

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9408, n9409, n9410, n9411, n9412, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10798;

  AND2_X1 U4988 ( .A1(n7221), .A2(n8915), .ZN(n8887) );
  INV_X2 U4990 ( .A(n6025), .ZN(n4927) );
  INV_X1 U4991 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5019) );
  INV_X2 U4993 ( .A(n10798), .ZN(n4925) );
  INV_X1 U4994 ( .A(n5968), .ZN(n5534) );
  NOR2_X1 U4995 ( .A1(n6632), .A2(n5284), .ZN(n5282) );
  INV_X1 U4996 ( .A(n8887), .ZN(n5034) );
  INV_X1 U4997 ( .A(n6881), .ZN(n6988) );
  INV_X1 U4998 ( .A(n7050), .ZN(n6015) );
  OR2_X1 U4999 ( .A1(n6279), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6296) );
  OAI22_X1 U5000 ( .A1(n9003), .A2(n9002), .B1(n9001), .B2(n9000), .ZN(n9030)
         );
  INV_X1 U5001 ( .A(n6401), .ZN(n8723) );
  INV_X1 U5002 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6232) );
  OR2_X1 U5004 ( .A1(n7448), .A2(n6981), .ZN(n10782) );
  OR3_X2 U5005 ( .A1(n8245), .A2(n8244), .A3(n8243), .ZN(n8246) );
  NOR2_X4 U5006 ( .A1(n6255), .A2(n6186), .ZN(n6302) );
  NAND2_X2 U5009 ( .A1(n6635), .A2(n8855), .ZN(n9167) );
  XNOR2_X2 U5010 ( .A(n5540), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5542) );
  NAND2_X2 U5011 ( .A1(n6200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6201) );
  NAND2_X2 U5012 ( .A1(n5049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6199) );
  XNOR2_X2 U5013 ( .A(n5708), .B(P1_IR_REG_30__SCAN_IN), .ZN(n10238) );
  NAND4_X1 U5014 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n8929)
         );
  NAND4_X1 U5015 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n6617)
         );
  INV_X4 U5016 ( .A(n6801), .ZN(n4926) );
  NAND4_X2 U5017 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n6724)
         );
  INV_X4 U5018 ( .A(n5836), .ZN(n5757) );
  OAI21_X1 U5019 ( .B1(n7036), .B2(n5582), .A(n5581), .ZN(n5584) );
  INV_X4 U5020 ( .A(n5701), .ZN(n7036) );
  AND3_X1 U5021 ( .A1(n6652), .A2(n6615), .A3(n6653), .ZN(n5338) );
  NAND2_X1 U5022 ( .A1(n9757), .A2(n5503), .ZN(n7004) );
  AND2_X1 U5023 ( .A1(n8276), .A2(n8275), .ZN(n10199) );
  NAND2_X1 U5024 ( .A1(n8232), .A2(n8231), .ZN(n9904) );
  NAND2_X1 U5025 ( .A1(n9019), .A2(n9020), .ZN(n9042) );
  XNOR2_X1 U5026 ( .A(n8268), .B(n8267), .ZN(n8529) );
  NAND2_X1 U5027 ( .A1(n5015), .A2(n5014), .ZN(n8684) );
  NAND2_X1 U5028 ( .A1(n6078), .A2(n6077), .ZN(n10013) );
  AND2_X1 U5029 ( .A1(n5512), .A2(n8863), .ZN(n5297) );
  AND2_X1 U5030 ( .A1(n5476), .A2(n5506), .ZN(n5007) );
  NAND2_X1 U5031 ( .A1(n5397), .A2(n5395), .ZN(n6120) );
  NAND2_X1 U5032 ( .A1(n6076), .A2(n5671), .ZN(n6089) );
  OAI21_X1 U5033 ( .B1(n6059), .B2(n6058), .A(n5665), .ZN(n6074) );
  NAND2_X1 U5034 ( .A1(n5105), .A2(n4987), .ZN(n7918) );
  OR2_X1 U5035 ( .A1(n7881), .A2(n7880), .ZN(n5105) );
  AND2_X1 U5036 ( .A1(n8463), .A2(n8333), .ZN(n7653) );
  NAND2_X1 U5037 ( .A1(n5848), .A2(n5847), .ZN(n7615) );
  OAI21_X1 U5038 ( .B1(n5424), .B2(n5256), .A(n5254), .ZN(n5918) );
  NAND2_X1 U5039 ( .A1(n5303), .A2(n5832), .ZN(n7691) );
  NAND2_X1 U5040 ( .A1(n5804), .A2(n5803), .ZN(n7418) );
  AND2_X1 U5041 ( .A1(n5119), .A2(n5118), .ZN(n10535) );
  OAI21_X1 U5042 ( .B1(n5779), .B2(n5778), .A(n5780), .ZN(n7046) );
  AOI21_X1 U5043 ( .B1(n7351), .B2(n7350), .A(n7349), .ZN(n10519) );
  AND2_X1 U5044 ( .A1(n5363), .A2(n4947), .ZN(n10628) );
  AND4_X1 U5045 ( .A1(n6220), .A2(n6219), .A3(n6221), .A4(n6222), .ZN(n8515)
         );
  NAND2_X1 U5046 ( .A1(n6364), .A2(n9717), .ZN(n6380) );
  INV_X1 U5047 ( .A(n6365), .ZN(n6364) );
  NAND2_X1 U5048 ( .A1(n7009), .A2(n7036), .ZN(n6274) );
  XNOR2_X1 U5049 ( .A(n6598), .B(n6597), .ZN(n8771) );
  INV_X1 U5050 ( .A(n8505), .ZN(n10692) );
  NAND2_X1 U5051 ( .A1(n7050), .A2(n5700), .ZN(n5997) );
  XNOR2_X1 U5052 ( .A(n6659), .B(n6658), .ZN(n8145) );
  NAND2_X1 U5053 ( .A1(n7387), .A2(n6951), .ZN(n8505) );
  CLKBUF_X1 U5054 ( .A(n6605), .Z(n8585) );
  CLKBUF_X3 U5055 ( .A(n6606), .Z(n9417) );
  OR2_X1 U5056 ( .A1(n6725), .A2(n6153), .ZN(n6154) );
  NAND2_X1 U5057 ( .A1(n5381), .A2(n5126), .ZN(n7050) );
  AND2_X1 U5058 ( .A1(n6153), .A2(n6951), .ZN(n10607) );
  CLKBUF_X1 U5059 ( .A(n6153), .Z(n9886) );
  XNOR2_X1 U5060 ( .A(n5538), .B(n5535), .ZN(n5574) );
  XNOR2_X1 U5061 ( .A(n5710), .B(n5707), .ZN(n5712) );
  XNOR2_X1 U5062 ( .A(n6656), .B(n6655), .ZN(n8516) );
  XNOR2_X1 U5063 ( .A(n5550), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U5064 ( .A1(n7025), .A2(n7026), .ZN(n7336) );
  NAND2_X2 U5065 ( .A1(n7036), .A2(P1_U3086), .ZN(n7238) );
  NAND4_X1 U5066 ( .A1(n5474), .A2(n4942), .A3(n5523), .A4(n5510), .ZN(n5709)
         );
  INV_X2 U5067 ( .A(n9409), .ZN(n9415) );
  OR2_X1 U5068 ( .A1(n5551), .A2(n10233), .ZN(n5998) );
  NOR2_X2 U5069 ( .A1(n7036), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10241) );
  AND2_X1 U5070 ( .A1(n5533), .A2(n5535), .ZN(n5474) );
  AND4_X1 U5071 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n5510)
         );
  AND2_X1 U5072 ( .A1(n6184), .A2(n6232), .ZN(n5482) );
  AND3_X1 U5073 ( .A1(n5018), .A2(n6594), .A3(n6195), .ZN(n5498) );
  AND4_X1 U5074 ( .A1(n5529), .A2(n5530), .A3(n5532), .A4(n5531), .ZN(n5533)
         );
  XNOR2_X1 U5075 ( .A(n6213), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7192) );
  INV_X1 U5076 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6427) );
  NOR2_X2 U5077 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5737) );
  NOR2_X1 U5078 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6187) );
  NOR2_X1 U5079 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6188) );
  NOR2_X1 U5080 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5473) );
  INV_X1 U5081 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5101) );
  INV_X1 U5082 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6271) );
  INV_X1 U5083 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6286) );
  INV_X1 U5084 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5020) );
  INV_X1 U5085 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6388) );
  INV_X1 U5086 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6415) );
  INV_X1 U5087 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5223) );
  NAND2_X1 U5088 ( .A1(n7226), .A2(n7362), .ZN(n7460) );
  INV_X2 U5089 ( .A(n5475), .ZN(n7226) );
  AOI21_X2 U5090 ( .B1(n8634), .B2(n8568), .A(n4985), .ZN(n8697) );
  NAND2_X2 U5091 ( .A1(n6605), .A2(n6606), .ZN(n7009) );
  XNOR2_X2 U5092 ( .A(n6199), .B(n6198), .ZN(n6204) );
  NAND2_X1 U5093 ( .A1(n5192), .A2(n8369), .ZN(n8370) );
  AND2_X1 U5094 ( .A1(n7971), .A2(n7970), .ZN(n7973) );
  OAI21_X1 U5095 ( .B1(n8549), .B2(n5489), .A(n5487), .ZN(n8555) );
  AOI21_X1 U5096 ( .B1(n5490), .B2(n5488), .A(n8553), .ZN(n5487) );
  INV_X1 U5097 ( .A(n5490), .ZN(n5489) );
  OR2_X1 U5098 ( .A1(n8733), .A2(n8721), .ZN(n8764) );
  NOR2_X1 U5099 ( .A1(n5361), .A2(n6247), .ZN(n5360) );
  AND2_X1 U5100 ( .A1(n5502), .A2(n6196), .ZN(n5501) );
  NOR2_X1 U5101 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5502) );
  INV_X1 U5102 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6208) );
  INV_X1 U5103 ( .A(n8443), .ZN(n5208) );
  BUF_X4 U5104 ( .A(n7036), .Z(n5700) );
  INV_X1 U5105 ( .A(n5725), .ZN(n5768) );
  AND2_X1 U5106 ( .A1(n5376), .A2(n5375), .ZN(n5522) );
  NOR2_X1 U5107 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5376) );
  NOR2_X1 U5108 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5375) );
  INV_X1 U5109 ( .A(n5255), .ZN(n5254) );
  OAI21_X1 U5110 ( .B1(n5423), .B2(n5256), .A(n5915), .ZN(n5255) );
  OR2_X1 U5111 ( .A1(n9099), .A2(n6547), .ZN(n5343) );
  NAND2_X1 U5112 ( .A1(n7009), .A2(n5701), .ZN(n6244) );
  INV_X1 U5113 ( .A(n5351), .ZN(n5103) );
  OR2_X1 U5114 ( .A1(n9928), .A2(n9941), .ZN(n6715) );
  INV_X1 U5115 ( .A(n5768), .ZN(n8230) );
  INV_X1 U5116 ( .A(n5997), .ZN(n8273) );
  MUX2_X1 U5117 ( .A(n8793), .B(n8792), .S(n8887), .Z(n8800) );
  OAI211_X1 U5118 ( .C1(n8815), .C2(n8805), .A(n8804), .B(n8811), .ZN(n8806)
         );
  NAND2_X1 U5119 ( .A1(n8857), .A2(n9184), .ZN(n5230) );
  NAND2_X1 U5120 ( .A1(n8358), .A2(n5194), .ZN(n5193) );
  NOR2_X1 U5121 ( .A1(n5196), .A2(n5195), .ZN(n5194) );
  NAND2_X1 U5122 ( .A1(n8365), .A2(n8400), .ZN(n5196) );
  NAND2_X1 U5123 ( .A1(n5211), .A2(n5213), .ZN(n8377) );
  AND2_X1 U5124 ( .A1(n9985), .A2(n5214), .ZN(n5213) );
  NAND2_X1 U5125 ( .A1(n4973), .A2(n8375), .ZN(n5214) );
  NAND2_X1 U5126 ( .A1(n5188), .A2(n8425), .ZN(n5187) );
  OAI21_X1 U5127 ( .B1(n8383), .B2(n8382), .A(n8400), .ZN(n5188) );
  INV_X1 U5128 ( .A(SI_25_), .ZN(n9657) );
  NAND2_X1 U5129 ( .A1(n9904), .A2(n9899), .ZN(n5009) );
  NAND2_X1 U5130 ( .A1(n6120), .A2(n6119), .ZN(n5688) );
  INV_X1 U5131 ( .A(SI_19_), .ZN(n9557) );
  INV_X1 U5132 ( .A(SI_8_), .ZN(n9683) );
  NAND2_X1 U5133 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  AND2_X1 U5134 ( .A1(n8546), .A2(n8620), .ZN(n8547) );
  OR2_X1 U5135 ( .A1(n8897), .A2(n8896), .ZN(n8902) );
  INV_X1 U5136 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6195) );
  OR2_X1 U5137 ( .A1(n9287), .A2(n9293), .ZN(n8883) );
  NAND2_X1 U5138 ( .A1(n9121), .A2(n5290), .ZN(n5289) );
  NOR2_X1 U5139 ( .A1(n8878), .A2(n5291), .ZN(n5290) );
  INV_X1 U5140 ( .A(n8874), .ZN(n5291) );
  NAND2_X1 U5141 ( .A1(n5287), .A2(n9259), .ZN(n5286) );
  OAI21_X1 U5142 ( .B1(n7069), .B2(P2_D_REG_0__SCAN_IN), .A(n7084), .ZN(n6668)
         );
  OR2_X1 U5143 ( .A1(n7069), .A2(n6679), .ZN(n6972) );
  AND2_X1 U5144 ( .A1(n5353), .A2(n5498), .ZN(n5351) );
  AND2_X1 U5145 ( .A1(n5497), .A2(n6689), .ZN(n5353) );
  NAND2_X2 U5146 ( .A1(n6730), .A2(n6154), .ZN(n6744) );
  AND2_X1 U5147 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  NOR2_X1 U5148 ( .A1(n9904), .A2(n8262), .ZN(n8434) );
  AOI21_X1 U5149 ( .B1(n8402), .B2(n8399), .A(n8398), .ZN(n8404) );
  AOI21_X1 U5150 ( .B1(n9904), .B2(n8400), .A(n8396), .ZN(n8397) );
  NAND2_X1 U5151 ( .A1(n9989), .A2(n4954), .ZN(n9969) );
  OR2_X1 U5152 ( .A1(n9471), .A2(n10111), .ZN(n8415) );
  OR2_X1 U5153 ( .A1(n10142), .A2(n10132), .ZN(n8367) );
  NAND2_X1 U5154 ( .A1(n10072), .A2(n8487), .ZN(n5083) );
  NOR2_X1 U5155 ( .A1(n8209), .A2(n8254), .ZN(n5079) );
  NAND2_X1 U5156 ( .A1(n7418), .A2(n7479), .ZN(n8318) );
  NAND2_X1 U5157 ( .A1(n8448), .A2(n8298), .ZN(n5159) );
  OAI21_X1 U5158 ( .B1(n8225), .B2(n9646), .A(n8224), .ZN(n8268) );
  OR2_X1 U5159 ( .A1(n8223), .A2(n8222), .ZN(n8224) );
  NAND2_X1 U5160 ( .A1(n6074), .A2(n6073), .ZN(n6076) );
  OAI21_X1 U5161 ( .B1(n5558), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5549) );
  AOI21_X1 U5162 ( .B1(n5418), .B2(n5420), .A(n6045), .ZN(n5415) );
  INV_X1 U5163 ( .A(n5812), .ZN(n5261) );
  NAND2_X1 U5164 ( .A1(n5266), .A2(n5843), .ZN(n5265) );
  NAND2_X1 U5165 ( .A1(n5481), .A2(n5480), .ZN(n5479) );
  AND2_X1 U5166 ( .A1(n7726), .A2(n7633), .ZN(n5500) );
  NAND2_X1 U5167 ( .A1(n8563), .A2(n8659), .ZN(n8631) );
  NAND2_X1 U5168 ( .A1(n5484), .A2(n8658), .ZN(n8563) );
  NOR2_X1 U5169 ( .A1(n8899), .A2(n8728), .ZN(n8729) );
  OR2_X1 U5170 ( .A1(n7698), .A2(n5120), .ZN(n5119) );
  NOR2_X1 U5171 ( .A1(n5121), .A2(n7709), .ZN(n5120) );
  INV_X1 U5172 ( .A(n7700), .ZN(n5121) );
  OAI21_X1 U5173 ( .B1(n9102), .B2(n6536), .A(n6535), .ZN(n9099) );
  AND2_X1 U5174 ( .A1(n5511), .A2(n8813), .ZN(n5293) );
  AND2_X1 U5175 ( .A1(n5356), .A2(n4946), .ZN(n5355) );
  NAND2_X1 U5177 ( .A1(n6616), .A2(n9340), .ZN(n5340) );
  INV_X1 U5178 ( .A(n8921), .ZN(n9293) );
  INV_X2 U5179 ( .A(n6274), .ZN(n6562) );
  INV_X1 U5180 ( .A(n9340), .ZN(n9323) );
  AND2_X1 U5181 ( .A1(n5501), .A2(n6208), .ZN(n5048) );
  XNOR2_X1 U5182 ( .A(n6209), .B(n6208), .ZN(n6605) );
  NAND2_X1 U5183 ( .A1(n6212), .A2(n6211), .ZN(n6606) );
  NAND2_X1 U5184 ( .A1(n5115), .A2(n5114), .ZN(n6212) );
  NAND2_X1 U5185 ( .A1(n6197), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5114) );
  AND2_X1 U5186 ( .A1(n8403), .A2(n9781), .ZN(n5414) );
  OAI21_X1 U5187 ( .B1(n8402), .B2(n8399), .A(n8401), .ZN(n5216) );
  AND2_X1 U5188 ( .A1(n8437), .A2(n8406), .ZN(n8407) );
  NAND2_X1 U5189 ( .A1(n6123), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U5190 ( .A1(n8393), .A2(n8392), .ZN(n8281) );
  OAI21_X1 U5191 ( .B1(n9963), .B2(n5167), .A(n5163), .ZN(n6151) );
  NAND2_X1 U5192 ( .A1(n9936), .A2(n6132), .ZN(n5167) );
  INV_X1 U5193 ( .A(n5164), .ZN(n5163) );
  OAI21_X1 U5194 ( .B1(n5310), .B2(n5165), .A(n6142), .ZN(n5164) );
  NOR2_X1 U5195 ( .A1(n6151), .A2(n6706), .ZN(n6701) );
  AOI21_X1 U5196 ( .B1(n9924), .B2(n5850), .A(n6150), .ZN(n9938) );
  OAI21_X1 U5197 ( .B1(n5370), .B2(n5177), .A(n5175), .ZN(n9967) );
  INV_X1 U5198 ( .A(n5387), .ZN(n5177) );
  AOI21_X1 U5199 ( .B1(n5176), .B2(n5387), .A(n4964), .ZN(n5175) );
  NOR2_X1 U5200 ( .A1(n4967), .A2(n5388), .ZN(n5387) );
  AND2_X1 U5201 ( .A1(n5372), .A2(n4945), .ZN(n5178) );
  INV_X1 U5202 ( .A(n7060), .ZN(n6022) );
  OR2_X1 U5203 ( .A1(n9431), .A2(n9771), .ZN(n8472) );
  NOR2_X1 U5204 ( .A1(n9431), .A2(n8035), .ZN(n8016) );
  NAND2_X1 U5205 ( .A1(n10690), .A2(n4950), .ZN(n7370) );
  NAND2_X1 U5206 ( .A1(n5558), .A2(n5557), .ZN(n6951) );
  NAND2_X1 U5207 ( .A1(n5127), .A2(n5128), .ZN(n5126) );
  NAND2_X1 U5208 ( .A1(n5697), .A2(n4932), .ZN(n5381) );
  NAND2_X1 U5209 ( .A1(n5382), .A2(n4966), .ZN(n5128) );
  NAND2_X1 U5210 ( .A1(n5703), .A2(n5702), .ZN(n9928) );
  NAND2_X1 U5211 ( .A1(n8583), .A2(n8273), .ZN(n5703) );
  NAND2_X1 U5212 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5710) );
  AOI21_X1 U5213 ( .B1(n5408), .B2(n5411), .A(n5407), .ZN(n5406) );
  NAND2_X1 U5214 ( .A1(n5918), .A2(n5408), .ZN(n5405) );
  INV_X1 U5215 ( .A(n5947), .ZN(n5407) );
  NAND2_X1 U5216 ( .A1(n5863), .A2(n5425), .ZN(n5424) );
  INV_X1 U5217 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5227) );
  NAND3_X1 U5218 ( .A1(n6688), .A2(n6687), .A3(n6686), .ZN(n7198) );
  NOR2_X1 U5219 ( .A1(n8587), .A2(n5486), .ZN(n5485) );
  INV_X1 U5220 ( .A(n8571), .ZN(n5486) );
  AND2_X1 U5221 ( .A1(n6176), .A2(n6175), .ZN(n9934) );
  XNOR2_X1 U5222 ( .A(n6705), .B(n8387), .ZN(n6167) );
  INV_X1 U5223 ( .A(n8452), .ZN(n5210) );
  INV_X1 U5224 ( .A(n8817), .ZN(n5040) );
  AOI21_X1 U5225 ( .B1(n5037), .B2(n8818), .A(n8887), .ZN(n5036) );
  INV_X1 U5226 ( .A(n8816), .ZN(n5037) );
  NAND2_X1 U5227 ( .A1(n9211), .A2(n8833), .ZN(n5235) );
  AOI211_X1 U5228 ( .C1(n8836), .C2(n4929), .A(n4974), .B(n5023), .ZN(n5021)
         );
  INV_X1 U5229 ( .A(n8355), .ZN(n5202) );
  NAND2_X1 U5230 ( .A1(n8363), .A2(n5198), .ZN(n5197) );
  AND2_X1 U5231 ( .A1(n8364), .A2(n8406), .ZN(n5198) );
  NAND2_X1 U5232 ( .A1(n8360), .A2(n5199), .ZN(n8361) );
  OR2_X1 U5233 ( .A1(n8858), .A2(n5229), .ZN(n5027) );
  MUX2_X1 U5234 ( .A(n8854), .B(n8853), .S(n8887), .Z(n8858) );
  AOI21_X1 U5235 ( .B1(n5231), .B2(n4959), .A(n5029), .ZN(n5028) );
  INV_X1 U5236 ( .A(n8865), .ZN(n5029) );
  NAND2_X1 U5237 ( .A1(n8872), .A2(n9118), .ZN(n5032) );
  NAND2_X1 U5238 ( .A1(n8379), .A2(n8421), .ZN(n5191) );
  INV_X1 U5239 ( .A(n8882), .ZN(n5238) );
  OAI21_X1 U5240 ( .B1(n5031), .B2(n5030), .A(n5240), .ZN(n5239) );
  NAND2_X1 U5241 ( .A1(n9107), .A2(n8876), .ZN(n5030) );
  AND2_X1 U5242 ( .A1(n8880), .A2(n8881), .ZN(n5240) );
  AOI21_X1 U5243 ( .B1(n8868), .B2(n9135), .A(n5032), .ZN(n5031) );
  INV_X1 U5244 ( .A(n5429), .ZN(n6574) );
  NAND2_X1 U5245 ( .A1(n5187), .A2(n5186), .ZN(n8389) );
  MUX2_X1 U5246 ( .A(n8428), .B(n8279), .S(n8400), .Z(n8280) );
  NAND2_X1 U5247 ( .A1(n5083), .A2(n5299), .ZN(n8418) );
  INV_X1 U5248 ( .A(n8406), .ZN(n8400) );
  NAND2_X1 U5249 ( .A1(n8290), .A2(n7554), .ZN(n8244) );
  NAND2_X1 U5250 ( .A1(n7885), .A2(n7886), .ZN(n7928) );
  OR2_X1 U5251 ( .A1(n6504), .A2(n6503), .ZN(n6506) );
  OR2_X1 U5252 ( .A1(n9348), .A2(n9183), .ZN(n8850) );
  NOR2_X1 U5253 ( .A1(n5280), .A2(n5038), .ZN(n5276) );
  OAI21_X1 U5254 ( .B1(n8819), .B2(n5280), .A(n8824), .ZN(n5279) );
  AOI21_X1 U5255 ( .B1(n5332), .B2(n5330), .A(n5329), .ZN(n5328) );
  INV_X1 U5256 ( .A(n5336), .ZN(n5330) );
  NOR2_X1 U5257 ( .A1(n7838), .A2(n5296), .ZN(n5295) );
  INV_X1 U5258 ( .A(n8795), .ZN(n5296) );
  OR2_X1 U5259 ( .A1(n7775), .A2(n8926), .ZN(n5334) );
  NAND2_X1 U5260 ( .A1(n6278), .A2(n6277), .ZN(n5335) );
  INV_X1 U5261 ( .A(n8771), .ZN(n7221) );
  INV_X1 U5262 ( .A(n5350), .ZN(n5349) );
  NOR2_X1 U5263 ( .A1(n5347), .A2(n5350), .ZN(n6663) );
  NAND2_X1 U5264 ( .A1(n5351), .A2(n5348), .ZN(n5347) );
  INV_X1 U5265 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5348) );
  INV_X1 U5266 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6689) );
  INV_X1 U5267 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5497) );
  INV_X1 U5268 ( .A(n6849), .ZN(n5448) );
  AND2_X1 U5269 ( .A1(n5446), .A2(n6852), .ZN(n5445) );
  NAND2_X1 U5270 ( .A1(n6849), .A2(n5447), .ZN(n5446) );
  AND2_X1 U5271 ( .A1(n5440), .A2(n5509), .ZN(n5052) );
  NOR2_X1 U5272 ( .A1(n9968), .A2(n9962), .ZN(n9940) );
  OR2_X1 U5273 ( .A1(n9947), .A2(n9926), .ZN(n8426) );
  NOR2_X1 U5274 ( .A1(n9995), .A2(n5144), .ZN(n5143) );
  INV_X1 U5275 ( .A(n5145), .ZN(n5144) );
  NOR2_X1 U5276 ( .A1(n4968), .A2(n5172), .ZN(n5171) );
  AND2_X1 U5277 ( .A1(n6011), .A2(n5173), .ZN(n5172) );
  INV_X1 U5278 ( .A(n5991), .ZN(n5173) );
  INV_X1 U5279 ( .A(n8256), .ZN(n5169) );
  OR2_X1 U5280 ( .A1(n10153), .A2(n10088), .ZN(n8256) );
  NOR2_X1 U5281 ( .A1(n5149), .A2(n10153), .ZN(n5148) );
  INV_X1 U5282 ( .A(n5150), .ZN(n5149) );
  OR2_X1 U5283 ( .A1(n10166), .A2(n10156), .ZN(n8359) );
  NOR2_X1 U5284 ( .A1(n8117), .A2(n5153), .ZN(n5152) );
  INV_X1 U5285 ( .A(n5154), .ZN(n5153) );
  INV_X1 U5286 ( .A(n8345), .ZN(n8471) );
  NAND2_X1 U5287 ( .A1(n7691), .A2(n7610), .ZN(n8240) );
  INV_X1 U5288 ( .A(n10628), .ZN(n6752) );
  INV_X1 U5289 ( .A(n5383), .ZN(n5382) );
  OAI21_X1 U5290 ( .B1(n5696), .B2(P1_IR_REG_28__SCAN_IN), .A(n5698), .ZN(
        n5383) );
  NAND2_X1 U5291 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(n5699), .ZN(n5698) );
  OR2_X1 U5292 ( .A1(n5574), .A2(P1_B_REG_SCAN_IN), .ZN(n5543) );
  AOI21_X1 U5293 ( .B1(n5398), .B2(n5400), .A(n5396), .ZN(n5395) );
  NAND2_X1 U5294 ( .A1(n6089), .A2(n5398), .ZN(n5397) );
  INV_X1 U5295 ( .A(n5682), .ZN(n5396) );
  INV_X1 U5296 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U5297 ( .A1(n5130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U5298 ( .A1(n5534), .A2(n5474), .ZN(n5130) );
  INV_X1 U5299 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5548) );
  INV_X1 U5300 ( .A(n5419), .ZN(n5418) );
  OAI21_X1 U5301 ( .B1(n5421), .B2(n5420), .A(n5656), .ZN(n5419) );
  AOI21_X1 U5302 ( .B1(n5932), .B2(n5410), .A(n5409), .ZN(n5408) );
  INV_X1 U5303 ( .A(n5635), .ZN(n5409) );
  INV_X1 U5304 ( .A(n5631), .ZN(n5410) );
  NOR2_X1 U5305 ( .A1(n5894), .A2(n5428), .ZN(n5423) );
  INV_X1 U5306 ( .A(n5608), .ZN(n5403) );
  AND2_X1 U5307 ( .A1(n5301), .A2(n5300), .ZN(n5602) );
  OR2_X1 U5308 ( .A1(n5700), .A2(n5302), .ZN(n5301) );
  NAND2_X1 U5309 ( .A1(n5700), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U5310 ( .A1(n5595), .A2(n5012), .ZN(n5011) );
  NAND2_X1 U5311 ( .A1(n5700), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5595) );
  OR2_X1 U5312 ( .A1(n5700), .A2(n5596), .ZN(n5012) );
  NAND2_X1 U5313 ( .A1(n8558), .A2(n8559), .ZN(n5484) );
  NAND2_X1 U5314 ( .A1(n8684), .A2(n8683), .ZN(n8611) );
  XNOR2_X1 U5315 ( .A(n9186), .B(n9333), .ZN(n8740) );
  OR2_X1 U5316 ( .A1(n6316), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U5317 ( .A1(n8631), .A2(n8632), .ZN(n8634) );
  INV_X1 U5318 ( .A(n8555), .ZN(n8557) );
  NAND2_X1 U5319 ( .A1(n5016), .A2(n4988), .ZN(n8539) );
  OAI21_X1 U5320 ( .B1(n5006), .B2(n5003), .A(n4936), .ZN(n5496) );
  INV_X1 U5321 ( .A(n8192), .ZN(n5003) );
  NAND2_X1 U5322 ( .A1(n5002), .A2(n8192), .ZN(n5001) );
  AND2_X1 U5323 ( .A1(n8905), .A2(n8906), .ZN(n5245) );
  AND2_X1 U5324 ( .A1(n5273), .A2(n8736), .ZN(n5272) );
  OR2_X1 U5325 ( .A1(n8734), .A2(n8906), .ZN(n5273) );
  AOI211_X1 U5326 ( .C1(n8737), .C2(n8733), .A(n8771), .B(n8908), .ZN(n8734)
         );
  AND2_X1 U5327 ( .A1(n5241), .A2(n8909), .ZN(n5043) );
  AND2_X1 U5328 ( .A1(n5249), .A2(n5242), .ZN(n5241) );
  NAND2_X1 U5329 ( .A1(n5248), .A2(n5243), .ZN(n5242) );
  OR2_X1 U5330 ( .A1(n8900), .A2(n5244), .ZN(n5044) );
  NAND2_X1 U5331 ( .A1(n5248), .A2(n8906), .ZN(n5244) );
  INV_X1 U5332 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6191) );
  NOR2_X1 U5333 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5018) );
  OR2_X1 U5334 ( .A1(n6261), .A2(n6205), .ZN(n5268) );
  INV_X1 U5335 ( .A(n7572), .ZN(n6202) );
  OAI21_X1 U5336 ( .B1(n9417), .B2(n6205), .A(n5113), .ZN(n5112) );
  NAND2_X1 U5337 ( .A1(n9417), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5113) );
  INV_X1 U5338 ( .A(n10538), .ZN(n5118) );
  NAND2_X1 U5339 ( .A1(n10554), .A2(n10555), .ZN(n10553) );
  NAND2_X1 U5340 ( .A1(n10553), .A2(n5394), .ZN(n7706) );
  NAND2_X1 U5341 ( .A1(n7707), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U5342 ( .A1(n7882), .A2(n7883), .ZN(n7919) );
  NAND2_X1 U5343 ( .A1(n8081), .A2(n8082), .ZN(n8935) );
  NAND2_X1 U5344 ( .A1(n8935), .A2(n5221), .ZN(n8956) );
  OR2_X1 U5345 ( .A1(n8939), .A2(n6363), .ZN(n5221) );
  AND2_X1 U5346 ( .A1(n5109), .A2(n5108), .ZN(n10574) );
  NAND2_X1 U5347 ( .A1(n8952), .A2(n8951), .ZN(n5108) );
  NAND2_X1 U5348 ( .A1(n8954), .A2(n8953), .ZN(n5109) );
  NAND2_X1 U5349 ( .A1(n9013), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9019) );
  OR2_X1 U5350 ( .A1(n9281), .A2(n9285), .ZN(n6645) );
  OR2_X1 U5351 ( .A1(n9295), .A2(n8570), .ZN(n9081) );
  NAND2_X1 U5352 ( .A1(n5289), .A2(n8739), .ZN(n9092) );
  INV_X1 U5353 ( .A(n6249), .ZN(n6585) );
  INV_X1 U5354 ( .A(n8765), .ZN(n9107) );
  NAND2_X1 U5355 ( .A1(n6512), .A2(n9640), .ZN(n6527) );
  INV_X1 U5356 ( .A(n6513), .ZN(n6512) );
  OR2_X1 U5357 ( .A1(n9385), .A2(n9315), .ZN(n8863) );
  NAND2_X1 U5358 ( .A1(n5315), .A2(n5317), .ZN(n9126) );
  AOI21_X1 U5359 ( .B1(n9168), .B2(n5318), .A(n4992), .ZN(n5317) );
  NAND2_X1 U5360 ( .A1(n5324), .A2(n9203), .ZN(n5323) );
  INV_X1 U5361 ( .A(n6453), .ZN(n5322) );
  NAND2_X1 U5362 ( .A1(n6631), .A2(n5285), .ZN(n5283) );
  NAND2_X1 U5363 ( .A1(n6633), .A2(n5286), .ZN(n5285) );
  NAND2_X1 U5364 ( .A1(n6376), .A2(n6375), .ZN(n8828) );
  INV_X1 U5365 ( .A(n8821), .ZN(n5280) );
  AND2_X1 U5366 ( .A1(n8818), .A2(n8809), .ZN(n8754) );
  OR2_X1 U5367 ( .A1(n7950), .A2(n7975), .ZN(n8813) );
  NAND2_X1 U5368 ( .A1(n6622), .A2(n6621), .ZN(n5294) );
  NAND2_X1 U5369 ( .A1(n6330), .A2(n6329), .ZN(n6343) );
  INV_X1 U5370 ( .A(n6331), .ZN(n6330) );
  NOR2_X1 U5371 ( .A1(n6292), .A2(n5337), .ZN(n5336) );
  INV_X1 U5372 ( .A(n6277), .ZN(n5337) );
  AND2_X1 U5373 ( .A1(n8795), .A2(n8794), .ZN(n8746) );
  NOR2_X1 U5374 ( .A1(n7587), .A2(n7513), .ZN(n5357) );
  AND2_X1 U5375 ( .A1(n8785), .A2(n8781), .ZN(n8742) );
  NAND2_X1 U5376 ( .A1(n6584), .A2(n6583), .ZN(n8726) );
  NAND2_X1 U5377 ( .A1(n6511), .A2(n6510), .ZN(n8873) );
  INV_X1 U5378 ( .A(n9314), .ZN(n9334) );
  INV_X1 U5379 ( .A(n7210), .ZN(n7213) );
  OR2_X1 U5380 ( .A1(n7230), .A2(n5034), .ZN(n9314) );
  NAND2_X1 U5381 ( .A1(n8771), .A2(n7908), .ZN(n10785) );
  NAND2_X1 U5382 ( .A1(n7230), .A2(n8887), .ZN(n9316) );
  NAND2_X1 U5383 ( .A1(n6604), .A2(n6680), .ZN(n9340) );
  NAND2_X1 U5384 ( .A1(n6666), .A2(n6688), .ZN(n7069) );
  XNOR2_X1 U5385 ( .A(n8516), .B(P2_B_REG_SCAN_IN), .ZN(n6660) );
  AND2_X1 U5386 ( .A1(n7198), .A2(n7086), .ZN(n7206) );
  OR2_X1 U5387 ( .A1(n6654), .A2(n9406), .ZN(n6656) );
  INV_X1 U5388 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U5389 ( .A1(n6596), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6600) );
  INV_X1 U5390 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U5391 ( .A1(n6600), .A2(n6599), .ZN(n6602) );
  INV_X1 U5392 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6309) );
  OR2_X1 U5393 ( .A1(n6079), .A2(n9438), .ZN(n6095) );
  NAND2_X1 U5394 ( .A1(n5455), .A2(n6922), .ZN(n5453) );
  NAND2_X1 U5395 ( .A1(n5064), .A2(n5454), .ZN(n5451) );
  NAND2_X1 U5396 ( .A1(n6922), .A2(n9496), .ZN(n5452) );
  INV_X1 U5397 ( .A(n6738), .ZN(n6881) );
  NAND2_X1 U5398 ( .A1(n5461), .A2(n5456), .ZN(n5455) );
  NAND2_X1 U5399 ( .A1(n5457), .A2(n9496), .ZN(n5456) );
  INV_X1 U5400 ( .A(n9495), .ZN(n5461) );
  INV_X1 U5401 ( .A(n9435), .ZN(n5457) );
  INV_X1 U5402 ( .A(n7244), .ZN(n5062) );
  OR2_X1 U5403 ( .A1(n5834), .A2(n7687), .ZN(n5852) );
  NAND2_X1 U5404 ( .A1(n9525), .A2(n9524), .ZN(n5454) );
  INV_X1 U5405 ( .A(n7292), .ZN(n5468) );
  INV_X1 U5406 ( .A(n6771), .ZN(n5465) );
  NAND2_X1 U5407 ( .A1(n5207), .A2(n5208), .ZN(n5206) );
  AND3_X1 U5408 ( .A1(n8277), .A2(n4928), .A3(n8499), .ZN(n8439) );
  NOR2_X1 U5409 ( .A1(n10376), .A2(n10375), .ZN(n10374) );
  NOR2_X1 U5410 ( .A1(n10374), .A2(n5090), .ZN(n10387) );
  AND2_X1 U5411 ( .A1(n10378), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5090) );
  OR2_X1 U5412 ( .A1(n10387), .A2(n10386), .ZN(n5089) );
  XNOR2_X1 U5413 ( .A(n9858), .B(n9857), .ZN(n10461) );
  NOR2_X1 U5414 ( .A1(n10440), .A2(n5091), .ZN(n9858) );
  AND2_X1 U5415 ( .A1(n10439), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5091) );
  NOR2_X1 U5416 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  AND2_X1 U5417 ( .A1(n6146), .A2(n9914), .ZN(n9924) );
  NAND2_X1 U5418 ( .A1(n8278), .A2(n8420), .ZN(n8387) );
  OAI22_X1 U5419 ( .A1(n9967), .A2(n6118), .B1(n10111), .B2(n5142), .ZN(n9963)
         );
  NAND2_X1 U5420 ( .A1(n9989), .A2(n8412), .ZN(n9971) );
  AND2_X1 U5421 ( .A1(n8412), .A2(n8409), .ZN(n9985) );
  AOI21_X1 U5422 ( .B1(n6072), .B2(n5373), .A(n4965), .ZN(n5372) );
  INV_X1 U5423 ( .A(n6057), .ZN(n5373) );
  NOR2_X1 U5424 ( .A1(n10025), .A2(n10033), .ZN(n5371) );
  OR2_X1 U5425 ( .A1(n10148), .A2(n10139), .ZN(n10042) );
  OR2_X1 U5426 ( .A1(n6035), .A2(n9507), .ZN(n6049) );
  NAND2_X1 U5427 ( .A1(n6164), .A2(n8482), .ZN(n10072) );
  NAND2_X1 U5428 ( .A1(n5074), .A2(n5072), .ZN(n6164) );
  AOI21_X1 U5429 ( .B1(n5075), .B2(n5076), .A(n5073), .ZN(n5072) );
  NAND2_X1 U5430 ( .A1(n8208), .A2(n5991), .ZN(n10077) );
  AND2_X1 U5431 ( .A1(n8359), .A2(n8233), .ZN(n8354) );
  NAND2_X1 U5432 ( .A1(n9780), .A2(n9426), .ZN(n5367) );
  NAND2_X1 U5433 ( .A1(n8024), .A2(n5368), .ZN(n5366) );
  NOR2_X1 U5434 ( .A1(n5965), .A2(n5369), .ZN(n5368) );
  INV_X1 U5435 ( .A(n5946), .ZN(n5369) );
  NAND2_X1 U5436 ( .A1(n8132), .A2(n8141), .ZN(n8131) );
  AND4_X1 U5437 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n9427)
         );
  AND2_X1 U5438 ( .A1(n8342), .A2(n8338), .ZN(n7801) );
  NAND2_X1 U5439 ( .A1(n5305), .A2(n7651), .ZN(n5304) );
  AND2_X1 U5440 ( .A1(n5306), .A2(n8333), .ZN(n5305) );
  NAND2_X1 U5441 ( .A1(n5883), .A2(n5882), .ZN(n7672) );
  OAI21_X1 U5442 ( .B1(n5070), .B2(n8464), .A(n8292), .ZN(n7652) );
  NOR2_X1 U5443 ( .A1(n7402), .A2(n8461), .ZN(n5070) );
  INV_X1 U5444 ( .A(n10703), .ZN(n10089) );
  OR2_X1 U5445 ( .A1(n7691), .A2(n7596), .ZN(n7597) );
  NAND2_X1 U5446 ( .A1(n5158), .A2(n5797), .ZN(n7369) );
  AND2_X1 U5447 ( .A1(n5772), .A2(n5771), .ZN(n10689) );
  NOR2_X1 U5448 ( .A1(n10661), .A2(n10662), .ZN(n10690) );
  OR2_X1 U5449 ( .A1(n10626), .A2(n6752), .ZN(n10661) );
  OR2_X1 U5450 ( .A1(n8436), .A2(n10245), .ZN(n10703) );
  NAND2_X1 U5451 ( .A1(n8529), .A2(n8273), .ZN(n8232) );
  INV_X1 U5452 ( .A(n10659), .ZN(n10698) );
  XNOR2_X1 U5453 ( .A(n8272), .B(n8271), .ZN(n9405) );
  OAI21_X1 U5454 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8272) );
  XNOR2_X1 U5455 ( .A(n5693), .B(n6576), .ZN(n8583) );
  NAND2_X1 U5456 ( .A1(n6575), .A2(n5429), .ZN(n5693) );
  NAND2_X1 U5457 ( .A1(n5697), .A2(n5696), .ZN(n6173) );
  XNOR2_X1 U5458 ( .A(n6134), .B(SI_27_), .ZN(n9414) );
  NAND2_X1 U5459 ( .A1(n6575), .A2(n6133), .ZN(n6134) );
  NAND2_X1 U5460 ( .A1(n5697), .A2(n5695), .ZN(n5539) );
  OAI21_X1 U5461 ( .B1(n6089), .B2(n5400), .A(n5398), .ZN(n6105) );
  NAND2_X1 U5462 ( .A1(n6091), .A2(n5677), .ZN(n6103) );
  NAND2_X1 U5463 ( .A1(n5526), .A2(n5525), .ZN(n5558) );
  NAND2_X1 U5464 ( .A1(n5417), .A2(n5655), .ZN(n6032) );
  XNOR2_X1 U5465 ( .A(n5554), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6153) );
  INV_X1 U5466 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5065) );
  AND2_X1 U5467 ( .A1(n5640), .A2(n5639), .ZN(n5947) );
  INV_X1 U5468 ( .A(n5408), .ZN(n5252) );
  NAND2_X1 U5469 ( .A1(n5424), .A2(n5253), .ZN(n5250) );
  AND2_X1 U5470 ( .A1(n5631), .A2(n5630), .ZN(n5915) );
  NAND2_X1 U5471 ( .A1(n5259), .A2(n5257), .ZN(n5859) );
  NAND2_X1 U5472 ( .A1(n5265), .A2(n5258), .ZN(n5257) );
  INV_X1 U5473 ( .A(n5263), .ZN(n5258) );
  NAND2_X1 U5474 ( .A1(n5262), .A2(n5616), .ZN(n5844) );
  NAND2_X1 U5475 ( .A1(n5815), .A2(n5266), .ZN(n5262) );
  NAND2_X1 U5476 ( .A1(n5815), .A2(n5613), .ZN(n5829) );
  OR2_X1 U5477 ( .A1(n5602), .A2(n5601), .ZN(n5604) );
  AND2_X1 U5478 ( .A1(n5608), .A2(n5607), .ZN(n5798) );
  NAND2_X1 U5479 ( .A1(n5767), .A2(n5600), .ZN(n5779) );
  NAND2_X1 U5480 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NOR2_X1 U5481 ( .A1(n10233), .A2(n5101), .ZN(n5100) );
  NAND2_X1 U5482 ( .A1(n5737), .A2(n5473), .ZN(n5102) );
  AND2_X1 U5483 ( .A1(n4995), .A2(n5479), .ZN(n8057) );
  INV_X1 U5484 ( .A(n7304), .ZN(n7305) );
  INV_X1 U5485 ( .A(n9219), .ZN(n9183) );
  OR2_X1 U5486 ( .A1(n8572), .A2(n9293), .ZN(n8573) );
  INV_X1 U5487 ( .A(n9261), .ZN(n8644) );
  NAND2_X1 U5488 ( .A1(n7743), .A2(n7742), .ZN(n7971) );
  INV_X1 U5489 ( .A(n8929), .ZN(n7513) );
  OAI211_X1 U5490 ( .C1(n7009), .C2(n7350), .A(n6234), .B(n6233), .ZN(n7467)
         );
  INV_X1 U5491 ( .A(n9292), .ZN(n8922) );
  INV_X1 U5492 ( .A(n9133), .ZN(n9300) );
  NAND4_X1 U5493 ( .A1(n6270), .A2(n6269), .A3(n6268), .A4(n6267), .ZN(n8927)
         );
  XNOR2_X1 U5494 ( .A(n5112), .B(n5110), .ZN(n7189) );
  NOR2_X1 U5495 ( .A1(n7354), .A2(n7355), .ZN(n7698) );
  NAND2_X1 U5496 ( .A1(n10550), .A2(n4991), .ZN(n7812) );
  XNOR2_X1 U5497 ( .A(n7919), .B(n5389), .ZN(n7922) );
  NAND2_X1 U5498 ( .A1(n7925), .A2(n7924), .ZN(n7985) );
  XNOR2_X1 U5499 ( .A(n8070), .B(n5391), .ZN(n8074) );
  AOI22_X1 U5500 ( .A1(n8069), .A2(n8068), .B1(n8067), .B2(n8072), .ZN(n8934)
         );
  NOR2_X1 U5501 ( .A1(n9050), .A2(n9033), .ZN(n9034) );
  NOR2_X1 U5502 ( .A1(n7015), .A2(n7014), .ZN(n10566) );
  AOI21_X1 U5503 ( .B1(n9038), .B2(n10579), .A(n5124), .ZN(n5123) );
  OAI21_X1 U5504 ( .B1(n9039), .B2(n9064), .A(n5125), .ZN(n5124) );
  AOI21_X1 U5505 ( .B1(n10564), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9036), .ZN(
        n5125) );
  INV_X1 U5506 ( .A(n5340), .ZN(n5339) );
  NAND2_X1 U5507 ( .A1(n5343), .A2(n6548), .ZN(n9088) );
  INV_X1 U5508 ( .A(n9325), .ZN(n9182) );
  NAND2_X1 U5509 ( .A1(n6406), .A2(n6405), .ZN(n9254) );
  OR2_X1 U5510 ( .A1(n7289), .A2(n6401), .ZN(n6406) );
  AND2_X1 U5511 ( .A1(n6392), .A2(n6391), .ZN(n9266) );
  OR2_X1 U5512 ( .A1(n7241), .A2(n6244), .ZN(n6392) );
  NAND2_X1 U5513 ( .A1(n6362), .A2(n6361), .ZN(n10766) );
  AND4_X1 U5514 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(n7761)
         );
  INV_X1 U5515 ( .A(n9274), .ZN(n9192) );
  INV_X1 U5516 ( .A(n5314), .ZN(n7362) );
  INV_X2 U5517 ( .A(n10782), .ZN(n10791) );
  NAND2_X1 U5518 ( .A1(n5338), .A2(n5340), .ZN(n6982) );
  AND2_X1 U5519 ( .A1(n5048), .A2(n5047), .ZN(n5046) );
  NAND2_X1 U5520 ( .A1(n9757), .A2(n6946), .ZN(n5435) );
  NAND2_X1 U5521 ( .A1(n5938), .A2(n5937), .ZN(n9431) );
  OR2_X1 U5522 ( .A1(n7241), .A2(n5997), .ZN(n5938) );
  AND2_X1 U5523 ( .A1(n6010), .A2(n6009), .ZN(n10074) );
  NAND2_X1 U5524 ( .A1(n6048), .A2(n6047), .ZN(n10142) );
  NAND2_X1 U5525 ( .A1(n5971), .A2(n5970), .ZN(n10171) );
  NAND2_X1 U5526 ( .A1(n6000), .A2(n5999), .ZN(n10159) );
  INV_X1 U5527 ( .A(n9779), .ZN(n9546) );
  NAND2_X1 U5528 ( .A1(n6966), .A2(n10245), .ZN(n9772) );
  AND3_X1 U5529 ( .A1(n5978), .A2(n5977), .A3(n5976), .ZN(n10163) );
  AND2_X1 U5530 ( .A1(n6964), .A2(n6950), .ZN(n9768) );
  INV_X1 U5531 ( .A(n10111), .ZN(n9501) );
  INV_X1 U5532 ( .A(n9991), .ZN(n10027) );
  INV_X1 U5533 ( .A(n10074), .ZN(n9786) );
  OR2_X1 U5534 ( .A1(n5758), .A2(n9817), .ZN(n5735) );
  OR2_X1 U5535 ( .A1(n5758), .A2(n7158), .ZN(n5721) );
  OR2_X1 U5536 ( .A1(n5759), .A2(n5713), .ZN(n5714) );
  NAND2_X1 U5537 ( .A1(n5757), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5716) );
  OR2_X1 U5538 ( .A1(n5758), .A2(n10605), .ZN(n5715) );
  NAND2_X1 U5539 ( .A1(n5097), .A2(n5096), .ZN(n5095) );
  AOI21_X1 U5540 ( .B1(n10585), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n10478), .ZN(
        n5096) );
  NAND2_X1 U5541 ( .A1(n10595), .A2(n10477), .ZN(n5097) );
  OR2_X1 U5542 ( .A1(n10369), .A2(n8506), .ZN(n10496) );
  OR2_X1 U5543 ( .A1(n6714), .A2(n6715), .ZN(n9903) );
  OAI21_X1 U5544 ( .B1(n9903), .B2(n5132), .A(n5131), .ZN(n5137) );
  NAND2_X1 U5545 ( .A1(n10199), .A2(n8399), .ZN(n5132) );
  INV_X1 U5546 ( .A(n5141), .ZN(n5131) );
  AND2_X1 U5547 ( .A1(n9928), .A2(n9782), .ZN(n6700) );
  AND2_X1 U5548 ( .A1(n10707), .A2(n7387), .ZN(n10674) );
  NAND2_X1 U5549 ( .A1(n9934), .A2(n5080), .ZN(n6182) );
  INV_X1 U5550 ( .A(n5081), .ZN(n5080) );
  OAI21_X1 U5551 ( .B1(n9923), .B2(n10183), .A(n6180), .ZN(n5081) );
  NAND4_X1 U5552 ( .A1(n5084), .A2(n4942), .A3(n5510), .A4(n5523), .ZN(n10234)
         );
  AND2_X1 U5553 ( .A1(n5533), .A2(n5085), .ZN(n5084) );
  AND2_X1 U5554 ( .A1(n5535), .A2(n5707), .ZN(n5085) );
  NOR2_X2 U5555 ( .A1(n7198), .A2(n7011), .ZN(P2_U3893) );
  OAI21_X1 U5556 ( .B1(n8766), .B2(n8775), .A(n8774), .ZN(n8767) );
  MUX2_X1 U5557 ( .A(n8803), .B(n8798), .S(n8887), .Z(n8801) );
  AND2_X1 U5558 ( .A1(n8813), .A2(n8797), .ZN(n8798) );
  NAND2_X1 U5559 ( .A1(n5035), .A2(n5033), .ZN(n5041) );
  OAI21_X1 U5560 ( .B1(n5039), .B2(n5038), .A(n5036), .ZN(n5042) );
  AOI21_X1 U5561 ( .B1(n4951), .B2(n8809), .A(n5034), .ZN(n5033) );
  NAND2_X1 U5562 ( .A1(n5233), .A2(n5034), .ZN(n5232) );
  NAND2_X1 U5563 ( .A1(n5235), .A2(n8887), .ZN(n5234) );
  NAND2_X1 U5564 ( .A1(n8837), .A2(n9266), .ZN(n5233) );
  NAND2_X1 U5565 ( .A1(n8838), .A2(n9212), .ZN(n5023) );
  NAND2_X1 U5566 ( .A1(n5022), .A2(n8843), .ZN(n8849) );
  NAND2_X1 U5567 ( .A1(n5022), .A2(n4963), .ZN(n8848) );
  INV_X1 U5568 ( .A(n8844), .ZN(n5024) );
  NAND2_X1 U5569 ( .A1(n5201), .A2(n5200), .ZN(n8360) );
  AND2_X1 U5570 ( .A1(n8354), .A2(n8353), .ZN(n5200) );
  NAND2_X1 U5571 ( .A1(n5203), .A2(n5202), .ZN(n5201) );
  AND2_X1 U5572 ( .A1(n8482), .A2(n8359), .ZN(n5199) );
  INV_X1 U5573 ( .A(n8857), .ZN(n5228) );
  INV_X1 U5574 ( .A(n9129), .ZN(n5026) );
  NOR2_X1 U5575 ( .A1(n5215), .A2(n4956), .ZN(n5212) );
  INV_X1 U5576 ( .A(n8375), .ZN(n5215) );
  NAND2_X1 U5577 ( .A1(n8384), .A2(n8400), .ZN(n5186) );
  NAND2_X1 U5578 ( .A1(n8380), .A2(n8406), .ZN(n5189) );
  NAND2_X1 U5579 ( .A1(n5191), .A2(n8400), .ZN(n5190) );
  INV_X1 U5580 ( .A(n8621), .ZN(n5488) );
  NAND2_X1 U5581 ( .A1(n8886), .A2(n8887), .ZN(n8889) );
  NAND2_X1 U5582 ( .A1(n5236), .A2(n8885), .ZN(n8890) );
  NAND2_X1 U5583 ( .A1(n5239), .A2(n5237), .ZN(n5236) );
  NOR2_X1 U5584 ( .A1(n9089), .A2(n5238), .ZN(n5237) );
  INV_X1 U5585 ( .A(n9514), .ZN(n5447) );
  INV_X1 U5586 ( .A(n8255), .ZN(n5385) );
  INV_X1 U5587 ( .A(n6012), .ZN(n5384) );
  NOR2_X1 U5588 ( .A1(n5986), .A2(n5985), .ZN(n6001) );
  AND2_X1 U5589 ( .A1(n7958), .A2(n9791), .ZN(n8345) );
  NOR2_X1 U5590 ( .A1(n10135), .A2(n10013), .ZN(n5145) );
  NAND3_X1 U5591 ( .A1(n6581), .A2(n6580), .A3(n6579), .ZN(n8223) );
  INV_X1 U5592 ( .A(SI_28_), .ZN(n9571) );
  NOR2_X1 U5593 ( .A1(n6013), .A2(n5422), .ZN(n5421) );
  INV_X1 U5594 ( .A(n5652), .ZN(n5422) );
  OAI211_X1 U5595 ( .C1(n5579), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5580), .ZN(n5586) );
  NAND2_X1 U5596 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  INV_X1 U5597 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5578) );
  INV_X1 U5598 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9710) );
  AND2_X1 U5599 ( .A1(n8055), .A2(n7747), .ZN(n5478) );
  INV_X1 U5600 ( .A(n5004), .ZN(n5002) );
  NOR2_X1 U5601 ( .A1(n8598), .A2(n5494), .ZN(n5493) );
  INV_X1 U5602 ( .A(n8532), .ZN(n5494) );
  NOR2_X1 U5603 ( .A1(n8898), .A2(n5247), .ZN(n5243) );
  NAND2_X1 U5604 ( .A1(n8907), .A2(n5247), .ZN(n5249) );
  AOI21_X1 U5605 ( .B1(n8898), .B2(n8899), .A(n8887), .ZN(n5248) );
  INV_X1 U5606 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U5607 ( .A1(n7703), .A2(n4953), .ZN(n7704) );
  NAND2_X1 U5608 ( .A1(n7708), .A2(n4957), .ZN(n7710) );
  NAND2_X1 U5609 ( .A1(n10545), .A2(n5218), .ZN(n7822) );
  NAND2_X1 U5610 ( .A1(n7707), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U5611 ( .A1(n10570), .A2(n8959), .ZN(n8990) );
  INV_X1 U5612 ( .A(n6548), .ZN(n5342) );
  AND2_X1 U5613 ( .A1(n5517), .A2(n9081), .ZN(n8881) );
  OR2_X1 U5614 ( .A1(n6493), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6495) );
  NOR2_X1 U5615 ( .A1(n9166), .A2(n5321), .ZN(n5316) );
  INV_X1 U5616 ( .A(n5323), .ZN(n5318) );
  NAND2_X1 U5617 ( .A1(n6458), .A2(n9708), .ZN(n6469) );
  INV_X1 U5618 ( .A(n6459), .ZN(n6458) );
  INV_X1 U5619 ( .A(n5287), .ZN(n5284) );
  NOR2_X1 U5620 ( .A1(n9244), .A2(n5288), .ZN(n5287) );
  INV_X1 U5621 ( .A(n6627), .ZN(n5288) );
  OR2_X1 U5622 ( .A1(n9254), .A2(n8644), .ZN(n9211) );
  INV_X1 U5623 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9717) );
  AND2_X1 U5624 ( .A1(n6654), .A2(n5501), .ZN(n6210) );
  OAI21_X1 U5625 ( .B1(n6663), .B2(n9406), .A(P2_IR_REG_27__SCAN_IN), .ZN(
        n5115) );
  OAI21_X1 U5626 ( .B1(n6360), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6373) );
  OR2_X1 U5627 ( .A1(n6349), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6360) );
  OR2_X1 U5628 ( .A1(n6339), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6349) );
  NOR2_X1 U5629 ( .A1(n5852), .A2(n5851), .ZN(n5869) );
  NAND2_X1 U5630 ( .A1(n6791), .A2(n6790), .ZN(n5059) );
  OAI21_X1 U5631 ( .B1(n7474), .B2(n7475), .A(n7476), .ZN(n6791) );
  OR2_X1 U5632 ( .A1(n6743), .A2(n6930), .ZN(n6749) );
  INV_X1 U5633 ( .A(n6759), .ZN(n6810) );
  NOR2_X1 U5634 ( .A1(n8281), .A2(n8280), .ZN(n8395) );
  MUX2_X1 U5635 ( .A(n8431), .B(n8429), .S(n8400), .Z(n8394) );
  NOR2_X1 U5636 ( .A1(n5010), .A2(n5008), .ZN(n8438) );
  NAND2_X1 U5637 ( .A1(n4928), .A2(n5009), .ZN(n5008) );
  AOI22_X1 U5638 ( .A1(n8435), .A2(n8497), .B1(n8433), .B2(n8434), .ZN(n5010)
         );
  AND2_X1 U5639 ( .A1(n9904), .A2(n8262), .ZN(n8432) );
  OR2_X1 U5640 ( .A1(n6714), .A2(n7243), .ZN(n8393) );
  OR2_X1 U5641 ( .A1(n8283), .A2(n5166), .ZN(n5165) );
  INV_X1 U5642 ( .A(n6132), .ZN(n5166) );
  OR2_X1 U5643 ( .A1(n9928), .A2(n9938), .ZN(n8278) );
  NAND2_X1 U5644 ( .A1(n9928), .A2(n9938), .ZN(n8420) );
  INV_X1 U5645 ( .A(n6086), .ZN(n5388) );
  INV_X1 U5646 ( .A(n5178), .ZN(n5176) );
  OR2_X1 U5647 ( .A1(n6095), .A2(n6094), .ZN(n6110) );
  AND2_X1 U5648 ( .A1(n6001), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6018) );
  INV_X1 U5649 ( .A(n10086), .ZN(n5073) );
  NOR2_X1 U5650 ( .A1(n10159), .A2(n10166), .ZN(n5150) );
  INV_X1 U5651 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5985) );
  OR2_X1 U5652 ( .A1(n5973), .A2(n5972), .ZN(n5986) );
  NOR2_X1 U5653 ( .A1(n5939), .A2(n9425), .ZN(n5957) );
  NOR2_X1 U5654 ( .A1(n5914), .A2(n5183), .ZN(n5182) );
  INV_X1 U5655 ( .A(n5893), .ZN(n5183) );
  INV_X1 U5656 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5906) );
  OR2_X1 U5657 ( .A1(n5907), .A2(n5906), .ZN(n5924) );
  NOR2_X1 U5658 ( .A1(n7672), .A2(n7658), .ZN(n5154) );
  OR2_X1 U5659 ( .A1(n6157), .A2(n8244), .ZN(n8464) );
  NAND2_X1 U5660 ( .A1(n10628), .A2(n5746), .ZN(n8451) );
  AND2_X1 U5661 ( .A1(n5382), .A2(n5474), .ZN(n5129) );
  AND2_X1 U5662 ( .A1(n8297), .A2(n8457), .ZN(n10696) );
  AND2_X1 U5663 ( .A1(n5701), .A2(n7050), .ZN(n5725) );
  AND2_X1 U5664 ( .A1(n6725), .A2(n9886), .ZN(n8406) );
  XNOR2_X1 U5665 ( .A(n8223), .B(n8222), .ZN(n8225) );
  NAND2_X1 U5666 ( .A1(n6133), .A2(n9654), .ZN(n5429) );
  NAND2_X1 U5667 ( .A1(n5688), .A2(n5430), .ZN(n6133) );
  AND2_X1 U5668 ( .A1(n5687), .A2(n5431), .ZN(n5430) );
  INV_X1 U5669 ( .A(n5690), .ZN(n5431) );
  AND2_X1 U5670 ( .A1(n5687), .A2(n5686), .ZN(n6119) );
  AND2_X1 U5671 ( .A1(n5682), .A2(n5681), .ZN(n6102) );
  INV_X1 U5672 ( .A(n5677), .ZN(n5400) );
  INV_X1 U5673 ( .A(n5399), .ZN(n5398) );
  OAI21_X1 U5674 ( .B1(n6088), .B2(n5400), .A(n6102), .ZN(n5399) );
  NAND2_X1 U5675 ( .A1(n6089), .A2(n6088), .ZN(n6091) );
  AND2_X1 U5676 ( .A1(n5671), .A2(n5670), .ZN(n6073) );
  NOR2_X1 U5677 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5524) );
  NAND2_X1 U5678 ( .A1(n4993), .A2(n5655), .ZN(n5420) );
  INV_X1 U5679 ( .A(SI_18_), .ZN(n9652) );
  NOR2_X1 U5680 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5066) );
  XNOR2_X1 U5681 ( .A(n5646), .B(n5645), .ZN(n5981) );
  INV_X1 U5682 ( .A(SI_17_), .ZN(n5645) );
  INV_X1 U5683 ( .A(SI_14_), .ZN(n9671) );
  INV_X1 U5684 ( .A(SI_13_), .ZN(n9674) );
  INV_X1 U5685 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5900) );
  OAI21_X1 U5686 ( .B1(n5616), .B2(n5264), .A(n4975), .ZN(n5263) );
  INV_X1 U5687 ( .A(n5843), .ZN(n5264) );
  NOR2_X1 U5688 ( .A1(n5828), .A2(n5267), .ZN(n5266) );
  OR2_X1 U5689 ( .A1(n6469), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U5690 ( .A1(n6477), .A2(n9710), .ZN(n6493) );
  INV_X1 U5691 ( .A(n6478), .ZN(n6477) );
  NAND2_X1 U5692 ( .A1(n8056), .A2(n8055), .ZN(n5477) );
  AND2_X1 U5693 ( .A1(n8693), .A2(n8566), .ZN(n8635) );
  AND2_X1 U5694 ( .A1(n8632), .A2(n8562), .ZN(n8659) );
  NAND2_X1 U5695 ( .A1(n4997), .A2(n5005), .ZN(n5004) );
  INV_X1 U5696 ( .A(n8190), .ZN(n5005) );
  NOR2_X1 U5697 ( .A1(n8679), .A2(n5491), .ZN(n5490) );
  INV_X1 U5698 ( .A(n8551), .ZN(n5491) );
  NAND2_X1 U5699 ( .A1(n8549), .A2(n8621), .ZN(n8623) );
  OR2_X1 U5700 ( .A1(n6539), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U5701 ( .A1(n8534), .A2(n8833), .ZN(n5495) );
  AOI21_X1 U5702 ( .B1(n6231), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7176), .ZN(
        n7025) );
  NAND2_X1 U5703 ( .A1(n10513), .A2(n4940), .ZN(n7338) );
  NAND2_X1 U5704 ( .A1(n7338), .A2(n7339), .ZN(n7708) );
  NAND2_X1 U5705 ( .A1(n7342), .A2(n7343), .ZN(n7703) );
  XNOR2_X1 U5706 ( .A(n7704), .B(n5220), .ZN(n10534) );
  NAND2_X1 U5707 ( .A1(n10534), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10533) );
  INV_X1 U5708 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U5709 ( .A(n7710), .B(n5220), .ZN(n10531) );
  NOR2_X1 U5710 ( .A1(n10535), .A2(n5116), .ZN(n10552) );
  NOR2_X1 U5711 ( .A1(n5117), .A2(n5220), .ZN(n5116) );
  INV_X1 U5712 ( .A(n7701), .ZN(n5117) );
  NAND2_X1 U5713 ( .A1(n10546), .A2(n10547), .ZN(n10545) );
  XNOR2_X1 U5714 ( .A(n7822), .B(n7816), .ZN(n7712) );
  NAND2_X1 U5715 ( .A1(n7712), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U5716 ( .A1(n7825), .A2(n7826), .ZN(n7885) );
  XNOR2_X1 U5717 ( .A(n7928), .B(n7921), .ZN(n7887) );
  NAND2_X1 U5718 ( .A1(n7887), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U5719 ( .A1(n8079), .A2(n8080), .ZN(n8081) );
  NAND2_X1 U5720 ( .A1(n8938), .A2(n5390), .ZN(n8967) );
  OR2_X1 U5721 ( .A1(n8939), .A2(n8075), .ZN(n5390) );
  NAND2_X1 U5722 ( .A1(n8957), .A2(n8958), .ZN(n10571) );
  NAND2_X1 U5723 ( .A1(n10571), .A2(n10572), .ZN(n10570) );
  XNOR2_X1 U5724 ( .A(n8990), .B(n8978), .ZN(n8960) );
  XNOR2_X1 U5725 ( .A(n9018), .B(n9028), .ZN(n9013) );
  NAND2_X1 U5726 ( .A1(n9011), .A2(n5219), .ZN(n9018) );
  OR2_X1 U5727 ( .A1(n9012), .A2(n9236), .ZN(n5219) );
  NAND2_X1 U5728 ( .A1(n6645), .A2(n6641), .ZN(n9073) );
  INV_X1 U5729 ( .A(n8881), .ZN(n9098) );
  OR2_X1 U5730 ( .A1(n6509), .A2(n6508), .ZN(n9112) );
  OR2_X1 U5731 ( .A1(n6495), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6513) );
  AND2_X1 U5732 ( .A1(n8850), .A2(n8847), .ZN(n9200) );
  NAND2_X1 U5733 ( .A1(n6434), .A2(n6433), .ZN(n6446) );
  INV_X1 U5734 ( .A(n6435), .ZN(n6434) );
  NAND2_X1 U5735 ( .A1(n6407), .A2(n9742), .ZN(n6420) );
  INV_X1 U5736 ( .A(n6408), .ZN(n6407) );
  OR2_X1 U5737 ( .A1(n6393), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U5738 ( .A1(n4986), .A2(n5287), .ZN(n9241) );
  NAND2_X1 U5739 ( .A1(n5275), .A2(n5278), .ZN(n6626) );
  INV_X1 U5740 ( .A(n5279), .ZN(n5278) );
  AND2_X1 U5741 ( .A1(n8834), .A2(n6400), .ZN(n9259) );
  NAND2_X1 U5742 ( .A1(n6379), .A2(n6378), .ZN(n6393) );
  INV_X1 U5743 ( .A(n6380), .ZN(n6379) );
  NAND2_X1 U5744 ( .A1(n5346), .A2(n5344), .ZN(n8096) );
  NOR2_X1 U5745 ( .A1(n5345), .A2(n4955), .ZN(n5344) );
  INV_X1 U5746 ( .A(n8149), .ZN(n5345) );
  NAND2_X1 U5747 ( .A1(n5346), .A2(n8149), .ZN(n8093) );
  AOI21_X1 U5748 ( .B1(n5328), .B2(n5333), .A(n4971), .ZN(n5325) );
  AND2_X1 U5749 ( .A1(n8790), .A2(n8787), .ZN(n8744) );
  AND2_X1 U5750 ( .A1(n8786), .A2(n8782), .ZN(n8779) );
  NAND2_X1 U5751 ( .A1(n7499), .A2(n8742), .ZN(n7498) );
  OR2_X1 U5752 ( .A1(n8515), .A2(n7509), .ZN(n8775) );
  AND2_X1 U5753 ( .A1(n8906), .A2(n7645), .ZN(n6977) );
  OR2_X1 U5754 ( .A1(n8887), .A2(n6976), .ZN(n7453) );
  NAND2_X1 U5755 ( .A1(n6667), .A2(n7081), .ZN(n7452) );
  OR2_X1 U5756 ( .A1(n7069), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U5757 ( .A1(n6419), .A2(n6418), .ZN(n8840) );
  AND4_X1 U5758 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n7579)
         );
  AND2_X1 U5759 ( .A1(n6665), .A2(n6664), .ZN(n6688) );
  XNOR2_X1 U5760 ( .A(n6690), .B(n6689), .ZN(n7966) );
  NAND2_X1 U5761 ( .A1(n5498), .A2(n5497), .ZN(n5352) );
  INV_X1 U5762 ( .A(n6810), .ZN(n6993) );
  AND2_X1 U5763 ( .A1(n6943), .A2(n6942), .ZN(n6944) );
  NAND2_X1 U5764 ( .A1(n5059), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U5765 ( .A1(n5055), .A2(n5058), .ZN(n6800) );
  INV_X1 U5766 ( .A(n5059), .ZN(n5055) );
  INV_X1 U5767 ( .A(n5441), .ZN(n5440) );
  OAI21_X1 U5768 ( .B1(n6866), .B2(n5442), .A(n6865), .ZN(n5441) );
  NAND2_X1 U5769 ( .A1(n5445), .A2(n5448), .ZN(n5442) );
  NOR2_X1 U5770 ( .A1(n6866), .A2(n5444), .ZN(n5443) );
  INV_X1 U5771 ( .A(n5445), .ZN(n5444) );
  OR2_X1 U5772 ( .A1(n9528), .A2(n9523), .ZN(n5459) );
  XNOR2_X1 U5773 ( .A(n6762), .B(n6930), .ZN(n6763) );
  INV_X1 U5774 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5851) );
  OAI21_X1 U5775 ( .B1(n5059), .B2(n5057), .A(n5056), .ZN(n7789) );
  NAND2_X1 U5776 ( .A1(n5058), .A2(n6799), .ZN(n5056) );
  NOR2_X1 U5777 ( .A1(n5058), .A2(n6799), .ZN(n5057) );
  NAND2_X1 U5778 ( .A1(n9443), .A2(n9444), .ZN(n5471) );
  OR2_X1 U5779 ( .A1(n9443), .A2(n9444), .ZN(n5472) );
  AOI21_X1 U5780 ( .B1(n8041), .B2(n7999), .A(n5437), .ZN(n5436) );
  INV_X1 U5781 ( .A(n8042), .ZN(n5437) );
  AND2_X1 U5782 ( .A1(n5746), .A2(n6881), .ZN(n6751) );
  NAND2_X1 U5783 ( .A1(n5051), .A2(n5050), .ZN(n9539) );
  NOR2_X1 U5784 ( .A1(n5508), .A2(n4941), .ZN(n5050) );
  OR2_X1 U5785 ( .A1(n6963), .A2(n6962), .ZN(n9759) );
  NOR2_X1 U5786 ( .A1(n8432), .A2(n8431), .ZN(n8497) );
  NAND2_X1 U5787 ( .A1(n8508), .A2(n6726), .ZN(n8436) );
  AND2_X1 U5788 ( .A1(n5089), .A2(n5088), .ZN(n10400) );
  NAND2_X1 U5789 ( .A1(n10393), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U5790 ( .A1(n10398), .A2(n5093), .ZN(n10414) );
  AND2_X1 U5791 ( .A1(n10406), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5093) );
  OR2_X1 U5792 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  INV_X1 U5793 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7687) );
  AND2_X1 U5794 ( .A1(n10415), .A2(n5092), .ZN(n7126) );
  NAND2_X1 U5795 ( .A1(n7123), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5092) );
  OR2_X1 U5796 ( .A1(n5919), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5936) );
  AND2_X1 U5797 ( .A1(n6141), .A2(n6140), .ZN(n9926) );
  OAI21_X1 U5798 ( .B1(n9952), .B2(n9936), .A(n5071), .ZN(n6705) );
  AOI21_X1 U5799 ( .B1(n5310), .B2(n8382), .A(n8386), .ZN(n5071) );
  INV_X1 U5800 ( .A(n9940), .ZN(n9958) );
  INV_X1 U5801 ( .A(n8283), .ZN(n9964) );
  NAND2_X1 U5802 ( .A1(n10020), .A2(n4949), .ZN(n9968) );
  AND2_X1 U5803 ( .A1(n9985), .A2(n9986), .ZN(n5298) );
  OAI21_X1 U5804 ( .B1(n10072), .B2(n8485), .A(n5082), .ZN(n10026) );
  AOI21_X1 U5805 ( .B1(n5299), .B2(n5195), .A(n8411), .ZN(n5082) );
  NAND2_X1 U5806 ( .A1(n8135), .A2(n5146), .ZN(n10055) );
  NOR2_X1 U5807 ( .A1(n5147), .A2(n10148), .ZN(n5146) );
  INV_X1 U5808 ( .A(n5148), .ZN(n5147) );
  NOR2_X1 U5809 ( .A1(n10055), .A2(n10142), .ZN(n10020) );
  INV_X1 U5810 ( .A(n5083), .ZN(n10041) );
  AOI21_X1 U5811 ( .B1(n5171), .B2(n5174), .A(n5169), .ZN(n5168) );
  INV_X1 U5812 ( .A(n6011), .ZN(n5174) );
  INV_X1 U5813 ( .A(n5079), .ZN(n5075) );
  AOI21_X1 U5814 ( .B1(n5079), .B2(n5078), .A(n5077), .ZN(n5076) );
  INV_X1 U5815 ( .A(n8359), .ZN(n5077) );
  NAND2_X1 U5816 ( .A1(n8135), .A2(n8218), .ZN(n10080) );
  NAND2_X1 U5817 ( .A1(n8135), .A2(n5150), .ZN(n10078) );
  NAND2_X1 U5818 ( .A1(n8029), .A2(n4958), .ZN(n5309) );
  NAND2_X1 U5819 ( .A1(n5309), .A2(n5307), .ZN(n8013) );
  NOR2_X1 U5820 ( .A1(n8253), .A2(n5308), .ZN(n5307) );
  INV_X1 U5821 ( .A(n8472), .ZN(n5308) );
  OAI21_X1 U5822 ( .B1(n7953), .B2(n8250), .A(n5931), .ZN(n8025) );
  NAND2_X1 U5823 ( .A1(n7655), .A2(n4933), .ZN(n8035) );
  NAND2_X1 U5824 ( .A1(n7655), .A2(n5152), .ZN(n7955) );
  OAI21_X1 U5825 ( .B1(n7663), .B2(n5181), .A(n5179), .ZN(n7953) );
  AOI21_X1 U5826 ( .B1(n5182), .B2(n5180), .A(n4962), .ZN(n5179) );
  INV_X1 U5827 ( .A(n5182), .ZN(n5181) );
  INV_X1 U5828 ( .A(n5892), .ZN(n5180) );
  NAND2_X1 U5829 ( .A1(n7651), .A2(n8333), .ZN(n7664) );
  NAND2_X1 U5830 ( .A1(n7655), .A2(n8005), .ZN(n7668) );
  NOR2_X1 U5831 ( .A1(n7615), .A2(n7597), .ZN(n7655) );
  INV_X1 U5832 ( .A(n8240), .ZN(n8327) );
  AND4_X1 U5833 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n7601)
         );
  NAND2_X1 U5834 ( .A1(n7406), .A2(n7485), .ZN(n7596) );
  AND2_X1 U5835 ( .A1(n8320), .A2(n8319), .ZN(n8242) );
  NAND2_X1 U5836 ( .A1(n7368), .A2(n5811), .ZN(n7405) );
  NOR2_X1 U5837 ( .A1(n7370), .A2(n7418), .ZN(n7406) );
  NAND2_X1 U5838 ( .A1(n6163), .A2(n8448), .ZN(n7402) );
  NAND2_X1 U5839 ( .A1(n8316), .A2(n8318), .ZN(n8239) );
  NOR2_X1 U5840 ( .A1(n5777), .A2(n5157), .ZN(n5156) );
  INV_X1 U5841 ( .A(n5762), .ZN(n5157) );
  NAND2_X1 U5842 ( .A1(n9797), .A2(n10691), .ZN(n5160) );
  INV_X1 U5843 ( .A(n6161), .ZN(n10652) );
  NAND2_X1 U5844 ( .A1(n8304), .A2(n8451), .ZN(n10632) );
  AND2_X1 U5845 ( .A1(n6739), .A2(n10193), .ZN(n10185) );
  INV_X1 U5846 ( .A(n6731), .ZN(n10616) );
  OAI21_X1 U5847 ( .B1(n10199), .B2(n8399), .A(n10192), .ZN(n5141) );
  NOR2_X1 U5848 ( .A1(n9903), .A2(n5135), .ZN(n5134) );
  NAND2_X1 U5849 ( .A1(n10199), .A2(n5136), .ZN(n5135) );
  NOR2_X1 U5850 ( .A1(n9904), .A2(n10095), .ZN(n5136) );
  NAND2_X1 U5851 ( .A1(n6136), .A2(n6135), .ZN(n9947) );
  OR2_X1 U5852 ( .A1(n10688), .A2(n10692), .ZN(n10750) );
  AND4_X1 U5853 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n7610)
         );
  AND4_X1 U5854 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n7688)
         );
  AND4_X1 U5855 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n7479)
         );
  NAND2_X1 U5856 ( .A1(n5575), .A2(n10232), .ZN(n7383) );
  XNOR2_X1 U5857 ( .A(n8225), .B(SI_29_), .ZN(n9411) );
  XNOR2_X1 U5858 ( .A(n5528), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7052) );
  INV_X1 U5859 ( .A(n6951), .ZN(n8441) );
  AND2_X1 U5860 ( .A1(n5613), .A2(n5612), .ZN(n5812) );
  AOI21_X1 U5861 ( .B1(n5798), .B2(n5404), .A(n5403), .ZN(n5401) );
  INV_X1 U5862 ( .A(n5604), .ZN(n5404) );
  CLKBUF_X1 U5863 ( .A(n5783), .Z(n5784) );
  INV_X1 U5864 ( .A(n5011), .ZN(n5598) );
  NAND2_X1 U5865 ( .A1(n5765), .A2(n5764), .ZN(n5767) );
  AND2_X1 U5866 ( .A1(n7634), .A2(n7633), .ZN(n7727) );
  NAND2_X1 U5867 ( .A1(n8697), .A2(n8571), .ZN(n8586) );
  NAND2_X1 U5868 ( .A1(n8533), .A2(n8532), .ZN(n8597) );
  INV_X1 U5869 ( .A(n9266), .ZN(n10778) );
  INV_X1 U5870 ( .A(n5484), .ZN(n5483) );
  NAND2_X1 U5871 ( .A1(n6484), .A2(n6483), .ZN(n9137) );
  AND2_X1 U5872 ( .A1(n7227), .A2(n7252), .ZN(n5017) );
  NAND2_X1 U5873 ( .A1(n5007), .A2(n5477), .ZN(n8191) );
  AND2_X1 U5874 ( .A1(n8634), .A2(n8635), .ZN(n8696) );
  OR2_X1 U5875 ( .A1(n8535), .A2(n8644), .ZN(n8536) );
  NAND2_X1 U5876 ( .A1(n5006), .A2(n5004), .ZN(n8193) );
  AND2_X1 U5877 ( .A1(n8623), .A2(n5490), .ZN(n8677) );
  NAND2_X1 U5878 ( .A1(n8623), .A2(n8551), .ZN(n8678) );
  OAI21_X1 U5879 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8107) );
  NAND2_X1 U5880 ( .A1(n7214), .A2(n9267), .ZN(n8689) );
  NAND2_X1 U5881 ( .A1(n8539), .A2(n9232), .ZN(n5014) );
  OAI21_X1 U5882 ( .B1(n8539), .B2(n9232), .A(n8649), .ZN(n5015) );
  INV_X1 U5883 ( .A(n8712), .ZN(n8685) );
  NAND2_X1 U5884 ( .A1(n5496), .A2(n5492), .ZN(n8707) );
  AND2_X1 U5885 ( .A1(n8708), .A2(n5495), .ZN(n5492) );
  AND2_X1 U5886 ( .A1(n5496), .A2(n5495), .ZN(n8709) );
  INV_X1 U5887 ( .A(n8691), .ZN(n8706) );
  INV_X1 U5888 ( .A(n8654), .ZN(n8715) );
  NAND2_X1 U5889 ( .A1(n5246), .A2(n5245), .ZN(n5045) );
  XNOR2_X1 U5890 ( .A(n6595), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9056) );
  XNOR2_X1 U5891 ( .A(n6603), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8915) );
  INV_X1 U5892 ( .A(n9285), .ZN(n8920) );
  NAND2_X1 U5893 ( .A1(n6559), .A2(n6558), .ZN(n8921) );
  NAND4_X1 U5894 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n8924)
         );
  NAND4_X1 U5895 ( .A1(n6321), .A2(n6320), .A3(n6319), .A4(n6318), .ZN(n7941)
         );
  OR2_X1 U5896 ( .A1(n6327), .A2(n6237), .ZN(n6238) );
  OR2_X1 U5897 ( .A1(n7572), .A2(n6226), .ZN(n6227) );
  OR2_X1 U5898 ( .A1(n6249), .A2(n7260), .ZN(n6230) );
  OR2_X1 U5899 ( .A1(n6249), .A2(n7490), .ZN(n5269) );
  AND2_X1 U5900 ( .A1(n5112), .A2(n5110), .ZN(n5111) );
  INV_X1 U5901 ( .A(n5119), .ZN(n10537) );
  INV_X1 U5902 ( .A(n7706), .ZN(n7815) );
  AND2_X1 U5903 ( .A1(n5107), .A2(n5106), .ZN(n7881) );
  NAND2_X1 U5904 ( .A1(n7810), .A2(n7816), .ZN(n5106) );
  NAND2_X1 U5905 ( .A1(n7812), .A2(n7811), .ZN(n5107) );
  OAI22_X1 U5906 ( .A1(n7922), .A2(n7948), .B1(n7921), .B2(n7920), .ZN(n7925)
         );
  AOI21_X1 U5907 ( .B1(n7918), .B2(n7917), .A(n5104), .ZN(n7984) );
  AND2_X1 U5908 ( .A1(n7916), .A2(n7921), .ZN(n5104) );
  OAI22_X1 U5909 ( .A1(n8074), .A2(n8073), .B1(n8072), .B2(n8071), .ZN(n8077)
         );
  NAND2_X1 U5910 ( .A1(n8077), .A2(n8076), .ZN(n8938) );
  OAI21_X1 U5911 ( .B1(n8934), .B2(n8933), .A(n4998), .ZN(n8954) );
  XNOR2_X1 U5912 ( .A(n8956), .B(n8952), .ZN(n8936) );
  OAI22_X1 U5913 ( .A1(n10574), .A2(n10573), .B1(n8955), .B2(n8965), .ZN(n8980) );
  OAI21_X1 U5914 ( .B1(n9040), .B2(n9207), .A(n9052), .ZN(n9041) );
  AND2_X1 U5915 ( .A1(n7576), .A2(n6591), .ZN(n9279) );
  NAND2_X1 U5916 ( .A1(n6564), .A2(n6563), .ZN(n9281) );
  NAND2_X1 U5917 ( .A1(n6550), .A2(n6549), .ZN(n9287) );
  AND2_X1 U5918 ( .A1(n6534), .A2(n6533), .ZN(n9292) );
  NAND2_X1 U5919 ( .A1(n6538), .A2(n6537), .ZN(n9295) );
  NAND2_X1 U5920 ( .A1(n9121), .A2(n8874), .ZN(n9108) );
  AND2_X1 U5921 ( .A1(n6519), .A2(n6518), .ZN(n9133) );
  NAND2_X1 U5922 ( .A1(n6525), .A2(n6524), .ZN(n9301) );
  NAND2_X1 U5923 ( .A1(n9158), .A2(n8863), .ZN(n9151) );
  NAND2_X1 U5924 ( .A1(n6492), .A2(n6491), .ZN(n9320) );
  NAND2_X1 U5925 ( .A1(n5319), .A2(n5323), .ZN(n9169) );
  NAND2_X1 U5926 ( .A1(n6454), .A2(n5320), .ZN(n5319) );
  NAND2_X1 U5927 ( .A1(n6468), .A2(n6467), .ZN(n9177) );
  NAND2_X1 U5928 ( .A1(n6454), .A2(n6453), .ZN(n9180) );
  NAND2_X1 U5929 ( .A1(n6445), .A2(n6444), .ZN(n9348) );
  AOI21_X1 U5930 ( .B1(n8166), .B2(n8819), .A(n5280), .ZN(n5277) );
  NAND2_X1 U5931 ( .A1(n5294), .A2(n8813), .ZN(n8151) );
  INV_X1 U5932 ( .A(n7941), .ZN(n7852) );
  NAND2_X1 U5933 ( .A1(n7767), .A2(n8795), .ZN(n7837) );
  NAND2_X1 U5934 ( .A1(n5327), .A2(n5332), .ZN(n7835) );
  NAND2_X1 U5935 ( .A1(n7781), .A2(n5336), .ZN(n5327) );
  NAND2_X1 U5936 ( .A1(n5331), .A2(n6277), .ZN(n7770) );
  OR2_X1 U5937 ( .A1(n7781), .A2(n6278), .ZN(n5331) );
  NAND2_X1 U5938 ( .A1(n7463), .A2(n7458), .ZN(n5362) );
  INV_X1 U5939 ( .A(n9155), .ZN(n9170) );
  OR2_X1 U5940 ( .A1(n9194), .A2(n7487), .ZN(n9274) );
  INV_X1 U5941 ( .A(n10785), .ZN(n10777) );
  AND2_X1 U5942 ( .A1(n8887), .A2(n6977), .ZN(n7506) );
  INV_X1 U5943 ( .A(n9265), .ZN(n9253) );
  OR2_X1 U5944 ( .A1(n6401), .A2(n7041), .ZN(n6245) );
  AND2_X1 U5945 ( .A1(n10791), .A2(n10777), .ZN(n9331) );
  AOI21_X1 U5946 ( .B1(n9405), .B2(n8723), .A(n8720), .ZN(n9366) );
  AOI21_X1 U5947 ( .B1(n8529), .B2(n8723), .A(n4996), .ZN(n9369) );
  INV_X1 U5948 ( .A(n8873), .ZN(n9377) );
  NAND2_X1 U5949 ( .A1(n6476), .A2(n6475), .ZN(n9385) );
  INV_X1 U5950 ( .A(n8840), .ZN(n9404) );
  NAND2_X1 U5951 ( .A1(n6326), .A2(n6325), .ZN(n7950) );
  OR2_X1 U5952 ( .A1(n6274), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6216) );
  AND2_X1 U5953 ( .A1(n7966), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7086) );
  NAND2_X1 U5954 ( .A1(n6654), .A2(n5048), .ZN(n6200) );
  INV_X1 U5955 ( .A(n6688), .ZN(n8204) );
  INV_X1 U5956 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6658) );
  INV_X1 U5957 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7910) );
  INV_X1 U5958 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6597) );
  INV_X1 U5959 ( .A(n10565), .ZN(n8965) );
  OR2_X1 U5960 ( .A1(n6312), .A2(n6311), .ZN(n7884) );
  NAND2_X1 U5961 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U5962 ( .A1(n9513), .A2(n9514), .ZN(n9420) );
  NAND2_X1 U5963 ( .A1(n5061), .A2(n8041), .ZN(n7998) );
  NAND2_X1 U5964 ( .A1(n6813), .A2(n6812), .ZN(n5061) );
  NAND2_X1 U5965 ( .A1(n6017), .A2(n6016), .ZN(n10153) );
  INV_X1 U5966 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9459) );
  CLKBUF_X1 U5967 ( .A(n9454), .Z(n9455) );
  AND2_X1 U5968 ( .A1(n6131), .A2(n6130), .ZN(n10103) );
  AND2_X1 U5969 ( .A1(n5453), .A2(n5450), .ZN(n5449) );
  INV_X1 U5970 ( .A(n9466), .ZN(n5450) );
  OR2_X1 U5971 ( .A1(n5469), .A2(n6774), .ZN(n7291) );
  NAND2_X1 U5972 ( .A1(n7245), .A2(n6771), .ZN(n5469) );
  AND2_X1 U5973 ( .A1(n6085), .A2(n6084), .ZN(n9991) );
  AOI21_X1 U5974 ( .B1(n5454), .B2(n5458), .A(n5455), .ZN(n9498) );
  NOR2_X1 U5975 ( .A1(n9523), .A2(n5460), .ZN(n5458) );
  AND2_X1 U5976 ( .A1(n5067), .A2(n5068), .ZN(n10700) );
  INV_X1 U5977 ( .A(n5069), .ZN(n5067) );
  AND2_X1 U5978 ( .A1(n5761), .A2(n5760), .ZN(n5068) );
  INV_X1 U5979 ( .A(n7056), .ZN(n10702) );
  AND2_X1 U5980 ( .A1(n6028), .A2(n6027), .ZN(n10054) );
  NAND2_X1 U5981 ( .A1(n5470), .A2(n5471), .ZN(n9505) );
  AND4_X1 U5982 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n9771)
         );
  INV_X1 U5983 ( .A(n9759), .ZN(n9774) );
  INV_X1 U5984 ( .A(n5454), .ZN(n9528) );
  AND2_X1 U5985 ( .A1(n5466), .A2(n5464), .ZN(n5463) );
  NAND2_X1 U5986 ( .A1(n6774), .A2(n5468), .ZN(n5466) );
  AND2_X1 U5987 ( .A1(n6955), .A2(n10718), .ZN(n9779) );
  NAND2_X1 U5988 ( .A1(n6966), .A2(n9810), .ZN(n9770) );
  OAI21_X1 U5989 ( .B1(n5412), .B2(n5206), .A(n4934), .ZN(n5205) );
  INV_X1 U5990 ( .A(n10054), .ZN(n10088) );
  INV_X1 U5991 ( .A(n10700), .ZN(n9798) );
  OR3_X1 U5992 ( .A1(n7052), .A2(P1_U3086), .A3(n6729), .ZN(n9799) );
  INV_X1 U5993 ( .A(n5089), .ZN(n10385) );
  AND2_X1 U5994 ( .A1(n7053), .A2(n7111), .ZN(n10585) );
  NOR2_X1 U5995 ( .A1(n10428), .A2(n5087), .ZN(n7265) );
  AND2_X1 U5996 ( .A1(n7273), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U5997 ( .A1(n7265), .A2(n7266), .ZN(n9854) );
  NOR2_X1 U5998 ( .A1(n10484), .A2(n10483), .ZN(n10482) );
  NAND2_X1 U5999 ( .A1(n9854), .A2(n5086), .ZN(n10484) );
  OR2_X1 U6000 ( .A1(n9855), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5086) );
  NOR2_X1 U6001 ( .A1(n10459), .A2(n9859), .ZN(n9862) );
  OR2_X1 U6002 ( .A1(n9907), .A2(n9906), .ZN(n10099) );
  OR2_X1 U6003 ( .A1(n6145), .A2(n6144), .ZN(n9914) );
  OR2_X1 U6004 ( .A1(n6701), .A2(n6152), .ZN(n9923) );
  NAND2_X1 U6005 ( .A1(n5162), .A2(n6132), .ZN(n9935) );
  NAND2_X1 U6006 ( .A1(n9963), .A2(n8283), .ZN(n5162) );
  INV_X1 U6007 ( .A(n5311), .ZN(n9937) );
  AND2_X1 U6008 ( .A1(n6117), .A2(n6116), .ZN(n10111) );
  NAND2_X1 U6009 ( .A1(n6122), .A2(n6121), .ZN(n9962) );
  NAND2_X1 U6010 ( .A1(n6087), .A2(n6086), .ZN(n9984) );
  NAND2_X1 U6011 ( .A1(n5370), .A2(n5178), .ZN(n6087) );
  AND2_X1 U6012 ( .A1(n6071), .A2(n6070), .ZN(n10126) );
  NAND2_X1 U6013 ( .A1(n5370), .A2(n5372), .ZN(n10014) );
  AND2_X1 U6014 ( .A1(n6056), .A2(n6055), .ZN(n10132) );
  NAND2_X1 U6015 ( .A1(n5374), .A2(n6057), .ZN(n10019) );
  NAND2_X1 U6016 ( .A1(n10032), .A2(n10043), .ZN(n5374) );
  AND2_X1 U6017 ( .A1(n6042), .A2(n6041), .ZN(n10139) );
  NAND2_X1 U6018 ( .A1(n5386), .A2(n6012), .ZN(n10064) );
  NAND2_X1 U6019 ( .A1(n10077), .A2(n6011), .ZN(n5386) );
  AND3_X1 U6020 ( .A1(n5990), .A2(n5989), .A3(n5988), .ZN(n10156) );
  NAND2_X1 U6021 ( .A1(n8131), .A2(n8481), .ZN(n8206) );
  NOR2_X1 U6022 ( .A1(n8141), .A2(n5365), .ZN(n5364) );
  INV_X1 U6023 ( .A(n5367), .ZN(n5365) );
  NAND2_X1 U6024 ( .A1(n5366), .A2(n5367), .ZN(n8142) );
  AND2_X1 U6025 ( .A1(n5304), .A2(n8341), .ZN(n7800) );
  NAND2_X1 U6026 ( .A1(n5184), .A2(n5893), .ZN(n7798) );
  NAND2_X1 U6027 ( .A1(n7663), .A2(n5892), .ZN(n5184) );
  INV_X1 U6028 ( .A(n10674), .ZN(n10010) );
  AND2_X1 U6029 ( .A1(n10690), .A2(n10689), .ZN(n7316) );
  NAND2_X1 U6030 ( .A1(n7066), .A2(n8273), .ZN(n5303) );
  INV_X1 U6031 ( .A(n7321), .ZN(n7393) );
  NAND2_X1 U6032 ( .A1(n5138), .A2(n5133), .ZN(n10196) );
  NAND2_X1 U6033 ( .A1(n9903), .A2(n5139), .ZN(n5138) );
  AOI21_X1 U6034 ( .B1(n5141), .B2(n5140), .A(n5134), .ZN(n5133) );
  AND2_X1 U6035 ( .A1(n8403), .A2(n5140), .ZN(n5139) );
  AND2_X1 U6036 ( .A1(n9912), .A2(n9916), .ZN(n6718) );
  NAND2_X1 U6037 ( .A1(n10758), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5379) );
  INV_X1 U6038 ( .A(n9962), .ZN(n10211) );
  INV_X1 U6039 ( .A(n10013), .ZN(n10221) );
  OR3_X1 U6040 ( .A1(n7052), .A2(n6957), .A3(P1_U3086), .ZN(n10362) );
  NAND2_X1 U6041 ( .A1(n10234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  INV_X1 U6042 ( .A(n5712), .ZN(n10242) );
  XNOR2_X1 U6043 ( .A(n6174), .B(P1_IR_REG_28__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U6044 ( .A1(n5539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5540) );
  INV_X1 U6045 ( .A(n6725), .ZN(n8508) );
  AOI21_X1 U6046 ( .B1(n5253), .B2(n5256), .A(n5252), .ZN(n5251) );
  NAND2_X1 U6047 ( .A1(n5933), .A2(n5932), .ZN(n5935) );
  OR2_X1 U6048 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U6049 ( .A1(n5896), .A2(n5627), .ZN(n5916) );
  NAND2_X1 U6050 ( .A1(n5424), .A2(n5427), .ZN(n5895) );
  NAND2_X1 U6051 ( .A1(n5799), .A2(n5798), .ZN(n5801) );
  NAND2_X1 U6052 ( .A1(n5780), .A2(n5604), .ZN(n5799) );
  NAND2_X1 U6053 ( .A1(n5099), .A2(n5098), .ZN(n5770) );
  NAND2_X1 U6054 ( .A1(n10233), .A2(n5101), .ZN(n5098) );
  NAND2_X1 U6055 ( .A1(n5102), .A2(n5100), .ZN(n5099) );
  OR2_X1 U6056 ( .A1(n5122), .A2(n9035), .ZN(P2_U3200) );
  OAI21_X1 U6057 ( .B1(n9037), .B2(n9044), .A(n5123), .ZN(n5122) );
  NOR2_X1 U6058 ( .A1(n5339), .A2(n5341), .ZN(n8521) );
  NOR2_X1 U6059 ( .A1(n5514), .A2(n6984), .ZN(n6985) );
  AOI21_X1 U6060 ( .B1(n7004), .B2(n7003), .A(n7002), .ZN(n7005) );
  OR2_X1 U6061 ( .A1(n10475), .A2(n5094), .ZN(P1_U3261) );
  OR2_X1 U6062 ( .A1(n10476), .A2(n5095), .ZN(n5094) );
  AOI21_X1 U6063 ( .B1(n9903), .B2(n8403), .A(n5137), .ZN(n10096) );
  NAND2_X1 U6064 ( .A1(n10756), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6065 ( .A1(n6182), .A2(n10757), .ZN(n5313) );
  NAND2_X1 U6066 ( .A1(n5380), .A2(n5377), .ZN(P1_U3518) );
  INV_X1 U6067 ( .A(n5378), .ZN(n5377) );
  NAND2_X1 U6068 ( .A1(n6182), .A2(n10761), .ZN(n5380) );
  OAI21_X1 U6069 ( .B1(n6183), .B2(n10220), .A(n5379), .ZN(n5378) );
  NAND2_X1 U6070 ( .A1(n10199), .A2(n8433), .ZN(n4928) );
  INV_X2 U6071 ( .A(n4926), .ZN(n6927) );
  INV_X1 U6072 ( .A(n9936), .ZN(n5310) );
  AND2_X1 U6073 ( .A1(n5234), .A2(n5232), .ZN(n4929) );
  NAND2_X1 U6074 ( .A1(n5711), .A2(n5712), .ZN(n5836) );
  NAND2_X1 U6075 ( .A1(n10020), .A2(n5145), .ZN(n4930) );
  INV_X1 U6076 ( .A(n8487), .ZN(n5195) );
  NAND2_X1 U6077 ( .A1(n5956), .A2(n5955), .ZN(n8017) );
  AND2_X1 U6078 ( .A1(n5483), .A2(n8658), .ZN(n4931) );
  NAND2_X1 U6079 ( .A1(n5451), .A2(n5453), .ZN(n9464) );
  AND2_X1 U6080 ( .A1(n5696), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4932) );
  INV_X1 U6081 ( .A(n5333), .ZN(n5332) );
  OAI21_X1 U6082 ( .B1(n6292), .B2(n5335), .A(n5334), .ZN(n5333) );
  AND2_X1 U6083 ( .A1(n5152), .A2(n7958), .ZN(n4933) );
  AND3_X1 U6084 ( .A1(n8442), .A2(n8441), .A3(n4981), .ZN(n4934) );
  INV_X1 U6085 ( .A(n8349), .ZN(n8251) );
  AND2_X1 U6086 ( .A1(n8284), .A2(n8373), .ZN(n10025) );
  AND2_X1 U6087 ( .A1(n7531), .A2(n7530), .ZN(n4935) );
  AND2_X1 U6088 ( .A1(n5254), .A2(n5932), .ZN(n5253) );
  XNOR2_X1 U6089 ( .A(n6734), .B(n6744), .ZN(n6750) );
  AND2_X1 U6090 ( .A1(n5493), .A2(n5001), .ZN(n4936) );
  NAND2_X1 U6091 ( .A1(n5051), .A2(n5053), .ZN(n4937) );
  OR2_X1 U6092 ( .A1(n7729), .A2(n7728), .ZN(n4938) );
  NAND2_X1 U6093 ( .A1(n6107), .A2(n6106), .ZN(n9471) );
  INV_X1 U6094 ( .A(n9471), .ZN(n5142) );
  INV_X1 U6095 ( .A(n10549), .ZN(n7707) );
  AND2_X1 U6096 ( .A1(n5000), .A2(n6800), .ZN(n4939) );
  NAND2_X1 U6097 ( .A1(n5062), .A2(n6768), .ZN(n7245) );
  INV_X1 U6098 ( .A(n5013), .ZN(n8542) );
  NAND2_X2 U6099 ( .A1(n10238), .A2(n10242), .ZN(n5758) );
  NAND4_X1 U6100 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n6739)
         );
  AND3_X1 U6101 ( .A1(n5473), .A2(n5101), .A3(n5737), .ZN(n5769) );
  OR2_X1 U6102 ( .A1(n7337), .A2(n10516), .ZN(n4940) );
  INV_X1 U6103 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5705) );
  INV_X1 U6104 ( .A(n8818), .ZN(n5038) );
  NAND2_X1 U6105 ( .A1(n5459), .A2(n9435), .ZN(n9434) );
  XOR2_X1 U6106 ( .A(n6875), .B(n6777), .Z(n4941) );
  AND3_X1 U6107 ( .A1(n5706), .A2(n5705), .A3(n5699), .ZN(n4942) );
  NAND2_X1 U6108 ( .A1(n6703), .A2(n6702), .ZN(n6714) );
  AND2_X1 U6109 ( .A1(n5867), .A2(n5866), .ZN(n8005) );
  NOR2_X1 U6110 ( .A1(n7187), .A2(n5111), .ZN(n4943) );
  AND2_X1 U6111 ( .A1(n9287), .A2(n8921), .ZN(n4944) );
  NAND2_X1 U6112 ( .A1(n8558), .A2(n8658), .ZN(n8604) );
  OR2_X1 U6113 ( .A1(n10013), .A2(n10027), .ZN(n4945) );
  OR2_X1 U6114 ( .A1(n7579), .A2(n10680), .ZN(n4946) );
  OR2_X1 U6115 ( .A1(n7040), .A2(n5997), .ZN(n4947) );
  NOR2_X1 U6116 ( .A1(n7021), .A2(n7022), .ZN(n4948) );
  NAND2_X1 U6117 ( .A1(n5482), .A2(n6231), .ZN(n6255) );
  INV_X1 U6118 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U6119 ( .A1(n5349), .A2(n5351), .ZN(n6661) );
  NAND2_X1 U6120 ( .A1(n6231), .A2(n6232), .ZN(n6242) );
  NAND2_X1 U6121 ( .A1(n6061), .A2(n6060), .ZN(n10135) );
  NAND2_X1 U6122 ( .A1(n5905), .A2(n5904), .ZN(n8117) );
  AND2_X1 U6123 ( .A1(n5143), .A2(n5142), .ZN(n4949) );
  AND2_X1 U6124 ( .A1(n7321), .A2(n10689), .ZN(n4950) );
  NAND2_X1 U6125 ( .A1(n5511), .A2(n8818), .ZN(n4951) );
  NAND2_X1 U6126 ( .A1(n5984), .A2(n5983), .ZN(n10166) );
  AND2_X1 U6127 ( .A1(n5027), .A2(n5028), .ZN(n4952) );
  OR2_X1 U6128 ( .A1(n7709), .A2(n7340), .ZN(n4953) );
  AND2_X1 U6129 ( .A1(n8376), .A2(n8412), .ZN(n4954) );
  INV_X1 U6130 ( .A(n9995), .ZN(n10216) );
  NOR2_X1 U6131 ( .A1(n10743), .A2(n8163), .ZN(n4955) );
  AND2_X1 U6132 ( .A1(n8414), .A2(n8406), .ZN(n4956) );
  OR2_X1 U6133 ( .A1(n7709), .A2(n7335), .ZN(n4957) );
  AND2_X1 U6134 ( .A1(n8251), .A2(n8339), .ZN(n4958) );
  OR2_X1 U6135 ( .A1(n9168), .A2(n5228), .ZN(n4959) );
  NAND2_X1 U6136 ( .A1(n6034), .A2(n6033), .ZN(n10148) );
  AND2_X1 U6137 ( .A1(n5313), .A2(n5312), .ZN(n4960) );
  AND2_X1 U6138 ( .A1(n5311), .A2(n5310), .ZN(n4961) );
  AND2_X1 U6139 ( .A1(n8117), .A2(n8051), .ZN(n4962) );
  NAND2_X1 U6140 ( .A1(n5922), .A2(n5921), .ZN(n10180) );
  INV_X1 U6141 ( .A(n7838), .ZN(n5329) );
  AND2_X1 U6142 ( .A1(n5024), .A2(n8843), .ZN(n4963) );
  AND2_X1 U6143 ( .A1(n8352), .A2(n8481), .ZN(n8141) );
  INV_X1 U6144 ( .A(n8141), .ZN(n5078) );
  INV_X1 U6145 ( .A(n5428), .ZN(n5427) );
  NOR2_X1 U6146 ( .A1(n9995), .A2(n10005), .ZN(n4964) );
  NOR2_X1 U6147 ( .A1(n10135), .A2(n10045), .ZN(n4965) );
  INV_X1 U6148 ( .A(n9797), .ZN(n10654) );
  OR2_X1 U6149 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(n10233), .ZN(n4966) );
  INV_X1 U6150 ( .A(n10033), .ZN(n10043) );
  AND2_X1 U6151 ( .A1(n8367), .A2(n8368), .ZN(n10033) );
  AND2_X1 U6152 ( .A1(n9995), .A2(n10005), .ZN(n4967) );
  OR2_X1 U6153 ( .A1(n5385), .A2(n5384), .ZN(n4968) );
  INV_X1 U6154 ( .A(n8485), .ZN(n5299) );
  NAND2_X1 U6155 ( .A1(n5587), .A2(n5185), .ZN(n4969) );
  INV_X1 U6156 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U6157 ( .A1(n8771), .A2(n7468), .ZN(n4970) );
  AND2_X1 U6158 ( .A1(n7905), .A2(n7761), .ZN(n4971) );
  NAND3_X1 U6159 ( .A1(n6302), .A2(n6194), .A3(n5498), .ZN(n4972) );
  AND2_X1 U6160 ( .A1(n10015), .A2(n8372), .ZN(n4973) );
  AND2_X1 U6161 ( .A1(n8471), .A2(n8339), .ZN(n8250) );
  AND2_X1 U6162 ( .A1(n4929), .A2(n9259), .ZN(n4974) );
  OR2_X1 U6163 ( .A1(n5618), .A2(SI_9_), .ZN(n4975) );
  INV_X1 U6164 ( .A(n5321), .ZN(n5320) );
  OR2_X1 U6165 ( .A1(n6466), .A2(n5322), .ZN(n5321) );
  NAND2_X1 U6166 ( .A1(n5462), .A2(n7292), .ZN(n5467) );
  INV_X1 U6167 ( .A(n5701), .ZN(n5579) );
  AND2_X1 U6168 ( .A1(n5451), .A2(n5449), .ZN(n9465) );
  NAND2_X1 U6169 ( .A1(n6216), .A2(n6217), .ZN(n5314) );
  AND2_X1 U6170 ( .A1(n5028), .A2(n5026), .ZN(n4976) );
  NOR2_X1 U6171 ( .A1(n5292), .A2(n8877), .ZN(n4977) );
  NOR2_X1 U6172 ( .A1(n4944), .A2(n5342), .ZN(n4978) );
  INV_X1 U6173 ( .A(n5229), .ZN(n5231) );
  OAI211_X1 U6174 ( .C1(n9168), .C2(n5230), .A(n8861), .B(n8862), .ZN(n5229)
         );
  INV_X1 U6175 ( .A(n5932), .ZN(n5411) );
  AND2_X1 U6176 ( .A1(n5635), .A2(n5634), .ZN(n5932) );
  AND2_X1 U6177 ( .A1(n8403), .A2(n9899), .ZN(n8437) );
  AND2_X1 U6178 ( .A1(n7801), .A2(n8341), .ZN(n4979) );
  AND2_X1 U6179 ( .A1(n6891), .A2(n5471), .ZN(n4980) );
  INV_X1 U6180 ( .A(n5508), .ZN(n5053) );
  NAND2_X1 U6181 ( .A1(n5208), .A2(n8407), .ZN(n4981) );
  INV_X1 U6182 ( .A(n5758), .ZN(n5850) );
  INV_X1 U6183 ( .A(n7921), .ZN(n5389) );
  INV_X1 U6184 ( .A(n8072), .ZN(n5391) );
  INV_X1 U6185 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5302) );
  OAI21_X1 U6186 ( .B1(n9513), .B2(n5448), .A(n5445), .ZN(n9474) );
  INV_X1 U6187 ( .A(n9232), .ZN(n9204) );
  AND2_X1 U6188 ( .A1(n5438), .A2(n6818), .ZN(n4982) );
  AND2_X1 U6189 ( .A1(n10020), .A2(n5143), .ZN(n4983) );
  AND2_X1 U6190 ( .A1(n10020), .A2(n6177), .ZN(n4984) );
  INV_X1 U6191 ( .A(n7192), .ZN(n5110) );
  NOR2_X1 U6192 ( .A1(n8567), .A2(n8693), .ZN(n4985) );
  OR2_X1 U6193 ( .A1(n9257), .A2(n9259), .ZN(n4986) );
  NAND2_X1 U6194 ( .A1(n6624), .A2(n8818), .ZN(n8166) );
  NAND2_X1 U6195 ( .A1(n5439), .A2(n5440), .ZN(n9486) );
  INV_X1 U6196 ( .A(n5277), .ZN(n8176) );
  NAND2_X1 U6197 ( .A1(n5170), .A2(n5168), .ZN(n10050) );
  INV_X1 U6198 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5047) );
  NOR2_X1 U6199 ( .A1(n8136), .A2(n10171), .ZN(n8135) );
  NAND2_X1 U6200 ( .A1(n8193), .A2(n8192), .ZN(n8533) );
  AND4_X1 U6201 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n9426)
         );
  OR2_X1 U6202 ( .A1(n7879), .A2(n7884), .ZN(n4987) );
  NAND2_X1 U6203 ( .A1(n8538), .A2(n9247), .ZN(n4988) );
  NAND2_X1 U6204 ( .A1(n8135), .A2(n5148), .ZN(n5151) );
  INV_X1 U6205 ( .A(n9496), .ZN(n5460) );
  AND2_X1 U6206 ( .A1(n4986), .A2(n6627), .ZN(n4989) );
  AND2_X1 U6207 ( .A1(n5309), .A2(n8472), .ZN(n4990) );
  INV_X1 U6208 ( .A(n5627), .ZN(n5256) );
  OR2_X1 U6209 ( .A1(n7702), .A2(n7707), .ZN(n4991) );
  NOR2_X1 U6210 ( .A1(n9177), .A2(n9325), .ZN(n4992) );
  NAND2_X1 U6211 ( .A1(n8642), .A2(n8643), .ZN(n5016) );
  INV_X1 U6212 ( .A(n8054), .ZN(n8056) );
  NAND2_X1 U6213 ( .A1(n7973), .A2(n7972), .ZN(n8054) );
  OR2_X1 U6214 ( .A1(n6030), .A2(SI_20_), .ZN(n4993) );
  AND3_X1 U6215 ( .A1(n5510), .A2(n5523), .A3(n5065), .ZN(n4994) );
  AND2_X1 U6216 ( .A1(n8054), .A2(n7747), .ZN(n4995) );
  NAND2_X1 U6217 ( .A1(n6457), .A2(n6456), .ZN(n9186) );
  INV_X1 U6218 ( .A(n9186), .ZN(n5324) );
  INV_X1 U6219 ( .A(n10757), .ZN(n10756) );
  AND2_X1 U6220 ( .A1(n7427), .A2(n7426), .ZN(n7524) );
  NOR2_X1 U6221 ( .A1(n6274), .A2(n8722), .ZN(n4996) );
  OAI21_X1 U6222 ( .B1(n7244), .B2(n5063), .A(n5463), .ZN(n7328) );
  NAND2_X1 U6223 ( .A1(n5326), .A2(n5325), .ZN(n7752) );
  NAND2_X1 U6224 ( .A1(n5362), .A2(n6235), .ZN(n7497) );
  OR2_X1 U6225 ( .A1(n8108), .A2(n8195), .ZN(n4997) );
  INV_X1 U6226 ( .A(n6668), .ZN(n7220) );
  NAND2_X1 U6227 ( .A1(n5469), .A2(n6774), .ZN(n7290) );
  NAND2_X1 U6228 ( .A1(n6800), .A2(n6796), .ZN(n7685) );
  NAND2_X1 U6229 ( .A1(n6815), .A2(n6814), .ZN(n8041) );
  NAND2_X1 U6230 ( .A1(n7655), .A2(n5154), .ZN(n5155) );
  INV_X1 U6231 ( .A(n10754), .ZN(n10183) );
  OR2_X1 U6232 ( .A1(n8931), .A2(n8932), .ZN(n4998) );
  OR2_X1 U6233 ( .A1(n5354), .A2(n5352), .ZN(n4999) );
  AND2_X1 U6234 ( .A1(n6796), .A2(n6799), .ZN(n5000) );
  INV_X1 U6235 ( .A(n10095), .ZN(n5140) );
  INV_X1 U6236 ( .A(n6153), .ZN(n7387) );
  NAND2_X1 U6237 ( .A1(n7089), .A2(n7088), .ZN(n7090) );
  OR2_X1 U6238 ( .A1(n10688), .A2(n8441), .ZN(n10660) );
  INV_X1 U6239 ( .A(n10660), .ZN(n10192) );
  AND2_X1 U6240 ( .A1(n7148), .A2(n7152), .ZN(n7139) );
  NAND4_X1 U6241 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n5475)
         );
  NAND2_X1 U6242 ( .A1(n6602), .A2(n6601), .ZN(n8906) );
  INV_X1 U6243 ( .A(n8906), .ZN(n5247) );
  INV_X1 U6244 ( .A(n10529), .ZN(n5220) );
  NAND3_X1 U6245 ( .A1(n5007), .A2(n5477), .A3(n4997), .ZN(n5006) );
  NAND2_X1 U6246 ( .A1(n5011), .A2(SI_4_), .ZN(n5600) );
  XNOR2_X1 U6247 ( .A(n7362), .B(n5013), .ZN(n7225) );
  OAI21_X2 U6248 ( .B1(n6668), .B2(n4970), .A(n7222), .ZN(n5013) );
  NAND3_X1 U6249 ( .A1(n7227), .A2(n7252), .A3(n7228), .ZN(n7253) );
  OAI21_X1 U6250 ( .B1(n7228), .B2(n5017), .A(n7253), .ZN(n7229) );
  AND2_X4 U6251 ( .A1(n5020), .A2(n5019), .ZN(n6231) );
  NAND2_X1 U6252 ( .A1(n8839), .A2(n5021), .ZN(n5022) );
  NAND2_X1 U6253 ( .A1(n5027), .A2(n4976), .ZN(n5025) );
  NAND2_X1 U6254 ( .A1(n5025), .A2(n8866), .ZN(n8867) );
  NAND2_X1 U6255 ( .A1(n8515), .A2(n7509), .ZN(n7223) );
  NAND3_X1 U6256 ( .A1(n8808), .A2(n8807), .A3(n8809), .ZN(n5035) );
  NAND3_X1 U6257 ( .A1(n8808), .A2(n5040), .A3(n8807), .ZN(n5039) );
  NAND2_X1 U6258 ( .A1(n5042), .A2(n5041), .ZN(n8826) );
  NAND3_X1 U6259 ( .A1(n5045), .A2(n5044), .A3(n5043), .ZN(n8910) );
  NAND2_X1 U6260 ( .A1(n6654), .A2(n5046), .ZN(n5049) );
  NAND2_X1 U6261 ( .A1(n5439), .A2(n5052), .ZN(n5051) );
  AND2_X2 U6262 ( .A1(n9456), .A2(n6899), .ZN(n6904) );
  NAND2_X1 U6263 ( .A1(n5054), .A2(n9453), .ZN(n9456) );
  NAND2_X1 U6264 ( .A1(n9454), .A2(n9451), .ZN(n5054) );
  NAND2_X1 U6265 ( .A1(n5470), .A2(n4980), .ZN(n9454) );
  INV_X1 U6266 ( .A(n6795), .ZN(n5058) );
  NAND2_X1 U6267 ( .A1(n5436), .A2(n5060), .ZN(n8044) );
  NAND3_X1 U6268 ( .A1(n6813), .A2(n6812), .A3(n8041), .ZN(n5060) );
  NAND2_X1 U6269 ( .A1(n5467), .A2(n6768), .ZN(n5063) );
  NAND2_X1 U6270 ( .A1(n7328), .A2(n7326), .ZN(n6784) );
  NOR2_X2 U6271 ( .A1(n9523), .A2(n5452), .ZN(n5064) );
  AND2_X2 U6272 ( .A1(n6907), .A2(n6906), .ZN(n9523) );
  AND3_X1 U6273 ( .A1(n5510), .A2(n5066), .A3(n5523), .ZN(n5551) );
  NAND2_X1 U6274 ( .A1(n5510), .A2(n5523), .ZN(n5968) );
  NAND4_X1 U6275 ( .A1(n5510), .A2(n5523), .A3(n5066), .A4(n5524), .ZN(n5555)
         );
  NAND2_X1 U6276 ( .A1(n10700), .A2(n10662), .ZN(n8452) );
  OAI22_X1 U6277 ( .A1(n5758), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n5759), .B2(
        n7099), .ZN(n5069) );
  NAND2_X1 U6278 ( .A1(n10002), .A2(n5298), .ZN(n9989) );
  NAND2_X1 U6279 ( .A1(n9952), .A2(n8422), .ZN(n5311) );
  NAND2_X1 U6280 ( .A1(n8132), .A2(n5076), .ZN(n5074) );
  OAI21_X1 U6281 ( .B1(n8132), .B2(n5075), .A(n5076), .ZN(n10087) );
  NOR2_X2 U6282 ( .A1(n5354), .A2(n5103), .ZN(n6654) );
  NAND2_X1 U6283 ( .A1(n5129), .A2(n5534), .ZN(n5127) );
  NOR2_X1 U6284 ( .A1(n9903), .A2(n9904), .ZN(n9907) );
  INV_X1 U6285 ( .A(n5151), .ZN(n10065) );
  NAND2_X1 U6286 ( .A1(n5763), .A2(n5156), .ZN(n5161) );
  NAND2_X1 U6287 ( .A1(n7369), .A2(n8239), .ZN(n7368) );
  NAND3_X1 U6288 ( .A1(n5161), .A2(n5160), .A3(n5159), .ZN(n5158) );
  INV_X1 U6289 ( .A(n5159), .ZN(n8237) );
  NAND2_X1 U6290 ( .A1(n5161), .A2(n5160), .ZN(n7315) );
  NAND2_X1 U6291 ( .A1(n10702), .A2(n7393), .ZN(n8448) );
  NAND2_X1 U6292 ( .A1(n5763), .A2(n5762), .ZN(n10686) );
  NAND2_X1 U6293 ( .A1(n8208), .A2(n5171), .ZN(n5170) );
  NAND3_X1 U6294 ( .A1(n5185), .A2(n5587), .A3(SI_1_), .ZN(n5724) );
  NAND2_X1 U6295 ( .A1(n5585), .A2(n5586), .ZN(n5185) );
  NAND2_X1 U6296 ( .A1(n5190), .A2(n5189), .ZN(n8383) );
  NAND4_X1 U6297 ( .A1(n5197), .A2(n8366), .A3(n10033), .A4(n5193), .ZN(n5192)
         );
  OR2_X1 U6298 ( .A1(n7046), .A2(n5997), .ZN(n5787) );
  OAI21_X1 U6299 ( .B1(n8350), .B2(n8349), .A(n5204), .ZN(n5203) );
  INV_X1 U6300 ( .A(n8351), .ZN(n5204) );
  AOI21_X1 U6301 ( .B1(n8444), .B2(n8445), .A(n5205), .ZN(n8513) );
  NOR2_X1 U6302 ( .A1(n5412), .A2(n8404), .ZN(n8408) );
  INV_X1 U6303 ( .A(n8404), .ZN(n5207) );
  NAND2_X1 U6304 ( .A1(n5209), .A2(n8448), .ZN(n8308) );
  NAND3_X1 U6305 ( .A1(n8297), .A2(n8298), .A3(n5210), .ZN(n5209) );
  NAND2_X1 U6306 ( .A1(n8298), .A2(n8297), .ZN(n8456) );
  NAND2_X1 U6307 ( .A1(n7321), .A2(n7056), .ZN(n8298) );
  NAND2_X1 U6308 ( .A1(n8371), .A2(n5212), .ZN(n5211) );
  NAND2_X1 U6309 ( .A1(n5216), .A2(n5414), .ZN(n5413) );
  AOI21_X2 U6310 ( .B1(n5217), .B2(n8395), .A(n8394), .ZN(n8402) );
  INV_X1 U6311 ( .A(n8391), .ZN(n5217) );
  NAND3_X1 U6312 ( .A1(n5779), .A2(n5798), .A3(n5778), .ZN(n5402) );
  AND2_X1 U6313 ( .A1(n5599), .A2(n5600), .ZN(n5764) );
  NAND2_X1 U6314 ( .A1(n5752), .A2(n5594), .ZN(n5765) );
  INV_X1 U6315 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5226) );
  INV_X1 U6316 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5225) );
  NAND3_X1 U6317 ( .A1(n5223), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5222) );
  NAND3_X1 U6318 ( .A1(n5227), .A2(n5226), .A3(n5225), .ZN(n5224) );
  NAND2_X1 U6319 ( .A1(n9254), .A2(n8644), .ZN(n8837) );
  NAND2_X1 U6320 ( .A1(n8902), .A2(n8901), .ZN(n5246) );
  NAND2_X1 U6321 ( .A1(n5250), .A2(n5251), .ZN(n5948) );
  NAND2_X1 U6322 ( .A1(n5424), .A2(n5423), .ZN(n5896) );
  NAND2_X1 U6323 ( .A1(n5813), .A2(n5812), .ZN(n5815) );
  NAND2_X1 U6324 ( .A1(n5813), .A2(n5260), .ZN(n5259) );
  INV_X1 U6325 ( .A(n5613), .ZN(n5267) );
  NOR2_X1 U6326 ( .A1(n5261), .A2(n5263), .ZN(n5260) );
  OAI211_X1 U6327 ( .C1(n8826), .C2(n8825), .A(n8824), .B(n8823), .ZN(n8832)
         );
  INV_X1 U6328 ( .A(n8902), .ZN(n8900) );
  INV_X1 U6329 ( .A(n6231), .ZN(n5393) );
  NAND2_X1 U6330 ( .A1(n5413), .A2(n8499), .ZN(n5412) );
  MUX2_X1 U6331 ( .A(n8311), .B(n8310), .S(n8400), .Z(n8317) );
  OR2_X1 U6332 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  AND2_X1 U6333 ( .A1(n9922), .A2(n6718), .ZN(n6719) );
  NAND2_X1 U6334 ( .A1(n9969), .A2(n8421), .ZN(n9953) );
  NAND2_X1 U6335 ( .A1(n8013), .A2(n8288), .ZN(n8132) );
  NAND2_X1 U6336 ( .A1(n6165), .A2(n8373), .ZN(n10003) );
  NAND2_X1 U6337 ( .A1(n6302), .A2(n6194), .ZN(n5354) );
  NAND2_X1 U6338 ( .A1(n9940), .A2(n10207), .ZN(n9941) );
  NAND2_X1 U6339 ( .A1(n6248), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6340 ( .A1(n6202), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6341 ( .A1(n5314), .A2(n5475), .ZN(n8774) );
  OAI21_X2 U6342 ( .B1(n8735), .B2(n8906), .A(n5272), .ZN(n5274) );
  NAND2_X1 U6343 ( .A1(n5274), .A2(n8910), .ZN(n8911) );
  NAND2_X1 U6344 ( .A1(n6624), .A2(n5276), .ZN(n5275) );
  NAND2_X1 U6345 ( .A1(n5283), .A2(n5281), .ZN(n9197) );
  NAND2_X1 U6346 ( .A1(n9257), .A2(n5282), .ZN(n5281) );
  NAND2_X1 U6347 ( .A1(n9197), .A2(n6634), .ZN(n9198) );
  NAND2_X1 U6348 ( .A1(n5289), .A2(n4977), .ZN(n9082) );
  INV_X1 U6349 ( .A(n5517), .ZN(n5292) );
  NAND2_X1 U6350 ( .A1(n5294), .A2(n5293), .ZN(n8090) );
  NAND2_X1 U6351 ( .A1(n7767), .A2(n5295), .ZN(n7753) );
  NAND2_X2 U6352 ( .A1(n6619), .A2(n8746), .ZN(n7767) );
  NOR2_X2 U6353 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  NAND2_X1 U6354 ( .A1(n9158), .A2(n5297), .ZN(n6637) );
  OR2_X2 U6355 ( .A1(n9156), .A2(n9159), .ZN(n9158) );
  NAND2_X1 U6356 ( .A1(n5304), .A2(n4979), .ZN(n7799) );
  INV_X1 U6357 ( .A(n8247), .ZN(n5306) );
  NAND2_X1 U6358 ( .A1(n7959), .A2(n8250), .ZN(n8029) );
  NAND2_X1 U6359 ( .A1(n6454), .A2(n5316), .ZN(n5315) );
  NAND2_X1 U6360 ( .A1(n7781), .A2(n5328), .ZN(n5326) );
  NAND2_X1 U6361 ( .A1(n6982), .A2(n6696), .ZN(n6699) );
  NAND2_X1 U6362 ( .A1(n6652), .A2(n6615), .ZN(n5341) );
  NAND2_X1 U6363 ( .A1(n5343), .A2(n4978), .ZN(n6561) );
  NAND2_X1 U6364 ( .A1(n8154), .A2(n8148), .ZN(n5346) );
  NAND3_X1 U6365 ( .A1(n6302), .A2(n6196), .A3(n6194), .ZN(n5350) );
  INV_X1 U6366 ( .A(n6235), .ZN(n5361) );
  NAND2_X1 U6367 ( .A1(n5358), .A2(n5356), .ZN(n7511) );
  NAND2_X1 U6368 ( .A1(n5358), .A2(n5355), .ZN(n6259) );
  AOI21_X1 U6369 ( .B1(n5360), .B2(n8772), .A(n5357), .ZN(n5356) );
  OR2_X1 U6370 ( .A1(n7463), .A2(n5359), .ZN(n5358) );
  INV_X1 U6371 ( .A(n5360), .ZN(n5359) );
  NAND2_X1 U6372 ( .A1(n7359), .A2(n8741), .ZN(n6225) );
  NAND2_X1 U6373 ( .A1(n8774), .A2(n7460), .ZN(n8741) );
  INV_X1 U6374 ( .A(n5745), .ZN(n5363) );
  NAND2_X1 U6375 ( .A1(n5366), .A2(n5364), .ZN(n8140) );
  NAND2_X1 U6376 ( .A1(n8024), .A2(n5946), .ZN(n8012) );
  NAND2_X1 U6377 ( .A1(n10032), .A2(n5371), .ZN(n5370) );
  MUX2_X1 U6378 ( .A(n6226), .B(P2_REG1_REG_2__SCAN_IN), .S(n7350), .Z(n7022)
         );
  XNOR2_X2 U6379 ( .A(n5392), .B(n6232), .ZN(n7350) );
  NAND2_X1 U6380 ( .A1(n5402), .A2(n5401), .ZN(n5813) );
  NAND2_X1 U6381 ( .A1(n5405), .A2(n5406), .ZN(n5950) );
  NAND2_X1 U6382 ( .A1(n5918), .A2(n5631), .ZN(n5933) );
  NAND2_X1 U6383 ( .A1(n5996), .A2(n5421), .ZN(n5417) );
  NAND2_X1 U6384 ( .A1(n5996), .A2(n5652), .ZN(n6014) );
  OAI21_X1 U6385 ( .B1(n5996), .B2(n5420), .A(n5418), .ZN(n6046) );
  NAND2_X1 U6386 ( .A1(n5416), .A2(n5415), .ZN(n5659) );
  NAND2_X1 U6387 ( .A1(n5996), .A2(n5418), .ZN(n5416) );
  NAND2_X1 U6388 ( .A1(n5863), .A2(n5624), .ZN(n5878) );
  NOR2_X1 U6389 ( .A1(n5877), .A2(n5426), .ZN(n5425) );
  INV_X1 U6390 ( .A(n5624), .ZN(n5426) );
  NOR2_X1 U6391 ( .A1(n5625), .A2(SI_11_), .ZN(n5428) );
  NAND2_X1 U6392 ( .A1(n5688), .A2(n5687), .ZN(n5691) );
  INV_X1 U6393 ( .A(n7004), .ZN(n6987) );
  NAND2_X1 U6394 ( .A1(n5432), .A2(n6971), .ZN(P1_U3214) );
  NAND2_X1 U6395 ( .A1(n5433), .A2(n9768), .ZN(n5432) );
  NAND2_X1 U6396 ( .A1(n5434), .A2(n7004), .ZN(n5433) );
  NAND2_X1 U6397 ( .A1(n5435), .A2(n6945), .ZN(n5434) );
  INV_X1 U6398 ( .A(n7998), .ZN(n5438) );
  NAND2_X1 U6399 ( .A1(n9513), .A2(n5443), .ZN(n5439) );
  INV_X1 U6400 ( .A(n6774), .ZN(n5462) );
  NAND2_X1 U6401 ( .A1(n5465), .A2(n5467), .ZN(n5464) );
  NAND2_X1 U6402 ( .A1(n9446), .A2(n5472), .ZN(n5470) );
  NAND4_X1 U6403 ( .A1(n5473), .A2(n5101), .A3(n5737), .A4(n5518), .ZN(n5783)
         );
  NAND2_X1 U6404 ( .A1(n5534), .A2(n5533), .ZN(n5537) );
  NAND2_X1 U6405 ( .A1(n7224), .A2(n5475), .ZN(n7227) );
  NAND2_X4 U6406 ( .A1(n6204), .A2(n6206), .ZN(n7572) );
  INV_X2 U6407 ( .A(n6203), .ZN(n6206) );
  INV_X1 U6408 ( .A(n8539), .ZN(n8651) );
  NAND2_X1 U6409 ( .A1(n8611), .A2(n5516), .ZN(n8548) );
  NAND3_X1 U6410 ( .A1(n5479), .A2(n5478), .A3(n8054), .ZN(n5476) );
  NAND2_X1 U6411 ( .A1(n5479), .A2(n8054), .ZN(n7974) );
  INV_X1 U6412 ( .A(n7972), .ZN(n5480) );
  INV_X1 U6413 ( .A(n7973), .ZN(n5481) );
  NAND2_X1 U6414 ( .A1(n8697), .A2(n5485), .ZN(n8588) );
  NAND2_X1 U6415 ( .A1(n8588), .A2(n8573), .ZN(n8576) );
  INV_X1 U6416 ( .A(n5496), .ZN(n8596) );
  NAND3_X1 U6417 ( .A1(n6302), .A2(n6194), .A3(n6195), .ZN(n6455) );
  NAND3_X1 U6418 ( .A1(n5499), .A2(n7738), .A3(n4938), .ZN(n7740) );
  NAND2_X1 U6419 ( .A1(n7634), .A2(n5500), .ZN(n5499) );
  AND2_X1 U6420 ( .A1(n4938), .A2(n5499), .ZN(n7739) );
  INV_X1 U6421 ( .A(n7740), .ZN(n7743) );
  INV_X1 U6422 ( .A(n5740), .ZN(n5742) );
  OR2_X1 U6423 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  OR2_X1 U6424 ( .A1(n7050), .A2(n5727), .ZN(n5728) );
  NOR2_X1 U6425 ( .A1(n7452), .A2(n6668), .ZN(n6974) );
  NAND2_X2 U6426 ( .A1(n6626), .A2(n8830), .ZN(n9257) );
  NOR2_X1 U6427 ( .A1(n6701), .A2(n6700), .ZN(n6704) );
  NAND2_X1 U6428 ( .A1(n10203), .A2(n10757), .ZN(n6722) );
  NOR2_X1 U6429 ( .A1(n8741), .A2(n7223), .ZN(n7456) );
  OAI21_X1 U6430 ( .B1(n10131), .B2(n6183), .A(n4960), .ZN(P1_U3550) );
  INV_X1 U6431 ( .A(n6261), .ZN(n6587) );
  NAND2_X2 U6432 ( .A1(n6207), .A2(n6206), .ZN(n6249) );
  NAND2_X2 U6433 ( .A1(n6207), .A2(n6203), .ZN(n6261) );
  OR2_X1 U6434 ( .A1(n6724), .A2(n6731), .ZN(n5730) );
  OR2_X1 U6435 ( .A1(n5712), .A2(n10238), .ZN(n5759) );
  OAI21_X1 U6436 ( .B1(n10653), .B2(n4926), .A(n6753), .ZN(n6754) );
  OR2_X1 U6437 ( .A1(n6210), .A2(n9406), .ZN(n6209) );
  OR2_X1 U6438 ( .A1(n7539), .A2(n5997), .ZN(n6000) );
  OR2_X1 U6439 ( .A1(n7289), .A2(n5997), .ZN(n5956) );
  OR2_X1 U6440 ( .A1(n7195), .A2(n5997), .ZN(n5922) );
  OR2_X1 U6441 ( .A1(n7160), .A2(n5997), .ZN(n5905) );
  OAI22_X1 U6442 ( .A1(n9167), .A2(n9168), .B1(n9391), .B2(n9325), .ZN(n9156)
         );
  AND2_X1 U6443 ( .A1(n6692), .A2(n6691), .ZN(n10792) );
  NOR2_X1 U6444 ( .A1(n6945), .A2(n6944), .ZN(n5503) );
  AND2_X1 U6445 ( .A1(n6998), .A2(n9768), .ZN(n5504) );
  AND2_X1 U6446 ( .A1(n8340), .A2(n8333), .ZN(n5505) );
  INV_X1 U6447 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6294) );
  INV_X1 U6448 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8147) );
  OR2_X1 U6449 ( .A1(n8106), .A2(n8163), .ZN(n5506) );
  NAND2_X1 U6450 ( .A1(n6957), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5507) );
  AND2_X1 U6451 ( .A1(n6872), .A2(n6871), .ZN(n5508) );
  INV_X1 U6452 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6329) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5582) );
  INV_X1 U6454 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5596) );
  AND2_X1 U6455 ( .A1(n7505), .A2(n9267), .ZN(n9194) );
  INV_X1 U6456 ( .A(n9194), .ZN(n9269) );
  NAND2_X1 U6457 ( .A1(n6490), .A2(n6489), .ZN(n9146) );
  NAND2_X1 U6458 ( .A1(n9488), .A2(n9487), .ZN(n5509) );
  OR2_X1 U6459 ( .A1(n10735), .A2(n7747), .ZN(n5511) );
  INV_X1 U6460 ( .A(n9904), .ZN(n8399) );
  OR2_X1 U6461 ( .A1(n9320), .A2(n9134), .ZN(n5512) );
  NAND2_X1 U6462 ( .A1(n7429), .A2(n7579), .ZN(n7543) );
  INV_X1 U6463 ( .A(n7543), .ZN(n7526) );
  AND2_X1 U6464 ( .A1(n6801), .A2(n6752), .ZN(n5513) );
  NAND2_X2 U6465 ( .A1(n7388), .A2(n10718), .ZN(n10707) );
  AND2_X1 U6466 ( .A1(n8726), .A2(n9331), .ZN(n5514) );
  NOR4_X1 U6467 ( .A1(n9159), .A2(n9184), .A3(n9217), .A4(n8758), .ZN(n5515)
         );
  INV_X1 U6468 ( .A(n10020), .ZN(n10034) );
  AND3_X1 U6469 ( .A1(n8617), .A2(n8610), .A3(n8619), .ZN(n5516) );
  INV_X1 U6470 ( .A(n9506), .ZN(n6891) );
  NAND2_X1 U6471 ( .A1(n9295), .A2(n8570), .ZN(n5517) );
  NAND2_X1 U6472 ( .A1(n5691), .A2(n5690), .ZN(n6575) );
  INV_X1 U6473 ( .A(n6575), .ZN(n5692) );
  INV_X1 U6474 ( .A(n10632), .ZN(n8235) );
  INV_X1 U6475 ( .A(n8894), .ZN(n8891) );
  NAND2_X1 U6476 ( .A1(n9285), .A2(n5034), .ZN(n8888) );
  NAND2_X1 U6477 ( .A1(n8889), .A2(n8888), .ZN(n8894) );
  NOR2_X1 U6478 ( .A1(n8733), .A2(n9369), .ZN(n8728) );
  NOR2_X1 U6479 ( .A1(n8904), .A2(n5034), .ZN(n8905) );
  AND2_X1 U6480 ( .A1(n8898), .A2(n8738), .ZN(n8901) );
  NOR2_X1 U6481 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6196) );
  INV_X1 U6482 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6185) );
  INV_X1 U6483 ( .A(n6750), .ZN(n6745) );
  INV_X1 U6484 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5694) );
  INV_X1 U6485 ( .A(n9103), .ZN(n8570) );
  INV_X1 U6486 ( .A(n9146), .ZN(n8559) );
  INV_X1 U6487 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6184) );
  OR2_X1 U6488 ( .A1(n9904), .A2(n8406), .ZN(n8401) );
  INV_X1 U6489 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5972) );
  INV_X1 U6490 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U6491 ( .A1(n7524), .A2(n7523), .ZN(n7532) );
  INV_X1 U6492 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9708) );
  INV_X1 U6493 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6594) );
  AND2_X1 U6494 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5789) );
  INV_X1 U6495 ( .A(n7247), .ZN(n6768) );
  INV_X1 U6496 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5923) );
  NOR2_X1 U6497 ( .A1(n6049), .A2(n9459), .ZN(n6062) );
  INV_X1 U6498 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U6499 ( .A1(n4928), .A2(n8397), .ZN(n8398) );
  AND2_X1 U6500 ( .A1(n5869), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5884) );
  INV_X1 U6501 ( .A(n10135), .ZN(n6177) );
  INV_X1 U6502 ( .A(n8293), .ZN(n8463) );
  INV_X1 U6503 ( .A(n5555), .ZN(n5526) );
  NAND2_X1 U6504 ( .A1(n6576), .A2(n5692), .ZN(n6580) );
  INV_X1 U6505 ( .A(SI_26_), .ZN(n9658) );
  NAND2_X1 U6506 ( .A1(n8550), .A2(n9315), .ZN(n8551) );
  OR2_X1 U6507 ( .A1(n5034), .A2(n6977), .ZN(n7197) );
  INV_X1 U6508 ( .A(n6631), .ZN(n6632) );
  AND2_X1 U6509 ( .A1(n8726), .A2(n9386), .ZN(n6694) );
  INV_X1 U6510 ( .A(n7999), .ZN(n6818) );
  OR2_X1 U6511 ( .A1(n5924), .A2(n5923), .ZN(n5939) );
  NAND2_X1 U6512 ( .A1(n5884), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5907) );
  AND2_X1 U6513 ( .A1(n6110), .A2(n6096), .ZN(n9996) );
  NAND2_X1 U6514 ( .A1(n6018), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6035) );
  INV_X1 U6515 ( .A(n8135), .ZN(n8211) );
  AND2_X1 U6516 ( .A1(n5544), .A2(n5543), .ZN(n5545) );
  AND2_X1 U6517 ( .A1(n5677), .A2(n5676), .ZN(n6088) );
  NAND2_X1 U6518 ( .A1(n5553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5554) );
  OR2_X1 U6519 ( .A1(n5902), .A2(n5901), .ZN(n5919) );
  NAND2_X1 U6520 ( .A1(n8531), .A2(n9262), .ZN(n8532) );
  NAND2_X1 U6521 ( .A1(n6526), .A2(n9720), .ZN(n6539) );
  NAND2_X1 U6522 ( .A1(n7232), .A2(n7231), .ZN(n8700) );
  INV_X1 U6523 ( .A(n7821), .ZN(n7816) );
  INV_X1 U6524 ( .A(n7009), .ZN(n7014) );
  OR2_X1 U6525 ( .A1(n6565), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8522) );
  OAI21_X1 U6526 ( .B1(n6647), .B2(n6646), .A(n8896), .ZN(n6648) );
  INV_X1 U6527 ( .A(n9326), .ZN(n9134) );
  INV_X1 U6528 ( .A(n9212), .ZN(n9230) );
  NAND2_X1 U6529 ( .A1(n7513), .A2(n7585), .ZN(n8785) );
  INV_X1 U6530 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6983) );
  OR3_X1 U6531 ( .A1(n7506), .A2(n10777), .A3(n6651), .ZN(n7486) );
  INV_X1 U6532 ( .A(n8824), .ZN(n8756) );
  INV_X1 U6533 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6198) );
  INV_X1 U6534 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9425) );
  INV_X1 U6535 ( .A(n6757), .ZN(n7141) );
  OR2_X1 U6536 ( .A1(n9754), .A2(n9755), .ZN(n6934) );
  AND4_X1 U6537 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n9517)
         );
  NAND2_X1 U6538 ( .A1(n4927), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5720) );
  INV_X1 U6539 ( .A(n10245), .ZN(n9810) );
  INV_X1 U6540 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7330) );
  OR2_X1 U6541 ( .A1(n10369), .A2(n10245), .ZN(n10451) );
  INV_X1 U6542 ( .A(n10607), .ZN(n9978) );
  NAND2_X1 U6543 ( .A1(n8296), .A2(n8304), .ZN(n10651) );
  NAND2_X1 U6544 ( .A1(n6725), .A2(n8234), .ZN(n10688) );
  INV_X1 U6545 ( .A(n8354), .ZN(n8209) );
  OR2_X1 U6546 ( .A1(n8436), .A2(n9810), .ZN(n10701) );
  OR2_X1 U6547 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  INV_X1 U6548 ( .A(n8700), .ZN(n8710) );
  AND2_X1 U6549 ( .A1(n6572), .A2(n6571), .ZN(n9285) );
  INV_X1 U6550 ( .A(n10566), .ZN(n9008) );
  INV_X1 U6551 ( .A(n10563), .ZN(n10564) );
  INV_X1 U6552 ( .A(n9064), .ZN(n10578) );
  NAND2_X1 U6553 ( .A1(n6649), .A2(n6648), .ZN(n8527) );
  INV_X1 U6554 ( .A(n9316), .ZN(n9335) );
  INV_X1 U6555 ( .A(n9267), .ZN(n9188) );
  NAND2_X1 U6556 ( .A1(n7213), .A2(n7212), .ZN(n9267) );
  INV_X1 U6557 ( .A(n9269), .ZN(n9189) );
  OR2_X1 U6558 ( .A1(n6974), .A2(n6973), .ZN(n7448) );
  AND2_X1 U6559 ( .A1(n7486), .A2(n7282), .ZN(n10787) );
  INV_X1 U6560 ( .A(n10787), .ZN(n10775) );
  OR2_X1 U6561 ( .A1(n7211), .A2(n7215), .ZN(n6691) );
  OAI21_X1 U6562 ( .B1(n10207), .B2(n9779), .A(n6969), .ZN(n6970) );
  AND2_X1 U6563 ( .A1(n6101), .A2(n6100), .ZN(n9974) );
  AND4_X1 U6564 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n6822)
         );
  INV_X1 U6565 ( .A(n10496), .ZN(n10587) );
  INV_X1 U6566 ( .A(n10451), .ZN(n10595) );
  INV_X1 U6567 ( .A(n10492), .ZN(n10591) );
  INV_X1 U6568 ( .A(n10670), .ZN(n10081) );
  AND2_X1 U6569 ( .A1(n10707), .A2(n10713), .ZN(n10016) );
  INV_X1 U6570 ( .A(n9915), .ZN(n10709) );
  NAND2_X1 U6571 ( .A1(n8405), .A2(n6166), .ZN(n10659) );
  INV_X1 U6572 ( .A(n10606), .ZN(n10193) );
  INV_X1 U6573 ( .A(n10750), .ZN(n10663) );
  NAND2_X1 U6574 ( .A1(n10655), .A2(n10665), .ZN(n10754) );
  INV_X1 U6575 ( .A(n5572), .ZN(n10231) );
  INV_X1 U6576 ( .A(n6729), .ZN(n6957) );
  INV_X1 U6577 ( .A(n7086), .ZN(n7011) );
  NAND2_X1 U6578 ( .A1(n7209), .A2(n7208), .ZN(n8691) );
  INV_X1 U6579 ( .A(n8689), .ZN(n8719) );
  OR2_X1 U6580 ( .A1(P2_U3150), .A2(n7017), .ZN(n10563) );
  NAND2_X1 U6581 ( .A1(n7489), .A2(n7488), .ZN(n9265) );
  INV_X1 U6582 ( .A(n9331), .ZN(n9362) );
  NOR2_X1 U6583 ( .A1(n6694), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U6584 ( .A1(n6693), .A2(n7213), .ZN(n9403) );
  NAND2_X1 U6585 ( .A1(n7206), .A2(n7069), .ZN(n7080) );
  INV_X1 U6586 ( .A(n7927), .ZN(n7987) );
  INV_X1 U6587 ( .A(n6970), .ZN(n6971) );
  INV_X1 U6588 ( .A(n9768), .ZN(n9541) );
  INV_X1 U6589 ( .A(n9926), .ZN(n9954) );
  INV_X1 U6590 ( .A(n9974), .ZN(n10005) );
  INV_X1 U6591 ( .A(n6822), .ZN(n9792) );
  INV_X1 U6592 ( .A(n7610), .ZN(n9795) );
  INV_X1 U6593 ( .A(n10585), .ZN(n10491) );
  INV_X1 U6594 ( .A(n10016), .ZN(n10094) );
  OR2_X1 U6595 ( .A1(n10362), .A2(n6954), .ZN(n10718) );
  AND2_X2 U6596 ( .A1(n6181), .A2(n5576), .ZN(n10757) );
  INV_X1 U6597 ( .A(n9947), .ZN(n10207) );
  NAND2_X1 U6598 ( .A1(n10761), .A2(n10663), .ZN(n10220) );
  INV_X1 U6599 ( .A(n10761), .ZN(n10758) );
  AND2_X2 U6600 ( .A1(n6181), .A2(n7383), .ZN(n10761) );
  NOR2_X1 U6601 ( .A1(n10362), .A2(n10231), .ZN(n10269) );
  INV_X1 U6602 ( .A(n10241), .ZN(n7593) );
  INV_X2 U6603 ( .A(n9799), .ZN(P1_U3973) );
  NAND2_X1 U6604 ( .A1(n6722), .A2(n6721), .ZN(P1_U3551) );
  INV_X2 U6605 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U6606 ( .A(n5783), .ZN(n5523) );
  NOR2_X1 U6607 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5521) );
  NOR2_X1 U6608 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5520) );
  NOR2_X1 U6609 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5519) );
  INV_X1 U6610 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6611 ( .A1(n5549), .A2(n5548), .ZN(n5527) );
  NAND2_X1 U6612 ( .A1(n5527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5528) );
  NOR2_X1 U6613 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5532) );
  NOR2_X1 U6614 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5531) );
  NOR2_X1 U6615 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5530) );
  NOR2_X1 U6616 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5529) );
  INV_X1 U6617 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5535) );
  OR2_X1 U6618 ( .A1(n5697), .A2(n5695), .ZN(n5536) );
  NAND2_X1 U6619 ( .A1(n5539), .A2(n5536), .ZN(n5546) );
  NAND2_X1 U6620 ( .A1(n5537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5538) );
  NOR2_X1 U6621 ( .A1(n5546), .A2(n5574), .ZN(n5541) );
  NAND2_X2 U6622 ( .A1(n5541), .A2(n5542), .ZN(n6729) );
  NAND3_X1 U6623 ( .A1(n5546), .A2(P1_B_REG_SCAN_IN), .A3(n5574), .ZN(n5544)
         );
  NAND2_X1 U6624 ( .A1(n5542), .A2(n5545), .ZN(n5572) );
  INV_X1 U6625 ( .A(n5546), .ZN(n8129) );
  OAI22_X1 U6626 ( .A1(n5572), .A2(P1_D_REG_1__SCAN_IN), .B1(n5542), .B2(n8129), .ZN(n6948) );
  INV_X1 U6627 ( .A(n6948), .ZN(n5547) );
  NOR2_X1 U6628 ( .A1(n10362), .A2(n5547), .ZN(n10360) );
  XNOR2_X1 U6629 ( .A(n5549), .B(n5548), .ZN(n6725) );
  NAND2_X1 U6630 ( .A1(n5558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5550) );
  INV_X1 U6631 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6632 ( .A1(n5998), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U6633 ( .A1(n5555), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5556) );
  MUX2_X1 U6634 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5556), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5557) );
  OR2_X1 U6635 ( .A1(n8436), .A2(n10692), .ZN(n7384) );
  INV_X1 U6636 ( .A(n6726), .ZN(n8234) );
  OR2_X1 U6637 ( .A1(n10688), .A2(n9978), .ZN(n6954) );
  NOR4_X1 U6638 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5562) );
  NOR4_X1 U6639 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5561) );
  NOR4_X1 U6640 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5560) );
  NOR4_X1 U6641 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5559) );
  NAND4_X1 U6642 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n5568)
         );
  NOR2_X1 U6643 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n5566) );
  NOR4_X1 U6644 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5565) );
  NOR4_X1 U6645 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5564) );
  NOR4_X1 U6646 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5563) );
  NAND4_X1 U6647 ( .A1(n5566), .A2(n5565), .A3(n5564), .A4(n5563), .ZN(n5567)
         );
  NOR2_X1 U6648 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  NOR2_X1 U6649 ( .A1(n5572), .A2(n5569), .ZN(n6947) );
  INV_X1 U6650 ( .A(n6947), .ZN(n5570) );
  AND3_X1 U6651 ( .A1(n7384), .A2(n6954), .A3(n5570), .ZN(n5571) );
  AND2_X1 U6652 ( .A1(n10360), .A2(n5571), .ZN(n6181) );
  INV_X1 U6653 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6654 ( .A1(n10231), .A2(n5573), .ZN(n5575) );
  INV_X1 U6655 ( .A(n5574), .ZN(n8010) );
  OR2_X1 U6656 ( .A1(n5542), .A2(n8010), .ZN(n10232) );
  INV_X1 U6657 ( .A(n7383), .ZN(n5576) );
  NAND2_X1 U6658 ( .A1(n10757), .A2(n10663), .ZN(n10131) );
  MUX2_X1 U6659 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5701), .Z(n5577) );
  NAND2_X1 U6660 ( .A1(n5577), .A2(SI_2_), .ZN(n5589) );
  OAI21_X1 U6661 ( .B1(n5577), .B2(SI_2_), .A(n5589), .ZN(n5741) );
  INV_X1 U6662 ( .A(n5741), .ZN(n5588) );
  INV_X1 U6663 ( .A(n5586), .ZN(n5583) );
  NAND2_X1 U6664 ( .A1(n5579), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U6665 ( .A1(n5583), .A2(n5584), .ZN(n5587) );
  INV_X1 U6666 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U6667 ( .A1(n5724), .A2(n5587), .ZN(n5740) );
  NAND2_X1 U6668 ( .A1(n5588), .A2(n5740), .ZN(n5743) );
  NAND2_X1 U6669 ( .A1(n5743), .A2(n5589), .ZN(n5750) );
  MUX2_X1 U6670 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7036), .Z(n5590) );
  NAND2_X1 U6671 ( .A1(n5590), .A2(SI_3_), .ZN(n5594) );
  INV_X1 U6672 ( .A(n5590), .ZN(n5592) );
  INV_X1 U6673 ( .A(SI_3_), .ZN(n5591) );
  NAND2_X1 U6674 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  AND2_X1 U6675 ( .A1(n5594), .A2(n5593), .ZN(n5749) );
  NAND2_X1 U6676 ( .A1(n5750), .A2(n5749), .ZN(n5752) );
  INV_X1 U6677 ( .A(SI_4_), .ZN(n5597) );
  NAND2_X1 U6678 ( .A1(n5598), .A2(n5597), .ZN(n5599) );
  INV_X1 U6679 ( .A(SI_5_), .ZN(n5601) );
  NAND2_X1 U6680 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  AND2_X1 U6681 ( .A1(n5604), .A2(n5603), .ZN(n5778) );
  MUX2_X1 U6682 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5700), .Z(n5605) );
  NAND2_X1 U6683 ( .A1(n5605), .A2(SI_6_), .ZN(n5608) );
  INV_X1 U6684 ( .A(n5605), .ZN(n5606) );
  INV_X1 U6685 ( .A(SI_6_), .ZN(n9685) );
  NAND2_X1 U6686 ( .A1(n5606), .A2(n9685), .ZN(n5607) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5700), .Z(n5609) );
  NAND2_X1 U6688 ( .A1(n5609), .A2(SI_7_), .ZN(n5613) );
  INV_X1 U6689 ( .A(n5609), .ZN(n5611) );
  INV_X1 U6690 ( .A(SI_7_), .ZN(n5610) );
  NAND2_X1 U6691 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  MUX2_X1 U6692 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5700), .Z(n5614) );
  XNOR2_X1 U6693 ( .A(n5614), .B(SI_8_), .ZN(n5828) );
  INV_X1 U6694 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U6695 ( .A1(n5615), .A2(n9683), .ZN(n5616) );
  MUX2_X1 U6696 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7036), .Z(n5618) );
  INV_X1 U6697 ( .A(SI_9_), .ZN(n5617) );
  XNOR2_X1 U6698 ( .A(n5618), .B(n5617), .ZN(n5843) );
  MUX2_X1 U6699 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7036), .Z(n5619) );
  NAND2_X1 U6700 ( .A1(n5619), .A2(SI_10_), .ZN(n5624) );
  INV_X1 U6701 ( .A(n5619), .ZN(n5621) );
  INV_X1 U6702 ( .A(SI_10_), .ZN(n5620) );
  NAND2_X1 U6703 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U6704 ( .A1(n5624), .A2(n5622), .ZN(n5860) );
  INV_X1 U6705 ( .A(n5860), .ZN(n5623) );
  NAND2_X1 U6706 ( .A1(n5859), .A2(n5623), .ZN(n5863) );
  MUX2_X1 U6707 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7036), .Z(n5625) );
  XNOR2_X1 U6708 ( .A(n5625), .B(SI_11_), .ZN(n5877) );
  MUX2_X1 U6709 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7036), .Z(n5626) );
  NAND2_X1 U6710 ( .A1(n5626), .A2(SI_12_), .ZN(n5627) );
  OAI21_X1 U6711 ( .B1(n5626), .B2(SI_12_), .A(n5627), .ZN(n5894) );
  MUX2_X1 U6712 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5700), .Z(n5628) );
  NAND2_X1 U6713 ( .A1(n5628), .A2(SI_13_), .ZN(n5631) );
  INV_X1 U6714 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U6715 ( .A1(n5629), .A2(n9674), .ZN(n5630) );
  MUX2_X1 U6716 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5700), .Z(n5632) );
  NAND2_X1 U6717 ( .A1(n5632), .A2(SI_14_), .ZN(n5635) );
  INV_X1 U6718 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U6719 ( .A1(n5633), .A2(n9671), .ZN(n5634) );
  MUX2_X1 U6720 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5700), .Z(n5636) );
  NAND2_X1 U6721 ( .A1(n5636), .A2(SI_15_), .ZN(n5640) );
  INV_X1 U6722 ( .A(n5636), .ZN(n5638) );
  INV_X1 U6723 ( .A(SI_15_), .ZN(n5637) );
  NAND2_X1 U6724 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U6725 ( .A1(n5950), .A2(n5640), .ZN(n5967) );
  MUX2_X1 U6726 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5700), .Z(n5641) );
  XNOR2_X1 U6727 ( .A(n5641), .B(SI_16_), .ZN(n5966) );
  INV_X1 U6728 ( .A(n5641), .ZN(n5643) );
  INV_X1 U6729 ( .A(SI_16_), .ZN(n5642) );
  NAND2_X1 U6730 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  OAI21_X1 U6731 ( .B1(n5967), .B2(n5966), .A(n5644), .ZN(n5980) );
  MUX2_X1 U6732 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5700), .Z(n5646) );
  NOR2_X1 U6733 ( .A1(n5646), .A2(SI_17_), .ZN(n5647) );
  AOI21_X1 U6734 ( .B1(n5980), .B2(n5981), .A(n5647), .ZN(n5992) );
  MUX2_X1 U6735 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5700), .Z(n5648) );
  NAND2_X1 U6736 ( .A1(n5648), .A2(SI_18_), .ZN(n5652) );
  INV_X1 U6737 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U6738 ( .A1(n5649), .A2(n9652), .ZN(n5650) );
  NAND2_X1 U6739 ( .A1(n5652), .A2(n5650), .ZN(n5993) );
  INV_X1 U6740 ( .A(n5993), .ZN(n5651) );
  NAND2_X1 U6741 ( .A1(n5992), .A2(n5651), .ZN(n5996) );
  MUX2_X1 U6742 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n5700), .Z(n5653) );
  XNOR2_X1 U6743 ( .A(n5653), .B(SI_19_), .ZN(n6013) );
  INV_X1 U6744 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U6745 ( .A1(n5654), .A2(n9557), .ZN(n5655) );
  MUX2_X1 U6746 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5700), .Z(n6030) );
  NAND2_X1 U6747 ( .A1(n6030), .A2(SI_20_), .ZN(n5656) );
  MUX2_X1 U6748 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5700), .Z(n5657) );
  XNOR2_X1 U6749 ( .A(n5657), .B(SI_21_), .ZN(n6045) );
  NAND2_X1 U6750 ( .A1(n5657), .A2(SI_21_), .ZN(n5658) );
  NAND2_X1 U6751 ( .A1(n5659), .A2(n5658), .ZN(n6059) );
  INV_X1 U6752 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5660) );
  MUX2_X1 U6753 ( .A(n7910), .B(n5660), .S(n5700), .Z(n5662) );
  INV_X1 U6754 ( .A(SI_22_), .ZN(n5661) );
  NAND2_X1 U6755 ( .A1(n5662), .A2(n5661), .ZN(n5665) );
  INV_X1 U6756 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U6757 ( .A1(n5663), .A2(SI_22_), .ZN(n5664) );
  NAND2_X1 U6758 ( .A1(n5665), .A2(n5664), .ZN(n6058) );
  INV_X1 U6759 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5667) );
  INV_X1 U6760 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5666) );
  MUX2_X1 U6761 ( .A(n5667), .B(n5666), .S(n5700), .Z(n5668) );
  INV_X1 U6762 ( .A(SI_23_), .ZN(n9559) );
  NAND2_X1 U6763 ( .A1(n5668), .A2(n9559), .ZN(n5671) );
  INV_X1 U6764 ( .A(n5668), .ZN(n5669) );
  NAND2_X1 U6765 ( .A1(n5669), .A2(SI_23_), .ZN(n5670) );
  INV_X1 U6766 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8518) );
  INV_X1 U6767 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5672) );
  MUX2_X1 U6768 ( .A(n8518), .B(n5672), .S(n5700), .Z(n5674) );
  INV_X1 U6769 ( .A(SI_24_), .ZN(n5673) );
  NAND2_X1 U6770 ( .A1(n5674), .A2(n5673), .ZN(n5677) );
  INV_X1 U6771 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U6772 ( .A1(n5675), .A2(SI_24_), .ZN(n5676) );
  INV_X1 U6773 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5678) );
  MUX2_X1 U6774 ( .A(n8147), .B(n5678), .S(n5700), .Z(n5679) );
  NAND2_X1 U6775 ( .A1(n5679), .A2(n9657), .ZN(n5682) );
  INV_X1 U6776 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U6777 ( .A1(n5680), .A2(SI_25_), .ZN(n5681) );
  INV_X1 U6778 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8203) );
  INV_X1 U6779 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5683) );
  MUX2_X1 U6780 ( .A(n8203), .B(n5683), .S(n5700), .Z(n5684) );
  NAND2_X1 U6781 ( .A1(n5684), .A2(n9658), .ZN(n5687) );
  INV_X1 U6782 ( .A(n5684), .ZN(n5685) );
  NAND2_X1 U6783 ( .A1(n5685), .A2(SI_26_), .ZN(n5686) );
  INV_X1 U6784 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9416) );
  INV_X1 U6785 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5689) );
  MUX2_X1 U6786 ( .A(n9416), .B(n5689), .S(n5700), .Z(n5690) );
  MUX2_X1 U6787 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7036), .Z(n6577) );
  XNOR2_X1 U6788 ( .A(n6577), .B(n9571), .ZN(n6576) );
  NAND2_X1 U6789 ( .A1(n5695), .A2(n5694), .ZN(n5704) );
  NAND2_X1 U6790 ( .A1(n5704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5696) );
  INV_X1 U6791 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6792 ( .A1(n8230), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5702) );
  INV_X1 U6793 ( .A(n5704), .ZN(n5706) );
  INV_X1 U6794 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5707) );
  NAND2_X2 U6795 ( .A1(n10238), .A2(n5712), .ZN(n6025) );
  NAND2_X1 U6796 ( .A1(n4927), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5717) );
  INV_X1 U6797 ( .A(n10238), .ZN(n5711) );
  INV_X1 U6798 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10605) );
  INV_X1 U6799 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5713) );
  INV_X1 U6800 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10365) );
  NOR2_X1 U6801 ( .A1(n5701), .A2(n9697), .ZN(n5718) );
  XNOR2_X1 U6802 ( .A(n5718), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10250) );
  MUX2_X1 U6803 ( .A(n10365), .B(n10250), .S(n7050), .Z(n10606) );
  NAND2_X1 U6804 ( .A1(n5757), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5722) );
  INV_X1 U6805 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7158) );
  INV_X1 U6806 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7096) );
  OR2_X1 U6807 ( .A1(n5759), .A2(n7096), .ZN(n5719) );
  INV_X1 U6808 ( .A(SI_1_), .ZN(n9691) );
  NAND2_X1 U6809 ( .A1(n4969), .A2(n9691), .ZN(n5723) );
  AND2_X1 U6810 ( .A1(n5724), .A2(n5723), .ZN(n6214) );
  INV_X1 U6811 ( .A(n6214), .ZN(n8520) );
  NAND2_X1 U6812 ( .A1(n5725), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6813 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5726) );
  XNOR2_X1 U6814 ( .A(n5726), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9805) );
  INV_X1 U6815 ( .A(n9805), .ZN(n5727) );
  OAI211_X2 U6816 ( .C1(n5997), .C2(n8520), .A(n5729), .B(n5728), .ZN(n6731)
         );
  XNOR2_X1 U6817 ( .A(n6724), .B(n6731), .ZN(n10187) );
  OAI21_X1 U6818 ( .B1(n10185), .B2(n10187), .A(n5730), .ZN(n10625) );
  NAND2_X1 U6819 ( .A1(n4927), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5736) );
  INV_X1 U6820 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9817) );
  INV_X1 U6821 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5731) );
  OR2_X1 U6822 ( .A1(n5836), .A2(n5731), .ZN(n5734) );
  INV_X1 U6823 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5732) );
  OR2_X1 U6824 ( .A1(n5759), .A2(n5732), .ZN(n5733) );
  NAND4_X1 U6825 ( .A1(n5736), .A2(n5735), .A3(n5734), .A4(n5733), .ZN(n5746)
         );
  INV_X1 U6826 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7037) );
  OR2_X1 U6827 ( .A1(n5737), .A2(n10233), .ZN(n5739) );
  INV_X1 U6828 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U6829 ( .A1(n5739), .A2(n5738), .ZN(n5753) );
  OAI21_X1 U6830 ( .B1(n5739), .B2(n5738), .A(n5753), .ZN(n7114) );
  OAI22_X1 U6831 ( .A1(n5768), .A2(n7037), .B1(n7050), .B2(n7114), .ZN(n5745)
         );
  NAND2_X1 U6832 ( .A1(n5742), .A2(n5741), .ZN(n5744) );
  NAND2_X1 U6833 ( .A1(n5744), .A2(n5743), .ZN(n7040) );
  INV_X1 U6834 ( .A(n5746), .ZN(n10653) );
  NAND2_X1 U6835 ( .A1(n6752), .A2(n10653), .ZN(n8304) );
  NAND2_X1 U6836 ( .A1(n10625), .A2(n10632), .ZN(n5748) );
  NAND2_X1 U6837 ( .A1(n10653), .A2(n10628), .ZN(n5747) );
  NAND2_X1 U6838 ( .A1(n5748), .A2(n5747), .ZN(n10649) );
  OR2_X1 U6839 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  NAND2_X1 U6840 ( .A1(n5752), .A2(n5751), .ZN(n7041) );
  OR2_X1 U6841 ( .A1(n7041), .A2(n5997), .ZN(n5756) );
  NAND2_X1 U6842 ( .A1(n5753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U6843 ( .A(n5754), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U6844 ( .A1(n8230), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6015), .B2(
        n9833), .ZN(n5755) );
  NAND2_X2 U6845 ( .A1(n5756), .A2(n5755), .ZN(n10662) );
  INV_X1 U6846 ( .A(n10662), .ZN(n10669) );
  NAND2_X1 U6847 ( .A1(n5757), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5761) );
  INV_X1 U6848 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7118) );
  OR2_X1 U6849 ( .A1(n6025), .A2(n7118), .ZN(n5760) );
  INV_X1 U6850 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U6851 ( .A1(n10669), .A2(n9798), .ZN(n8454) );
  NAND2_X1 U6852 ( .A1(n8454), .A2(n8452), .ZN(n6161) );
  NAND2_X1 U6853 ( .A1(n10649), .A2(n6161), .ZN(n5763) );
  NAND2_X1 U6854 ( .A1(n10700), .A2(n10669), .ZN(n5762) );
  OR2_X1 U6855 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NAND2_X1 U6856 ( .A1(n5767), .A2(n5766), .ZN(n7044) );
  OR2_X1 U6857 ( .A1(n7044), .A2(n5997), .ZN(n5772) );
  INV_X2 U6858 ( .A(n5768), .ZN(n8274) );
  NOR2_X1 U6859 ( .A1(n5770), .A2(n5769), .ZN(n10594) );
  AOI22_X1 U6860 ( .A1(n8274), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6015), .B2(
        n10594), .ZN(n5771) );
  NAND2_X1 U6861 ( .A1(n5757), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5776) );
  XNOR2_X1 U6862 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10719) );
  OR2_X1 U6863 ( .A1(n5758), .A2(n10719), .ZN(n5775) );
  INV_X1 U6864 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10706) );
  OR2_X1 U6865 ( .A1(n6025), .A2(n10706), .ZN(n5774) );
  INV_X1 U6866 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7101) );
  OR2_X1 U6867 ( .A1(n5759), .A2(n7101), .ZN(n5773) );
  NAND4_X1 U6868 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n9797)
         );
  AND2_X1 U6869 ( .A1(n10689), .A2(n10654), .ZN(n5777) );
  NOR2_X1 U6870 ( .A1(n5769), .A2(n10233), .ZN(n5781) );
  MUX2_X1 U6871 ( .A(n10233), .B(n5781), .S(P1_IR_REG_5__SCAN_IN), .Z(n5782)
         );
  INV_X1 U6872 ( .A(n5782), .ZN(n5785) );
  AND2_X1 U6873 ( .A1(n5785), .A2(n5784), .ZN(n10378) );
  AOI22_X1 U6874 ( .A1(n8274), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6015), .B2(
        n10378), .ZN(n5786) );
  AND2_X2 U6875 ( .A1(n5787), .A2(n5786), .ZN(n7321) );
  NAND2_X1 U6876 ( .A1(n5757), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5796) );
  INV_X1 U6877 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5788) );
  OR2_X1 U6878 ( .A1(n5759), .A2(n5788), .ZN(n5795) );
  NAND2_X1 U6879 ( .A1(n5789), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5805) );
  INV_X1 U6880 ( .A(n5789), .ZN(n5791) );
  INV_X1 U6881 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6882 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NAND2_X1 U6883 ( .A1(n5805), .A2(n5792), .ZN(n7389) );
  OR2_X1 U6884 ( .A1(n5758), .A2(n7389), .ZN(n5794) );
  INV_X1 U6885 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7390) );
  OR2_X1 U6886 ( .A1(n6025), .A2(n7390), .ZN(n5793) );
  NAND4_X1 U6887 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n7056)
         );
  NAND2_X1 U6888 ( .A1(n7321), .A2(n10702), .ZN(n5797) );
  OR2_X1 U6889 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  NAND2_X1 U6890 ( .A1(n5801), .A2(n5800), .ZN(n7048) );
  OR2_X1 U6891 ( .A1(n7048), .A2(n5997), .ZN(n5804) );
  NAND2_X1 U6892 ( .A1(n5784), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U6893 ( .A(n5802), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U6894 ( .A1(n8274), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6015), .B2(
        n10393), .ZN(n5803) );
  NAND2_X1 U6895 ( .A1(n5757), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5810) );
  INV_X1 U6896 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7103) );
  OR2_X1 U6897 ( .A1(n7060), .A2(n7103), .ZN(n5809) );
  NOR2_X1 U6898 ( .A1(n5805), .A2(n7330), .ZN(n5819) );
  INV_X1 U6899 ( .A(n5819), .ZN(n5821) );
  NAND2_X1 U6900 ( .A1(n5805), .A2(n7330), .ZN(n5806) );
  NAND2_X1 U6901 ( .A1(n5821), .A2(n5806), .ZN(n7415) );
  OR2_X1 U6902 ( .A1(n5758), .A2(n7415), .ZN(n5808) );
  INV_X1 U6903 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7113) );
  OR2_X1 U6904 ( .A1(n6025), .A2(n7113), .ZN(n5807) );
  OR2_X1 U6905 ( .A1(n7418), .A2(n7479), .ZN(n8316) );
  INV_X1 U6906 ( .A(n7479), .ZN(n7296) );
  OR2_X1 U6907 ( .A1(n7418), .A2(n7296), .ZN(n5811) );
  OR2_X1 U6908 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U6909 ( .A1(n5815), .A2(n5814), .ZN(n7055) );
  OR2_X1 U6910 ( .A1(n7055), .A2(n5997), .ZN(n5818) );
  OR2_X1 U6911 ( .A1(n5784), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U6912 ( .A1(n5830), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5816) );
  XNOR2_X1 U6913 ( .A(n5816), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U6914 ( .A1(n8274), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6015), .B2(
        n10406), .ZN(n5817) );
  NAND2_X1 U6915 ( .A1(n5818), .A2(n5817), .ZN(n7445) );
  NAND2_X1 U6916 ( .A1(n5757), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5826) );
  INV_X1 U6917 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7105) );
  OR2_X1 U6918 ( .A1(n7060), .A2(n7105), .ZN(n5825) );
  NAND2_X1 U6919 ( .A1(n5819), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5834) );
  INV_X1 U6920 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U6921 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND2_X1 U6922 ( .A1(n5834), .A2(n5822), .ZN(n7480) );
  OR2_X1 U6923 ( .A1(n5758), .A2(n7480), .ZN(n5824) );
  INV_X1 U6924 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7407) );
  OR2_X1 U6925 ( .A1(n6025), .A2(n7407), .ZN(n5823) );
  OR2_X1 U6926 ( .A1(n7445), .A2(n7688), .ZN(n8320) );
  AND2_X1 U6927 ( .A1(n7445), .A2(n7688), .ZN(n8313) );
  INV_X1 U6928 ( .A(n8313), .ZN(n8319) );
  INV_X1 U6929 ( .A(n8242), .ZN(n7552) );
  NAND2_X1 U6930 ( .A1(n7405), .A2(n7552), .ZN(n7404) );
  INV_X1 U6931 ( .A(n7688), .ZN(n9796) );
  OR2_X1 U6932 ( .A1(n7445), .A2(n9796), .ZN(n5827) );
  NAND2_X1 U6933 ( .A1(n7404), .A2(n5827), .ZN(n7595) );
  XNOR2_X1 U6934 ( .A(n5829), .B(n5828), .ZN(n7066) );
  NOR2_X1 U6935 ( .A1(n5830), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5846) );
  OR2_X1 U6936 ( .A1(n5846), .A2(n10233), .ZN(n5831) );
  XNOR2_X1 U6937 ( .A(n5831), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7123) );
  AOI22_X1 U6938 ( .A1(n8274), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6015), .B2(
        n7123), .ZN(n5832) );
  NAND2_X1 U6939 ( .A1(n6022), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5841) );
  INV_X1 U6940 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5833) );
  OR2_X1 U6941 ( .A1(n6025), .A2(n5833), .ZN(n5840) );
  NAND2_X1 U6942 ( .A1(n5834), .A2(n7687), .ZN(n5835) );
  NAND2_X1 U6943 ( .A1(n5852), .A2(n5835), .ZN(n7689) );
  OR2_X1 U6944 ( .A1(n5758), .A2(n7689), .ZN(n5839) );
  INV_X1 U6945 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5837) );
  OR2_X1 U6946 ( .A1(n5836), .A2(n5837), .ZN(n5838) );
  XNOR2_X1 U6947 ( .A(n7691), .B(n9795), .ZN(n8331) );
  INV_X1 U6948 ( .A(n8331), .ZN(n7599) );
  NAND2_X1 U6949 ( .A1(n7595), .A2(n7599), .ZN(n7594) );
  OR2_X1 U6950 ( .A1(n7691), .A2(n9795), .ZN(n5842) );
  NAND2_X1 U6951 ( .A1(n7594), .A2(n5842), .ZN(n7558) );
  XNOR2_X1 U6952 ( .A(n5844), .B(n5843), .ZN(n7073) );
  NAND2_X1 U6953 ( .A1(n7073), .A2(n8273), .ZN(n5848) );
  INV_X1 U6954 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6955 ( .A1(n5846), .A2(n5845), .ZN(n5902) );
  NAND2_X1 U6956 ( .A1(n5902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U6957 ( .A(n5864), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7271) );
  AOI22_X1 U6958 ( .A1(n8274), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6015), .B2(
        n7271), .ZN(n5847) );
  NAND2_X1 U6959 ( .A1(n5757), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5857) );
  INV_X1 U6960 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5849) );
  OR2_X1 U6961 ( .A1(n7060), .A2(n5849), .ZN(n5856) );
  INV_X1 U6962 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7560) );
  OR2_X1 U6963 ( .A1(n6025), .A2(n7560), .ZN(n5855) );
  INV_X1 U6964 ( .A(n5869), .ZN(n5870) );
  NAND2_X1 U6965 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U6966 ( .A1(n5870), .A2(n5853), .ZN(n7792) );
  OR2_X1 U6967 ( .A1(n5758), .A2(n7792), .ZN(n5854) );
  OR2_X1 U6968 ( .A1(n7615), .A2(n7601), .ZN(n8290) );
  NAND2_X1 U6969 ( .A1(n7615), .A2(n7601), .ZN(n8292) );
  NAND2_X1 U6970 ( .A1(n8290), .A2(n8292), .ZN(n8329) );
  NAND2_X1 U6971 ( .A1(n7558), .A2(n8329), .ZN(n7557) );
  INV_X1 U6972 ( .A(n7601), .ZN(n9794) );
  OR2_X1 U6973 ( .A1(n7615), .A2(n9794), .ZN(n5858) );
  NAND2_X1 U6974 ( .A1(n7557), .A2(n5858), .ZN(n7649) );
  INV_X1 U6975 ( .A(n5859), .ZN(n5861) );
  NAND2_X1 U6976 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U6977 ( .A1(n5863), .A2(n5862), .ZN(n7072) );
  OR2_X1 U6978 ( .A1(n7072), .A2(n5997), .ZN(n5867) );
  INV_X1 U6979 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6980 ( .A1(n5864), .A2(n5899), .ZN(n5865) );
  NAND2_X1 U6981 ( .A1(n5865), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U6982 ( .A(n5879), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U6983 ( .A1(n8274), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10502), 
        .B2(n6015), .ZN(n5866) );
  NAND2_X1 U6984 ( .A1(n6022), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5875) );
  INV_X1 U6985 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5868) );
  OR2_X1 U6986 ( .A1(n5836), .A2(n5868), .ZN(n5874) );
  INV_X1 U6987 ( .A(n5884), .ZN(n5886) );
  INV_X1 U6988 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U6989 ( .A1(n5870), .A2(n8000), .ZN(n5871) );
  NAND2_X1 U6990 ( .A1(n5886), .A2(n5871), .ZN(n8001) );
  OR2_X1 U6991 ( .A1(n5758), .A2(n8001), .ZN(n5873) );
  INV_X1 U6992 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7656) );
  OR2_X1 U6993 ( .A1(n6025), .A2(n7656), .ZN(n5872) );
  NAND4_X1 U6994 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n9793)
         );
  AND2_X1 U6995 ( .A1(n8005), .A2(n9793), .ZN(n8293) );
  INV_X1 U6996 ( .A(n8005), .ZN(n7658) );
  INV_X1 U6997 ( .A(n9793), .ZN(n8047) );
  NAND2_X1 U6998 ( .A1(n7658), .A2(n8047), .ZN(n8333) );
  INV_X1 U6999 ( .A(n7653), .ZN(n8245) );
  NAND2_X1 U7000 ( .A1(n7649), .A2(n8245), .ZN(n7648) );
  NAND2_X1 U7001 ( .A1(n8005), .A2(n8047), .ZN(n5876) );
  NAND2_X1 U7002 ( .A1(n7648), .A2(n5876), .ZN(n7663) );
  XNOR2_X1 U7003 ( .A(n5878), .B(n5877), .ZN(n7134) );
  NAND2_X1 U7004 ( .A1(n7134), .A2(n8273), .ZN(n5883) );
  NAND2_X1 U7005 ( .A1(n5879), .A2(n5900), .ZN(n5880) );
  NAND2_X1 U7006 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7007 ( .A(n5881), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7273) );
  AOI22_X1 U7008 ( .A1(n7273), .A2(n6015), .B1(P2_DATAO_REG_11__SCAN_IN), .B2(
        n8274), .ZN(n5882) );
  NAND2_X1 U7009 ( .A1(n5757), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5891) );
  INV_X1 U7010 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7272) );
  OR2_X1 U7011 ( .A1(n7060), .A2(n7272), .ZN(n5890) );
  INV_X1 U7012 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7013 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7014 ( .A1(n5907), .A2(n5887), .ZN(n8048) );
  OR2_X1 U7015 ( .A1(n5758), .A2(n8048), .ZN(n5889) );
  INV_X1 U7016 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7670) );
  OR2_X1 U7017 ( .A1(n6025), .A2(n7670), .ZN(n5888) );
  NAND2_X1 U7018 ( .A1(n7672), .A2(n9792), .ZN(n5892) );
  OR2_X1 U7019 ( .A1(n7672), .A2(n9792), .ZN(n5893) );
  NAND2_X1 U7020 ( .A1(n5895), .A2(n5894), .ZN(n5897) );
  NAND2_X1 U7021 ( .A1(n5897), .A2(n5896), .ZN(n7160) );
  INV_X1 U7022 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5898) );
  NAND3_X1 U7023 ( .A1(n5900), .A2(n5899), .A3(n5898), .ZN(n5901) );
  NAND2_X1 U7024 ( .A1(n5919), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U7025 ( .A(n5903), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U7026 ( .A1(n8274), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6015), .B2(
        n9855), .ZN(n5904) );
  NAND2_X1 U7027 ( .A1(n5757), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5913) );
  INV_X1 U7028 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7268) );
  OR2_X1 U7029 ( .A1(n7060), .A2(n7268), .ZN(n5912) );
  NAND2_X1 U7030 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U7031 ( .A1(n5924), .A2(n5908), .ZN(n8122) );
  OR2_X1 U7032 ( .A1(n5758), .A2(n8122), .ZN(n5911) );
  INV_X1 U7033 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5909) );
  OR2_X1 U7034 ( .A1(n6025), .A2(n5909), .ZN(n5910) );
  INV_X1 U7035 ( .A(n9517), .ZN(n8051) );
  NOR2_X1 U7036 ( .A1(n8117), .A2(n8051), .ZN(n5914) );
  OR2_X1 U7037 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  NAND2_X1 U7038 ( .A1(n5918), .A2(n5917), .ZN(n7195) );
  NAND2_X1 U7039 ( .A1(n5936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7040 ( .A(n5920), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U7041 ( .A1(n6015), .A2(n10487), .B1(n8230), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5921) );
  INV_X1 U7042 ( .A(n10180), .ZN(n7958) );
  NAND2_X1 U7043 ( .A1(n6022), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5930) );
  INV_X1 U7044 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9853) );
  OR2_X1 U7045 ( .A1(n6025), .A2(n9853), .ZN(n5929) );
  NAND2_X1 U7046 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  NAND2_X1 U7047 ( .A1(n5939), .A2(n5925), .ZN(n9518) );
  OR2_X1 U7048 ( .A1(n5758), .A2(n9518), .ZN(n5928) );
  INV_X1 U7049 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7050 ( .A1(n5836), .A2(n5926), .ZN(n5927) );
  INV_X1 U7051 ( .A(n9427), .ZN(n9791) );
  NAND2_X1 U7052 ( .A1(n10180), .A2(n9427), .ZN(n8339) );
  OR2_X1 U7053 ( .A1(n10180), .A2(n9791), .ZN(n5931) );
  INV_X1 U7054 ( .A(n8025), .ZN(n5945) );
  NAND2_X1 U7055 ( .A1(n5935), .A2(n5934), .ZN(n7241) );
  OAI21_X1 U7056 ( .B1(n5936), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7057 ( .A(n5952), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U7058 ( .A1(n10439), .A2(n6015), .B1(n8230), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7059 ( .A1(n5757), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5944) );
  INV_X1 U7060 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8184) );
  OR2_X1 U7061 ( .A1(n7060), .A2(n8184), .ZN(n5943) );
  INV_X1 U7062 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8036) );
  OR2_X1 U7063 ( .A1(n6025), .A2(n8036), .ZN(n5942) );
  INV_X1 U7064 ( .A(n5957), .ZN(n5959) );
  NAND2_X1 U7065 ( .A1(n5939), .A2(n9425), .ZN(n5940) );
  NAND2_X1 U7066 ( .A1(n5959), .A2(n5940), .ZN(n9428) );
  OR2_X1 U7067 ( .A1(n5758), .A2(n9428), .ZN(n5941) );
  NAND2_X1 U7068 ( .A1(n9431), .A2(n9771), .ZN(n8287) );
  NAND2_X1 U7069 ( .A1(n8472), .A2(n8287), .ZN(n8349) );
  NAND2_X1 U7070 ( .A1(n5945), .A2(n8349), .ZN(n8024) );
  INV_X1 U7071 ( .A(n9771), .ZN(n9790) );
  NAND2_X1 U7072 ( .A1(n9431), .A2(n9790), .ZN(n5946) );
  NAND2_X1 U7073 ( .A1(n5950), .A2(n5949), .ZN(n7289) );
  INV_X1 U7074 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7075 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7076 ( .A1(n5953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7077 ( .A(n5954), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U7078 ( .A1(n10464), .A2(n6015), .B1(n8230), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7079 ( .A1(n5957), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5973) );
  INV_X1 U7080 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7081 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7082 ( .A1(n5973), .A2(n5960), .ZN(n9773) );
  OR2_X1 U7083 ( .A1(n9773), .A2(n5758), .ZN(n5964) );
  NAND2_X1 U7084 ( .A1(n5757), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7085 ( .A1(n4927), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5962) );
  INV_X1 U7086 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10457) );
  OR2_X1 U7087 ( .A1(n7060), .A2(n10457), .ZN(n5961) );
  INV_X1 U7088 ( .A(n9426), .ZN(n9789) );
  AND2_X1 U7089 ( .A1(n8017), .A2(n9789), .ZN(n5965) );
  XNOR2_X1 U7090 ( .A(n5967), .B(n5966), .ZN(n7311) );
  NAND2_X1 U7091 ( .A1(n7311), .A2(n8273), .ZN(n5971) );
  NAND2_X1 U7092 ( .A1(n5968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5969) );
  XNOR2_X1 U7093 ( .A(n5969), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U7094 ( .A1(n8274), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6015), .B2(
        n9874), .ZN(n5970) );
  NAND2_X1 U7095 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  AND2_X1 U7096 ( .A1(n5986), .A2(n5974), .ZN(n9481) );
  NAND2_X1 U7097 ( .A1(n9481), .A2(n5850), .ZN(n5978) );
  AOI22_X1 U7098 ( .A1(n6022), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n5757), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5977) );
  INV_X1 U7099 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7100 ( .A1(n6025), .A2(n5975), .ZN(n5976) );
  OR2_X1 U7101 ( .A1(n10171), .A2(n10163), .ZN(n8352) );
  NAND2_X1 U7102 ( .A1(n10171), .A2(n10163), .ZN(n8481) );
  INV_X1 U7103 ( .A(n10163), .ZN(n9788) );
  NAND2_X1 U7104 ( .A1(n10171), .A2(n9788), .ZN(n5979) );
  NAND2_X1 U7105 ( .A1(n8140), .A2(n5979), .ZN(n8210) );
  XNOR2_X1 U7106 ( .A(n5980), .B(n5981), .ZN(n7567) );
  NAND2_X1 U7107 ( .A1(n7567), .A2(n8273), .ZN(n5984) );
  OR2_X1 U7108 ( .A1(n4994), .A2(n10233), .ZN(n5982) );
  XNOR2_X1 U7109 ( .A(n5982), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9890) );
  AOI22_X1 U7110 ( .A1(n8274), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6015), .B2(
        n9890), .ZN(n5983) );
  INV_X1 U7111 ( .A(n6001), .ZN(n6003) );
  NAND2_X1 U7112 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7113 ( .A1(n6003), .A2(n5987), .ZN(n9490) );
  OR2_X1 U7114 ( .A1(n9490), .A2(n5758), .ZN(n5990) );
  AOI22_X1 U7115 ( .A1(n6022), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5757), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5989) );
  INV_X1 U7116 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8213) );
  OR2_X1 U7117 ( .A1(n6025), .A2(n8213), .ZN(n5988) );
  NAND2_X1 U7118 ( .A1(n10166), .A2(n10156), .ZN(n8233) );
  NAND2_X1 U7119 ( .A1(n8210), .A2(n8209), .ZN(n8208) );
  INV_X1 U7120 ( .A(n10156), .ZN(n9787) );
  NAND2_X1 U7121 ( .A1(n10166), .A2(n9787), .ZN(n5991) );
  INV_X1 U7122 ( .A(n5992), .ZN(n5994) );
  NAND2_X1 U7123 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  NAND2_X1 U7124 ( .A1(n5996), .A2(n5995), .ZN(n7539) );
  XNOR2_X1 U7125 ( .A(n5998), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U7126 ( .A1(n8274), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6015), .B2(
        n10477), .ZN(n5999) );
  INV_X1 U7127 ( .A(n6018), .ZN(n6020) );
  INV_X1 U7128 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7129 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  AND2_X1 U7130 ( .A1(n6020), .A2(n6004), .ZN(n10082) );
  NAND2_X1 U7131 ( .A1(n10082), .A2(n5850), .ZN(n6010) );
  INV_X1 U7132 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7133 ( .A1(n5757), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7134 ( .A1(n4927), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6005) );
  OAI211_X1 U7135 ( .C1(n7060), .C2(n6007), .A(n6006), .B(n6005), .ZN(n6008)
         );
  INV_X1 U7136 ( .A(n6008), .ZN(n6009) );
  OR2_X1 U7137 ( .A1(n10159), .A2(n9786), .ZN(n6011) );
  NAND2_X1 U7138 ( .A1(n10159), .A2(n9786), .ZN(n6012) );
  XNOR2_X1 U7139 ( .A(n6014), .B(n6013), .ZN(n7620) );
  NAND2_X1 U7140 ( .A1(n7620), .A2(n8273), .ZN(n6017) );
  AOI22_X1 U7141 ( .A1(n8230), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9886), .B2(
        n6015), .ZN(n6016) );
  INV_X1 U7142 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7143 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7144 ( .A1(n6035), .A2(n6021), .ZN(n10067) );
  OR2_X1 U7145 ( .A1(n10067), .A2(n5758), .ZN(n6028) );
  INV_X1 U7146 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U7147 ( .A1(n6022), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7148 ( .A1(n5757), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6023) );
  OAI211_X1 U7149 ( .C1(n6025), .C2(n10068), .A(n6024), .B(n6023), .ZN(n6026)
         );
  INV_X1 U7150 ( .A(n6026), .ZN(n6027) );
  NAND2_X1 U7151 ( .A1(n10153), .A2(n10088), .ZN(n8255) );
  INV_X1 U7152 ( .A(SI_20_), .ZN(n6029) );
  XNOR2_X1 U7153 ( .A(n6030), .B(n6029), .ZN(n6031) );
  XNOR2_X1 U7154 ( .A(n6032), .B(n6031), .ZN(n7695) );
  NAND2_X1 U7155 ( .A1(n7695), .A2(n8273), .ZN(n6034) );
  NAND2_X1 U7156 ( .A1(n8274), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6033) );
  INV_X1 U7157 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U7158 ( .A1(n6035), .A2(n9507), .ZN(n6036) );
  AND2_X1 U7159 ( .A1(n6049), .A2(n6036), .ZN(n10057) );
  NAND2_X1 U7160 ( .A1(n10057), .A2(n5850), .ZN(n6042) );
  INV_X1 U7161 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7162 ( .A1(n5757), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7163 ( .A1(n4927), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6037) );
  OAI211_X1 U7164 ( .C1(n7060), .C2(n6039), .A(n6038), .B(n6037), .ZN(n6040)
         );
  INV_X1 U7165 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7166 ( .A1(n10148), .A2(n10139), .ZN(n8365) );
  NAND2_X1 U7167 ( .A1(n10042), .A2(n8365), .ZN(n10051) );
  NAND2_X1 U7168 ( .A1(n10050), .A2(n10051), .ZN(n6044) );
  INV_X1 U7169 ( .A(n10139), .ZN(n9785) );
  OR2_X1 U7170 ( .A1(n10148), .A2(n9785), .ZN(n6043) );
  NAND2_X1 U7171 ( .A1(n6044), .A2(n6043), .ZN(n10032) );
  XNOR2_X1 U7172 ( .A(n6046), .B(n6045), .ZN(n7857) );
  NAND2_X1 U7173 ( .A1(n7857), .A2(n8273), .ZN(n6048) );
  NAND2_X1 U7174 ( .A1(n8274), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6047) );
  INV_X1 U7175 ( .A(n6062), .ZN(n6064) );
  NAND2_X1 U7176 ( .A1(n6049), .A2(n9459), .ZN(n6050) );
  NAND2_X1 U7177 ( .A1(n6064), .A2(n6050), .ZN(n10035) );
  OR2_X1 U7178 ( .A1(n10035), .A2(n5758), .ZN(n6056) );
  INV_X1 U7179 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7180 ( .A1(n5757), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7181 ( .A1(n4927), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7182 ( .C1(n7060), .C2(n6053), .A(n6052), .B(n6051), .ZN(n6054)
         );
  INV_X1 U7183 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7184 ( .A1(n10142), .A2(n10132), .ZN(n8368) );
  INV_X1 U7185 ( .A(n10132), .ZN(n9784) );
  OR2_X1 U7186 ( .A1(n10142), .A2(n9784), .ZN(n6057) );
  XNOR2_X1 U7187 ( .A(n6059), .B(n6058), .ZN(n7896) );
  NAND2_X1 U7188 ( .A1(n7896), .A2(n8273), .ZN(n6061) );
  NAND2_X1 U7189 ( .A1(n8274), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7190 ( .A1(n6062), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6079) );
  INV_X1 U7191 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7192 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  NAND2_X1 U7193 ( .A1(n6079), .A2(n6065), .ZN(n10021) );
  OR2_X1 U7194 ( .A1(n10021), .A2(n5758), .ZN(n6071) );
  INV_X1 U7195 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7196 ( .A1(n5757), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7197 ( .A1(n4927), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6066) );
  OAI211_X1 U7198 ( .C1(n7060), .C2(n6068), .A(n6067), .B(n6066), .ZN(n6069)
         );
  INV_X1 U7199 ( .A(n6069), .ZN(n6070) );
  OR2_X1 U7200 ( .A1(n10135), .A2(n10126), .ZN(n8284) );
  NAND2_X1 U7201 ( .A1(n10135), .A2(n10126), .ZN(n8373) );
  INV_X1 U7202 ( .A(n10025), .ZN(n6072) );
  INV_X1 U7203 ( .A(n10126), .ZN(n10045) );
  NAND2_X1 U7204 ( .A1(n6076), .A2(n6075), .ZN(n7964) );
  NAND2_X1 U7205 ( .A1(n7964), .A2(n8273), .ZN(n6078) );
  NAND2_X1 U7206 ( .A1(n8230), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6077) );
  INV_X1 U7207 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U7208 ( .A1(n6079), .A2(n9438), .ZN(n6080) );
  NAND2_X1 U7209 ( .A1(n6095), .A2(n6080), .ZN(n10007) );
  OR2_X1 U7210 ( .A1(n10007), .A2(n5758), .ZN(n6085) );
  INV_X1 U7211 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U7212 ( .A1(n5757), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7213 ( .A1(n4927), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6081) );
  OAI211_X1 U7214 ( .C1(n7060), .C2(n10129), .A(n6082), .B(n6081), .ZN(n6083)
         );
  INV_X1 U7215 ( .A(n6083), .ZN(n6084) );
  NAND2_X1 U7216 ( .A1(n10013), .A2(n10027), .ZN(n6086) );
  OR2_X1 U7217 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  NAND2_X1 U7218 ( .A1(n6091), .A2(n6090), .ZN(n8009) );
  NAND2_X1 U7219 ( .A1(n8009), .A2(n8273), .ZN(n6093) );
  NAND2_X1 U7220 ( .A1(n8274), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6092) );
  NAND2_X2 U7221 ( .A1(n6093), .A2(n6092), .ZN(n9995) );
  INV_X1 U7222 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7223 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7224 ( .A1(n9996), .A2(n5850), .ZN(n6101) );
  INV_X1 U7225 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U7226 ( .A1(n5757), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7227 ( .A1(n4927), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6097) );
  OAI211_X1 U7228 ( .C1(n7060), .C2(n10122), .A(n6098), .B(n6097), .ZN(n6099)
         );
  INV_X1 U7229 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U7230 ( .A1(n6105), .A2(n6104), .ZN(n8128) );
  NAND2_X1 U7231 ( .A1(n8128), .A2(n8273), .ZN(n6107) );
  NAND2_X1 U7232 ( .A1(n8230), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6106) );
  INV_X1 U7233 ( .A(n6110), .ZN(n6108) );
  NAND2_X1 U7234 ( .A1(n6108), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6125) );
  INV_X1 U7235 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7236 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  NAND2_X1 U7237 ( .A1(n6125), .A2(n6111), .ZN(n9467) );
  OR2_X1 U7238 ( .A1(n9467), .A2(n5758), .ZN(n6117) );
  INV_X1 U7239 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7240 ( .A1(n5757), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7241 ( .A1(n4927), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7242 ( .C1(n7060), .C2(n6114), .A(n6113), .B(n6112), .ZN(n6115)
         );
  INV_X1 U7243 ( .A(n6115), .ZN(n6116) );
  NOR2_X1 U7244 ( .A1(n9471), .A2(n9501), .ZN(n6118) );
  XNOR2_X1 U7245 ( .A(n6120), .B(n6119), .ZN(n8201) );
  NAND2_X1 U7246 ( .A1(n8201), .A2(n8273), .ZN(n6122) );
  NAND2_X1 U7247 ( .A1(n8274), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6121) );
  INV_X1 U7248 ( .A(n6125), .ZN(n6123) );
  INV_X1 U7249 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7250 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  NAND2_X1 U7251 ( .A1(n6145), .A2(n6126), .ZN(n9758) );
  OR2_X1 U7252 ( .A1(n9758), .A2(n5758), .ZN(n6131) );
  INV_X1 U7253 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U7254 ( .A1(n4927), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7255 ( .A1(n5757), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6127) );
  OAI211_X1 U7256 ( .C1(n7060), .C2(n10114), .A(n6128), .B(n6127), .ZN(n6129)
         );
  INV_X1 U7257 ( .A(n6129), .ZN(n6130) );
  NOR2_X1 U7258 ( .A1(n9962), .A2(n10103), .ZN(n8384) );
  INV_X1 U7259 ( .A(n8384), .ZN(n8425) );
  AND2_X1 U7260 ( .A1(n9962), .A2(n10103), .ZN(n8382) );
  INV_X1 U7261 ( .A(n8382), .ZN(n8422) );
  NAND2_X1 U7262 ( .A1(n8425), .A2(n8422), .ZN(n8283) );
  INV_X1 U7263 ( .A(n10103), .ZN(n9783) );
  NAND2_X1 U7264 ( .A1(n9962), .A2(n9783), .ZN(n6132) );
  NAND2_X1 U7265 ( .A1(n9414), .A2(n8273), .ZN(n6136) );
  NAND2_X1 U7266 ( .A1(n8274), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7267 ( .A(n6145), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U7268 ( .A1(n9943), .A2(n5850), .ZN(n6141) );
  INV_X1 U7269 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U7270 ( .A1(n5757), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7271 ( .A1(n4927), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6137) );
  OAI211_X1 U7272 ( .C1(n7060), .C2(n10107), .A(n6138), .B(n6137), .ZN(n6139)
         );
  INV_X1 U7273 ( .A(n6139), .ZN(n6140) );
  NAND2_X1 U7274 ( .A1(n9947), .A2(n9926), .ZN(n8419) );
  NAND2_X1 U7275 ( .A1(n8426), .A2(n8419), .ZN(n9936) );
  OR2_X1 U7276 ( .A1(n9947), .A2(n9954), .ZN(n6142) );
  INV_X1 U7277 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6965) );
  INV_X1 U7278 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6143) );
  OAI21_X1 U7279 ( .B1(n6145), .B2(n6965), .A(n6143), .ZN(n6146) );
  NAND2_X1 U7280 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6144) );
  INV_X1 U7281 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7282 ( .A1(n4927), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7283 ( .A1(n5757), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U7284 ( .C1(n7060), .C2(n6149), .A(n6148), .B(n6147), .ZN(n6150)
         );
  INV_X1 U7285 ( .A(n8387), .ZN(n6706) );
  AND2_X1 U7286 ( .A1(n6151), .A2(n6706), .ZN(n6152) );
  OR2_X1 U7287 ( .A1(n8436), .A2(n8505), .ZN(n8507) );
  OAI21_X1 U7288 ( .B1(n8505), .B2(n8234), .A(n6154), .ZN(n6155) );
  NAND2_X1 U7289 ( .A1(n8507), .A2(n6155), .ZN(n10655) );
  NAND2_X1 U7290 ( .A1(n8406), .A2(n6951), .ZN(n10665) );
  OR2_X1 U7291 ( .A1(n9995), .A2(n9974), .ZN(n8412) );
  NAND2_X1 U7292 ( .A1(n9995), .A2(n9974), .ZN(n8409) );
  NAND2_X1 U7293 ( .A1(n8368), .A2(n8365), .ZN(n6156) );
  AND2_X1 U7294 ( .A1(n6156), .A2(n8367), .ZN(n8411) );
  OR2_X1 U7295 ( .A1(n10153), .A2(n10054), .ZN(n10039) );
  AND2_X1 U7296 ( .A1(n10042), .A2(n10039), .ZN(n8364) );
  NAND2_X1 U7297 ( .A1(n8367), .A2(n8364), .ZN(n8485) );
  NOR2_X1 U7298 ( .A1(n7691), .A2(n7610), .ZN(n8326) );
  INV_X1 U7299 ( .A(n8326), .ZN(n7554) );
  NAND2_X1 U7300 ( .A1(n8240), .A2(n8319), .ZN(n6158) );
  AND2_X1 U7301 ( .A1(n8320), .A2(n8316), .ZN(n8314) );
  NOR2_X1 U7302 ( .A1(n6158), .A2(n8314), .ZN(n6157) );
  INV_X1 U7303 ( .A(n8318), .ZN(n7400) );
  OR2_X1 U7304 ( .A1(n6158), .A2(n7400), .ZN(n8461) );
  NOR2_X1 U7305 ( .A1(n6739), .A2(n10606), .ZN(n10186) );
  NAND2_X1 U7306 ( .A1(n10187), .A2(n10186), .ZN(n6160) );
  INV_X1 U7307 ( .A(n6724), .ZN(n10634) );
  NAND2_X1 U7308 ( .A1(n10634), .A2(n6731), .ZN(n6159) );
  NAND2_X1 U7309 ( .A1(n6160), .A2(n6159), .ZN(n10631) );
  NAND2_X1 U7310 ( .A1(n10631), .A2(n8451), .ZN(n8296) );
  NAND2_X1 U7311 ( .A1(n10651), .A2(n10652), .ZN(n10650) );
  NAND2_X1 U7312 ( .A1(n10650), .A2(n8452), .ZN(n10697) );
  NAND2_X1 U7313 ( .A1(n10689), .A2(n9797), .ZN(n8297) );
  INV_X1 U7314 ( .A(n10689), .ZN(n10691) );
  AND2_X1 U7315 ( .A1(n10691), .A2(n10654), .ZN(n8300) );
  INV_X1 U7316 ( .A(n8300), .ZN(n8457) );
  NAND2_X1 U7317 ( .A1(n10697), .A2(n10696), .ZN(n6162) );
  NAND2_X1 U7318 ( .A1(n6162), .A2(n8457), .ZN(n7317) );
  NAND2_X1 U7319 ( .A1(n7317), .A2(n8237), .ZN(n6163) );
  NAND2_X1 U7320 ( .A1(n7652), .A2(n7653), .ZN(n7651) );
  OR2_X1 U7321 ( .A1(n7672), .A2(n6822), .ZN(n8341) );
  NAND2_X1 U7322 ( .A1(n7672), .A2(n6822), .ZN(n8334) );
  NAND2_X1 U7323 ( .A1(n8341), .A2(n8334), .ZN(n8247) );
  OR2_X1 U7324 ( .A1(n8117), .A2(n9517), .ZN(n8342) );
  NAND2_X1 U7325 ( .A1(n8117), .A2(n9517), .ZN(n8338) );
  NAND2_X1 U7326 ( .A1(n7799), .A2(n8338), .ZN(n7959) );
  OR2_X1 U7327 ( .A1(n8017), .A2(n9426), .ZN(n8476) );
  NAND2_X1 U7328 ( .A1(n8017), .A2(n9426), .ZN(n8288) );
  NAND2_X1 U7329 ( .A1(n8476), .A2(n8288), .ZN(n8253) );
  XNOR2_X1 U7330 ( .A(n10159), .B(n9786), .ZN(n10086) );
  OR2_X1 U7331 ( .A1(n10159), .A2(n10074), .ZN(n8482) );
  NAND2_X1 U7332 ( .A1(n10153), .A2(n10054), .ZN(n8487) );
  NAND2_X1 U7333 ( .A1(n10026), .A2(n10025), .ZN(n6165) );
  OR2_X1 U7334 ( .A1(n10013), .A2(n9991), .ZN(n8374) );
  NAND2_X1 U7335 ( .A1(n10013), .A2(n9991), .ZN(n9986) );
  NAND2_X1 U7336 ( .A1(n8374), .A2(n9986), .ZN(n10015) );
  INV_X1 U7337 ( .A(n10015), .ZN(n10004) );
  NAND2_X1 U7338 ( .A1(n10003), .A2(n10004), .ZN(n10002) );
  NAND2_X1 U7339 ( .A1(n9471), .A2(n10111), .ZN(n8421) );
  NAND2_X1 U7340 ( .A1(n8415), .A2(n8421), .ZN(n9972) );
  NAND2_X1 U7341 ( .A1(n9964), .A2(n9953), .ZN(n9952) );
  NAND2_X1 U7342 ( .A1(n8508), .A2(n9886), .ZN(n8405) );
  NAND2_X1 U7343 ( .A1(n6726), .A2(n8441), .ZN(n6166) );
  OR2_X1 U7344 ( .A1(n6167), .A2(n10698), .ZN(n6176) );
  INV_X1 U7345 ( .A(n9914), .ZN(n6172) );
  INV_X1 U7346 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7347 ( .A1(n4927), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7348 ( .A1(n5757), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6168) );
  OAI211_X1 U7349 ( .C1(n7060), .C2(n6170), .A(n6169), .B(n6168), .ZN(n6171)
         );
  AOI21_X1 U7350 ( .B1(n6172), .B2(n5850), .A(n6171), .ZN(n7243) );
  OAI21_X1 U7351 ( .B1(n6173), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7352 ( .A1(n7243), .A2(n10703), .ZN(n6175) );
  INV_X1 U7353 ( .A(n10148), .ZN(n10060) );
  INV_X1 U7354 ( .A(n8017), .ZN(n9780) );
  INV_X1 U7355 ( .A(n7445), .ZN(n7485) );
  NAND2_X1 U7356 ( .A1(n10616), .A2(n10606), .ZN(n10626) );
  NAND2_X1 U7357 ( .A1(n9780), .A2(n8016), .ZN(n8136) );
  AOI21_X1 U7358 ( .B1(n9928), .B2(n9941), .A(n10660), .ZN(n6178) );
  NAND2_X1 U7359 ( .A1(n6178), .A2(n6715), .ZN(n9930) );
  OR2_X1 U7360 ( .A1(n9926), .A2(n10701), .ZN(n6179) );
  AND2_X1 U7361 ( .A1(n9930), .A2(n6179), .ZN(n6180) );
  INV_X1 U7362 ( .A(n9928), .ZN(n6183) );
  NAND3_X1 U7363 ( .A1(n6271), .A2(n6286), .A3(n6185), .ZN(n6186) );
  NOR2_X1 U7364 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6189) );
  NAND4_X1 U7365 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6427), .ZN(n6193)
         );
  NAND4_X1 U7366 ( .A1(n6191), .A2(n6388), .A3(n6190), .A4(n6415), .ZN(n6192)
         );
  INV_X1 U7367 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6197) );
  XNOR2_X2 U7368 ( .A(n6201), .B(n5047), .ZN(n6203) );
  AND2_X4 U7369 ( .A1(n6204), .A2(n6203), .ZN(n6248) );
  INV_X2 U7370 ( .A(n6204), .ZN(n6207) );
  INV_X1 U7371 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6205) );
  INV_X1 U7372 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7490) );
  INV_X1 U7373 ( .A(n6210), .ZN(n6211) );
  NAND2_X1 U7374 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6213) );
  OAI22_X1 U7375 ( .A1(n6244), .A2(n6214), .B1(n7192), .B2(n7009), .ZN(n6215)
         );
  INV_X1 U7376 ( .A(n6215), .ZN(n6217) );
  INV_X1 U7377 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10512) );
  OR2_X1 U7378 ( .A1(n6249), .A2(n10512), .ZN(n6222) );
  INV_X1 U7379 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6218) );
  OR2_X1 U7380 ( .A1(n6261), .A2(n6218), .ZN(n6221) );
  NAND2_X1 U7381 ( .A1(n6202), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7382 ( .A1(n6248), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7383 ( .A1(n5701), .A2(SI_0_), .ZN(n6223) );
  XNOR2_X1 U7384 ( .A(n6223), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9418) );
  MUX2_X1 U7385 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9418), .S(n7009), .Z(n7509) );
  INV_X1 U7386 ( .A(n7509), .ZN(n7284) );
  OR2_X1 U7387 ( .A1(n8515), .A2(n7284), .ZN(n7359) );
  NAND2_X1 U7388 ( .A1(n7226), .A2(n5314), .ZN(n6224) );
  NAND2_X1 U7389 ( .A1(n6225), .A2(n6224), .ZN(n7463) );
  INV_X1 U7390 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7260) );
  OR2_X1 U7391 ( .A1(n6261), .A2(n7473), .ZN(n6229) );
  NAND2_X1 U7392 ( .A1(n6248), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6228) );
  INV_X1 U7393 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7394 ( .A1(n6244), .A2(n7040), .ZN(n6234) );
  INV_X1 U7395 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7039) );
  OR2_X1 U7396 ( .A1(n6274), .A2(n7039), .ZN(n6233) );
  XNOR2_X2 U7397 ( .A(n6617), .B(n7467), .ZN(n8772) );
  INV_X1 U7398 ( .A(n8772), .ZN(n7458) );
  INV_X1 U7399 ( .A(n6617), .ZN(n7580) );
  INV_X1 U7400 ( .A(n7467), .ZN(n8768) );
  NAND2_X1 U7401 ( .A1(n7580), .A2(n8768), .ZN(n6235) );
  NAND2_X1 U7402 ( .A1(n6587), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6241) );
  INV_X1 U7403 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6236) );
  OR2_X1 U7404 ( .A1(n7572), .A2(n6236), .ZN(n6240) );
  OR2_X1 U7405 ( .A1(n6249), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6239) );
  INV_X1 U7406 ( .A(n6248), .ZN(n6327) );
  INV_X1 U7407 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7408 ( .A1(n6242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6243) );
  XNOR2_X1 U7409 ( .A(n6243), .B(n6184), .ZN(n7352) );
  INV_X1 U7410 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7042) );
  OR2_X1 U7411 ( .A1(n6274), .A2(n7042), .ZN(n6246) );
  OAI211_X1 U7412 ( .C1(n7009), .C2(n7352), .A(n6246), .B(n6245), .ZN(n7585)
         );
  NOR2_X1 U7413 ( .A1(n8929), .A2(n7585), .ZN(n6247) );
  INV_X1 U7414 ( .A(n7585), .ZN(n7587) );
  NAND2_X1 U7415 ( .A1(n6248), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6254) );
  INV_X1 U7416 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7335) );
  OR2_X1 U7417 ( .A1(n6261), .A2(n7335), .ZN(n6253) );
  INV_X2 U7418 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9620) );
  INV_X2 U7419 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9550) );
  NAND2_X1 U7420 ( .A1(n9620), .A2(n9550), .ZN(n6264) );
  NAND2_X1 U7421 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6250) );
  AND2_X1 U7422 ( .A1(n6264), .A2(n6250), .ZN(n7516) );
  OR2_X1 U7423 ( .A1(n6249), .A2(n7516), .ZN(n6252) );
  INV_X1 U7424 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7340) );
  OR2_X1 U7425 ( .A1(n7572), .A2(n7340), .ZN(n6251) );
  NAND2_X1 U7426 ( .A1(n6255), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6272) );
  XNOR2_X1 U7427 ( .A(n6272), .B(n6271), .ZN(n7699) );
  OR2_X1 U7428 ( .A1(n6274), .A2(n5596), .ZN(n6257) );
  OR2_X1 U7429 ( .A1(n6401), .A2(n7044), .ZN(n6256) );
  OAI211_X1 U7430 ( .C1(n7009), .C2(n7699), .A(n6257), .B(n6256), .ZN(n7428)
         );
  INV_X1 U7431 ( .A(n7428), .ZN(n10680) );
  NAND2_X1 U7432 ( .A1(n7579), .A2(n10680), .ZN(n6258) );
  NAND2_X1 U7433 ( .A1(n6259), .A2(n6258), .ZN(n7781) );
  NAND2_X1 U7434 ( .A1(n6248), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6270) );
  INV_X1 U7435 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6260) );
  OR2_X1 U7436 ( .A1(n6261), .A2(n6260), .ZN(n6269) );
  INV_X1 U7437 ( .A(n6264), .ZN(n6263) );
  NAND2_X1 U7438 ( .A1(n6263), .A2(n6262), .ZN(n6279) );
  NAND2_X1 U7439 ( .A1(n6264), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6265) );
  AND2_X1 U7440 ( .A1(n6279), .A2(n6265), .ZN(n7780) );
  OR2_X1 U7441 ( .A1(n6249), .A2(n7780), .ZN(n6268) );
  INV_X1 U7442 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7443 ( .A1(n7572), .A2(n6266), .ZN(n6267) );
  NAND2_X1 U7444 ( .A1(n6272), .A2(n6271), .ZN(n6273) );
  NAND2_X1 U7445 ( .A1(n6273), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  XNOR2_X1 U7446 ( .A(n6287), .B(n6286), .ZN(n10529) );
  OR2_X1 U7447 ( .A1(n6274), .A2(n5302), .ZN(n6276) );
  OR2_X1 U7448 ( .A1(n6401), .A2(n7046), .ZN(n6275) );
  OAI211_X1 U7449 ( .C1(n7009), .C2(n10529), .A(n6276), .B(n6275), .ZN(n7521)
         );
  NOR2_X1 U7450 ( .A1(n8927), .A2(n7521), .ZN(n6278) );
  NAND2_X1 U7451 ( .A1(n8927), .A2(n7521), .ZN(n6277) );
  NAND2_X1 U7452 ( .A1(n6248), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6285) );
  INV_X1 U7453 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7772) );
  OR2_X1 U7454 ( .A1(n6261), .A2(n7772), .ZN(n6284) );
  NAND2_X1 U7455 ( .A1(n6279), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6280) );
  AND2_X1 U7456 ( .A1(n6296), .A2(n6280), .ZN(n7773) );
  OR2_X1 U7457 ( .A1(n6249), .A2(n7773), .ZN(n6283) );
  INV_X1 U7458 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6281) );
  OR2_X1 U7459 ( .A1(n7572), .A2(n6281), .ZN(n6282) );
  NAND4_X1 U7460 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n8926)
         );
  NAND2_X1 U7461 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  NAND2_X1 U7462 ( .A1(n6288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6289) );
  XNOR2_X1 U7463 ( .A(n6289), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10549) );
  OR2_X1 U7464 ( .A1(n7048), .A2(n6401), .ZN(n6291) );
  NAND2_X1 U7465 ( .A1(n6562), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6290) );
  OAI211_X1 U7466 ( .C1(n7009), .C2(n7707), .A(n6291), .B(n6290), .ZN(n7775)
         );
  AND2_X1 U7467 ( .A1(n8926), .A2(n7775), .ZN(n6292) );
  NAND2_X1 U7468 ( .A1(n6248), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6301) );
  INV_X1 U7469 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6293) );
  OR2_X1 U7470 ( .A1(n6261), .A2(n6293), .ZN(n6300) );
  INV_X1 U7471 ( .A(n6296), .ZN(n6295) );
  NAND2_X1 U7472 ( .A1(n6295), .A2(n6294), .ZN(n6316) );
  NAND2_X1 U7473 ( .A1(n6296), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6297) );
  AND2_X1 U7474 ( .A1(n6316), .A2(n6297), .ZN(n7839) );
  OR2_X1 U7475 ( .A1(n6249), .A2(n7839), .ZN(n6299) );
  INV_X1 U7476 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7477 ( .A1(n7572), .A2(n7813), .ZN(n6298) );
  OR2_X1 U7478 ( .A1(n7055), .A2(n6401), .ZN(n6307) );
  NOR2_X1 U7479 ( .A1(n6302), .A2(n9406), .ZN(n6303) );
  MUX2_X1 U7480 ( .A(n9406), .B(n6303), .S(P2_IR_REG_7__SCAN_IN), .Z(n6305) );
  INV_X1 U7481 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6304) );
  AND2_X1 U7482 ( .A1(n6302), .A2(n6304), .ZN(n6310) );
  OR2_X1 U7483 ( .A1(n6305), .A2(n6310), .ZN(n7821) );
  AOI22_X1 U7484 ( .A1(n6562), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7014), .B2(
        n7816), .ZN(n6306) );
  NAND2_X1 U7485 ( .A1(n6307), .A2(n6306), .ZN(n7912) );
  OR2_X1 U7486 ( .A1(n7761), .A2(n7912), .ZN(n7754) );
  NAND2_X1 U7487 ( .A1(n7761), .A2(n7912), .ZN(n8802) );
  NAND2_X1 U7488 ( .A1(n7754), .A2(n8802), .ZN(n7838) );
  INV_X1 U7489 ( .A(n7912), .ZN(n7905) );
  NAND2_X1 U7490 ( .A1(n7066), .A2(n8723), .ZN(n6314) );
  NOR2_X1 U7491 ( .A1(n6310), .A2(n9406), .ZN(n6308) );
  MUX2_X1 U7492 ( .A(n9406), .B(n6308), .S(P2_IR_REG_8__SCAN_IN), .Z(n6312) );
  NAND2_X1 U7493 ( .A1(n6310), .A2(n6309), .ZN(n6339) );
  INV_X1 U7494 ( .A(n6339), .ZN(n6311) );
  INV_X1 U7495 ( .A(n7884), .ZN(n7820) );
  AOI22_X1 U7496 ( .A1(n6562), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7014), .B2(
        n7820), .ZN(n6313) );
  NAND2_X1 U7497 ( .A1(n6314), .A2(n6313), .ZN(n7876) );
  NAND2_X1 U7498 ( .A1(n6248), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6321) );
  INV_X1 U7499 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6315) );
  OR2_X1 U7500 ( .A1(n6261), .A2(n6315), .ZN(n6320) );
  NAND2_X1 U7501 ( .A1(n6316), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6317) );
  AND2_X1 U7502 ( .A1(n6331), .A2(n6317), .ZN(n7757) );
  OR2_X1 U7503 ( .A1(n6249), .A2(n7757), .ZN(n6319) );
  INV_X1 U7504 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7817) );
  OR2_X1 U7505 ( .A1(n7572), .A2(n7817), .ZN(n6318) );
  OR2_X1 U7506 ( .A1(n7876), .A2(n7852), .ZN(n8797) );
  NAND2_X1 U7507 ( .A1(n7876), .A2(n7852), .ZN(n8803) );
  NAND2_X1 U7508 ( .A1(n8797), .A2(n8803), .ZN(n7755) );
  NAND2_X1 U7509 ( .A1(n7752), .A2(n7755), .ZN(n6323) );
  OR2_X1 U7510 ( .A1(n7876), .A2(n7941), .ZN(n6322) );
  NAND2_X1 U7511 ( .A1(n6323), .A2(n6322), .ZN(n7847) );
  NAND2_X1 U7512 ( .A1(n7073), .A2(n8723), .ZN(n6326) );
  NAND2_X1 U7513 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6324) );
  XNOR2_X1 U7514 ( .A(n6324), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7921) );
  AOI22_X1 U7515 ( .A1(n6562), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7014), .B2(
        n7921), .ZN(n6325) );
  NAND2_X1 U7516 ( .A1(n6587), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6336) );
  INV_X1 U7517 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6328) );
  OR2_X1 U7518 ( .A1(n6327), .A2(n6328), .ZN(n6335) );
  NAND2_X1 U7519 ( .A1(n6331), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6332) );
  AND2_X1 U7520 ( .A1(n6343), .A2(n6332), .ZN(n7745) );
  OR2_X1 U7521 ( .A1(n6249), .A2(n7745), .ZN(n6334) );
  OR2_X1 U7522 ( .A1(n7572), .A2(n7948), .ZN(n6333) );
  INV_X1 U7523 ( .A(n8924), .ZN(n7975) );
  NAND2_X1 U7524 ( .A1(n7950), .A2(n7975), .ZN(n8811) );
  NAND2_X1 U7525 ( .A1(n8813), .A2(n8811), .ZN(n7848) );
  NAND2_X1 U7526 ( .A1(n7847), .A2(n7848), .ZN(n6338) );
  OR2_X1 U7527 ( .A1(n7950), .A2(n8924), .ZN(n6337) );
  NAND2_X1 U7528 ( .A1(n6338), .A2(n6337), .ZN(n8154) );
  OR2_X1 U7529 ( .A1(n7072), .A2(n6244), .ZN(n6342) );
  NAND2_X1 U7530 ( .A1(n6349), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6340) );
  XNOR2_X1 U7531 ( .A(n6340), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7927) );
  AOI22_X1 U7532 ( .A1(n6562), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7014), .B2(
        n7927), .ZN(n6341) );
  NAND2_X1 U7533 ( .A1(n6342), .A2(n6341), .ZN(n10735) );
  NAND2_X1 U7534 ( .A1(n6248), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6348) );
  INV_X1 U7535 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7923) );
  OR2_X1 U7536 ( .A1(n7572), .A2(n7923), .ZN(n6347) );
  OR2_X2 U7537 ( .A1(n6343), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7538 ( .A1(n6343), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6344) );
  AND2_X1 U7539 ( .A1(n6354), .A2(n6344), .ZN(n8152) );
  OR2_X1 U7540 ( .A1(n6249), .A2(n8152), .ZN(n6346) );
  OR2_X1 U7541 ( .A1(n6261), .A2(n7926), .ZN(n6345) );
  NAND4_X1 U7542 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n8923)
         );
  NAND2_X1 U7543 ( .A1(n10735), .A2(n8923), .ZN(n8148) );
  OR2_X1 U7544 ( .A1(n10735), .A2(n8923), .ZN(n8149) );
  NAND2_X1 U7545 ( .A1(n7134), .A2(n8723), .ZN(n6352) );
  NAND2_X1 U7546 ( .A1(n6360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U7547 ( .A(n6350), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8072) );
  AOI22_X1 U7548 ( .A1(n6562), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7014), .B2(
        n8072), .ZN(n6351) );
  NAND2_X1 U7549 ( .A1(n6352), .A2(n6351), .ZN(n10743) );
  NAND2_X1 U7550 ( .A1(n6248), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6359) );
  INV_X1 U7551 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6353) );
  OR2_X1 U7552 ( .A1(n6261), .A2(n6353), .ZN(n6358) );
  OR2_X2 U7553 ( .A1(n6354), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U7554 ( .A1(n6354), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6355) );
  AND2_X1 U7555 ( .A1(n6365), .A2(n6355), .ZN(n8060) );
  OR2_X1 U7556 ( .A1(n6249), .A2(n8060), .ZN(n6357) );
  INV_X1 U7557 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8073) );
  OR2_X1 U7558 ( .A1(n7572), .A2(n8073), .ZN(n6356) );
  NAND4_X1 U7559 ( .A1(n6359), .A2(n6358), .A3(n6357), .A4(n6356), .ZN(n8163)
         );
  NAND2_X1 U7560 ( .A1(n10743), .A2(n8163), .ZN(n8092) );
  NAND2_X1 U7561 ( .A1(n8096), .A2(n8092), .ZN(n8162) );
  OR2_X1 U7562 ( .A1(n7160), .A2(n6244), .ZN(n6362) );
  XNOR2_X1 U7563 ( .A(n6373), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8939) );
  AOI22_X1 U7564 ( .A1(n6562), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7014), .B2(
        n8939), .ZN(n6361) );
  NAND2_X1 U7565 ( .A1(n6248), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6370) );
  INV_X1 U7566 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6363) );
  OR2_X1 U7567 ( .A1(n6261), .A2(n6363), .ZN(n6369) );
  NAND2_X1 U7568 ( .A1(n6365), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6366) );
  AND2_X1 U7569 ( .A1(n6380), .A2(n6366), .ZN(n8165) );
  OR2_X1 U7570 ( .A1(n6249), .A2(n8165), .ZN(n6368) );
  INV_X1 U7571 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8075) );
  OR2_X1 U7572 ( .A1(n7572), .A2(n8075), .ZN(n6367) );
  NAND4_X1 U7573 ( .A1(n6370), .A2(n6369), .A3(n6368), .A4(n6367), .ZN(n8195)
         );
  OR2_X1 U7574 ( .A1(n10766), .A2(n8195), .ZN(n6625) );
  NAND2_X1 U7575 ( .A1(n8162), .A2(n6625), .ZN(n6371) );
  NAND2_X1 U7576 ( .A1(n10766), .A2(n8195), .ZN(n8109) );
  NAND2_X1 U7577 ( .A1(n6371), .A2(n8109), .ZN(n8171) );
  OR2_X1 U7578 ( .A1(n7195), .A2(n6401), .ZN(n6376) );
  INV_X1 U7579 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7580 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  NAND2_X1 U7581 ( .A1(n6374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6389) );
  XNOR2_X1 U7582 ( .A(n6389), .B(n6388), .ZN(n8968) );
  INV_X1 U7583 ( .A(n8968), .ZN(n8952) );
  AOI22_X1 U7584 ( .A1(n6562), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7014), .B2(
        n8952), .ZN(n6375) );
  NAND2_X1 U7585 ( .A1(n6248), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6386) );
  INV_X1 U7586 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6377) );
  OR2_X1 U7587 ( .A1(n6261), .A2(n6377), .ZN(n6385) );
  INV_X1 U7588 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7589 ( .A1(n6380), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6381) );
  AND2_X1 U7590 ( .A1(n6393), .A2(n6381), .ZN(n8194) );
  OR2_X1 U7591 ( .A1(n6249), .A2(n8194), .ZN(n6384) );
  INV_X1 U7592 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6382) );
  OR2_X1 U7593 ( .A1(n7572), .A2(n6382), .ZN(n6383) );
  NAND4_X1 U7594 ( .A1(n6386), .A2(n6385), .A3(n6384), .A4(n6383), .ZN(n9262)
         );
  XNOR2_X1 U7595 ( .A(n8828), .B(n9262), .ZN(n8824) );
  NAND2_X1 U7596 ( .A1(n8171), .A2(n8756), .ZN(n8170) );
  NAND2_X1 U7597 ( .A1(n8828), .A2(n9262), .ZN(n6387) );
  NAND2_X1 U7598 ( .A1(n8170), .A2(n6387), .ZN(n9260) );
  NAND2_X1 U7599 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U7600 ( .A1(n6390), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6403) );
  XNOR2_X1 U7601 ( .A(n6403), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U7602 ( .A1(n6562), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7014), .B2(
        n10565), .ZN(n6391) );
  NAND2_X1 U7603 ( .A1(n6248), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6399) );
  INV_X1 U7604 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8966) );
  OR2_X1 U7605 ( .A1(n7572), .A2(n8966), .ZN(n6398) );
  NAND2_X1 U7606 ( .A1(n6393), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6394) );
  AND2_X1 U7607 ( .A1(n6408), .A2(n6394), .ZN(n9268) );
  OR2_X1 U7608 ( .A1(n6249), .A2(n9268), .ZN(n6397) );
  INV_X1 U7609 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6395) );
  OR2_X1 U7610 ( .A1(n6261), .A2(n6395), .ZN(n6396) );
  NAND4_X1 U7611 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n9246)
         );
  NAND2_X1 U7612 ( .A1(n10778), .A2(n9246), .ZN(n8834) );
  OR2_X1 U7613 ( .A1(n10778), .A2(n9246), .ZN(n6400) );
  NAND2_X1 U7614 ( .A1(n9260), .A2(n9259), .ZN(n9258) );
  NAND2_X1 U7615 ( .A1(n9258), .A2(n8834), .ZN(n9245) );
  INV_X1 U7616 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7617 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  NAND2_X1 U7618 ( .A1(n6404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6416) );
  XNOR2_X1 U7619 ( .A(n6416), .B(n6415), .ZN(n8991) );
  INV_X1 U7620 ( .A(n8991), .ZN(n8978) );
  AOI22_X1 U7621 ( .A1(n6562), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8978), .B2(
        n7014), .ZN(n6405) );
  NAND2_X1 U7622 ( .A1(n6248), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6413) );
  INV_X1 U7623 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9251) );
  OR2_X1 U7624 ( .A1(n6261), .A2(n9251), .ZN(n6412) );
  NAND2_X1 U7625 ( .A1(n6408), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6409) );
  AND2_X1 U7626 ( .A1(n6420), .A2(n6409), .ZN(n9250) );
  OR2_X1 U7627 ( .A1(n6249), .A2(n9250), .ZN(n6411) );
  INV_X1 U7628 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8949) );
  OR2_X1 U7629 ( .A1(n7572), .A2(n8949), .ZN(n6410) );
  NAND4_X1 U7630 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .ZN(n9261)
         );
  NAND2_X1 U7631 ( .A1(n9211), .A2(n8837), .ZN(n9244) );
  NAND2_X1 U7632 ( .A1(n9245), .A2(n9244), .ZN(n9243) );
  NAND2_X1 U7633 ( .A1(n9254), .A2(n9261), .ZN(n6414) );
  NAND2_X1 U7634 ( .A1(n9243), .A2(n6414), .ZN(n9231) );
  NAND2_X1 U7635 ( .A1(n7311), .A2(n8723), .ZN(n6419) );
  NAND2_X1 U7636 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  NAND2_X1 U7637 ( .A1(n6417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6428) );
  XNOR2_X1 U7638 ( .A(n6428), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9012) );
  AOI22_X1 U7639 ( .A1(n6562), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9012), .B2(
        n7014), .ZN(n6418) );
  NAND2_X1 U7640 ( .A1(n6248), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6425) );
  INV_X1 U7641 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9236) );
  OR2_X1 U7642 ( .A1(n6261), .A2(n9236), .ZN(n6424) );
  OR2_X2 U7643 ( .A1(n6420), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7644 ( .A1(n6420), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6421) );
  AND2_X1 U7645 ( .A1(n6435), .A2(n6421), .ZN(n9235) );
  OR2_X1 U7646 ( .A1(n6249), .A2(n9235), .ZN(n6423) );
  INV_X1 U7647 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9360) );
  OR2_X1 U7648 ( .A1(n7572), .A2(n9360), .ZN(n6422) );
  NAND4_X1 U7649 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n9247)
         );
  XNOR2_X1 U7650 ( .A(n8840), .B(n9247), .ZN(n9212) );
  NAND2_X1 U7651 ( .A1(n9231), .A2(n9230), .ZN(n9229) );
  NAND2_X1 U7652 ( .A1(n8840), .A2(n9247), .ZN(n6426) );
  NAND2_X1 U7653 ( .A1(n9229), .A2(n6426), .ZN(n9218) );
  NAND2_X1 U7654 ( .A1(n7567), .A2(n8723), .ZN(n6432) );
  NAND2_X1 U7655 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  NAND2_X1 U7656 ( .A1(n6429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6430) );
  XNOR2_X1 U7657 ( .A(n6430), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9028) );
  AOI22_X1 U7658 ( .A1(n9028), .A2(n7014), .B1(n6562), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6431) );
  NAND2_X2 U7659 ( .A1(n6432), .A2(n6431), .ZN(n9355) );
  NAND2_X1 U7660 ( .A1(n6248), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6441) );
  INV_X1 U7661 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9224) );
  OR2_X1 U7662 ( .A1(n6261), .A2(n9224), .ZN(n6440) );
  INV_X1 U7663 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U7664 ( .A1(n6435), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6436) );
  AND2_X1 U7665 ( .A1(n6446), .A2(n6436), .ZN(n9223) );
  OR2_X1 U7666 ( .A1(n6249), .A2(n9223), .ZN(n6439) );
  INV_X1 U7667 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6437) );
  OR2_X1 U7668 ( .A1(n7572), .A2(n6437), .ZN(n6438) );
  NAND4_X1 U7669 ( .A1(n6441), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n9232)
         );
  XNOR2_X1 U7670 ( .A(n9355), .B(n9204), .ZN(n9217) );
  NAND2_X1 U7671 ( .A1(n9218), .A2(n9217), .ZN(n9216) );
  NAND2_X1 U7672 ( .A1(n9355), .A2(n9232), .ZN(n6442) );
  NAND2_X1 U7673 ( .A1(n9216), .A2(n6442), .ZN(n9201) );
  OR2_X1 U7674 ( .A1(n7539), .A2(n6244), .ZN(n6445) );
  NAND2_X1 U7675 ( .A1(n5354), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6443) );
  XNOR2_X1 U7676 ( .A(n6443), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9052) );
  AOI22_X1 U7677 ( .A1(n6562), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7014), .B2(
        n9052), .ZN(n6444) );
  OR2_X2 U7678 ( .A1(n6446), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7679 ( .A1(n6446), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U7680 ( .A1(n6459), .A2(n6447), .ZN(n9205) );
  NAND2_X1 U7681 ( .A1(n6585), .A2(n9205), .ZN(n6451) );
  INV_X1 U7682 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9207) );
  OR2_X1 U7683 ( .A1(n6261), .A2(n9207), .ZN(n6450) );
  INV_X1 U7684 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9396) );
  OR2_X1 U7685 ( .A1(n6327), .A2(n9396), .ZN(n6449) );
  INV_X1 U7686 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9352) );
  OR2_X1 U7687 ( .A1(n7572), .A2(n9352), .ZN(n6448) );
  NAND4_X1 U7688 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n9219)
         );
  OR2_X1 U7689 ( .A1(n9348), .A2(n9219), .ZN(n6452) );
  NAND2_X1 U7690 ( .A1(n9201), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U7691 ( .A1(n9348), .A2(n9219), .ZN(n6453) );
  NAND2_X1 U7692 ( .A1(n7620), .A2(n8723), .ZN(n6457) );
  NAND2_X1 U7693 ( .A1(n6455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6595) );
  AOI22_X1 U7694 ( .A1(n6562), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9056), .B2(
        n7014), .ZN(n6456) );
  NAND2_X1 U7695 ( .A1(n6459), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U7696 ( .A1(n6469), .A2(n6460), .ZN(n9187) );
  NAND2_X1 U7697 ( .A1(n6585), .A2(n9187), .ZN(n6465) );
  INV_X1 U7698 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6461) );
  OR2_X1 U7699 ( .A1(n6261), .A2(n6461), .ZN(n6464) );
  INV_X1 U7700 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9393) );
  OR2_X1 U7701 ( .A1(n6327), .A2(n9393), .ZN(n6463) );
  INV_X1 U7702 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9346) );
  OR2_X1 U7703 ( .A1(n7572), .A2(n9346), .ZN(n6462) );
  NAND4_X1 U7704 ( .A1(n6465), .A2(n6464), .A3(n6463), .A4(n6462), .ZN(n9333)
         );
  AND2_X1 U7705 ( .A1(n9186), .A2(n9333), .ZN(n6466) );
  NAND2_X1 U7706 ( .A1(n7695), .A2(n8723), .ZN(n6468) );
  NAND2_X1 U7707 ( .A1(n6562), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7708 ( .A1(n6469), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7709 ( .A1(n6478), .A2(n6470), .ZN(n9172) );
  NAND2_X1 U7710 ( .A1(n9172), .A2(n6585), .ZN(n6474) );
  NAND2_X1 U7711 ( .A1(n6587), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U7712 ( .A1(n6248), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U7713 ( .A1(n6202), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6471) );
  NAND4_X1 U7714 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n9325)
         );
  XNOR2_X1 U7715 ( .A(n9177), .B(n9182), .ZN(n9168) );
  NAND2_X1 U7716 ( .A1(n7857), .A2(n8723), .ZN(n6476) );
  NAND2_X1 U7717 ( .A1(n6562), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6475) );
  INV_X1 U7718 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U7719 ( .A1(n6478), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7720 ( .A1(n6493), .A2(n6479), .ZN(n9160) );
  NAND2_X1 U7721 ( .A1(n9160), .A2(n6585), .ZN(n6481) );
  AOI22_X1 U7722 ( .A1(n6587), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6248), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6480) );
  OAI211_X1 U7723 ( .C1(n7572), .C2(n6482), .A(n6481), .B(n6480), .ZN(n9336)
         );
  INV_X1 U7724 ( .A(n9336), .ZN(n9315) );
  NAND2_X1 U7725 ( .A1(n9385), .A2(n9315), .ZN(n8864) );
  NAND2_X1 U7726 ( .A1(n8863), .A2(n8864), .ZN(n9159) );
  NAND2_X1 U7727 ( .A1(n7964), .A2(n8723), .ZN(n6484) );
  NAND2_X1 U7728 ( .A1(n6562), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U7729 ( .A1(n6495), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U7730 ( .A1(n6513), .A2(n6485), .ZN(n9138) );
  NAND2_X1 U7731 ( .A1(n9138), .A2(n6585), .ZN(n6490) );
  INV_X1 U7732 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U7733 ( .A1(n6248), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7734 ( .A1(n6587), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6486) );
  OAI211_X1 U7735 ( .C1(n9312), .C2(n7572), .A(n6487), .B(n6486), .ZN(n6488)
         );
  INV_X1 U7736 ( .A(n6488), .ZN(n6489) );
  NAND2_X1 U7737 ( .A1(n9137), .A2(n9146), .ZN(n6502) );
  INV_X1 U7738 ( .A(n6502), .ZN(n6501) );
  NAND2_X1 U7739 ( .A1(n7896), .A2(n8723), .ZN(n6492) );
  NAND2_X1 U7740 ( .A1(n6562), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6491) );
  INV_X1 U7741 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U7742 ( .A1(n6493), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7743 ( .A1(n6495), .A2(n6494), .ZN(n9147) );
  NAND2_X1 U7744 ( .A1(n9147), .A2(n6585), .ZN(n6497) );
  AOI22_X1 U7745 ( .A1(n6587), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n6248), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6496) );
  OAI211_X1 U7746 ( .C1(n7572), .C2(n6498), .A(n6497), .B(n6496), .ZN(n9326)
         );
  OR2_X1 U7747 ( .A1(n9320), .A2(n9326), .ZN(n9127) );
  OR2_X1 U7748 ( .A1(n9137), .A2(n9146), .ZN(n6499) );
  AND2_X1 U7749 ( .A1(n9127), .A2(n6499), .ZN(n6500) );
  OR2_X1 U7750 ( .A1(n6501), .A2(n6500), .ZN(n6507) );
  INV_X1 U7751 ( .A(n6507), .ZN(n6504) );
  NAND2_X1 U7752 ( .A1(n9320), .A2(n9326), .ZN(n9129) );
  AND2_X1 U7753 ( .A1(n9129), .A2(n6502), .ZN(n6503) );
  AND2_X1 U7754 ( .A1(n9159), .A2(n6506), .ZN(n6505) );
  NAND2_X1 U7755 ( .A1(n9126), .A2(n6505), .ZN(n9113) );
  INV_X1 U7756 ( .A(n6506), .ZN(n6509) );
  OR2_X1 U7757 ( .A1(n9385), .A2(n9336), .ZN(n9143) );
  AND2_X1 U7758 ( .A1(n9143), .A2(n6507), .ZN(n6508) );
  NAND2_X1 U7759 ( .A1(n8009), .A2(n8723), .ZN(n6511) );
  NAND2_X1 U7760 ( .A1(n6562), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6510) );
  INV_X1 U7761 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U7762 ( .A1(n6513), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U7763 ( .A1(n6527), .A2(n6514), .ZN(n9122) );
  NAND2_X1 U7764 ( .A1(n9122), .A2(n6585), .ZN(n6519) );
  INV_X1 U7765 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U7766 ( .A1(n6587), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U7767 ( .A1(n6248), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6515) );
  OAI211_X1 U7768 ( .C1(n9308), .C2(n7572), .A(n6516), .B(n6515), .ZN(n6517)
         );
  INV_X1 U7769 ( .A(n6517), .ZN(n6518) );
  OR2_X1 U7770 ( .A1(n8873), .A2(n9300), .ZN(n6520) );
  AND2_X1 U7771 ( .A1(n9112), .A2(n6520), .ZN(n6521) );
  NAND2_X1 U7772 ( .A1(n9113), .A2(n6521), .ZN(n6523) );
  NAND2_X1 U7773 ( .A1(n8873), .A2(n9300), .ZN(n6522) );
  NAND2_X1 U7774 ( .A1(n6523), .A2(n6522), .ZN(n9102) );
  NAND2_X1 U7775 ( .A1(n8128), .A2(n8723), .ZN(n6525) );
  NAND2_X1 U7776 ( .A1(n6562), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6524) );
  INV_X1 U7777 ( .A(n6527), .ZN(n6526) );
  INV_X1 U7778 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U7779 ( .A1(n6527), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U7780 ( .A1(n6539), .A2(n6528), .ZN(n9105) );
  NAND2_X1 U7781 ( .A1(n9105), .A2(n6585), .ZN(n6534) );
  INV_X1 U7782 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U7783 ( .A1(n6587), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U7784 ( .A1(n6248), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6529) );
  OAI211_X1 U7785 ( .C1(n6531), .C2(n7572), .A(n6530), .B(n6529), .ZN(n6532)
         );
  INV_X1 U7786 ( .A(n6532), .ZN(n6533) );
  AND2_X1 U7787 ( .A1(n9301), .A2(n8922), .ZN(n6536) );
  OR2_X1 U7788 ( .A1(n9301), .A2(n8922), .ZN(n6535) );
  NAND2_X1 U7789 ( .A1(n8201), .A2(n8723), .ZN(n6538) );
  NAND2_X1 U7790 ( .A1(n6562), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7791 ( .A1(n6539), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U7792 ( .A1(n6552), .A2(n6540), .ZN(n9094) );
  NAND2_X1 U7793 ( .A1(n9094), .A2(n6585), .ZN(n6546) );
  INV_X1 U7794 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7795 ( .A1(n6587), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U7796 ( .A1(n6248), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6541) );
  OAI211_X1 U7797 ( .C1(n6543), .C2(n7572), .A(n6542), .B(n6541), .ZN(n6544)
         );
  INV_X1 U7798 ( .A(n6544), .ZN(n6545) );
  NAND2_X2 U7799 ( .A1(n6546), .A2(n6545), .ZN(n9103) );
  NOR2_X1 U7800 ( .A1(n9295), .A2(n9103), .ZN(n6547) );
  NAND2_X1 U7801 ( .A1(n9295), .A2(n9103), .ZN(n6548) );
  NAND2_X1 U7802 ( .A1(n9414), .A2(n8723), .ZN(n6550) );
  NAND2_X1 U7803 ( .A1(n6562), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6549) );
  INV_X1 U7804 ( .A(n6552), .ZN(n6551) );
  INV_X1 U7805 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U7806 ( .A1(n6551), .A2(n9703), .ZN(n6565) );
  NAND2_X1 U7807 ( .A1(n6552), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U7808 ( .A1(n6565), .A2(n6553), .ZN(n9084) );
  NAND2_X1 U7809 ( .A1(n9084), .A2(n6585), .ZN(n6559) );
  INV_X1 U7810 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7811 ( .A1(n6587), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7812 ( .A1(n6248), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6554) );
  OAI211_X1 U7813 ( .C1(n6556), .C2(n7572), .A(n6555), .B(n6554), .ZN(n6557)
         );
  INV_X1 U7814 ( .A(n6557), .ZN(n6558) );
  OR2_X1 U7815 ( .A1(n9287), .A2(n8921), .ZN(n6560) );
  NAND2_X1 U7816 ( .A1(n6561), .A2(n6560), .ZN(n9074) );
  NAND2_X1 U7817 ( .A1(n8583), .A2(n8723), .ZN(n6564) );
  NAND2_X1 U7818 ( .A1(n6562), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7819 ( .A1(n6565), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U7820 ( .A1(n8522), .A2(n6566), .ZN(n9075) );
  NAND2_X1 U7821 ( .A1(n9075), .A2(n6585), .ZN(n6572) );
  INV_X1 U7822 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U7823 ( .A1(n6587), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U7824 ( .A1(n6248), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6567) );
  OAI211_X1 U7825 ( .C1(n6569), .C2(n7572), .A(n6568), .B(n6567), .ZN(n6570)
         );
  INV_X1 U7826 ( .A(n6570), .ZN(n6571) );
  NOR2_X1 U7827 ( .A1(n9281), .A2(n8920), .ZN(n6573) );
  INV_X1 U7828 ( .A(n9281), .ZN(n8886) );
  OAI22_X1 U7829 ( .A1(n9074), .A2(n6573), .B1(n9285), .B2(n8886), .ZN(n6593)
         );
  NAND2_X1 U7830 ( .A1(n6574), .A2(n6576), .ZN(n6581) );
  INV_X1 U7831 ( .A(n6577), .ZN(n6578) );
  NAND2_X1 U7832 ( .A1(n6578), .A2(n9571), .ZN(n6579) );
  INV_X1 U7833 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6582) );
  INV_X1 U7834 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9412) );
  MUX2_X1 U7835 ( .A(n6582), .B(n9412), .S(n5701), .Z(n8222) );
  NAND2_X1 U7836 ( .A1(n9411), .A2(n8723), .ZN(n6584) );
  OR2_X1 U7837 ( .A1(n6274), .A2(n9412), .ZN(n6583) );
  INV_X1 U7838 ( .A(n8522), .ZN(n6586) );
  NAND2_X1 U7839 ( .A1(n6586), .A2(n6585), .ZN(n7576) );
  NAND2_X1 U7840 ( .A1(n6248), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U7841 ( .A1(n6587), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6588) );
  OAI211_X1 U7842 ( .C1(n7572), .C2(n6983), .A(n6589), .B(n6588), .ZN(n6590)
         );
  INV_X1 U7843 ( .A(n6590), .ZN(n6591) );
  XNOR2_X1 U7844 ( .A(n8726), .B(n9279), .ZN(n8896) );
  INV_X1 U7845 ( .A(n8896), .ZN(n6592) );
  XNOR2_X1 U7846 ( .A(n6593), .B(n6592), .ZN(n6616) );
  NAND2_X1 U7847 ( .A1(n6595), .A2(n6594), .ZN(n6596) );
  NAND2_X1 U7848 ( .A1(n6602), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6598) );
  OR2_X1 U7849 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  OR2_X1 U7850 ( .A1(n8771), .A2(n8906), .ZN(n6604) );
  NAND2_X1 U7851 ( .A1(n4972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7852 ( .A1(n8915), .A2(n9056), .ZN(n6680) );
  INV_X1 U7853 ( .A(n8585), .ZN(n8912) );
  INV_X1 U7854 ( .A(n9417), .ZN(n7028) );
  NAND2_X1 U7855 ( .A1(n8912), .A2(n7028), .ZN(n6607) );
  NAND2_X1 U7856 ( .A1(n7009), .A2(n6607), .ZN(n7230) );
  AND2_X1 U7857 ( .A1(n7009), .A2(P2_B_REG_SCAN_IN), .ZN(n6608) );
  NOR2_X1 U7858 ( .A1(n9316), .A2(n6608), .ZN(n9065) );
  INV_X1 U7859 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U7860 ( .A1(n6248), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6611) );
  INV_X1 U7861 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6609) );
  OR2_X1 U7862 ( .A1(n6261), .A2(n6609), .ZN(n6610) );
  OAI211_X1 U7863 ( .C1(n6612), .C2(n7572), .A(n6611), .B(n6610), .ZN(n6613)
         );
  INV_X1 U7864 ( .A(n6613), .ZN(n6614) );
  NAND2_X1 U7865 ( .A1(n7576), .A2(n6614), .ZN(n8919) );
  AOI22_X1 U7866 ( .A1(n8920), .A2(n9334), .B1(n9065), .B2(n8919), .ZN(n6615)
         );
  NAND2_X1 U7867 ( .A1(n7456), .A2(n8772), .ZN(n7461) );
  INV_X1 U7868 ( .A(n7460), .ZN(n8766) );
  NOR2_X1 U7869 ( .A1(n6617), .A2(n8768), .ZN(n6618) );
  AOI21_X1 U7870 ( .B1(n8772), .B2(n8766), .A(n6618), .ZN(n8777) );
  NAND2_X1 U7871 ( .A1(n7461), .A2(n8777), .ZN(n7499) );
  NAND2_X1 U7872 ( .A1(n8929), .A2(n7587), .ZN(n8781) );
  NAND2_X1 U7873 ( .A1(n7498), .A2(n8785), .ZN(n7515) );
  OR2_X1 U7874 ( .A1(n7579), .A2(n7428), .ZN(n8786) );
  NAND2_X1 U7875 ( .A1(n7579), .A2(n7428), .ZN(n8782) );
  NAND2_X1 U7876 ( .A1(n7515), .A2(n8779), .ZN(n7514) );
  NAND2_X1 U7877 ( .A1(n7514), .A2(n8782), .ZN(n7779) );
  INV_X1 U7878 ( .A(n8927), .ZN(n7535) );
  NAND2_X1 U7879 ( .A1(n7535), .A2(n7521), .ZN(n8790) );
  INV_X1 U7880 ( .A(n7521), .ZN(n10720) );
  NAND2_X1 U7881 ( .A1(n8927), .A2(n10720), .ZN(n8787) );
  NAND2_X1 U7882 ( .A1(n7779), .A2(n8744), .ZN(n7766) );
  NAND2_X1 U7883 ( .A1(n7766), .A2(n8790), .ZN(n6619) );
  INV_X1 U7884 ( .A(n8926), .ZN(n7843) );
  NAND2_X1 U7885 ( .A1(n7843), .A2(n7775), .ZN(n8795) );
  INV_X1 U7886 ( .A(n7775), .ZN(n10727) );
  NAND2_X1 U7887 ( .A1(n8926), .A2(n10727), .ZN(n8794) );
  AND2_X1 U7888 ( .A1(n8797), .A2(n7754), .ZN(n8810) );
  NAND2_X1 U7889 ( .A1(n7753), .A2(n8810), .ZN(n6620) );
  NAND2_X1 U7890 ( .A1(n6620), .A2(n8803), .ZN(n7854) );
  INV_X1 U7891 ( .A(n7854), .ZN(n6622) );
  INV_X1 U7892 ( .A(n7848), .ZN(n6621) );
  INV_X1 U7893 ( .A(n8923), .ZN(n7747) );
  INV_X1 U7894 ( .A(n8163), .ZN(n6623) );
  NAND2_X1 U7895 ( .A1(n10743), .A2(n6623), .ZN(n8809) );
  NAND2_X1 U7896 ( .A1(n10735), .A2(n7747), .ZN(n8804) );
  AND2_X1 U7897 ( .A1(n8809), .A2(n8804), .ZN(n8816) );
  NAND2_X1 U7898 ( .A1(n8090), .A2(n8816), .ZN(n6624) );
  OR2_X1 U7899 ( .A1(n10743), .A2(n6623), .ZN(n8818) );
  NAND2_X1 U7900 ( .A1(n6625), .A2(n8109), .ZN(n8819) );
  INV_X1 U7901 ( .A(n8195), .ZN(n8820) );
  OR2_X1 U7902 ( .A1(n10766), .A2(n8820), .ZN(n8821) );
  INV_X1 U7903 ( .A(n9262), .ZN(n8827) );
  OR2_X1 U7904 ( .A1(n8828), .A2(n8827), .ZN(n8830) );
  INV_X1 U7905 ( .A(n9246), .ZN(n8833) );
  NAND2_X1 U7906 ( .A1(n10778), .A2(n8833), .ZN(n6627) );
  INV_X1 U7907 ( .A(n9217), .ZN(n6628) );
  INV_X1 U7908 ( .A(n9247), .ZN(n8713) );
  OR2_X1 U7909 ( .A1(n8840), .A2(n8713), .ZN(n9213) );
  AND2_X1 U7910 ( .A1(n6628), .A2(n9213), .ZN(n6629) );
  AND2_X1 U7911 ( .A1(n9211), .A2(n6629), .ZN(n6633) );
  INV_X1 U7912 ( .A(n6629), .ZN(n6630) );
  OR2_X1 U7913 ( .A1(n6630), .A2(n9212), .ZN(n6631) );
  NAND2_X1 U7914 ( .A1(n9348), .A2(n9183), .ZN(n8847) );
  NAND2_X1 U7915 ( .A1(n9355), .A2(n9204), .ZN(n9196) );
  AND2_X1 U7916 ( .A1(n9200), .A2(n9196), .ZN(n6634) );
  NAND2_X1 U7917 ( .A1(n9198), .A2(n8850), .ZN(n9185) );
  NAND2_X1 U7918 ( .A1(n9185), .A2(n8740), .ZN(n6635) );
  INV_X1 U7919 ( .A(n9333), .ZN(n9203) );
  OR2_X1 U7920 ( .A1(n9186), .A2(n9203), .ZN(n8855) );
  INV_X1 U7921 ( .A(n9177), .ZN(n9391) );
  NAND2_X1 U7922 ( .A1(n9320), .A2(n9134), .ZN(n6636) );
  NAND2_X1 U7923 ( .A1(n6637), .A2(n6636), .ZN(n9136) );
  XNOR2_X1 U7924 ( .A(n9137), .B(n9146), .ZN(n9135) );
  AND2_X1 U7925 ( .A1(n9137), .A2(n8559), .ZN(n8869) );
  AOI21_X1 U7926 ( .B1(n9136), .B2(n9135), .A(n8869), .ZN(n9119) );
  XNOR2_X1 U7927 ( .A(n8873), .B(n9300), .ZN(n9118) );
  NAND2_X1 U7928 ( .A1(n9119), .A2(n9118), .ZN(n9121) );
  OR2_X1 U7929 ( .A1(n8873), .A2(n9133), .ZN(n8874) );
  NOR2_X1 U7930 ( .A1(n9301), .A2(n9292), .ZN(n8878) );
  NAND2_X1 U7931 ( .A1(n9301), .A2(n9292), .ZN(n8739) );
  AND2_X1 U7932 ( .A1(n8883), .A2(n9081), .ZN(n6644) );
  NAND2_X1 U7933 ( .A1(n9082), .A2(n6644), .ZN(n6638) );
  NAND2_X1 U7934 ( .A1(n9287), .A2(n9293), .ZN(n8884) );
  NAND2_X1 U7935 ( .A1(n6638), .A2(n8884), .ZN(n9072) );
  NAND2_X1 U7936 ( .A1(n9281), .A2(n9285), .ZN(n6641) );
  INV_X1 U7937 ( .A(n9073), .ZN(n6639) );
  NAND2_X1 U7938 ( .A1(n9072), .A2(n6639), .ZN(n6640) );
  NAND2_X1 U7939 ( .A1(n6640), .A2(n6641), .ZN(n8731) );
  NAND2_X1 U7940 ( .A1(n8731), .A2(n6592), .ZN(n6649) );
  INV_X1 U7941 ( .A(n8883), .ZN(n6642) );
  OAI211_X1 U7942 ( .C1(n6642), .C2(n5517), .A(n6641), .B(n8884), .ZN(n6643)
         );
  AOI21_X1 U7943 ( .B1(n9092), .B2(n6644), .A(n6643), .ZN(n6647) );
  INV_X1 U7944 ( .A(n6645), .ZN(n6646) );
  INV_X1 U7945 ( .A(n9056), .ZN(n7645) );
  INV_X1 U7946 ( .A(n8915), .ZN(n7908) );
  NAND2_X1 U7947 ( .A1(n7645), .A2(n8915), .ZN(n6975) );
  INV_X1 U7948 ( .A(n6975), .ZN(n6650) );
  NOR2_X1 U7949 ( .A1(n6977), .A2(n6650), .ZN(n6651) );
  INV_X1 U7950 ( .A(n7486), .ZN(n8155) );
  NAND2_X1 U7951 ( .A1(n8527), .A2(n8155), .ZN(n6652) );
  NAND2_X1 U7952 ( .A1(n8906), .A2(n9056), .ZN(n7468) );
  OR2_X1 U7953 ( .A1(n7468), .A2(n8915), .ZN(n7282) );
  INV_X1 U7954 ( .A(n7282), .ZN(n10733) );
  NAND2_X1 U7955 ( .A1(n8527), .A2(n10733), .ZN(n6653) );
  NAND2_X1 U7956 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  NAND2_X1 U7957 ( .A1(n6657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U7958 ( .A1(n6660), .A2(n8145), .ZN(n6666) );
  NAND2_X1 U7959 ( .A1(n6661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U7960 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6662), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6665) );
  INV_X1 U7961 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U7962 ( .A1(n8145), .A2(n8204), .ZN(n7081) );
  NAND2_X1 U7963 ( .A1(n8204), .A2(n8516), .ZN(n7084) );
  NOR2_X1 U7964 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6672) );
  NOR4_X1 U7965 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6671) );
  NOR4_X1 U7966 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6670) );
  NOR4_X1 U7967 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6669) );
  NAND4_X1 U7968 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6678)
         );
  NOR4_X1 U7969 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6676) );
  NOR4_X1 U7970 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6675) );
  NOR4_X1 U7971 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6674) );
  NOR4_X1 U7972 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6673) );
  NAND4_X1 U7973 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6677)
         );
  NOR2_X1 U7974 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  NAND2_X1 U7975 ( .A1(n6974), .A2(n6972), .ZN(n7211) );
  NOR2_X1 U7976 ( .A1(n6680), .A2(n8906), .ZN(n6681) );
  NAND2_X1 U7977 ( .A1(n8771), .A2(n6681), .ZN(n7204) );
  OR2_X1 U7978 ( .A1(n7211), .A2(n7204), .ZN(n6685) );
  NAND3_X1 U7979 ( .A1(n7452), .A2(n6668), .A3(n6972), .ZN(n7216) );
  INV_X1 U7980 ( .A(n7216), .ZN(n6683) );
  INV_X1 U7981 ( .A(n7468), .ZN(n7212) );
  OR2_X1 U7982 ( .A1(n10785), .A2(n7212), .ZN(n8174) );
  NAND3_X1 U7983 ( .A1(n5034), .A2(n10785), .A3(n7204), .ZN(n6682) );
  NAND2_X1 U7984 ( .A1(n8174), .A2(n6682), .ZN(n7196) );
  NAND2_X1 U7985 ( .A1(n6683), .A2(n7196), .ZN(n6684) );
  NAND2_X1 U7986 ( .A1(n6685), .A2(n6684), .ZN(n6693) );
  INV_X1 U7987 ( .A(n8145), .ZN(n6687) );
  INV_X1 U7988 ( .A(n8516), .ZN(n6686) );
  NAND2_X1 U7989 ( .A1(n4999), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U7990 ( .A1(n6693), .A2(n7206), .ZN(n6692) );
  NAND2_X1 U7991 ( .A1(n7206), .A2(n7506), .ZN(n7215) );
  INV_X2 U7992 ( .A(n10792), .ZN(n6696) );
  NAND2_X1 U7993 ( .A1(n7206), .A2(n10777), .ZN(n7210) );
  INV_X1 U7994 ( .A(n9403), .ZN(n9386) );
  INV_X1 U7995 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6695) );
  NOR2_X1 U7996 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  NAND2_X1 U7997 ( .A1(n6699), .A2(n6698), .ZN(P2_U3456) );
  INV_X1 U7998 ( .A(n9938), .ZN(n9782) );
  NAND2_X1 U7999 ( .A1(n9411), .A2(n8273), .ZN(n6703) );
  NAND2_X1 U8000 ( .A1(n8230), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U8001 ( .A1(n6714), .A2(n7243), .ZN(n8392) );
  XNOR2_X1 U8002 ( .A(n6704), .B(n8281), .ZN(n9911) );
  NAND2_X1 U8003 ( .A1(n9911), .A2(n10754), .ZN(n6720) );
  INV_X1 U8004 ( .A(n8420), .ZN(n8279) );
  AOI21_X1 U8005 ( .B1(n6706), .B2(n6705), .A(n8279), .ZN(n6707) );
  XNOR2_X1 U8006 ( .A(n8281), .B(n6707), .ZN(n6713) );
  INV_X1 U8007 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8008 ( .A1(n4927), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U8009 ( .A1(n5757), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6708) );
  OAI211_X1 U8010 ( .C1(n7060), .C2(n6710), .A(n6709), .B(n6708), .ZN(n9781)
         );
  INV_X1 U8011 ( .A(n9781), .ZN(n8262) );
  XNOR2_X1 U8012 ( .A(n6173), .B(n5699), .ZN(n10364) );
  AND2_X1 U8013 ( .A1(n10364), .A2(P1_B_REG_SCAN_IN), .ZN(n6711) );
  OR2_X1 U8014 ( .A1(n10703), .A2(n6711), .ZN(n9900) );
  OAI22_X1 U8015 ( .A1(n9938), .A2(n10701), .B1(n8262), .B2(n9900), .ZN(n6712)
         );
  AOI21_X1 U8016 ( .B1(n6713), .B2(n10659), .A(n6712), .ZN(n9922) );
  INV_X1 U8017 ( .A(n6714), .ZN(n6717) );
  INV_X1 U8018 ( .A(n6715), .ZN(n6716) );
  OAI211_X1 U8019 ( .C1(n6717), .C2(n6716), .A(n10192), .B(n9903), .ZN(n9912)
         );
  NAND2_X1 U8020 ( .A1(n6714), .A2(n10663), .ZN(n9916) );
  NAND2_X1 U8021 ( .A1(n6720), .A2(n6719), .ZN(n10203) );
  OR2_X1 U8022 ( .A1(n10757), .A2(n6170), .ZN(n6721) );
  NAND2_X1 U8023 ( .A1(n6951), .A2(n6726), .ZN(n6728) );
  INV_X1 U8024 ( .A(n6728), .ZN(n6723) );
  AND2_X2 U8025 ( .A1(n6723), .A2(n6729), .ZN(n6801) );
  NAND2_X1 U8026 ( .A1(n6724), .A2(n6801), .ZN(n6733) );
  NAND2_X1 U8027 ( .A1(n6725), .A2(n10692), .ZN(n6727) );
  NAND2_X1 U8028 ( .A1(n10607), .A2(n6726), .ZN(n8027) );
  NAND3_X1 U8029 ( .A1(n6727), .A2(n6729), .A3(n8027), .ZN(n6738) );
  NAND2_X2 U8030 ( .A1(n6738), .A2(n6744), .ZN(n6759) );
  NAND2_X1 U8031 ( .A1(n6759), .A2(n6731), .ZN(n6732) );
  NAND2_X1 U8032 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  NAND2_X1 U8033 ( .A1(n6759), .A2(n10193), .ZN(n6736) );
  NAND2_X1 U8034 ( .A1(n6739), .A2(n6801), .ZN(n6735) );
  NAND2_X1 U8035 ( .A1(n6736), .A2(n6735), .ZN(n6743) );
  INV_X1 U8036 ( .A(n6743), .ZN(n6737) );
  NAND2_X1 U8037 ( .A1(n6737), .A2(n5507), .ZN(n7089) );
  NAND2_X1 U8038 ( .A1(n6881), .A2(n6739), .ZN(n6742) );
  OAI22_X1 U8039 ( .A1(n4926), .A2(n10606), .B1(n6729), .B2(n10365), .ZN(n6740) );
  INV_X1 U8040 ( .A(n6740), .ZN(n6741) );
  NAND2_X1 U8041 ( .A1(n6742), .A2(n6741), .ZN(n7088) );
  CLKBUF_X3 U8042 ( .A(n6744), .Z(n6930) );
  NAND3_X1 U8043 ( .A1(n6745), .A2(n7090), .A3(n6749), .ZN(n6748) );
  NAND2_X1 U8044 ( .A1(n6881), .A2(n6724), .ZN(n6747) );
  NAND2_X1 U8045 ( .A1(n6801), .A2(n6731), .ZN(n6746) );
  NAND2_X1 U8046 ( .A1(n6747), .A2(n6746), .ZN(n7149) );
  NAND2_X1 U8047 ( .A1(n6748), .A2(n7149), .ZN(n7148) );
  NAND2_X1 U8048 ( .A1(n7090), .A2(n6749), .ZN(n7147) );
  NAND2_X1 U8049 ( .A1(n7147), .A2(n6750), .ZN(n7152) );
  NOR2_X1 U8050 ( .A1(n6751), .A2(n5513), .ZN(n6756) );
  NAND2_X1 U8051 ( .A1(n6752), .A2(n6759), .ZN(n6753) );
  INV_X2 U8052 ( .A(n6930), .ZN(n6777) );
  XNOR2_X1 U8053 ( .A(n6754), .B(n6777), .ZN(n6755) );
  NAND2_X1 U8054 ( .A1(n6755), .A2(n6756), .ZN(n6758) );
  OAI21_X1 U8055 ( .B1(n6756), .B2(n6755), .A(n6758), .ZN(n6757) );
  NAND2_X1 U8056 ( .A1(n7139), .A2(n7141), .ZN(n7140) );
  NAND2_X1 U8057 ( .A1(n7140), .A2(n6758), .ZN(n7167) );
  NAND2_X1 U8058 ( .A1(n6759), .A2(n10662), .ZN(n6761) );
  NAND2_X1 U8059 ( .A1(n9798), .A2(n6801), .ZN(n6760) );
  NAND2_X1 U8060 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  AOI22_X1 U8061 ( .A1(n6881), .A2(n9798), .B1(n6927), .B2(n10662), .ZN(n6764)
         );
  XNOR2_X1 U8062 ( .A(n6763), .B(n6764), .ZN(n7168) );
  NAND2_X1 U8063 ( .A1(n7167), .A2(n7168), .ZN(n7166) );
  INV_X1 U8064 ( .A(n6763), .ZN(n6765) );
  NAND2_X1 U8065 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  NAND2_X1 U8066 ( .A1(n7166), .A2(n6766), .ZN(n7244) );
  OAI22_X1 U8067 ( .A1(n10689), .A2(n6810), .B1(n10654), .B2(n4926), .ZN(n6767) );
  XNOR2_X1 U8068 ( .A(n6767), .B(n6930), .ZN(n6770) );
  OAI22_X1 U8069 ( .A1(n10689), .A2(n4926), .B1(n10654), .B2(n6988), .ZN(n6769) );
  XNOR2_X1 U8070 ( .A(n6770), .B(n6769), .ZN(n7247) );
  NAND2_X1 U8071 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  OAI22_X1 U8072 ( .A1(n7321), .A2(n6810), .B1(n10702), .B2(n4926), .ZN(n6772)
         );
  XNOR2_X1 U8073 ( .A(n6772), .B(n6930), .ZN(n6774) );
  AND2_X1 U8074 ( .A1(n6881), .A2(n7056), .ZN(n6773) );
  AOI21_X1 U8075 ( .B1(n7393), .B2(n6927), .A(n6773), .ZN(n7292) );
  NAND2_X1 U8076 ( .A1(n7418), .A2(n6993), .ZN(n6776) );
  OR2_X1 U8077 ( .A1(n7479), .A2(n4926), .ZN(n6775) );
  NAND2_X1 U8078 ( .A1(n6776), .A2(n6775), .ZN(n6778) );
  XNOR2_X1 U8079 ( .A(n6778), .B(n6777), .ZN(n6780) );
  NOR2_X1 U8080 ( .A1(n7479), .A2(n6988), .ZN(n6779) );
  AOI21_X1 U8081 ( .B1(n7418), .B2(n6927), .A(n6779), .ZN(n6781) );
  NAND2_X1 U8082 ( .A1(n6780), .A2(n6781), .ZN(n7326) );
  INV_X1 U8083 ( .A(n6780), .ZN(n6783) );
  INV_X1 U8084 ( .A(n6781), .ZN(n6782) );
  NAND2_X1 U8085 ( .A1(n6783), .A2(n6782), .ZN(n7327) );
  NAND2_X1 U8086 ( .A1(n6784), .A2(n7327), .ZN(n7474) );
  NAND2_X1 U8087 ( .A1(n7445), .A2(n6927), .ZN(n6786) );
  OR2_X1 U8088 ( .A1(n7688), .A2(n6988), .ZN(n6785) );
  NAND2_X1 U8089 ( .A1(n6786), .A2(n6785), .ZN(n7475) );
  NAND2_X1 U8090 ( .A1(n7445), .A2(n6993), .ZN(n6788) );
  OR2_X1 U8091 ( .A1(n7688), .A2(n4926), .ZN(n6787) );
  NAND2_X1 U8092 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  XNOR2_X1 U8093 ( .A(n6789), .B(n6930), .ZN(n7476) );
  NAND2_X1 U8094 ( .A1(n7474), .A2(n7475), .ZN(n6790) );
  NAND2_X1 U8095 ( .A1(n7691), .A2(n6759), .ZN(n6793) );
  OR2_X1 U8096 ( .A1(n7610), .A2(n4926), .ZN(n6792) );
  NAND2_X1 U8097 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  XNOR2_X1 U8098 ( .A(n6794), .B(n6930), .ZN(n6795) );
  NAND2_X1 U8099 ( .A1(n7691), .A2(n6927), .ZN(n6798) );
  OR2_X1 U8100 ( .A1(n7610), .A2(n6988), .ZN(n6797) );
  NAND2_X1 U8101 ( .A1(n6798), .A2(n6797), .ZN(n7686) );
  INV_X1 U8102 ( .A(n7686), .ZN(n6799) );
  NAND2_X1 U8103 ( .A1(n7615), .A2(n6993), .ZN(n6803) );
  OR2_X1 U8104 ( .A1(n7601), .A2(n4926), .ZN(n6802) );
  NAND2_X1 U8105 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  XNOR2_X1 U8106 ( .A(n6804), .B(n6930), .ZN(n6806) );
  NOR2_X1 U8107 ( .A1(n7601), .A2(n6988), .ZN(n6805) );
  AOI21_X1 U8108 ( .B1(n7615), .B2(n6927), .A(n6805), .ZN(n6807) );
  XNOR2_X1 U8109 ( .A(n6806), .B(n6807), .ZN(n7790) );
  NAND2_X1 U8110 ( .A1(n7789), .A2(n7790), .ZN(n7788) );
  INV_X1 U8111 ( .A(n6806), .ZN(n6808) );
  NAND2_X1 U8112 ( .A1(n6808), .A2(n6807), .ZN(n6809) );
  NAND2_X1 U8113 ( .A1(n7788), .A2(n6809), .ZN(n6815) );
  INV_X1 U8114 ( .A(n6815), .ZN(n6813) );
  OAI22_X1 U8115 ( .A1(n8005), .A2(n6810), .B1(n8047), .B2(n4926), .ZN(n6811)
         );
  XNOR2_X1 U8116 ( .A(n6811), .B(n6777), .ZN(n6814) );
  INV_X1 U8117 ( .A(n6814), .ZN(n6812) );
  OR2_X1 U8118 ( .A1(n8005), .A2(n4926), .ZN(n6817) );
  NAND2_X1 U8119 ( .A1(n6881), .A2(n9793), .ZN(n6816) );
  NAND2_X1 U8120 ( .A1(n6817), .A2(n6816), .ZN(n7999) );
  NAND2_X1 U8121 ( .A1(n7672), .A2(n6759), .ZN(n6820) );
  OR2_X1 U8122 ( .A1(n6822), .A2(n4926), .ZN(n6819) );
  NAND2_X1 U8123 ( .A1(n6820), .A2(n6819), .ZN(n6821) );
  XNOR2_X1 U8124 ( .A(n6821), .B(n6777), .ZN(n6825) );
  NOR2_X1 U8125 ( .A1(n6822), .A2(n6988), .ZN(n6823) );
  AOI21_X1 U8126 ( .B1(n7672), .B2(n6927), .A(n6823), .ZN(n6824) );
  NAND2_X1 U8127 ( .A1(n6825), .A2(n6824), .ZN(n6827) );
  OR2_X1 U8128 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  AND2_X1 U8129 ( .A1(n6827), .A2(n6826), .ZN(n8042) );
  NAND2_X1 U8130 ( .A1(n8044), .A2(n6827), .ZN(n8119) );
  NAND2_X1 U8131 ( .A1(n8117), .A2(n6759), .ZN(n6829) );
  OR2_X1 U8132 ( .A1(n9517), .A2(n4926), .ZN(n6828) );
  NAND2_X1 U8133 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  XNOR2_X1 U8134 ( .A(n6830), .B(n6930), .ZN(n6832) );
  NOR2_X1 U8135 ( .A1(n9517), .A2(n6988), .ZN(n6831) );
  AOI21_X1 U8136 ( .B1(n8117), .B2(n6927), .A(n6831), .ZN(n6833) );
  XNOR2_X1 U8137 ( .A(n6832), .B(n6833), .ZN(n8120) );
  NAND2_X1 U8138 ( .A1(n8119), .A2(n8120), .ZN(n8118) );
  INV_X1 U8139 ( .A(n6832), .ZN(n6834) );
  NAND2_X1 U8140 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  NAND2_X1 U8141 ( .A1(n8118), .A2(n6835), .ZN(n9513) );
  NAND2_X1 U8142 ( .A1(n10180), .A2(n6759), .ZN(n6837) );
  OR2_X1 U8143 ( .A1(n9427), .A2(n4926), .ZN(n6836) );
  NAND2_X1 U8144 ( .A1(n6837), .A2(n6836), .ZN(n6838) );
  XNOR2_X1 U8145 ( .A(n6838), .B(n6930), .ZN(n6845) );
  NAND2_X1 U8146 ( .A1(n10180), .A2(n6927), .ZN(n6840) );
  OR2_X1 U8147 ( .A1(n9427), .A2(n6988), .ZN(n6839) );
  NAND2_X1 U8148 ( .A1(n6840), .A2(n6839), .ZN(n6846) );
  NAND2_X1 U8149 ( .A1(n6845), .A2(n6846), .ZN(n9514) );
  NAND2_X1 U8150 ( .A1(n9431), .A2(n6759), .ZN(n6842) );
  OR2_X1 U8151 ( .A1(n9771), .A2(n4926), .ZN(n6841) );
  NAND2_X1 U8152 ( .A1(n6842), .A2(n6841), .ZN(n6843) );
  XNOR2_X1 U8153 ( .A(n6843), .B(n6777), .ZN(n9422) );
  NOR2_X1 U8154 ( .A1(n9771), .A2(n6988), .ZN(n6844) );
  AOI21_X1 U8155 ( .B1(n9431), .B2(n6927), .A(n6844), .ZN(n9421) );
  INV_X1 U8156 ( .A(n6845), .ZN(n6848) );
  INV_X1 U8157 ( .A(n6846), .ZN(n6847) );
  AND2_X1 U8158 ( .A1(n6848), .A2(n6847), .ZN(n9419) );
  AOI21_X1 U8159 ( .B1(n9422), .B2(n9421), .A(n9419), .ZN(n6849) );
  INV_X1 U8160 ( .A(n9422), .ZN(n6851) );
  INV_X1 U8161 ( .A(n9421), .ZN(n6850) );
  NAND2_X1 U8162 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  NAND2_X1 U8163 ( .A1(n10171), .A2(n6759), .ZN(n6854) );
  OR2_X1 U8164 ( .A1(n10163), .A2(n4926), .ZN(n6853) );
  NAND2_X1 U8165 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  XNOR2_X1 U8166 ( .A(n6855), .B(n6777), .ZN(n9478) );
  NOR2_X1 U8167 ( .A1(n10163), .A2(n6988), .ZN(n6856) );
  AOI21_X1 U8168 ( .B1(n10171), .B2(n6927), .A(n6856), .ZN(n9477) );
  NOR2_X1 U8169 ( .A1(n9426), .A2(n6988), .ZN(n6857) );
  AOI21_X1 U8170 ( .B1(n8017), .B2(n6927), .A(n6857), .ZN(n9767) );
  NAND2_X1 U8171 ( .A1(n8017), .A2(n6759), .ZN(n6859) );
  OR2_X1 U8172 ( .A1(n9426), .A2(n4926), .ZN(n6858) );
  NAND2_X1 U8173 ( .A1(n6859), .A2(n6858), .ZN(n6860) );
  XNOR2_X1 U8174 ( .A(n6860), .B(n6777), .ZN(n9475) );
  OAI22_X1 U8175 ( .A1(n9478), .A2(n9477), .B1(n9767), .B2(n9475), .ZN(n6866)
         );
  NAND2_X1 U8176 ( .A1(n9475), .A2(n9767), .ZN(n6862) );
  INV_X1 U8177 ( .A(n9477), .ZN(n6861) );
  NAND2_X1 U8178 ( .A1(n6862), .A2(n6861), .ZN(n6864) );
  INV_X1 U8179 ( .A(n6862), .ZN(n6863) );
  AOI22_X1 U8180 ( .A1(n9478), .A2(n6864), .B1(n6863), .B2(n9477), .ZN(n6865)
         );
  NAND2_X1 U8181 ( .A1(n10166), .A2(n6759), .ZN(n6868) );
  NAND2_X1 U8182 ( .A1(n9787), .A2(n6927), .ZN(n6867) );
  NAND2_X1 U8183 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  XNOR2_X1 U8184 ( .A(n6869), .B(n6777), .ZN(n9488) );
  NOR2_X1 U8185 ( .A1(n10156), .A2(n6988), .ZN(n6870) );
  AOI21_X1 U8186 ( .B1(n10166), .B2(n6927), .A(n6870), .ZN(n9487) );
  INV_X1 U8187 ( .A(n9488), .ZN(n6872) );
  INV_X1 U8188 ( .A(n9487), .ZN(n6871) );
  NAND2_X1 U8189 ( .A1(n10159), .A2(n6759), .ZN(n6874) );
  NAND2_X1 U8190 ( .A1(n9786), .A2(n6927), .ZN(n6873) );
  NAND2_X1 U8191 ( .A1(n6874), .A2(n6873), .ZN(n6875) );
  NAND2_X1 U8192 ( .A1(n10159), .A2(n6927), .ZN(n6877) );
  NAND2_X1 U8193 ( .A1(n9786), .A2(n6881), .ZN(n6876) );
  NAND2_X1 U8194 ( .A1(n6877), .A2(n6876), .ZN(n9538) );
  NAND2_X1 U8195 ( .A1(n9539), .A2(n9538), .ZN(n9537) );
  NAND2_X1 U8196 ( .A1(n4937), .A2(n4941), .ZN(n9542) );
  NAND2_X1 U8197 ( .A1(n9537), .A2(n9542), .ZN(n9446) );
  NAND2_X1 U8198 ( .A1(n10153), .A2(n6993), .ZN(n6879) );
  NAND2_X1 U8199 ( .A1(n10088), .A2(n6927), .ZN(n6878) );
  NAND2_X1 U8200 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  XNOR2_X1 U8201 ( .A(n6880), .B(n6930), .ZN(n9443) );
  NAND2_X1 U8202 ( .A1(n10153), .A2(n6927), .ZN(n6883) );
  NAND2_X1 U8203 ( .A1(n10088), .A2(n6881), .ZN(n6882) );
  NAND2_X1 U8204 ( .A1(n6883), .A2(n6882), .ZN(n9444) );
  NAND2_X1 U8205 ( .A1(n10148), .A2(n6993), .ZN(n6885) );
  OR2_X1 U8206 ( .A1(n10139), .A2(n4926), .ZN(n6884) );
  NAND2_X1 U8207 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  XNOR2_X1 U8208 ( .A(n6886), .B(n6777), .ZN(n6889) );
  NOR2_X1 U8209 ( .A1(n10139), .A2(n6988), .ZN(n6887) );
  AOI21_X1 U8210 ( .B1(n10148), .B2(n6927), .A(n6887), .ZN(n6888) );
  NAND2_X1 U8211 ( .A1(n6889), .A2(n6888), .ZN(n9451) );
  OR2_X1 U8212 ( .A1(n6889), .A2(n6888), .ZN(n6890) );
  NAND2_X1 U8213 ( .A1(n9451), .A2(n6890), .ZN(n9506) );
  NAND2_X1 U8214 ( .A1(n10142), .A2(n6993), .ZN(n6893) );
  NAND2_X1 U8215 ( .A1(n9784), .A2(n6927), .ZN(n6892) );
  NAND2_X1 U8216 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  XNOR2_X1 U8217 ( .A(n6894), .B(n6777), .ZN(n6897) );
  NOR2_X1 U8218 ( .A1(n10132), .A2(n6988), .ZN(n6895) );
  AOI21_X1 U8219 ( .B1(n10142), .B2(n6801), .A(n6895), .ZN(n6896) );
  NAND2_X1 U8220 ( .A1(n6897), .A2(n6896), .ZN(n6899) );
  OR2_X1 U8221 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  AND2_X1 U8222 ( .A1(n6899), .A2(n6898), .ZN(n9453) );
  NAND2_X1 U8223 ( .A1(n10135), .A2(n6993), .ZN(n6901) );
  OR2_X1 U8224 ( .A1(n10126), .A2(n4926), .ZN(n6900) );
  NAND2_X1 U8225 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  XNOR2_X1 U8226 ( .A(n6902), .B(n6930), .ZN(n6905) );
  NAND2_X1 U8227 ( .A1(n6904), .A2(n6905), .ZN(n9525) );
  NOR2_X1 U8228 ( .A1(n10126), .A2(n6988), .ZN(n6903) );
  AOI21_X1 U8229 ( .B1(n10135), .B2(n6801), .A(n6903), .ZN(n9524) );
  INV_X1 U8230 ( .A(n6904), .ZN(n6907) );
  INV_X1 U8231 ( .A(n6905), .ZN(n6906) );
  NAND2_X1 U8232 ( .A1(n10013), .A2(n6993), .ZN(n6909) );
  NAND2_X1 U8233 ( .A1(n10027), .A2(n6927), .ZN(n6908) );
  NAND2_X1 U8234 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  XNOR2_X1 U8235 ( .A(n6910), .B(n6777), .ZN(n6913) );
  NOR2_X1 U8236 ( .A1(n9991), .A2(n6988), .ZN(n6911) );
  AOI21_X1 U8237 ( .B1(n10013), .B2(n6801), .A(n6911), .ZN(n6912) );
  NAND2_X1 U8238 ( .A1(n6913), .A2(n6912), .ZN(n9496) );
  OR2_X1 U8239 ( .A1(n6913), .A2(n6912), .ZN(n6914) );
  AND2_X1 U8240 ( .A1(n9496), .A2(n6914), .ZN(n9435) );
  NAND2_X1 U8241 ( .A1(n9995), .A2(n6993), .ZN(n6916) );
  NAND2_X1 U8242 ( .A1(n10005), .A2(n6927), .ZN(n6915) );
  NAND2_X1 U8243 ( .A1(n6916), .A2(n6915), .ZN(n6917) );
  XNOR2_X1 U8244 ( .A(n6917), .B(n6777), .ZN(n6920) );
  NOR2_X1 U8245 ( .A1(n9974), .A2(n6988), .ZN(n6918) );
  AOI21_X1 U8246 ( .B1(n9995), .B2(n6801), .A(n6918), .ZN(n6919) );
  NAND2_X1 U8247 ( .A1(n6920), .A2(n6919), .ZN(n6922) );
  OR2_X1 U8248 ( .A1(n6920), .A2(n6919), .ZN(n6921) );
  NAND2_X1 U8249 ( .A1(n6922), .A2(n6921), .ZN(n9495) );
  NAND2_X1 U8250 ( .A1(n9471), .A2(n6993), .ZN(n6924) );
  NAND2_X1 U8251 ( .A1(n9501), .A2(n6927), .ZN(n6923) );
  NAND2_X1 U8252 ( .A1(n6924), .A2(n6923), .ZN(n6925) );
  XNOR2_X1 U8253 ( .A(n6925), .B(n6930), .ZN(n6933) );
  OAI22_X1 U8254 ( .A1(n5142), .A2(n4926), .B1(n10111), .B2(n6988), .ZN(n6932)
         );
  XNOR2_X1 U8255 ( .A(n6933), .B(n6932), .ZN(n9466) );
  NOR2_X1 U8256 ( .A1(n10103), .A2(n6988), .ZN(n6926) );
  AOI21_X1 U8257 ( .B1(n9962), .B2(n6801), .A(n6926), .ZN(n6941) );
  NAND2_X1 U8258 ( .A1(n9962), .A2(n6993), .ZN(n6929) );
  NAND2_X1 U8259 ( .A1(n9783), .A2(n6927), .ZN(n6928) );
  NAND2_X1 U8260 ( .A1(n6929), .A2(n6928), .ZN(n6931) );
  XNOR2_X1 U8261 ( .A(n6931), .B(n6930), .ZN(n6943) );
  XOR2_X1 U8262 ( .A(n6941), .B(n6943), .Z(n9754) );
  NOR2_X1 U8263 ( .A1(n6933), .A2(n6932), .ZN(n9755) );
  OR2_X2 U8264 ( .A1(n9465), .A2(n6934), .ZN(n9757) );
  NAND2_X1 U8265 ( .A1(n9947), .A2(n6993), .ZN(n6936) );
  OR2_X1 U8266 ( .A1(n9926), .A2(n4926), .ZN(n6935) );
  NAND2_X1 U8267 ( .A1(n6936), .A2(n6935), .ZN(n6937) );
  XNOR2_X1 U8268 ( .A(n6937), .B(n6777), .ZN(n6940) );
  NOR2_X1 U8269 ( .A1(n9926), .A2(n6988), .ZN(n6938) );
  AOI21_X1 U8270 ( .B1(n9947), .B2(n6801), .A(n6938), .ZN(n6939) );
  NAND2_X1 U8271 ( .A1(n6940), .A2(n6939), .ZN(n6998) );
  OAI21_X1 U8272 ( .B1(n6940), .B2(n6939), .A(n6998), .ZN(n6945) );
  INV_X1 U8273 ( .A(n6941), .ZN(n6942) );
  INV_X1 U8274 ( .A(n6944), .ZN(n6946) );
  OR2_X1 U8275 ( .A1(n6948), .A2(n6947), .ZN(n7382) );
  NOR2_X1 U8276 ( .A1(n7382), .A2(n7383), .ZN(n6956) );
  INV_X1 U8277 ( .A(n10362), .ZN(n6949) );
  AND2_X1 U8278 ( .A1(n6956), .A2(n6949), .ZN(n6964) );
  AND2_X1 U8279 ( .A1(n10750), .A2(n8436), .ZN(n6950) );
  INV_X1 U8280 ( .A(n6964), .ZN(n6953) );
  OR2_X1 U8281 ( .A1(n10688), .A2(n6951), .ZN(n6952) );
  OR2_X1 U8282 ( .A1(n6953), .A2(n6952), .ZN(n6955) );
  INV_X1 U8283 ( .A(n6956), .ZN(n6961) );
  NAND2_X1 U8284 ( .A1(n6961), .A2(n10750), .ZN(n6960) );
  NOR2_X1 U8285 ( .A1(n7052), .A2(n6957), .ZN(n6958) );
  AND2_X1 U8286 ( .A1(n6958), .A2(n7384), .ZN(n6959) );
  AOI21_X1 U8287 ( .B1(n6960), .B2(n6959), .A(P1_U3086), .ZN(n6963) );
  AND2_X1 U8288 ( .A1(n8441), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7696) );
  AND2_X1 U8289 ( .A1(n6961), .A2(n7696), .ZN(n6962) );
  INV_X1 U8290 ( .A(n8507), .ZN(n10603) );
  AND2_X1 U8291 ( .A1(n6964), .A2(n10603), .ZN(n6966) );
  OAI22_X1 U8292 ( .A1(n10103), .A2(n9772), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6965), .ZN(n6968) );
  NOR2_X1 U8293 ( .A1(n9938), .A2(n9770), .ZN(n6967) );
  AOI211_X1 U8294 ( .C1(n9943), .C2(n9759), .A(n6968), .B(n6967), .ZN(n6969)
         );
  NAND2_X1 U8295 ( .A1(n7206), .A2(n6972), .ZN(n6973) );
  OAI21_X1 U8296 ( .B1(n7221), .B2(n7282), .A(n7220), .ZN(n6978) );
  NOR2_X1 U8297 ( .A1(n6975), .A2(n8906), .ZN(n6976) );
  NAND2_X1 U8298 ( .A1(n7453), .A2(n7197), .ZN(n7449) );
  NAND2_X1 U8299 ( .A1(n6978), .A2(n7449), .ZN(n6980) );
  NAND2_X1 U8300 ( .A1(n7452), .A2(n7453), .ZN(n6979) );
  NAND2_X1 U8301 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  NAND2_X1 U8302 ( .A1(n6982), .A2(n10791), .ZN(n6986) );
  NOR2_X1 U8303 ( .A1(n10791), .A2(n6983), .ZN(n6984) );
  NAND2_X1 U8304 ( .A1(n6986), .A2(n6985), .ZN(P2_U3488) );
  NAND2_X1 U8305 ( .A1(n6987), .A2(n9768), .ZN(n7007) );
  NAND2_X1 U8306 ( .A1(n9928), .A2(n6801), .ZN(n6990) );
  OR2_X1 U8307 ( .A1(n9938), .A2(n6988), .ZN(n6989) );
  NAND2_X1 U8308 ( .A1(n6990), .A2(n6989), .ZN(n6991) );
  XNOR2_X1 U8309 ( .A(n6991), .B(n6777), .ZN(n6995) );
  NOR2_X1 U8310 ( .A1(n9938), .A2(n4926), .ZN(n6992) );
  AOI21_X1 U8311 ( .B1(n9928), .B2(n6993), .A(n6992), .ZN(n6994) );
  XNOR2_X1 U8312 ( .A(n6995), .B(n6994), .ZN(n7006) );
  AND2_X1 U8313 ( .A1(n7006), .A2(n5504), .ZN(n7003) );
  INV_X1 U8314 ( .A(n9772), .ZN(n9529) );
  NAND2_X1 U8315 ( .A1(n9954), .A2(n9529), .ZN(n6997) );
  AOI22_X1 U8316 ( .A1(n9924), .A2(n9759), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6996) );
  OAI211_X1 U8317 ( .C1(n7243), .C2(n9770), .A(n6997), .B(n6996), .ZN(n7000)
         );
  NOR3_X1 U8318 ( .A1(n7006), .A2(n9541), .A3(n6998), .ZN(n6999) );
  AOI211_X1 U8319 ( .C1(n9928), .C2(n9546), .A(n7000), .B(n6999), .ZN(n7001)
         );
  INV_X1 U8320 ( .A(n7001), .ZN(n7002) );
  OAI21_X1 U8321 ( .B1(n7007), .B2(n7006), .A(n7005), .ZN(P1_U3220) );
  NAND2_X1 U8322 ( .A1(n7198), .A2(n5034), .ZN(n7008) );
  NAND2_X1 U8323 ( .A1(n7008), .A2(n7966), .ZN(n7013) );
  NAND2_X1 U8324 ( .A1(n7009), .A2(n7013), .ZN(n7010) );
  NAND2_X1 U8325 ( .A1(n7010), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U8326 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  MUX2_X1 U8327 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9417), .Z(n7351) );
  XNOR2_X1 U8328 ( .A(n7351), .B(n7350), .ZN(n7012) );
  MUX2_X1 U8329 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n9417), .Z(n10507) );
  INV_X1 U8330 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7023) );
  NOR2_X1 U8331 ( .A1(n10507), .A2(n7023), .ZN(n7188) );
  NOR2_X1 U8332 ( .A1(n7189), .A2(n7188), .ZN(n7187) );
  NAND2_X1 U8333 ( .A1(P2_U3893), .A2(n8585), .ZN(n10536) );
  NOR2_X1 U8334 ( .A1(n4943), .A2(n7012), .ZN(n7349) );
  AOI211_X1 U8335 ( .C1(n7012), .C2(n4943), .A(n10536), .B(n7349), .ZN(n7035)
         );
  NAND2_X1 U8336 ( .A1(n7013), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7019) );
  INV_X2 U8337 ( .A(P2_U3893), .ZN(n8930) );
  MUX2_X1 U8338 ( .A(n7019), .B(n8930), .S(n8912), .Z(n7015) );
  NOR2_X1 U8339 ( .A1(n9008), .A2(n7350), .ZN(n7034) );
  INV_X1 U8340 ( .A(n7966), .ZN(n7016) );
  NOR2_X1 U8341 ( .A1(n7198), .A2(n7016), .ZN(n7017) );
  INV_X1 U8342 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7018) );
  OAI22_X1 U8343 ( .A1(n10563), .A2(n7018), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7260), .ZN(n7033) );
  OR2_X1 U8344 ( .A1(n7019), .A2(n8585), .ZN(n7027) );
  NOR2_X2 U8345 ( .A1(n7027), .A2(n7028), .ZN(n10579) );
  INV_X1 U8346 ( .A(n10579), .ZN(n7031) );
  NAND2_X1 U8347 ( .A1(n7023), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7020) );
  AOI22_X1 U8348 ( .A1(n7192), .A2(n7020), .B1(n6231), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n7181) );
  AND2_X1 U8349 ( .A1(n7181), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7179) );
  AOI21_X1 U8350 ( .B1(n6231), .B2(P2_REG1_REG_0__SCAN_IN), .A(n7179), .ZN(
        n7021) );
  AOI21_X1 U8351 ( .B1(n7022), .B2(n7021), .A(n4948), .ZN(n7030) );
  INV_X1 U8352 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7473) );
  MUX2_X1 U8353 ( .A(n7473), .B(P2_REG2_REG_2__SCAN_IN), .S(n7350), .Z(n7026)
         );
  NAND2_X1 U8354 ( .A1(n7023), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7024) );
  AOI22_X1 U8355 ( .A1(n7192), .A2(n7024), .B1(n6231), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n7178) );
  AND2_X1 U8356 ( .A1(n7178), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7176) );
  AOI21_X1 U8357 ( .B1(n7026), .B2(n7025), .A(n7336), .ZN(n7029) );
  INV_X1 U8358 ( .A(n7027), .ZN(n10509) );
  NAND2_X1 U8359 ( .A1(n10509), .A2(n7028), .ZN(n9064) );
  OAI22_X1 U8360 ( .A1(n7031), .A2(n7030), .B1(n7029), .B2(n9064), .ZN(n7032)
         );
  OR4_X1 U8361 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(P2_U3184)
         );
  OAI222_X1 U8362 ( .A1(P1_U3086), .A2(n7114), .B1(n7238), .B2(n7040), .C1(
        n7037), .C2(n7593), .ZN(P1_U3353) );
  AOI22_X1 U8363 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9833), .B1(n10241), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n7038) );
  OAI21_X1 U8364 ( .B1(n7041), .B2(n7238), .A(n7038), .ZN(P1_U3352) );
  NOR2_X1 U8365 ( .A1(n5701), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9409) );
  OAI222_X1 U8366 ( .A1(n4925), .A2(n7040), .B1(n7350), .B2(P2_U3151), .C1(
        n7039), .C2(n9415), .ZN(P2_U3293) );
  OAI222_X1 U8367 ( .A1(n9415), .A2(n7042), .B1(n7352), .B2(P2_U3151), .C1(
        n4925), .C2(n7041), .ZN(P2_U3292) );
  AOI22_X1 U8368 ( .A1(n10594), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10241), .ZN(n7043) );
  OAI21_X1 U8369 ( .B1(n7044), .B2(n7238), .A(n7043), .ZN(P1_U3351) );
  OAI222_X1 U8370 ( .A1(n4925), .A2(n8520), .B1(n5110), .B2(P2_U3151), .C1(
        n5582), .C2(n9415), .ZN(P2_U3294) );
  OAI222_X1 U8371 ( .A1(n4925), .A2(n7046), .B1(n9415), .B2(n5302), .C1(
        P2_U3151), .C2(n10529), .ZN(P2_U3290) );
  OAI222_X1 U8372 ( .A1(n9415), .A2(n5596), .B1(n7699), .B2(P2_U3151), .C1(
        n4925), .C2(n7044), .ZN(P2_U3291) );
  INV_X1 U8373 ( .A(n10378), .ZN(n7121) );
  INV_X1 U8374 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7045) );
  OAI222_X1 U8375 ( .A1(P1_U3086), .A2(n7121), .B1(n7238), .B2(n7046), .C1(
        n7045), .C2(n7593), .ZN(P1_U3350) );
  AOI22_X1 U8376 ( .A1(n10393), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10241), .ZN(n7047) );
  OAI21_X1 U8377 ( .B1(n7048), .B2(n7238), .A(n7047), .ZN(P1_U3349) );
  INV_X1 U8378 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7064) );
  OAI222_X1 U8379 ( .A1(n4925), .A2(n7048), .B1(n9415), .B2(n7064), .C1(
        P2_U3151), .C2(n7707), .ZN(P2_U3289) );
  INV_X1 U8380 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7049) );
  OAI222_X1 U8381 ( .A1(n4925), .A2(n7055), .B1(n7821), .B2(P2_U3151), .C1(
        n7049), .C2(n9415), .ZN(P2_U3288) );
  OR2_X1 U8382 ( .A1(n7052), .A2(n8436), .ZN(n7051) );
  AND2_X1 U8383 ( .A1(n7051), .A2(n7050), .ZN(n7112) );
  INV_X1 U8384 ( .A(n7112), .ZN(n7053) );
  NAND2_X1 U8385 ( .A1(n7052), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8509) );
  NAND2_X1 U8386 ( .A1(n10362), .A2(n8509), .ZN(n7111) );
  NOR2_X1 U8387 ( .A1(n10585), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8388 ( .A(n10406), .ZN(n7106) );
  INV_X1 U8389 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7054) );
  OAI222_X1 U8390 ( .A1(P1_U3086), .A2(n7106), .B1(n7238), .B2(n7055), .C1(
        n7054), .C2(n7593), .ZN(P1_U3348) );
  NAND2_X1 U8391 ( .A1(P1_U3973), .A2(n7056), .ZN(n7057) );
  OAI21_X1 U8392 ( .B1(P1_U3973), .B2(n5302), .A(n7057), .ZN(P1_U3559) );
  INV_X1 U8393 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7062) );
  INV_X1 U8394 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U8395 ( .A1(n4927), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7059) );
  NAND2_X1 U8396 ( .A1(n5757), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7058) );
  OAI211_X1 U8397 ( .C1(n7060), .C2(n10097), .A(n7059), .B(n7058), .ZN(n8433)
         );
  NAND2_X1 U8398 ( .A1(P1_U3973), .A2(n8433), .ZN(n7061) );
  OAI21_X1 U8399 ( .B1(P1_U3973), .B2(n7062), .A(n7061), .ZN(P1_U3585) );
  NAND2_X1 U8400 ( .A1(n7296), .A2(P1_U3973), .ZN(n7063) );
  OAI21_X1 U8401 ( .B1(P1_U3973), .B2(n7064), .A(n7063), .ZN(P1_U3560) );
  INV_X1 U8402 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U8403 ( .A1(n8051), .A2(P1_U3973), .ZN(n7065) );
  OAI21_X1 U8404 ( .B1(n7146), .B2(P1_U3973), .A(n7065), .ZN(P1_U3566) );
  INV_X1 U8405 ( .A(n7123), .ZN(n10420) );
  INV_X1 U8406 ( .A(n7066), .ZN(n7067) );
  INV_X1 U8407 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7094) );
  OAI222_X1 U8408 ( .A1(n10420), .A2(P1_U3086), .B1(n7238), .B2(n7067), .C1(
        n7593), .C2(n7094), .ZN(P1_U3347) );
  INV_X1 U8409 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7068) );
  OAI222_X1 U8410 ( .A1(n9415), .A2(n7068), .B1(n4925), .B2(n7067), .C1(
        P2_U3151), .C2(n7884), .ZN(P2_U3287) );
  AND2_X1 U8411 ( .A1(n7080), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8412 ( .A1(n7080), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8413 ( .A1(n7080), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8414 ( .A1(n7080), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8415 ( .A1(n7080), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8416 ( .A1(n7080), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8417 ( .A1(n7080), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8418 ( .A1(n7080), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8419 ( .A1(n7080), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8420 ( .A1(n7080), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8421 ( .A1(n7080), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8422 ( .A1(n7080), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8423 ( .A1(n7080), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AOI22_X1 U8424 ( .A1(n10502), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10241), .ZN(n7070) );
  OAI21_X1 U8425 ( .B1(n7072), .B2(n7238), .A(n7070), .ZN(P1_U3345) );
  INV_X1 U8426 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7071) );
  OAI222_X1 U8427 ( .A1(n4925), .A2(n7072), .B1(n7987), .B2(P2_U3151), .C1(
        n7071), .C2(n9415), .ZN(P2_U3285) );
  INV_X1 U8428 ( .A(n7073), .ZN(n7076) );
  INV_X1 U8429 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7074) );
  OAI222_X1 U8430 ( .A1(n4925), .A2(n7076), .B1(n5389), .B2(P2_U3151), .C1(
        n7074), .C2(n9415), .ZN(P2_U3286) );
  INV_X1 U8431 ( .A(n7271), .ZN(n7130) );
  INV_X1 U8432 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7075) );
  OAI222_X1 U8433 ( .A1(P1_U3086), .A2(n7130), .B1(n7238), .B2(n7076), .C1(
        n7075), .C2(n7593), .ZN(P1_U3346) );
  INV_X1 U8434 ( .A(n10688), .ZN(n10602) );
  NOR2_X1 U8435 ( .A1(n10634), .A2(n10703), .ZN(n10610) );
  INV_X1 U8436 ( .A(n10186), .ZN(n7077) );
  NAND2_X1 U8437 ( .A1(n6739), .A2(n10606), .ZN(n8450) );
  AND2_X1 U8438 ( .A1(n7077), .A2(n8450), .ZN(n10604) );
  AOI21_X1 U8439 ( .B1(n10698), .B2(n10183), .A(n10604), .ZN(n7078) );
  AOI211_X1 U8440 ( .C1(n10602), .C2(n10193), .A(n10610), .B(n7078), .ZN(n7162) );
  NAND2_X1 U8441 ( .A1(n10756), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7079) );
  OAI21_X1 U8442 ( .B1(n7162), .B2(n10756), .A(n7079), .ZN(P1_U3522) );
  INV_X1 U8443 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7083) );
  INV_X1 U8444 ( .A(n7081), .ZN(n7082) );
  AOI22_X1 U8445 ( .A1(n7080), .A2(n7083), .B1(n7086), .B2(n7082), .ZN(
        P2_U3377) );
  INV_X1 U8446 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7087) );
  INV_X1 U8447 ( .A(n7084), .ZN(n7085) );
  AOI22_X1 U8448 ( .A1(n7080), .A2(n7087), .B1(n7086), .B2(n7085), .ZN(
        P2_U3376) );
  NOR2_X1 U8449 ( .A1(n9759), .A2(P1_U3086), .ZN(n7159) );
  INV_X1 U8450 ( .A(n9770), .ZN(n9762) );
  AOI22_X1 U8451 ( .A1(n9762), .A2(n6724), .B1(n9546), .B2(n10193), .ZN(n7092)
         );
  OR2_X1 U8452 ( .A1(n7089), .A2(n7088), .ZN(n9812) );
  NAND3_X1 U8453 ( .A1(n9812), .A2(n9768), .A3(n7090), .ZN(n7091) );
  OAI211_X1 U8454 ( .C1(n7159), .C2(n10605), .A(n7092), .B(n7091), .ZN(
        P1_U3232) );
  NAND2_X1 U8455 ( .A1(n7941), .A2(P2_U3893), .ZN(n7093) );
  OAI21_X1 U8456 ( .B1(P2_U3893), .B2(n7094), .A(n7093), .ZN(P2_U3499) );
  AND2_X1 U8457 ( .A1(n7080), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8458 ( .A1(n7080), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8459 ( .A1(n7080), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8460 ( .A1(n7080), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8461 ( .A1(n7080), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8462 ( .A1(n7080), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8463 ( .A1(n7080), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8464 ( .A1(n7080), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8465 ( .A1(n7080), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8466 ( .A1(n7080), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8467 ( .A1(n7080), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8468 ( .A1(n7080), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8469 ( .A1(n7080), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8470 ( .A1(n7080), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8471 ( .A1(n7080), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8472 ( .A1(n7080), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8473 ( .A1(n7080), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  INV_X1 U8474 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U8475 ( .A1(n8163), .A2(P2_U3893), .ZN(n7095) );
  OAI21_X1 U8476 ( .B1(P2_U3893), .B2(n7135), .A(n7095), .ZN(P2_U3502) );
  XNOR2_X1 U8477 ( .A(n7114), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9823) );
  XNOR2_X1 U8478 ( .A(n9805), .B(n7096), .ZN(n9802) );
  AND2_X1 U8479 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9801) );
  NAND2_X1 U8480 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  NAND2_X1 U8481 ( .A1(n9805), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U8482 ( .A1(n9800), .A2(n7097), .ZN(n9822) );
  NAND2_X1 U8483 ( .A1(n9823), .A2(n9822), .ZN(n9821) );
  INV_X1 U8484 ( .A(n7114), .ZN(n9820) );
  NAND2_X1 U8485 ( .A1(n9820), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7098) );
  NAND2_X1 U8486 ( .A1(n9821), .A2(n7098), .ZN(n9838) );
  XNOR2_X1 U8487 ( .A(n9833), .B(n7099), .ZN(n9839) );
  NAND2_X1 U8488 ( .A1(n9838), .A2(n9839), .ZN(n9837) );
  NAND2_X1 U8489 ( .A1(n9833), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U8490 ( .A1(n9837), .A2(n7100), .ZN(n10592) );
  XNOR2_X1 U8491 ( .A(n10594), .B(n7101), .ZN(n10593) );
  NAND2_X1 U8492 ( .A1(n10592), .A2(n10593), .ZN(n10590) );
  NAND2_X1 U8493 ( .A1(n10594), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U8494 ( .A1(n10590), .A2(n7102), .ZN(n10372) );
  MUX2_X1 U8495 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5788), .S(n10378), .Z(n10373) );
  AND2_X1 U8496 ( .A1(n10372), .A2(n10373), .ZN(n10370) );
  AOI21_X1 U8497 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10378), .A(n10370), .ZN(
        n10390) );
  MUX2_X1 U8498 ( .A(n7103), .B(P1_REG1_REG_6__SCAN_IN), .S(n10393), .Z(n10389) );
  NOR2_X1 U8499 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  AOI21_X1 U8500 ( .B1(n10393), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10388), .ZN(
        n10403) );
  MUX2_X1 U8501 ( .A(n7105), .B(P1_REG1_REG_7__SCAN_IN), .S(n10406), .Z(n10402) );
  NOR2_X1 U8502 ( .A1(n10403), .A2(n10402), .ZN(n10401) );
  INV_X1 U8503 ( .A(n10401), .ZN(n7104) );
  OAI21_X1 U8504 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n10412) );
  INV_X1 U8505 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7107) );
  MUX2_X1 U8506 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7107), .S(n7123), .Z(n10411)
         );
  NAND2_X1 U8507 ( .A1(n10412), .A2(n10411), .ZN(n10410) );
  INV_X1 U8508 ( .A(n10410), .ZN(n7108) );
  AOI21_X1 U8509 ( .B1(n7123), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7108), .ZN(
        n7110) );
  AOI22_X1 U8510 ( .A1(n7271), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n5849), .B2(
        n7130), .ZN(n7109) );
  NAND2_X1 U8511 ( .A1(n7109), .A2(n7110), .ZN(n7270) );
  OAI21_X1 U8512 ( .B1(n7110), .B2(n7109), .A(n7270), .ZN(n7132) );
  NAND2_X1 U8513 ( .A1(n7112), .A2(n7111), .ZN(n10369) );
  OR2_X1 U8514 ( .A1(n10369), .A2(n10364), .ZN(n10492) );
  AND2_X1 U8515 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7794) );
  AOI21_X1 U8516 ( .B1(n10585), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7794), .ZN(
        n7129) );
  NAND2_X1 U8517 ( .A1(n10245), .A2(n10364), .ZN(n8506) );
  XNOR2_X1 U8518 ( .A(n7123), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n10413) );
  MUX2_X1 U8519 ( .A(n7113), .B(P1_REG2_REG_6__SCAN_IN), .S(n10393), .Z(n10386) );
  XNOR2_X1 U8520 ( .A(n7114), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9826) );
  INV_X1 U8521 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7115) );
  XNOR2_X1 U8522 ( .A(n9805), .B(n7115), .ZN(n9804) );
  AND2_X1 U8523 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9814) );
  NAND2_X1 U8524 ( .A1(n9804), .A2(n9814), .ZN(n9803) );
  NAND2_X1 U8525 ( .A1(n9805), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U8526 ( .A1(n9803), .A2(n7116), .ZN(n9825) );
  NAND2_X1 U8527 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  NAND2_X1 U8528 ( .A1(n9820), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7117) );
  NAND2_X1 U8529 ( .A1(n9824), .A2(n7117), .ZN(n9835) );
  XNOR2_X1 U8530 ( .A(n9833), .B(n7118), .ZN(n9836) );
  NAND2_X1 U8531 ( .A1(n9835), .A2(n9836), .ZN(n9834) );
  NAND2_X1 U8532 ( .A1(n9833), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7119) );
  NAND2_X1 U8533 ( .A1(n9834), .A2(n7119), .ZN(n10588) );
  XNOR2_X1 U8534 ( .A(n10594), .B(n10706), .ZN(n10589) );
  NAND2_X1 U8535 ( .A1(n10588), .A2(n10589), .ZN(n10586) );
  NAND2_X1 U8536 ( .A1(n10594), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7120) );
  AND2_X1 U8537 ( .A1(n10586), .A2(n7120), .ZN(n10376) );
  AOI22_X1 U8538 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7121), .B1(n10378), .B2(
        n7390), .ZN(n10375) );
  NAND2_X1 U8539 ( .A1(n10406), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7122) );
  OAI21_X1 U8540 ( .B1(n10406), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7122), .ZN(
        n10399) );
  NOR2_X1 U8541 ( .A1(n10400), .A2(n10399), .ZN(n10398) );
  NOR2_X1 U8542 ( .A1(n7271), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7124) );
  AOI21_X1 U8543 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7271), .A(n7124), .ZN(
        n7125) );
  NAND2_X1 U8544 ( .A1(n7125), .A2(n7126), .ZN(n7262) );
  OAI21_X1 U8545 ( .B1(n7126), .B2(n7125), .A(n7262), .ZN(n7127) );
  NAND2_X1 U8546 ( .A1(n10587), .A2(n7127), .ZN(n7128) );
  OAI211_X1 U8547 ( .C1(n10451), .C2(n7130), .A(n7129), .B(n7128), .ZN(n7131)
         );
  AOI21_X1 U8548 ( .B1(n7132), .B2(n10591), .A(n7131), .ZN(n7133) );
  INV_X1 U8549 ( .A(n7133), .ZN(P1_U3252) );
  INV_X1 U8550 ( .A(n7273), .ZN(n10434) );
  INV_X1 U8551 ( .A(n7134), .ZN(n7136) );
  OAI222_X1 U8552 ( .A1(n10434), .A2(P1_U3086), .B1(n7238), .B2(n7136), .C1(
        n7593), .C2(n7135), .ZN(P1_U3344) );
  INV_X1 U8553 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7137) );
  OAI222_X1 U8554 ( .A1(n9415), .A2(n7137), .B1(n4925), .B2(n7136), .C1(
        P2_U3151), .C2(n5391), .ZN(P2_U3284) );
  INV_X1 U8555 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U8556 ( .A1(n8195), .A2(P2_U3893), .ZN(n7138) );
  OAI21_X1 U8557 ( .B1(P2_U3893), .B2(n7161), .A(n7138), .ZN(P2_U3503) );
  OAI21_X1 U8558 ( .B1(n7139), .B2(n7141), .A(n7140), .ZN(n7142) );
  NAND2_X1 U8559 ( .A1(n7142), .A2(n9768), .ZN(n7145) );
  OAI22_X1 U8560 ( .A1(n9772), .A2(n10634), .B1(n9779), .B2(n10628), .ZN(n7143) );
  AOI21_X1 U8561 ( .B1(n9762), .B2(n9798), .A(n7143), .ZN(n7144) );
  OAI211_X1 U8562 ( .C1(n7159), .C2(n9817), .A(n7145), .B(n7144), .ZN(P1_U3237) );
  INV_X1 U8563 ( .A(n8939), .ZN(n8931) );
  OAI222_X1 U8564 ( .A1(n4925), .A2(n7160), .B1(n9415), .B2(n7146), .C1(
        P2_U3151), .C2(n8931), .ZN(P2_U3283) );
  INV_X1 U8565 ( .A(n7149), .ZN(n7153) );
  XOR2_X1 U8566 ( .A(n7147), .B(n6750), .Z(n7150) );
  OAI21_X1 U8567 ( .B1(n7150), .B2(n7149), .A(n7148), .ZN(n7151) );
  OAI21_X1 U8568 ( .B1(n7153), .B2(n7152), .A(n7151), .ZN(n7154) );
  NAND2_X1 U8569 ( .A1(n7154), .A2(n9768), .ZN(n7157) );
  INV_X1 U8570 ( .A(n6739), .ZN(n10188) );
  OAI22_X1 U8571 ( .A1(n9772), .A2(n10188), .B1(n9779), .B2(n10616), .ZN(n7155) );
  AOI21_X1 U8572 ( .B1(n9762), .B2(n5746), .A(n7155), .ZN(n7156) );
  OAI211_X1 U8573 ( .C1(n7159), .C2(n7158), .A(n7157), .B(n7156), .ZN(P1_U3222) );
  INV_X1 U8574 ( .A(n9855), .ZN(n7277) );
  OAI222_X1 U8575 ( .A1(n7277), .A2(P1_U3086), .B1(n7593), .B2(n7161), .C1(
        n7160), .C2(n7238), .ZN(P1_U3343) );
  INV_X1 U8576 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7164) );
  OR2_X1 U8577 ( .A1(n7162), .A2(n10758), .ZN(n7163) );
  OAI21_X1 U8578 ( .B1(n10761), .B2(n7164), .A(n7163), .ZN(P1_U3453) );
  NAND2_X1 U8579 ( .A1(n10027), .A2(P1_U3973), .ZN(n7165) );
  OAI21_X1 U8580 ( .B1(P1_U3973), .B2(n5667), .A(n7165), .ZN(P1_U3577) );
  OAI21_X1 U8581 ( .B1(n7168), .B2(n7167), .A(n7166), .ZN(n7173) );
  OAI22_X1 U8582 ( .A1(n10653), .A2(n9772), .B1(n9770), .B2(n10654), .ZN(n7172) );
  NAND2_X1 U8583 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9830) );
  INV_X1 U8584 ( .A(n9830), .ZN(n7169) );
  AOI21_X1 U8585 ( .B1(n9546), .B2(n10662), .A(n7169), .ZN(n7170) );
  OAI21_X1 U8586 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n9774), .A(n7170), .ZN(
        n7171) );
  AOI211_X1 U8587 ( .C1(n7173), .C2(n9768), .A(n7172), .B(n7171), .ZN(n7174)
         );
  INV_X1 U8588 ( .A(n7174), .ZN(P1_U3218) );
  INV_X1 U8589 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7175) );
  OAI222_X1 U8590 ( .A1(n4925), .A2(n7195), .B1(n8968), .B2(P2_U3151), .C1(
        n7175), .C2(n9415), .ZN(P2_U3282) );
  INV_X1 U8591 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7186) );
  INV_X1 U8592 ( .A(n7176), .ZN(n7177) );
  OAI21_X1 U8593 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n7178), .A(n7177), .ZN(
        n7183) );
  INV_X1 U8594 ( .A(n7179), .ZN(n7180) );
  OAI21_X1 U8595 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n7181), .A(n7180), .ZN(
        n7182) );
  AOI22_X1 U8596 ( .A1(n10578), .A2(n7183), .B1(n10579), .B2(n7182), .ZN(n7185) );
  NAND2_X1 U8597 ( .A1(P2_U3151), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7184) );
  OAI211_X1 U8598 ( .C1(n7186), .C2(n10563), .A(n7185), .B(n7184), .ZN(n7191)
         );
  AOI211_X1 U8599 ( .C1(n7189), .C2(n7188), .A(n10536), .B(n7187), .ZN(n7190)
         );
  AOI211_X1 U8600 ( .C1(n10566), .C2(n7192), .A(n7191), .B(n7190), .ZN(n7193)
         );
  INV_X1 U8601 ( .A(n7193), .ZN(P2_U3183) );
  INV_X1 U8602 ( .A(n10487), .ZN(n9852) );
  INV_X1 U8603 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7194) );
  OAI222_X1 U8604 ( .A1(P1_U3086), .A2(n9852), .B1(n7238), .B2(n7195), .C1(
        n7194), .C2(n7593), .ZN(P1_U3342) );
  NAND2_X1 U8605 ( .A1(n7211), .A2(n7196), .ZN(n7201) );
  AND3_X1 U8606 ( .A1(n7198), .A2(n7966), .A3(n7197), .ZN(n7200) );
  INV_X1 U8607 ( .A(n7204), .ZN(n7199) );
  NAND2_X1 U8608 ( .A1(n7216), .A2(n7199), .ZN(n7207) );
  NAND3_X1 U8609 ( .A1(n7201), .A2(n7200), .A3(n7207), .ZN(n7203) );
  INV_X1 U8610 ( .A(n7215), .ZN(n8913) );
  AND2_X1 U8611 ( .A1(n7216), .A2(n8913), .ZN(n7202) );
  AOI21_X2 U8612 ( .B1(n7203), .B2(P2_STATE_REG_SCAN_IN), .A(n7202), .ZN(n8654) );
  NOR2_X1 U8613 ( .A1(n8715), .A2(P2_U3151), .ZN(n7261) );
  AND2_X1 U8614 ( .A1(n8775), .A2(n7223), .ZN(n8745) );
  INV_X1 U8615 ( .A(n8745), .ZN(n7218) );
  NAND2_X1 U8616 ( .A1(n5034), .A2(n10785), .ZN(n7205) );
  OAI21_X1 U8617 ( .B1(n7211), .B2(n7205), .A(n7204), .ZN(n7209) );
  AND2_X1 U8618 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  OR2_X1 U8619 ( .A1(n7211), .A2(n7210), .ZN(n7214) );
  NOR2_X1 U8620 ( .A1(n7216), .A2(n7215), .ZN(n7232) );
  NAND2_X1 U8621 ( .A1(n7232), .A2(n7230), .ZN(n8712) );
  OAI22_X1 U8622 ( .A1(n8719), .A2(n7284), .B1(n7226), .B2(n8712), .ZN(n7217)
         );
  AOI21_X1 U8623 ( .B1(n7218), .B2(n8706), .A(n7217), .ZN(n7219) );
  OAI21_X1 U8624 ( .B1(n7261), .B2(n10512), .A(n7219), .ZN(P2_U3172) );
  NAND2_X1 U8625 ( .A1(n7221), .A2(n8906), .ZN(n7222) );
  OAI21_X1 U8626 ( .B1(n7509), .B2(n5013), .A(n7223), .ZN(n7228) );
  INV_X1 U8627 ( .A(n7225), .ZN(n7224) );
  NAND2_X1 U8628 ( .A1(n7226), .A2(n7225), .ZN(n7252) );
  NAND2_X1 U8629 ( .A1(n7229), .A2(n8706), .ZN(n7236) );
  INV_X1 U8630 ( .A(n7230), .ZN(n7231) );
  NAND2_X1 U8631 ( .A1(n8685), .A2(n6617), .ZN(n7233) );
  OAI21_X1 U8632 ( .B1(n8515), .B2(n8700), .A(n7233), .ZN(n7234) );
  AOI21_X1 U8633 ( .B1(n7362), .B2(n8689), .A(n7234), .ZN(n7235) );
  OAI211_X1 U8634 ( .C1(n7261), .C2(n7490), .A(n7236), .B(n7235), .ZN(P2_U3162) );
  AOI22_X1 U8635 ( .A1(n10439), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10241), .ZN(n7237) );
  OAI21_X1 U8636 ( .B1(n7241), .B2(n7238), .A(n7237), .ZN(P1_U3341) );
  NAND2_X1 U8637 ( .A1(n9501), .A2(P1_U3973), .ZN(n7239) );
  OAI21_X1 U8638 ( .B1(P1_U3973), .B2(n8147), .A(n7239), .ZN(P1_U3579) );
  INV_X1 U8639 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7240) );
  OAI222_X1 U8640 ( .A1(n4925), .A2(n7241), .B1(n8965), .B2(P2_U3151), .C1(
        n7240), .C2(n9415), .ZN(P2_U3281) );
  NAND2_X1 U8641 ( .A1(n9799), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7242) );
  OAI21_X1 U8642 ( .B1(n7243), .B2(n9799), .A(n7242), .ZN(P1_U3583) );
  INV_X1 U8643 ( .A(n7245), .ZN(n7246) );
  AOI211_X1 U8644 ( .C1(n7247), .C2(n7244), .A(n9541), .B(n7246), .ZN(n7251)
         );
  OAI22_X1 U8645 ( .A1(n10700), .A2(n9772), .B1(n9770), .B2(n10702), .ZN(n7250) );
  AND2_X1 U8646 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10584) );
  AOI21_X1 U8647 ( .B1(n9546), .B2(n10691), .A(n10584), .ZN(n7248) );
  OAI21_X1 U8648 ( .B1(n9774), .B2(n10719), .A(n7248), .ZN(n7249) );
  OR3_X1 U8649 ( .A1(n7251), .A2(n7250), .A3(n7249), .ZN(P1_U3230) );
  XNOR2_X1 U8650 ( .A(n7467), .B(n5013), .ZN(n7300) );
  XNOR2_X1 U8651 ( .A(n7300), .B(n6617), .ZN(n7255) );
  NAND2_X1 U8652 ( .A1(n7253), .A2(n7252), .ZN(n7254) );
  NAND2_X1 U8653 ( .A1(n7254), .A2(n7255), .ZN(n7302) );
  OAI21_X1 U8654 ( .B1(n7255), .B2(n7254), .A(n7302), .ZN(n7256) );
  NAND2_X1 U8655 ( .A1(n7256), .A2(n8706), .ZN(n7259) );
  OAI22_X1 U8656 ( .A1(n7513), .A2(n8712), .B1(n7226), .B2(n8700), .ZN(n7257)
         );
  AOI21_X1 U8657 ( .B1(n7467), .B2(n8689), .A(n7257), .ZN(n7258) );
  OAI211_X1 U8658 ( .C1(n7261), .C2(n7260), .A(n7259), .B(n7258), .ZN(P2_U3177) );
  AOI22_X1 U8659 ( .A1(n9855), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n5909), .B2(
        n7277), .ZN(n7266) );
  OAI21_X1 U8660 ( .B1(n7271), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7262), .ZN(
        n10499) );
  NAND2_X1 U8661 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10502), .ZN(n7263) );
  OAI21_X1 U8662 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10502), .A(n7263), .ZN(
        n10498) );
  NOR2_X1 U8663 ( .A1(n10499), .A2(n10498), .ZN(n10497) );
  AOI21_X1 U8664 ( .B1(n10502), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10497), .ZN(
        n10429) );
  NAND2_X1 U8665 ( .A1(n7273), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U8666 ( .B1(n7273), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7264), .ZN(
        n10430) );
  NOR2_X1 U8667 ( .A1(n10429), .A2(n10430), .ZN(n10428) );
  OAI21_X1 U8668 ( .B1(n7266), .B2(n7265), .A(n9854), .ZN(n7267) );
  INV_X1 U8669 ( .A(n7267), .ZN(n7281) );
  AOI22_X1 U8670 ( .A1(n9855), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7268), .B2(
        n7277), .ZN(n7275) );
  INV_X1 U8671 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7269) );
  MUX2_X1 U8672 ( .A(n7269), .B(P1_REG1_REG_10__SCAN_IN), .S(n10502), .Z(
        n10494) );
  OAI21_X1 U8673 ( .B1(n7271), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7270), .ZN(
        n10495) );
  NOR2_X1 U8674 ( .A1(n10494), .A2(n10495), .ZN(n10493) );
  AOI21_X1 U8675 ( .B1(n10502), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10493), .ZN(
        n10425) );
  MUX2_X1 U8676 ( .A(n7272), .B(P1_REG1_REG_11__SCAN_IN), .S(n7273), .Z(n10426) );
  NOR2_X1 U8677 ( .A1(n10425), .A2(n10426), .ZN(n10424) );
  AOI21_X1 U8678 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n7273), .A(n10424), .ZN(
        n7274) );
  NAND2_X1 U8679 ( .A1(n7275), .A2(n7274), .ZN(n9844) );
  OAI21_X1 U8680 ( .B1(n7275), .B2(n7274), .A(n9844), .ZN(n7279) );
  AND2_X1 U8681 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8124) );
  AOI21_X1 U8682 ( .B1(n10585), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8124), .ZN(
        n7276) );
  OAI21_X1 U8683 ( .B1(n7277), .B2(n10451), .A(n7276), .ZN(n7278) );
  AOI21_X1 U8684 ( .B1(n7279), .B2(n10591), .A(n7278), .ZN(n7280) );
  OAI21_X1 U8685 ( .B1(n7281), .B2(n10496), .A(n7280), .ZN(P1_U3255) );
  INV_X1 U8686 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7286) );
  NOR2_X1 U8687 ( .A1(n10775), .A2(n9340), .ZN(n7283) );
  OAI222_X1 U8688 ( .A1(n7284), .A2(n10785), .B1(n8745), .B2(n7283), .C1(n9316), .C2(n7226), .ZN(n9363) );
  NAND2_X1 U8689 ( .A1(n9363), .A2(n6696), .ZN(n7285) );
  OAI21_X1 U8690 ( .B1(n7286), .B2(n6696), .A(n7285), .ZN(P2_U3390) );
  INV_X1 U8691 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7287) );
  OAI222_X1 U8692 ( .A1(n4925), .A2(n7289), .B1(n8991), .B2(P2_U3151), .C1(
        n7287), .C2(n9415), .ZN(P2_U3280) );
  INV_X1 U8693 ( .A(n10464), .ZN(n9857) );
  INV_X1 U8694 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7288) );
  OAI222_X1 U8695 ( .A1(P1_U3086), .A2(n9857), .B1(n7238), .B2(n7289), .C1(
        n7288), .C2(n7593), .ZN(P1_U3340) );
  NAND2_X1 U8696 ( .A1(n7291), .A2(n7290), .ZN(n7293) );
  XNOR2_X1 U8697 ( .A(n7293), .B(n7292), .ZN(n7299) );
  NAND2_X1 U8698 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10382) );
  INV_X1 U8699 ( .A(n10382), .ZN(n7295) );
  OAI22_X1 U8700 ( .A1(n9774), .A2(n7389), .B1(n9772), .B2(n10654), .ZN(n7294)
         );
  AOI211_X1 U8701 ( .C1(n9762), .C2(n7296), .A(n7295), .B(n7294), .ZN(n7298)
         );
  NAND2_X1 U8702 ( .A1(n9546), .A2(n7393), .ZN(n7297) );
  OAI211_X1 U8703 ( .C1(n7299), .C2(n9541), .A(n7298), .B(n7297), .ZN(P1_U3227) );
  NAND2_X1 U8704 ( .A1(n7580), .A2(n7300), .ZN(n7301) );
  NAND2_X1 U8705 ( .A1(n7302), .A2(n7301), .ZN(n7303) );
  XNOR2_X1 U8706 ( .A(n7585), .B(n8542), .ZN(n7425) );
  XNOR2_X1 U8707 ( .A(n7425), .B(n8929), .ZN(n7304) );
  AOI21_X1 U8708 ( .B1(n7303), .B2(n7304), .A(n8691), .ZN(n7307) );
  INV_X1 U8709 ( .A(n7303), .ZN(n7306) );
  NAND2_X1 U8710 ( .A1(n7306), .A2(n7305), .ZN(n7427) );
  NAND2_X1 U8711 ( .A1(n7307), .A2(n7427), .ZN(n7310) );
  INV_X1 U8712 ( .A(n7579), .ZN(n8928) );
  NOR2_X1 U8713 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9550), .ZN(n10524) );
  OAI22_X1 U8714 ( .A1(n8719), .A2(n7587), .B1(n7580), .B2(n8700), .ZN(n7308)
         );
  AOI211_X1 U8715 ( .C1(n8685), .C2(n8928), .A(n10524), .B(n7308), .ZN(n7309)
         );
  OAI211_X1 U8716 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8654), .A(n7310), .B(
        n7309), .ZN(P2_U3158) );
  INV_X1 U8717 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7312) );
  INV_X1 U8718 ( .A(n7311), .ZN(n7314) );
  INV_X1 U8719 ( .A(n9012), .ZN(n9000) );
  OAI222_X1 U8720 ( .A1(n9415), .A2(n7312), .B1(n4925), .B2(n7314), .C1(
        P2_U3151), .C2(n9000), .ZN(P2_U3279) );
  INV_X1 U8721 ( .A(n9874), .ZN(n9851) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7313) );
  OAI222_X1 U8723 ( .A1(n9851), .A2(P1_U3086), .B1(n7238), .B2(n7314), .C1(
        n7313), .C2(n7593), .ZN(P1_U3339) );
  XNOR2_X1 U8724 ( .A(n7315), .B(n8237), .ZN(n7397) );
  OAI211_X1 U8725 ( .C1(n7316), .C2(n7321), .A(n10192), .B(n7370), .ZN(n7395)
         );
  OAI21_X1 U8726 ( .B1(n10654), .B2(n10701), .A(n7395), .ZN(n7319) );
  XOR2_X1 U8727 ( .A(n8237), .B(n7317), .Z(n7318) );
  OAI22_X1 U8728 ( .A1(n7318), .A2(n10698), .B1(n7479), .B2(n10703), .ZN(n7381) );
  AOI211_X1 U8729 ( .C1(n7397), .C2(n10754), .A(n7319), .B(n7381), .ZN(n7325)
         );
  INV_X1 U8730 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7320) );
  OAI22_X1 U8731 ( .A1(n10220), .A2(n7321), .B1(n10761), .B2(n7320), .ZN(n7322) );
  INV_X1 U8732 ( .A(n7322), .ZN(n7323) );
  OAI21_X1 U8733 ( .B1(n7325), .B2(n10758), .A(n7323), .ZN(P1_U3468) );
  INV_X1 U8734 ( .A(n10131), .ZN(n7865) );
  AOI22_X1 U8735 ( .A1(n7865), .A2(n7393), .B1(n10756), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7324) );
  OAI21_X1 U8736 ( .B1(n7325), .B2(n10756), .A(n7324), .ZN(P1_U3527) );
  NAND2_X1 U8737 ( .A1(n7327), .A2(n7326), .ZN(n7329) );
  XOR2_X1 U8738 ( .A(n7329), .B(n7328), .Z(n7334) );
  NOR2_X1 U8739 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7330), .ZN(n10395) );
  OAI22_X1 U8740 ( .A1(n9774), .A2(n7415), .B1(n9772), .B2(n10702), .ZN(n7331)
         );
  AOI211_X1 U8741 ( .C1(n9762), .C2(n9796), .A(n10395), .B(n7331), .ZN(n7333)
         );
  NAND2_X1 U8742 ( .A1(n9546), .A2(n7418), .ZN(n7332) );
  OAI211_X1 U8743 ( .C1(n7334), .C2(n9541), .A(n7333), .B(n7332), .ZN(P1_U3239) );
  INV_X1 U8744 ( .A(n7699), .ZN(n7709) );
  INV_X1 U8745 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7348) );
  MUX2_X1 U8746 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7335), .S(n7699), .Z(n7339)
         );
  AOI21_X1 U8747 ( .B1(n7350), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7336), .ZN(
        n7337) );
  INV_X1 U8748 ( .A(n7352), .ZN(n10516) );
  XNOR2_X1 U8749 ( .A(n7337), .B(n7352), .ZN(n10514) );
  NAND2_X1 U8750 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n10514), .ZN(n10513) );
  OAI21_X1 U8751 ( .B1(n7339), .B2(n7338), .A(n7708), .ZN(n7345) );
  MUX2_X1 U8752 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7340), .S(n7699), .Z(n7343)
         );
  AOI21_X1 U8753 ( .B1(n7350), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4948), .ZN(
        n7341) );
  XNOR2_X1 U8754 ( .A(n7341), .B(n7352), .ZN(n10521) );
  NAND2_X1 U8755 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n10521), .ZN(n10520) );
  OAI21_X1 U8756 ( .B1(n7341), .B2(n10516), .A(n10520), .ZN(n7342) );
  OAI21_X1 U8757 ( .B1(n7343), .B2(n7342), .A(n7703), .ZN(n7344) );
  AOI22_X1 U8758 ( .A1(n10578), .A2(n7345), .B1(n10579), .B2(n7344), .ZN(n7347) );
  NOR2_X1 U8759 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9620), .ZN(n7434) );
  INV_X1 U8760 ( .A(n7434), .ZN(n7346) );
  OAI211_X1 U8761 ( .C1(n7348), .C2(n10563), .A(n7347), .B(n7346), .ZN(n7357)
         );
  MUX2_X1 U8762 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9417), .Z(n7700) );
  XNOR2_X1 U8763 ( .A(n7700), .B(n7699), .ZN(n7355) );
  MUX2_X1 U8764 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9417), .Z(n7353) );
  XOR2_X1 U8765 ( .A(n7352), .B(n7353), .Z(n10518) );
  NAND2_X1 U8766 ( .A1(n10519), .A2(n10518), .ZN(n10517) );
  OAI21_X1 U8767 ( .B1(n7353), .B2(n7352), .A(n10517), .ZN(n7354) );
  AOI211_X1 U8768 ( .C1(n7355), .C2(n7354), .A(n10536), .B(n7698), .ZN(n7356)
         );
  AOI211_X1 U8769 ( .C1(n10566), .C2(n7709), .A(n7357), .B(n7356), .ZN(n7358)
         );
  INV_X1 U8770 ( .A(n7358), .ZN(P2_U3186) );
  XNOR2_X1 U8771 ( .A(n8741), .B(n7359), .ZN(n7493) );
  OAI22_X1 U8772 ( .A1(n7580), .A2(n9316), .B1(n8515), .B2(n9314), .ZN(n7361)
         );
  AOI21_X1 U8773 ( .B1(n7223), .B2(n8741), .A(n7456), .ZN(n7496) );
  NOR2_X1 U8774 ( .A1(n7496), .A2(n10787), .ZN(n7360) );
  AOI211_X1 U8775 ( .C1(n9340), .C2(n7493), .A(n7361), .B(n7360), .ZN(n7367)
         );
  AOI22_X1 U8776 ( .A1(n9331), .A2(n7362), .B1(n10782), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7363) );
  OAI21_X1 U8777 ( .B1(n7367), .B2(n10782), .A(n7363), .ZN(P2_U3460) );
  INV_X1 U8778 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7364) );
  OAI22_X1 U8779 ( .A1(n5314), .A2(n9403), .B1(n6696), .B2(n7364), .ZN(n7365)
         );
  INV_X1 U8780 ( .A(n7365), .ZN(n7366) );
  OAI21_X1 U8781 ( .B1(n7367), .B2(n10792), .A(n7366), .ZN(P2_U3393) );
  OAI21_X1 U8782 ( .B1(n7369), .B2(n8239), .A(n7368), .ZN(n7422) );
  INV_X1 U8783 ( .A(n7418), .ZN(n7376) );
  INV_X1 U8784 ( .A(n7370), .ZN(n7372) );
  INV_X1 U8785 ( .A(n7406), .ZN(n7371) );
  OAI211_X1 U8786 ( .C1(n7376), .C2(n7372), .A(n7371), .B(n10192), .ZN(n7420)
         );
  OAI21_X1 U8787 ( .B1(n10702), .B2(n10701), .A(n7420), .ZN(n7374) );
  XNOR2_X1 U8788 ( .A(n7402), .B(n8239), .ZN(n7373) );
  OAI22_X1 U8789 ( .A1(n7373), .A2(n10698), .B1(n7688), .B2(n10703), .ZN(n7414) );
  AOI211_X1 U8790 ( .C1(n10754), .C2(n7422), .A(n7374), .B(n7414), .ZN(n7380)
         );
  INV_X1 U8791 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7375) );
  OAI22_X1 U8792 ( .A1(n10220), .A2(n7376), .B1(n10761), .B2(n7375), .ZN(n7377) );
  INV_X1 U8793 ( .A(n7377), .ZN(n7378) );
  OAI21_X1 U8794 ( .B1(n7380), .B2(n10758), .A(n7378), .ZN(P1_U3471) );
  AOI22_X1 U8795 ( .A1(n7865), .A2(n7418), .B1(n10756), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7379) );
  OAI21_X1 U8796 ( .B1(n7380), .B2(n10756), .A(n7379), .ZN(P1_U3528) );
  INV_X1 U8797 ( .A(n7381), .ZN(n7399) );
  NOR2_X1 U8798 ( .A1(n10362), .A2(n7382), .ZN(n7386) );
  AND2_X1 U8799 ( .A1(n7384), .A2(n7383), .ZN(n7385) );
  NAND2_X1 U8800 ( .A1(n7386), .A2(n7385), .ZN(n7388) );
  INV_X2 U8801 ( .A(n10707), .ZN(n10714) );
  NAND2_X1 U8802 ( .A1(n10655), .A2(n8027), .ZN(n10713) );
  OR2_X1 U8803 ( .A1(n7388), .A2(n10607), .ZN(n9915) );
  NAND2_X1 U8804 ( .A1(n10709), .A2(n10663), .ZN(n10670) );
  OAI22_X1 U8805 ( .A1(n10707), .A2(n7390), .B1(n7389), .B2(n10718), .ZN(n7392) );
  INV_X1 U8806 ( .A(n10701), .ZN(n8133) );
  NAND2_X1 U8807 ( .A1(n10707), .A2(n8133), .ZN(n10085) );
  NOR2_X1 U8808 ( .A1(n10085), .A2(n10654), .ZN(n7391) );
  AOI211_X1 U8809 ( .C1(n10081), .C2(n7393), .A(n7392), .B(n7391), .ZN(n7394)
         );
  OAI21_X1 U8810 ( .B1(n10010), .B2(n7395), .A(n7394), .ZN(n7396) );
  AOI21_X1 U8811 ( .B1(n7397), .B2(n10016), .A(n7396), .ZN(n7398) );
  OAI21_X1 U8812 ( .B1(n7399), .B2(n10714), .A(n7398), .ZN(P1_U3288) );
  INV_X1 U8813 ( .A(n8239), .ZN(n7401) );
  AOI21_X1 U8814 ( .B1(n7402), .B2(n7401), .A(n7400), .ZN(n7553) );
  XNOR2_X1 U8815 ( .A(n7553), .B(n8242), .ZN(n7403) );
  OAI22_X1 U8816 ( .A1(n7403), .A2(n10698), .B1(n7610), .B2(n10703), .ZN(n7439) );
  INV_X1 U8817 ( .A(n7439), .ZN(n7413) );
  OAI21_X1 U8818 ( .B1(n7405), .B2(n7552), .A(n7404), .ZN(n7441) );
  OAI211_X1 U8819 ( .C1(n7485), .C2(n7406), .A(n10192), .B(n7596), .ZN(n7438)
         );
  OAI22_X1 U8820 ( .A1(n10707), .A2(n7407), .B1(n7480), .B2(n10718), .ZN(n7409) );
  NOR2_X1 U8821 ( .A1(n10085), .A2(n7479), .ZN(n7408) );
  AOI211_X1 U8822 ( .C1(n10081), .C2(n7445), .A(n7409), .B(n7408), .ZN(n7410)
         );
  OAI21_X1 U8823 ( .B1(n7438), .B2(n10010), .A(n7410), .ZN(n7411) );
  AOI21_X1 U8824 ( .B1(n7441), .B2(n10016), .A(n7411), .ZN(n7412) );
  OAI21_X1 U8825 ( .B1(n7413), .B2(n10714), .A(n7412), .ZN(P1_U3286) );
  INV_X1 U8826 ( .A(n7414), .ZN(n7424) );
  OAI22_X1 U8827 ( .A1(n10707), .A2(n7113), .B1(n7415), .B2(n10718), .ZN(n7417) );
  NOR2_X1 U8828 ( .A1(n10085), .A2(n10702), .ZN(n7416) );
  AOI211_X1 U8829 ( .C1(n10081), .C2(n7418), .A(n7417), .B(n7416), .ZN(n7419)
         );
  OAI21_X1 U8830 ( .B1(n7420), .B2(n10010), .A(n7419), .ZN(n7421) );
  AOI21_X1 U8831 ( .B1(n7422), .B2(n10016), .A(n7421), .ZN(n7423) );
  OAI21_X1 U8832 ( .B1(n7424), .B2(n10714), .A(n7423), .ZN(P1_U3287) );
  NAND2_X1 U8833 ( .A1(n7425), .A2(n8929), .ZN(n7426) );
  XNOR2_X1 U8834 ( .A(n7428), .B(n5013), .ZN(n7429) );
  INV_X1 U8835 ( .A(n7429), .ZN(n7430) );
  NAND2_X1 U8836 ( .A1(n7430), .A2(n8928), .ZN(n7431) );
  AND2_X1 U8837 ( .A1(n7543), .A2(n7431), .ZN(n7522) );
  NAND2_X1 U8838 ( .A1(n7524), .A2(n7522), .ZN(n7542) );
  OAI21_X1 U8839 ( .B1(n7524), .B2(n7522), .A(n7542), .ZN(n7432) );
  NAND2_X1 U8840 ( .A1(n7432), .A2(n8706), .ZN(n7436) );
  OAI22_X1 U8841 ( .A1(n8719), .A2(n10680), .B1(n7535), .B2(n8712), .ZN(n7433)
         );
  AOI211_X1 U8842 ( .C1(n8710), .C2(n8929), .A(n7434), .B(n7433), .ZN(n7435)
         );
  OAI211_X1 U8843 ( .C1(n7516), .C2(n8654), .A(n7436), .B(n7435), .ZN(P2_U3170) );
  AOI22_X1 U8844 ( .A1(n10477), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10241), .ZN(n7437) );
  OAI21_X1 U8845 ( .B1(n7539), .B2(n7238), .A(n7437), .ZN(P1_U3337) );
  OAI21_X1 U8846 ( .B1(n7479), .B2(n10701), .A(n7438), .ZN(n7440) );
  AOI211_X1 U8847 ( .C1(n10754), .C2(n7441), .A(n7440), .B(n7439), .ZN(n7447)
         );
  INV_X1 U8848 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7442) );
  OAI22_X1 U8849 ( .A1(n7485), .A2(n10220), .B1(n10761), .B2(n7442), .ZN(n7443) );
  INV_X1 U8850 ( .A(n7443), .ZN(n7444) );
  OAI21_X1 U8851 ( .B1(n7447), .B2(n10758), .A(n7444), .ZN(P1_U3474) );
  AOI22_X1 U8852 ( .A1(n7865), .A2(n7445), .B1(n10756), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7446) );
  OAI21_X1 U8853 ( .B1(n7447), .B2(n10756), .A(n7446), .ZN(P1_U3529) );
  INV_X1 U8854 ( .A(n7448), .ZN(n7455) );
  INV_X1 U8855 ( .A(n7449), .ZN(n7450) );
  NAND2_X1 U8856 ( .A1(n7220), .A2(n7450), .ZN(n7451) );
  OAI21_X1 U8857 ( .B1(n7453), .B2(n7452), .A(n7451), .ZN(n7454) );
  NAND2_X1 U8858 ( .A1(n7455), .A2(n7454), .ZN(n7505) );
  INV_X1 U8859 ( .A(n7456), .ZN(n7457) );
  NAND2_X1 U8860 ( .A1(n7457), .A2(n7460), .ZN(n7459) );
  MUX2_X1 U8861 ( .A(n7460), .B(n7459), .S(n7458), .Z(n7462) );
  NAND2_X1 U8862 ( .A1(n7462), .A2(n7461), .ZN(n10646) );
  INV_X1 U8863 ( .A(n10646), .ZN(n7470) );
  OR2_X1 U8864 ( .A1(n8771), .A2(n7468), .ZN(n7778) );
  XNOR2_X1 U8865 ( .A(n7463), .B(n8772), .ZN(n7465) );
  AOI22_X1 U8866 ( .A1(n5475), .A2(n9334), .B1(n9335), .B2(n8929), .ZN(n7464)
         );
  OAI21_X1 U8867 ( .B1(n7465), .B2(n9323), .A(n7464), .ZN(n7466) );
  AOI21_X1 U8868 ( .B1(n10646), .B2(n8155), .A(n7466), .ZN(n10643) );
  AND2_X1 U8869 ( .A1(n7467), .A2(n10777), .ZN(n10645) );
  AOI22_X1 U8870 ( .A1(n10645), .A2(n7468), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9188), .ZN(n7469) );
  OAI211_X1 U8871 ( .C1(n7470), .C2(n7778), .A(n10643), .B(n7469), .ZN(n7471)
         );
  NAND2_X1 U8872 ( .A1(n7471), .A2(n9269), .ZN(n7472) );
  OAI21_X1 U8873 ( .B1(n7473), .B2(n9269), .A(n7472), .ZN(P2_U3231) );
  XNOR2_X1 U8874 ( .A(n7476), .B(n7475), .ZN(n7477) );
  XNOR2_X1 U8875 ( .A(n7474), .B(n7477), .ZN(n7478) );
  NAND2_X1 U8876 ( .A1(n7478), .A2(n9768), .ZN(n7484) );
  NAND2_X1 U8877 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10407) );
  INV_X1 U8878 ( .A(n10407), .ZN(n7482) );
  OAI22_X1 U8879 ( .A1(n9774), .A2(n7480), .B1(n9772), .B2(n7479), .ZN(n7481)
         );
  AOI211_X1 U8880 ( .C1(n9762), .C2(n9795), .A(n7482), .B(n7481), .ZN(n7483)
         );
  OAI211_X1 U8881 ( .C1(n7485), .C2(n9779), .A(n7484), .B(n7483), .ZN(P1_U3213) );
  AND2_X1 U8882 ( .A1(n7486), .A2(n7778), .ZN(n7487) );
  INV_X1 U8883 ( .A(n7505), .ZN(n7489) );
  INV_X1 U8884 ( .A(n8174), .ZN(n7488) );
  OAI22_X1 U8885 ( .A1(n9265), .A2(n5314), .B1(n7490), .B2(n9267), .ZN(n7492)
         );
  OR2_X1 U8886 ( .A1(n9194), .A2(n9314), .ZN(n9175) );
  OR2_X1 U8887 ( .A1(n9194), .A2(n9316), .ZN(n9093) );
  OAI22_X1 U8888 ( .A1(n8515), .A2(n9175), .B1(n9093), .B2(n7580), .ZN(n7491)
         );
  AOI211_X1 U8889 ( .C1(P2_REG2_REG_1__SCAN_IN), .C2(n9189), .A(n7492), .B(
        n7491), .ZN(n7495) );
  OR2_X1 U8890 ( .A1(n9194), .A2(n9323), .ZN(n9155) );
  NAND2_X1 U8891 ( .A1(n7493), .A2(n9170), .ZN(n7494) );
  OAI211_X1 U8892 ( .C1(n7496), .C2(n9274), .A(n7495), .B(n7494), .ZN(P2_U3232) );
  XNOR2_X1 U8893 ( .A(n7497), .B(n8742), .ZN(n7581) );
  OAI21_X1 U8894 ( .B1(n7499), .B2(n8742), .A(n7498), .ZN(n7584) );
  NAND2_X1 U8895 ( .A1(n7584), .A2(n9192), .ZN(n7503) );
  OAI22_X1 U8896 ( .A1(n9265), .A2(n7587), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9267), .ZN(n7501) );
  OAI22_X1 U8897 ( .A1(n7579), .A2(n9093), .B1(n9175), .B2(n7580), .ZN(n7500)
         );
  AOI211_X1 U8898 ( .C1(P2_REG2_REG_3__SCAN_IN), .C2(n9189), .A(n7501), .B(
        n7500), .ZN(n7502) );
  OAI211_X1 U8899 ( .C1(n7581), .C2(n9155), .A(n7503), .B(n7502), .ZN(P2_U3230) );
  NAND2_X1 U8900 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n9188), .ZN(n7504) );
  OAI21_X1 U8901 ( .B1(n9269), .B2(n6218), .A(n7504), .ZN(n7508) );
  NOR4_X1 U8902 ( .A1(n8745), .A2(n7506), .A3(n10777), .A4(n7505), .ZN(n7507)
         );
  AOI211_X1 U8903 ( .C1(n9253), .C2(n7509), .A(n7508), .B(n7507), .ZN(n7510)
         );
  OAI21_X1 U8904 ( .B1(n7226), .B2(n9093), .A(n7510), .ZN(P2_U3233) );
  XOR2_X1 U8905 ( .A(n7511), .B(n8779), .Z(n7512) );
  OAI222_X1 U8906 ( .A1(n9314), .A2(n7513), .B1(n9316), .B2(n7535), .C1(n7512), 
        .C2(n9323), .ZN(n10681) );
  INV_X1 U8907 ( .A(n10681), .ZN(n7520) );
  OAI21_X1 U8908 ( .B1(n7515), .B2(n8779), .A(n7514), .ZN(n10683) );
  NOR2_X1 U8909 ( .A1(n9269), .A2(n7335), .ZN(n7518) );
  OAI22_X1 U8910 ( .A1(n9265), .A2(n10680), .B1(n7516), .B2(n9267), .ZN(n7517)
         );
  AOI211_X1 U8911 ( .C1(n10683), .C2(n9192), .A(n7518), .B(n7517), .ZN(n7519)
         );
  OAI21_X1 U8912 ( .B1(n7520), .B2(n9194), .A(n7519), .ZN(P2_U3229) );
  XNOR2_X1 U8913 ( .A(n7521), .B(n5013), .ZN(n7525) );
  XNOR2_X1 U8914 ( .A(n7525), .B(n8927), .ZN(n7544) );
  AND2_X1 U8915 ( .A1(n7522), .A2(n7544), .ZN(n7523) );
  NAND2_X1 U8916 ( .A1(n7535), .A2(n7525), .ZN(n7527) );
  NAND2_X1 U8917 ( .A1(n7544), .A2(n7526), .ZN(n7546) );
  AND2_X1 U8918 ( .A1(n7527), .A2(n7546), .ZN(n7531) );
  NAND2_X1 U8919 ( .A1(n7532), .A2(n7531), .ZN(n7528) );
  XNOR2_X1 U8920 ( .A(n7775), .B(n8542), .ZN(n7632) );
  XNOR2_X1 U8921 ( .A(n7632), .B(n8926), .ZN(n7529) );
  AOI21_X1 U8922 ( .B1(n7528), .B2(n7529), .A(n8691), .ZN(n7533) );
  INV_X1 U8923 ( .A(n7529), .ZN(n7530) );
  NAND2_X1 U8924 ( .A1(n7532), .A2(n4935), .ZN(n7634) );
  NAND2_X1 U8925 ( .A1(n7533), .A2(n7634), .ZN(n7538) );
  INV_X1 U8926 ( .A(n7761), .ZN(n8925) );
  INV_X1 U8927 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7534) );
  NOR2_X1 U8928 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7534), .ZN(n10558) );
  OAI22_X1 U8929 ( .A1(n8719), .A2(n10727), .B1(n7535), .B2(n8700), .ZN(n7536)
         );
  AOI211_X1 U8930 ( .C1(n8685), .C2(n8925), .A(n10558), .B(n7536), .ZN(n7537)
         );
  OAI211_X1 U8931 ( .C1(n7773), .C2(n8654), .A(n7538), .B(n7537), .ZN(P2_U3179) );
  INV_X1 U8932 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7540) );
  INV_X1 U8933 ( .A(n9052), .ZN(n9044) );
  OAI222_X1 U8934 ( .A1(n9415), .A2(n7540), .B1(n9044), .B2(P2_U3151), .C1(
        n4925), .C2(n7539), .ZN(P2_U3277) );
  NAND2_X1 U8935 ( .A1(n8930), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7541) );
  OAI21_X1 U8936 ( .B1(n9279), .B2(n8930), .A(n7541), .ZN(P2_U3520) );
  INV_X1 U8937 ( .A(n7542), .ZN(n7545) );
  NOR3_X1 U8938 ( .A1(n7545), .A2(n7526), .A3(n7544), .ZN(n7548) );
  NAND2_X1 U8939 ( .A1(n7532), .A2(n7546), .ZN(n7547) );
  OAI21_X1 U8940 ( .B1(n7548), .B2(n7547), .A(n8706), .ZN(n7551) );
  NOR2_X1 U8941 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6262), .ZN(n10540) );
  OAI22_X1 U8942 ( .A1(n8719), .A2(n10720), .B1(n7579), .B2(n8700), .ZN(n7549)
         );
  AOI211_X1 U8943 ( .C1(n8685), .C2(n8926), .A(n10540), .B(n7549), .ZN(n7550)
         );
  OAI211_X1 U8944 ( .C1(n7780), .C2(n8654), .A(n7551), .B(n7550), .ZN(P2_U3167) );
  OAI21_X1 U8945 ( .B1(n7553), .B2(n7552), .A(n8319), .ZN(n7600) );
  OAI21_X1 U8946 ( .B1(n7600), .B2(n8327), .A(n7554), .ZN(n7555) );
  XOR2_X1 U8947 ( .A(n8329), .B(n7555), .Z(n7556) );
  NOR2_X1 U8948 ( .A1(n7556), .A2(n10698), .ZN(n7611) );
  INV_X1 U8949 ( .A(n7611), .ZN(n7566) );
  OAI21_X1 U8950 ( .B1(n7558), .B2(n8329), .A(n7557), .ZN(n7613) );
  AOI211_X1 U8951 ( .C1(n7615), .C2(n7597), .A(n10660), .B(n7655), .ZN(n7559)
         );
  AOI21_X1 U8952 ( .B1(n10089), .B2(n9793), .A(n7559), .ZN(n7609) );
  NOR2_X1 U8953 ( .A1(n10085), .A2(n7610), .ZN(n7562) );
  OAI22_X1 U8954 ( .A1(n10707), .A2(n7560), .B1(n7792), .B2(n10718), .ZN(n7561) );
  AOI211_X1 U8955 ( .C1(n7615), .C2(n10081), .A(n7562), .B(n7561), .ZN(n7563)
         );
  OAI21_X1 U8956 ( .B1(n7609), .B2(n10010), .A(n7563), .ZN(n7564) );
  AOI21_X1 U8957 ( .B1(n10016), .B2(n7613), .A(n7564), .ZN(n7565) );
  OAI21_X1 U8958 ( .B1(n7566), .B2(n10714), .A(n7565), .ZN(P1_U3284) );
  INV_X1 U8959 ( .A(n7567), .ZN(n7591) );
  INV_X1 U8960 ( .A(n9028), .ZN(n9023) );
  INV_X1 U8961 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7568) );
  OAI222_X1 U8962 ( .A1(n4925), .A2(n7591), .B1(n9023), .B2(P2_U3151), .C1(
        n7568), .C2(n9415), .ZN(P2_U3278) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7578) );
  INV_X1 U8964 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U8965 ( .A1(n6248), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7571) );
  INV_X1 U8966 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7569) );
  OR2_X1 U8967 ( .A1(n6261), .A2(n7569), .ZN(n7570) );
  OAI211_X1 U8968 ( .C1(n7573), .C2(n7572), .A(n7571), .B(n7570), .ZN(n7574)
         );
  INV_X1 U8969 ( .A(n7574), .ZN(n7575) );
  NAND2_X1 U8970 ( .A1(n7576), .A2(n7575), .ZN(n9066) );
  NAND2_X1 U8971 ( .A1(n9066), .A2(P2_U3893), .ZN(n7577) );
  OAI21_X1 U8972 ( .B1(P2_U3893), .B2(n7578), .A(n7577), .ZN(P2_U3522) );
  OAI22_X1 U8973 ( .A1(n7580), .A2(n9314), .B1(n7579), .B2(n9316), .ZN(n7583)
         );
  NOR2_X1 U8974 ( .A1(n7581), .A2(n9323), .ZN(n7582) );
  AOI211_X1 U8975 ( .C1(n10775), .C2(n7584), .A(n7583), .B(n7582), .ZN(n7590)
         );
  AOI22_X1 U8976 ( .A1(n9331), .A2(n7585), .B1(n10782), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7586) );
  OAI21_X1 U8977 ( .B1(n7590), .B2(n10782), .A(n7586), .ZN(P2_U3462) );
  OAI22_X1 U8978 ( .A1(n7587), .A2(n9403), .B1(n6696), .B2(n6237), .ZN(n7588)
         );
  INV_X1 U8979 ( .A(n7588), .ZN(n7589) );
  OAI21_X1 U8980 ( .B1(n7590), .B2(n10792), .A(n7589), .ZN(P2_U3399) );
  INV_X1 U8981 ( .A(n9890), .ZN(n9879) );
  INV_X1 U8982 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7592) );
  OAI222_X1 U8983 ( .A1(n9879), .A2(P1_U3086), .B1(n7593), .B2(n7592), .C1(
        n7591), .C2(n7238), .ZN(P1_U3338) );
  OAI21_X1 U8984 ( .B1(n7595), .B2(n7599), .A(n7594), .ZN(n7629) );
  INV_X1 U8985 ( .A(n7691), .ZN(n7604) );
  INV_X1 U8986 ( .A(n7596), .ZN(n7598) );
  OAI211_X1 U8987 ( .C1(n7604), .C2(n7598), .A(n10192), .B(n7597), .ZN(n7627)
         );
  OAI21_X1 U8988 ( .B1(n7688), .B2(n10701), .A(n7627), .ZN(n7603) );
  XNOR2_X1 U8989 ( .A(n7600), .B(n7599), .ZN(n7602) );
  OAI22_X1 U8990 ( .A1(n7602), .A2(n10698), .B1(n7601), .B2(n10703), .ZN(n7622) );
  AOI211_X1 U8991 ( .C1(n10754), .C2(n7629), .A(n7603), .B(n7622), .ZN(n7608)
         );
  OAI22_X1 U8992 ( .A1(n7604), .A2(n10220), .B1(n10761), .B2(n5837), .ZN(n7605) );
  INV_X1 U8993 ( .A(n7605), .ZN(n7606) );
  OAI21_X1 U8994 ( .B1(n7608), .B2(n10758), .A(n7606), .ZN(P1_U3477) );
  AOI22_X1 U8995 ( .A1(n7691), .A2(n7865), .B1(n10756), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7607) );
  OAI21_X1 U8996 ( .B1(n7608), .B2(n10756), .A(n7607), .ZN(P1_U3530) );
  OAI21_X1 U8997 ( .B1(n7610), .B2(n10701), .A(n7609), .ZN(n7612) );
  AOI211_X1 U8998 ( .C1(n10754), .C2(n7613), .A(n7612), .B(n7611), .ZN(n7619)
         );
  AOI22_X1 U8999 ( .A1(n7615), .A2(n7865), .B1(n10756), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7614) );
  OAI21_X1 U9000 ( .B1(n7619), .B2(n10756), .A(n7614), .ZN(P1_U3531) );
  INV_X1 U9001 ( .A(n7615), .ZN(n7797) );
  INV_X1 U9002 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7616) );
  OAI22_X1 U9003 ( .A1(n7797), .A2(n10220), .B1(n10761), .B2(n7616), .ZN(n7617) );
  INV_X1 U9004 ( .A(n7617), .ZN(n7618) );
  OAI21_X1 U9005 ( .B1(n7619), .B2(n10758), .A(n7618), .ZN(P1_U3480) );
  INV_X1 U9006 ( .A(n7620), .ZN(n7646) );
  AOI22_X1 U9007 ( .A1(n9886), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10241), .ZN(n7621) );
  OAI21_X1 U9008 ( .B1(n7646), .B2(n7238), .A(n7621), .ZN(P1_U3336) );
  INV_X1 U9009 ( .A(n7622), .ZN(n7631) );
  INV_X1 U9010 ( .A(n7689), .ZN(n7623) );
  INV_X1 U9011 ( .A(n10718), .ZN(n10638) );
  AOI22_X1 U9012 ( .A1(n10714), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7623), .B2(
        n10638), .ZN(n7624) );
  OAI21_X1 U9013 ( .B1(n7688), .B2(n10085), .A(n7624), .ZN(n7625) );
  AOI21_X1 U9014 ( .B1(n7691), .B2(n10081), .A(n7625), .ZN(n7626) );
  OAI21_X1 U9015 ( .B1(n7627), .B2(n10010), .A(n7626), .ZN(n7628) );
  AOI21_X1 U9016 ( .B1(n7629), .B2(n10016), .A(n7628), .ZN(n7630) );
  OAI21_X1 U9017 ( .B1(n7631), .B2(n10714), .A(n7630), .ZN(P1_U3285) );
  NAND2_X1 U9018 ( .A1(n7632), .A2(n8926), .ZN(n7633) );
  XNOR2_X1 U9019 ( .A(n7912), .B(n8574), .ZN(n7635) );
  NAND2_X1 U9020 ( .A1(n7635), .A2(n7761), .ZN(n7728) );
  INV_X1 U9021 ( .A(n7635), .ZN(n7636) );
  NAND2_X1 U9022 ( .A1(n7636), .A2(n8925), .ZN(n7637) );
  AND2_X1 U9023 ( .A1(n7728), .A2(n7637), .ZN(n7724) );
  NAND2_X1 U9024 ( .A1(n7727), .A2(n7724), .ZN(n7730) );
  OAI21_X1 U9025 ( .B1(n7727), .B2(n7724), .A(n7730), .ZN(n7643) );
  OR2_X1 U9026 ( .A1(n8654), .A2(n7839), .ZN(n7641) );
  NOR2_X1 U9027 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6294), .ZN(n7714) );
  AOI21_X1 U9028 ( .B1(n8710), .B2(n8926), .A(n7714), .ZN(n7640) );
  NAND2_X1 U9029 ( .A1(n8689), .A2(n7912), .ZN(n7639) );
  NAND2_X1 U9030 ( .A1(n8685), .A2(n7941), .ZN(n7638) );
  NAND4_X1 U9031 ( .A1(n7641), .A2(n7640), .A3(n7639), .A4(n7638), .ZN(n7642)
         );
  AOI21_X1 U9032 ( .B1(n7643), .B2(n8706), .A(n7642), .ZN(n7644) );
  INV_X1 U9033 ( .A(n7644), .ZN(P2_U3153) );
  INV_X1 U9034 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7647) );
  OAI222_X1 U9035 ( .A1(n9415), .A2(n7647), .B1(n4925), .B2(n7646), .C1(
        P2_U3151), .C2(n7645), .ZN(P2_U3276) );
  OAI21_X1 U9036 ( .B1(n7649), .B2(n8245), .A(n7648), .ZN(n7650) );
  INV_X1 U9037 ( .A(n7650), .ZN(n7679) );
  OAI21_X1 U9038 ( .B1(n7653), .B2(n7652), .A(n7651), .ZN(n7654) );
  AOI222_X1 U9039 ( .A1(n10659), .A2(n7654), .B1(n9792), .B2(n10089), .C1(
        n9794), .C2(n8133), .ZN(n7678) );
  INV_X1 U9040 ( .A(n7678), .ZN(n7661) );
  OAI211_X1 U9041 ( .C1(n8005), .C2(n7655), .A(n10192), .B(n7668), .ZN(n7677)
         );
  OAI22_X1 U9042 ( .A1(n10707), .A2(n7656), .B1(n8001), .B2(n10718), .ZN(n7657) );
  AOI21_X1 U9043 ( .B1(n7658), .B2(n10081), .A(n7657), .ZN(n7659) );
  OAI21_X1 U9044 ( .B1(n7677), .B2(n10010), .A(n7659), .ZN(n7660) );
  AOI21_X1 U9045 ( .B1(n7661), .B2(n10707), .A(n7660), .ZN(n7662) );
  OAI21_X1 U9046 ( .B1(n7679), .B2(n10094), .A(n7662), .ZN(P1_U3283) );
  XNOR2_X1 U9047 ( .A(n7663), .B(n8247), .ZN(n10755) );
  INV_X1 U9048 ( .A(n10755), .ZN(n7676) );
  XNOR2_X1 U9049 ( .A(n7664), .B(n8247), .ZN(n7665) );
  OR2_X1 U9050 ( .A1(n7665), .A2(n10698), .ZN(n7667) );
  AOI22_X1 U9051 ( .A1(n8051), .A2(n10089), .B1(n8133), .B2(n9793), .ZN(n7666)
         );
  NAND2_X1 U9052 ( .A1(n7667), .A2(n7666), .ZN(n10753) );
  INV_X1 U9053 ( .A(n7672), .ZN(n10751) );
  INV_X1 U9054 ( .A(n7668), .ZN(n7669) );
  OAI211_X1 U9055 ( .C1(n10751), .C2(n7669), .A(n10192), .B(n5155), .ZN(n10749) );
  OAI22_X1 U9056 ( .A1(n10707), .A2(n7670), .B1(n8048), .B2(n10718), .ZN(n7671) );
  AOI21_X1 U9057 ( .B1(n7672), .B2(n10081), .A(n7671), .ZN(n7673) );
  OAI21_X1 U9058 ( .B1(n10749), .B2(n10010), .A(n7673), .ZN(n7674) );
  AOI21_X1 U9059 ( .B1(n10753), .B2(n10707), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9060 ( .B1(n7676), .B2(n10094), .A(n7675), .ZN(P1_U3282) );
  OAI211_X1 U9061 ( .C1(n7679), .C2(n10183), .A(n7678), .B(n7677), .ZN(n7683)
         );
  OAI22_X1 U9062 ( .A1(n8005), .A2(n10131), .B1(n10757), .B2(n7269), .ZN(n7680) );
  AOI21_X1 U9063 ( .B1(n7683), .B2(n10757), .A(n7680), .ZN(n7681) );
  INV_X1 U9064 ( .A(n7681), .ZN(P1_U3532) );
  OAI22_X1 U9065 ( .A1(n8005), .A2(n10220), .B1(n10761), .B2(n5868), .ZN(n7682) );
  AOI21_X1 U9066 ( .B1(n7683), .B2(n10761), .A(n7682), .ZN(n7684) );
  INV_X1 U9067 ( .A(n7684), .ZN(P1_U3483) );
  AOI21_X1 U9068 ( .B1(n7686), .B2(n7685), .A(n4939), .ZN(n7694) );
  NOR2_X1 U9069 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7687), .ZN(n10421) );
  OAI22_X1 U9070 ( .A1(n9774), .A2(n7689), .B1(n9772), .B2(n7688), .ZN(n7690)
         );
  AOI211_X1 U9071 ( .C1(n9762), .C2(n9794), .A(n10421), .B(n7690), .ZN(n7693)
         );
  NAND2_X1 U9072 ( .A1(n7691), .A2(n9546), .ZN(n7692) );
  OAI211_X1 U9073 ( .C1(n7694), .C2(n9541), .A(n7693), .B(n7692), .ZN(P1_U3221) );
  INV_X1 U9074 ( .A(n7695), .ZN(n7736) );
  AOI21_X1 U9075 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n10241), .A(n7696), .ZN(
        n7697) );
  OAI21_X1 U9076 ( .B1(n7736), .B2(n7238), .A(n7697), .ZN(P1_U3335) );
  MUX2_X1 U9077 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9417), .Z(n7809) );
  XNOR2_X1 U9078 ( .A(n7809), .B(n7816), .ZN(n7811) );
  MUX2_X1 U9079 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9417), .Z(n7702) );
  MUX2_X1 U9080 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9417), .Z(n7701) );
  XNOR2_X1 U9081 ( .A(n7701), .B(n10529), .ZN(n10538) );
  XNOR2_X1 U9082 ( .A(n7702), .B(n10549), .ZN(n10551) );
  NAND2_X1 U9083 ( .A1(n10552), .A2(n10551), .ZN(n10550) );
  XOR2_X1 U9084 ( .A(n7811), .B(n7812), .Z(n7720) );
  AOI22_X1 U9085 ( .A1(n10549), .A2(n6281), .B1(P2_REG1_REG_6__SCAN_IN), .B2(
        n7707), .ZN(n10555) );
  NAND2_X1 U9086 ( .A1(n7704), .A2(n10529), .ZN(n7705) );
  NAND2_X1 U9087 ( .A1(n7705), .A2(n10533), .ZN(n10554) );
  XNOR2_X1 U9088 ( .A(n7706), .B(n7821), .ZN(n7814) );
  XOR2_X1 U9089 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7814), .Z(n7718) );
  AOI22_X1 U9090 ( .A1(n10549), .A2(n7772), .B1(P2_REG2_REG_6__SCAN_IN), .B2(
        n7707), .ZN(n10547) );
  NAND2_X1 U9091 ( .A1(n7710), .A2(n10529), .ZN(n7711) );
  NAND2_X1 U9092 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n10531), .ZN(n10530) );
  NAND2_X1 U9093 ( .A1(n7711), .A2(n10530), .ZN(n10546) );
  OAI21_X1 U9094 ( .B1(n7712), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7823), .ZN(
        n7713) );
  NAND2_X1 U9095 ( .A1(n7713), .A2(n10578), .ZN(n7716) );
  AOI21_X1 U9096 ( .B1(n10564), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7714), .ZN(
        n7715) );
  OAI211_X1 U9097 ( .C1(n9008), .C2(n7821), .A(n7716), .B(n7715), .ZN(n7717)
         );
  AOI21_X1 U9098 ( .B1(n10579), .B2(n7718), .A(n7717), .ZN(n7719) );
  OAI21_X1 U9099 ( .B1(n7720), .B2(n10536), .A(n7719), .ZN(P2_U3189) );
  INV_X1 U9100 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7721) );
  NOR2_X1 U9101 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7721), .ZN(n7828) );
  NOR2_X1 U9102 ( .A1(n7761), .A2(n8700), .ZN(n7722) );
  AOI211_X1 U9103 ( .C1(n8685), .C2(n8924), .A(n7828), .B(n7722), .ZN(n7723)
         );
  OAI21_X1 U9104 ( .B1(n7757), .B2(n8654), .A(n7723), .ZN(n7733) );
  XNOR2_X1 U9105 ( .A(n7876), .B(n8574), .ZN(n7737) );
  XNOR2_X1 U9106 ( .A(n7737), .B(n7941), .ZN(n7725) );
  AND2_X1 U9107 ( .A1(n7724), .A2(n7725), .ZN(n7726) );
  INV_X1 U9108 ( .A(n7725), .ZN(n7729) );
  NAND3_X1 U9109 ( .A1(n7730), .A2(n7729), .A3(n7728), .ZN(n7731) );
  AOI21_X1 U9110 ( .B1(n7739), .B2(n7731), .A(n8691), .ZN(n7732) );
  AOI211_X1 U9111 ( .C1(n7876), .C2(n8689), .A(n7733), .B(n7732), .ZN(n7734)
         );
  INV_X1 U9112 ( .A(n7734), .ZN(P2_U3161) );
  INV_X1 U9113 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7735) );
  OAI222_X1 U9114 ( .A1(n4925), .A2(n7736), .B1(n8906), .B2(P2_U3151), .C1(
        n7735), .C2(n9415), .ZN(P2_U3275) );
  INV_X1 U9115 ( .A(n7950), .ZN(n7751) );
  NAND2_X1 U9116 ( .A1(n7737), .A2(n7852), .ZN(n7738) );
  XNOR2_X1 U9117 ( .A(n7950), .B(n8542), .ZN(n7969) );
  XNOR2_X1 U9118 ( .A(n7969), .B(n8924), .ZN(n7741) );
  AOI21_X1 U9119 ( .B1(n7740), .B2(n7741), .A(n8691), .ZN(n7744) );
  INV_X1 U9120 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U9121 ( .A1(n7744), .A2(n7971), .ZN(n7750) );
  INV_X1 U9122 ( .A(n7745), .ZN(n7849) );
  NOR2_X1 U9123 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6329), .ZN(n7889) );
  AOI21_X1 U9124 ( .B1(n8710), .B2(n7941), .A(n7889), .ZN(n7746) );
  OAI21_X1 U9125 ( .B1(n7747), .B2(n8712), .A(n7746), .ZN(n7748) );
  AOI21_X1 U9126 ( .B1(n7849), .B2(n8715), .A(n7748), .ZN(n7749) );
  OAI211_X1 U9127 ( .C1(n7751), .C2(n8719), .A(n7750), .B(n7749), .ZN(P2_U3171) );
  INV_X1 U9128 ( .A(n7755), .ZN(n8751) );
  XNOR2_X1 U9129 ( .A(n7752), .B(n8751), .ZN(n7869) );
  NAND2_X1 U9130 ( .A1(n7753), .A2(n7754), .ZN(n7756) );
  XNOR2_X1 U9131 ( .A(n7756), .B(n7755), .ZN(n7871) );
  NAND2_X1 U9132 ( .A1(n7871), .A2(n9192), .ZN(n7764) );
  INV_X1 U9133 ( .A(n9093), .ZN(n9171) );
  NAND2_X1 U9134 ( .A1(n9171), .A2(n8924), .ZN(n7760) );
  NOR2_X1 U9135 ( .A1(n9267), .A2(n7757), .ZN(n7758) );
  AOI21_X1 U9136 ( .B1(n9194), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7758), .ZN(
        n7759) );
  OAI211_X1 U9137 ( .C1(n7761), .C2(n9175), .A(n7760), .B(n7759), .ZN(n7762)
         );
  AOI21_X1 U9138 ( .B1(n9253), .B2(n7876), .A(n7762), .ZN(n7763) );
  OAI211_X1 U9139 ( .C1(n7869), .C2(n9155), .A(n7764), .B(n7763), .ZN(P2_U3225) );
  INV_X1 U9140 ( .A(n8790), .ZN(n7765) );
  NOR2_X1 U9141 ( .A1(n8746), .A2(n7765), .ZN(n7769) );
  INV_X1 U9142 ( .A(n7767), .ZN(n7768) );
  AOI21_X1 U9143 ( .B1(n7769), .B2(n7766), .A(n7768), .ZN(n10728) );
  XNOR2_X1 U9144 ( .A(n7770), .B(n8746), .ZN(n7771) );
  AOI222_X1 U9145 ( .A1(n9340), .A2(n7771), .B1(n8925), .B2(n9335), .C1(n8927), 
        .C2(n9334), .ZN(n10726) );
  MUX2_X1 U9146 ( .A(n7772), .B(n10726), .S(n9269), .Z(n7777) );
  INV_X1 U9147 ( .A(n7773), .ZN(n7774) );
  AOI22_X1 U9148 ( .A1(n9253), .A2(n7775), .B1(n9188), .B2(n7774), .ZN(n7776)
         );
  OAI211_X1 U9149 ( .C1(n10728), .C2(n9274), .A(n7777), .B(n7776), .ZN(
        P2_U3227) );
  NOR2_X1 U9150 ( .A1(n9189), .A2(n7778), .ZN(n8526) );
  OAI21_X1 U9151 ( .B1(n7779), .B2(n8744), .A(n7766), .ZN(n10723) );
  OAI22_X1 U9152 ( .A1(n9265), .A2(n10720), .B1(n7780), .B2(n9267), .ZN(n7786)
         );
  XNOR2_X1 U9153 ( .A(n7781), .B(n8744), .ZN(n7784) );
  NAND2_X1 U9154 ( .A1(n10723), .A2(n8155), .ZN(n7783) );
  AOI22_X1 U9155 ( .A1(n8928), .A2(n9334), .B1(n9335), .B2(n8926), .ZN(n7782)
         );
  OAI211_X1 U9156 ( .C1(n9323), .C2(n7784), .A(n7783), .B(n7782), .ZN(n10721)
         );
  MUX2_X1 U9157 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10721), .S(n9269), .Z(n7785)
         );
  AOI211_X1 U9158 ( .C1(n8526), .C2(n10723), .A(n7786), .B(n7785), .ZN(n7787)
         );
  INV_X1 U9159 ( .A(n7787), .ZN(P2_U3228) );
  OAI21_X1 U9160 ( .B1(n7790), .B2(n7789), .A(n7788), .ZN(n7791) );
  NAND2_X1 U9161 ( .A1(n7791), .A2(n9768), .ZN(n7796) );
  OAI22_X1 U9162 ( .A1(n9774), .A2(n7792), .B1(n9770), .B2(n8047), .ZN(n7793)
         );
  AOI211_X1 U9163 ( .C1(n9529), .C2(n9795), .A(n7794), .B(n7793), .ZN(n7795)
         );
  OAI211_X1 U9164 ( .C1(n7797), .C2(n9779), .A(n7796), .B(n7795), .ZN(P1_U3231) );
  INV_X1 U9165 ( .A(n7801), .ZN(n8248) );
  XNOR2_X1 U9166 ( .A(n7798), .B(n8248), .ZN(n7862) );
  OAI21_X1 U9167 ( .B1(n7801), .B2(n7800), .A(n7799), .ZN(n7802) );
  AOI222_X1 U9168 ( .A1(n10659), .A2(n7802), .B1(n9791), .B2(n10089), .C1(
        n9792), .C2(n8133), .ZN(n7859) );
  OAI22_X1 U9169 ( .A1(n10707), .A2(n5909), .B1(n8122), .B2(n10718), .ZN(n7803) );
  AOI21_X1 U9170 ( .B1(n8117), .B2(n10081), .A(n7803), .ZN(n7806) );
  AOI21_X1 U9171 ( .B1(n8117), .B2(n5155), .A(n10660), .ZN(n7804) );
  AND2_X1 U9172 ( .A1(n7804), .A2(n7955), .ZN(n7861) );
  NAND2_X1 U9173 ( .A1(n7861), .A2(n10674), .ZN(n7805) );
  OAI211_X1 U9174 ( .C1(n7859), .C2(n10714), .A(n7806), .B(n7805), .ZN(n7807)
         );
  AOI21_X1 U9175 ( .B1(n10016), .B2(n7862), .A(n7807), .ZN(n7808) );
  INV_X1 U9176 ( .A(n7808), .ZN(P1_U3281) );
  MUX2_X1 U9177 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9417), .Z(n7879) );
  XNOR2_X1 U9178 ( .A(n7879), .B(n7884), .ZN(n7880) );
  INV_X1 U9179 ( .A(n7809), .ZN(n7810) );
  XOR2_X1 U9180 ( .A(n7880), .B(n7881), .Z(n7834) );
  OAI22_X1 U9181 ( .A1(n7816), .A2(n7815), .B1(n7814), .B2(n7813), .ZN(n7819)
         );
  MUX2_X1 U9182 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7817), .S(n7884), .Z(n7818)
         );
  NAND2_X1 U9183 ( .A1(n7818), .A2(n7819), .ZN(n7882) );
  OAI21_X1 U9184 ( .B1(n7819), .B2(n7818), .A(n7882), .ZN(n7832) );
  AOI22_X1 U9185 ( .A1(n7820), .A2(n6315), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n7884), .ZN(n7826) );
  NAND2_X1 U9186 ( .A1(n7822), .A2(n7821), .ZN(n7824) );
  NAND2_X1 U9187 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  OAI21_X1 U9188 ( .B1(n7826), .B2(n7825), .A(n7885), .ZN(n7827) );
  NAND2_X1 U9189 ( .A1(n7827), .A2(n10578), .ZN(n7830) );
  AOI21_X1 U9190 ( .B1(n10564), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7828), .ZN(
        n7829) );
  OAI211_X1 U9191 ( .C1(n9008), .C2(n7884), .A(n7830), .B(n7829), .ZN(n7831)
         );
  AOI21_X1 U9192 ( .B1(n10579), .B2(n7832), .A(n7831), .ZN(n7833) );
  OAI21_X1 U9193 ( .B1(n7834), .B2(n10536), .A(n7833), .ZN(P2_U3190) );
  XNOR2_X1 U9194 ( .A(n7835), .B(n5329), .ZN(n7903) );
  INV_X1 U9195 ( .A(n7753), .ZN(n7836) );
  AOI21_X1 U9196 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7900) );
  NOR2_X1 U9197 ( .A1(n9265), .A2(n7905), .ZN(n7845) );
  NAND2_X1 U9198 ( .A1(n9171), .A2(n7941), .ZN(n7842) );
  NOR2_X1 U9199 ( .A1(n9267), .A2(n7839), .ZN(n7840) );
  AOI21_X1 U9200 ( .B1(n9194), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7840), .ZN(
        n7841) );
  OAI211_X1 U9201 ( .C1(n7843), .C2(n9175), .A(n7842), .B(n7841), .ZN(n7844)
         );
  AOI211_X1 U9202 ( .C1(n7900), .C2(n9192), .A(n7845), .B(n7844), .ZN(n7846)
         );
  OAI21_X1 U9203 ( .B1(n7903), .B2(n9155), .A(n7846), .ZN(P2_U3226) );
  XNOR2_X1 U9204 ( .A(n7847), .B(n6621), .ZN(n7943) );
  NAND2_X1 U9205 ( .A1(n9171), .A2(n8923), .ZN(n7851) );
  AOI22_X1 U9206 ( .A1(n9189), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9188), .B2(
        n7849), .ZN(n7850) );
  OAI211_X1 U9207 ( .C1(n7852), .C2(n9175), .A(n7851), .B(n7850), .ZN(n7853)
         );
  AOI21_X1 U9208 ( .B1(n9253), .B2(n7950), .A(n7853), .ZN(n7856) );
  XNOR2_X1 U9209 ( .A(n7854), .B(n6621), .ZN(n7945) );
  NAND2_X1 U9210 ( .A1(n7945), .A2(n9192), .ZN(n7855) );
  OAI211_X1 U9211 ( .C1(n7943), .C2(n9155), .A(n7856), .B(n7855), .ZN(P2_U3224) );
  INV_X1 U9212 ( .A(n7857), .ZN(n7898) );
  AOI22_X1 U9213 ( .A1(n6726), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10241), .ZN(n7858) );
  OAI21_X1 U9214 ( .B1(n7898), .B2(n7238), .A(n7858), .ZN(P1_U3334) );
  INV_X1 U9215 ( .A(n7859), .ZN(n7860) );
  AOI211_X1 U9216 ( .C1(n10754), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7867)
         );
  INV_X1 U9217 ( .A(n10220), .ZN(n7863) );
  AOI22_X1 U9218 ( .A1(n8117), .A2(n7863), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n10758), .ZN(n7864) );
  OAI21_X1 U9219 ( .B1(n7867), .B2(n10758), .A(n7864), .ZN(P1_U3489) );
  AOI22_X1 U9220 ( .A1(n8117), .A2(n7865), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n10756), .ZN(n7866) );
  OAI21_X1 U9221 ( .B1(n7867), .B2(n10756), .A(n7866), .ZN(P1_U3534) );
  AOI22_X1 U9222 ( .A1(n8925), .A2(n9334), .B1(n9335), .B2(n8924), .ZN(n7868)
         );
  OAI21_X1 U9223 ( .B1(n7869), .B2(n9323), .A(n7868), .ZN(n7870) );
  AOI21_X1 U9224 ( .B1(n10775), .B2(n7871), .A(n7870), .ZN(n7878) );
  INV_X1 U9225 ( .A(n7876), .ZN(n7873) );
  INV_X1 U9226 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7872) );
  OAI22_X1 U9227 ( .A1(n7873), .A2(n9403), .B1(n6696), .B2(n7872), .ZN(n7874)
         );
  INV_X1 U9228 ( .A(n7874), .ZN(n7875) );
  OAI21_X1 U9229 ( .B1(n7878), .B2(n10792), .A(n7875), .ZN(P2_U3414) );
  AOI22_X1 U9230 ( .A1(n7876), .A2(n9331), .B1(n10782), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7877) );
  OAI21_X1 U9231 ( .B1(n7878), .B2(n10782), .A(n7877), .ZN(P2_U3467) );
  MUX2_X1 U9232 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9417), .Z(n7915) );
  XNOR2_X1 U9233 ( .A(n7915), .B(n7921), .ZN(n7917) );
  XOR2_X1 U9234 ( .A(n7917), .B(n7918), .Z(n7895) );
  NAND2_X1 U9235 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7884), .ZN(n7883) );
  XOR2_X1 U9236 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7922), .Z(n7893) );
  NAND2_X1 U9237 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7884), .ZN(n7886) );
  OAI21_X1 U9238 ( .B1(n7887), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7929), .ZN(
        n7888) );
  NAND2_X1 U9239 ( .A1(n7888), .A2(n10578), .ZN(n7891) );
  AOI21_X1 U9240 ( .B1(n10564), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7889), .ZN(
        n7890) );
  OAI211_X1 U9241 ( .C1(n9008), .C2(n5389), .A(n7891), .B(n7890), .ZN(n7892)
         );
  AOI21_X1 U9242 ( .B1(n7893), .B2(n10579), .A(n7892), .ZN(n7894) );
  OAI21_X1 U9243 ( .B1(n7895), .B2(n10536), .A(n7894), .ZN(P2_U3191) );
  INV_X1 U9244 ( .A(n7896), .ZN(n7909) );
  AOI22_X1 U9245 ( .A1(n8508), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10241), .ZN(n7897) );
  OAI21_X1 U9246 ( .B1(n7909), .B2(n7238), .A(n7897), .ZN(P1_U3333) );
  INV_X1 U9247 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7899) );
  OAI222_X1 U9248 ( .A1(n9415), .A2(n7899), .B1(n4925), .B2(n7898), .C1(
        P2_U3151), .C2(n8771), .ZN(P2_U3274) );
  NAND2_X1 U9249 ( .A1(n7900), .A2(n10775), .ZN(n7902) );
  AOI22_X1 U9250 ( .A1(n9334), .A2(n8926), .B1(n7941), .B2(n9335), .ZN(n7901)
         );
  OAI211_X1 U9251 ( .C1(n9323), .C2(n7903), .A(n7902), .B(n7901), .ZN(n7911)
         );
  INV_X1 U9252 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7904) );
  OAI22_X1 U9253 ( .A1(n7905), .A2(n9403), .B1(n6696), .B2(n7904), .ZN(n7906)
         );
  AOI21_X1 U9254 ( .B1(n7911), .B2(n6696), .A(n7906), .ZN(n7907) );
  INV_X1 U9255 ( .A(n7907), .ZN(P2_U3411) );
  OAI222_X1 U9256 ( .A1(n9415), .A2(n7910), .B1(n4925), .B2(n7909), .C1(
        P2_U3151), .C2(n7908), .ZN(P2_U3273) );
  NAND2_X1 U9257 ( .A1(n7911), .A2(n10791), .ZN(n7914) );
  NAND2_X1 U9258 ( .A1(n9331), .A2(n7912), .ZN(n7913) );
  OAI211_X1 U9259 ( .C1(n10791), .C2(n7813), .A(n7914), .B(n7913), .ZN(
        P2_U3466) );
  MUX2_X1 U9260 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9417), .Z(n7982) );
  XNOR2_X1 U9261 ( .A(n7982), .B(n7987), .ZN(n7983) );
  INV_X1 U9262 ( .A(n7915), .ZN(n7916) );
  XOR2_X1 U9263 ( .A(n7983), .B(n7984), .Z(n7940) );
  INV_X1 U9264 ( .A(n7919), .ZN(n7920) );
  MUX2_X1 U9265 ( .A(n7923), .B(P2_REG1_REG_10__SCAN_IN), .S(n7927), .Z(n7924)
         );
  OAI21_X1 U9266 ( .B1(n7925), .B2(n7924), .A(n7985), .ZN(n7938) );
  INV_X1 U9267 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7926) );
  AOI22_X1 U9268 ( .A1(n7927), .A2(n7926), .B1(P2_REG2_REG_10__SCAN_IN), .B2(
        n7987), .ZN(n7932) );
  NAND2_X1 U9269 ( .A1(n7928), .A2(n5389), .ZN(n7930) );
  NAND2_X1 U9270 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NAND2_X1 U9271 ( .A1(n7932), .A2(n7931), .ZN(n7988) );
  OAI21_X1 U9272 ( .B1(n7932), .B2(n7931), .A(n7988), .ZN(n7933) );
  NAND2_X1 U9273 ( .A1(n7933), .A2(n10578), .ZN(n7936) );
  INV_X1 U9274 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U9275 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7934), .ZN(n7977) );
  AOI21_X1 U9276 ( .B1(n10564), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7977), .ZN(
        n7935) );
  OAI211_X1 U9277 ( .C1(n9008), .C2(n7987), .A(n7936), .B(n7935), .ZN(n7937)
         );
  AOI21_X1 U9278 ( .B1(n10579), .B2(n7938), .A(n7937), .ZN(n7939) );
  OAI21_X1 U9279 ( .B1(n7940), .B2(n10536), .A(n7939), .ZN(P2_U3192) );
  AOI22_X1 U9280 ( .A1(n9335), .A2(n8923), .B1(n7941), .B2(n9334), .ZN(n7942)
         );
  OAI21_X1 U9281 ( .B1(n7943), .B2(n9323), .A(n7942), .ZN(n7944) );
  AOI21_X1 U9282 ( .B1(n7945), .B2(n10775), .A(n7944), .ZN(n7952) );
  NOR2_X1 U9283 ( .A1(n6696), .A2(n6328), .ZN(n7946) );
  AOI21_X1 U9284 ( .B1(n9386), .B2(n7950), .A(n7946), .ZN(n7947) );
  OAI21_X1 U9285 ( .B1(n7952), .B2(n10792), .A(n7947), .ZN(P2_U3417) );
  INV_X1 U9286 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7948) );
  NOR2_X1 U9287 ( .A1(n10791), .A2(n7948), .ZN(n7949) );
  AOI21_X1 U9288 ( .B1(n7950), .B2(n9331), .A(n7949), .ZN(n7951) );
  OAI21_X1 U9289 ( .B1(n7952), .B2(n10782), .A(n7951), .ZN(P2_U3468) );
  XOR2_X1 U9290 ( .A(n8250), .B(n7953), .Z(n10184) );
  INV_X1 U9291 ( .A(n8035), .ZN(n7954) );
  AOI211_X1 U9292 ( .C1(n10180), .C2(n7955), .A(n10660), .B(n7954), .ZN(n10179) );
  INV_X1 U9293 ( .A(n9518), .ZN(n7956) );
  AOI22_X1 U9294 ( .A1(n10714), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7956), .B2(
        n10638), .ZN(n7957) );
  OAI21_X1 U9295 ( .B1(n7958), .B2(n10670), .A(n7957), .ZN(n7962) );
  OAI21_X1 U9296 ( .B1(n8250), .B2(n7959), .A(n8029), .ZN(n7960) );
  AOI222_X1 U9297 ( .A1(n10659), .A2(n7960), .B1(n9790), .B2(n10089), .C1(
        n8051), .C2(n8133), .ZN(n10182) );
  NOR2_X1 U9298 ( .A1(n10182), .A2(n10714), .ZN(n7961) );
  AOI211_X1 U9299 ( .C1(n10179), .C2(n10674), .A(n7962), .B(n7961), .ZN(n7963)
         );
  OAI21_X1 U9300 ( .B1(n10094), .B2(n10184), .A(n7963), .ZN(P1_U3280) );
  INV_X1 U9301 ( .A(n7964), .ZN(n7968) );
  NAND2_X1 U9302 ( .A1(n10241), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7965) );
  OAI211_X1 U9303 ( .C1(n7968), .C2(n7238), .A(n7965), .B(n8509), .ZN(P1_U3332) );
  OR2_X1 U9304 ( .A1(n7966), .A2(P2_U3151), .ZN(n8917) );
  NAND2_X1 U9305 ( .A1(n9409), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7967) );
  OAI211_X1 U9306 ( .C1(n7968), .C2(n4925), .A(n8917), .B(n7967), .ZN(P2_U3272) );
  NAND2_X1 U9307 ( .A1(n7969), .A2(n8924), .ZN(n7970) );
  XNOR2_X1 U9308 ( .A(n10735), .B(n8574), .ZN(n7972) );
  AOI21_X1 U9309 ( .B1(n8923), .B2(n7974), .A(n8057), .ZN(n7981) );
  NOR2_X1 U9310 ( .A1(n7975), .A2(n8700), .ZN(n7976) );
  AOI211_X1 U9311 ( .C1(n8685), .C2(n8163), .A(n7977), .B(n7976), .ZN(n7978)
         );
  OAI21_X1 U9312 ( .B1(n8152), .B2(n8654), .A(n7978), .ZN(n7979) );
  AOI21_X1 U9313 ( .B1(n10735), .B2(n8689), .A(n7979), .ZN(n7980) );
  OAI21_X1 U9314 ( .B1(n7981), .B2(n8691), .A(n7980), .ZN(P2_U3157) );
  MUX2_X1 U9315 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9417), .Z(n8066) );
  XNOR2_X1 U9316 ( .A(n8066), .B(n8072), .ZN(n8068) );
  OAI22_X1 U9317 ( .A1(n7984), .A2(n7983), .B1(n7982), .B2(n7987), .ZN(n8069)
         );
  XOR2_X1 U9318 ( .A(n8068), .B(n8069), .Z(n7997) );
  NAND2_X1 U9319 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7987), .ZN(n7986) );
  NAND2_X1 U9320 ( .A1(n7986), .A2(n7985), .ZN(n8070) );
  XOR2_X1 U9321 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8074), .Z(n7995) );
  NAND2_X1 U9322 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7987), .ZN(n7989) );
  NAND2_X1 U9323 ( .A1(n7989), .A2(n7988), .ZN(n8078) );
  XNOR2_X1 U9324 ( .A(n8078), .B(n8072), .ZN(n7990) );
  NAND2_X1 U9325 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n7990), .ZN(n8079) );
  OAI21_X1 U9326 ( .B1(n7990), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8079), .ZN(
        n7991) );
  NAND2_X1 U9327 ( .A1(n7991), .A2(n10578), .ZN(n7993) );
  INV_X1 U9328 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9625) );
  NOR2_X1 U9329 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9625), .ZN(n8061) );
  AOI21_X1 U9330 ( .B1(n10564), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8061), .ZN(
        n7992) );
  OAI211_X1 U9331 ( .C1(n9008), .C2(n5391), .A(n7993), .B(n7992), .ZN(n7994)
         );
  AOI21_X1 U9332 ( .B1(n7995), .B2(n10579), .A(n7994), .ZN(n7996) );
  OAI21_X1 U9333 ( .B1(n7997), .B2(n10536), .A(n7996), .ZN(P2_U3193) );
  AOI21_X1 U9334 ( .B1(n7999), .B2(n7998), .A(n4982), .ZN(n8008) );
  NOR2_X1 U9335 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8000), .ZN(n10504) );
  AOI21_X1 U9336 ( .B1(n9762), .B2(n9792), .A(n10504), .ZN(n8004) );
  INV_X1 U9337 ( .A(n8001), .ZN(n8002) );
  AOI22_X1 U9338 ( .A1(n9529), .A2(n9794), .B1(n8002), .B2(n9759), .ZN(n8003)
         );
  OAI211_X1 U9339 ( .C1(n8005), .C2(n9779), .A(n8004), .B(n8003), .ZN(n8006)
         );
  INV_X1 U9340 ( .A(n8006), .ZN(n8007) );
  OAI21_X1 U9341 ( .B1(n8008), .B2(n9541), .A(n8007), .ZN(P1_U3217) );
  INV_X1 U9342 ( .A(n8009), .ZN(n8517) );
  AOI22_X1 U9343 ( .A1(n8010), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10241), .ZN(n8011) );
  OAI21_X1 U9344 ( .B1(n8517), .B2(n7238), .A(n8011), .ZN(P1_U3331) );
  XNOR2_X1 U9345 ( .A(n8012), .B(n8253), .ZN(n10178) );
  INV_X1 U9346 ( .A(n8253), .ZN(n8014) );
  OAI21_X1 U9347 ( .B1(n4990), .B2(n8014), .A(n8013), .ZN(n8015) );
  AOI222_X1 U9348 ( .A1(n10659), .A2(n8015), .B1(n9788), .B2(n10089), .C1(
        n9790), .C2(n8133), .ZN(n10177) );
  INV_X1 U9349 ( .A(n10177), .ZN(n8022) );
  OR2_X1 U9350 ( .A1(n8016), .A2(n10660), .ZN(n8034) );
  AOI21_X1 U9351 ( .B1(n8016), .B2(n10192), .A(n10663), .ZN(n8018) );
  MUX2_X1 U9352 ( .A(n8034), .B(n8018), .S(n8017), .Z(n10176) );
  INV_X1 U9353 ( .A(n9773), .ZN(n8019) );
  AOI22_X1 U9354 ( .A1(n10714), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8019), .B2(
        n10638), .ZN(n8020) );
  OAI21_X1 U9355 ( .B1(n10176), .B2(n9915), .A(n8020), .ZN(n8021) );
  AOI21_X1 U9356 ( .B1(n8022), .B2(n10707), .A(n8021), .ZN(n8023) );
  OAI21_X1 U9357 ( .B1(n10094), .B2(n10178), .A(n8023), .ZN(P1_U3278) );
  NAND2_X1 U9358 ( .A1(n8025), .A2(n8251), .ZN(n8026) );
  NAND2_X1 U9359 ( .A1(n8024), .A2(n8026), .ZN(n8179) );
  INV_X1 U9360 ( .A(n8027), .ZN(n8028) );
  NAND2_X1 U9361 ( .A1(n10707), .A2(n8028), .ZN(n10619) );
  NAND2_X1 U9362 ( .A1(n8029), .A2(n8339), .ZN(n8030) );
  XNOR2_X1 U9363 ( .A(n8030), .B(n8251), .ZN(n8032) );
  OAI22_X1 U9364 ( .A1(n9426), .A2(n10703), .B1(n9427), .B2(n10701), .ZN(n8031) );
  AOI21_X1 U9365 ( .B1(n8032), .B2(n10659), .A(n8031), .ZN(n8033) );
  OAI21_X1 U9366 ( .B1(n8179), .B2(n10655), .A(n8033), .ZN(n8180) );
  NAND2_X1 U9367 ( .A1(n8180), .A2(n10707), .ZN(n8040) );
  AOI21_X1 U9368 ( .B1(n9431), .B2(n8035), .A(n8034), .ZN(n8181) );
  INV_X1 U9369 ( .A(n9431), .ZN(n8189) );
  NOR2_X1 U9370 ( .A1(n8189), .A2(n10670), .ZN(n8038) );
  OAI22_X1 U9371 ( .A1(n10707), .A2(n8036), .B1(n9428), .B2(n10718), .ZN(n8037) );
  AOI211_X1 U9372 ( .C1(n8181), .C2(n10674), .A(n8038), .B(n8037), .ZN(n8039)
         );
  OAI211_X1 U9373 ( .C1(n8179), .C2(n10619), .A(n8040), .B(n8039), .ZN(
        P1_U3279) );
  INV_X1 U9374 ( .A(n8041), .ZN(n8043) );
  NOR3_X1 U9375 ( .A1(n4982), .A2(n8043), .A3(n8042), .ZN(n8046) );
  INV_X1 U9376 ( .A(n8044), .ZN(n8045) );
  OAI21_X1 U9377 ( .B1(n8046), .B2(n8045), .A(n9768), .ZN(n8053) );
  NAND2_X1 U9378 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10436) );
  INV_X1 U9379 ( .A(n10436), .ZN(n8050) );
  OAI22_X1 U9380 ( .A1(n9774), .A2(n8048), .B1(n9772), .B2(n8047), .ZN(n8049)
         );
  AOI211_X1 U9381 ( .C1(n9762), .C2(n8051), .A(n8050), .B(n8049), .ZN(n8052)
         );
  OAI211_X1 U9382 ( .C1(n10751), .C2(n9779), .A(n8053), .B(n8052), .ZN(
        P1_U3236) );
  INV_X1 U9383 ( .A(n10743), .ZN(n8101) );
  XNOR2_X1 U9384 ( .A(n10743), .B(n8574), .ZN(n8105) );
  XNOR2_X1 U9385 ( .A(n8105), .B(n8163), .ZN(n8055) );
  INV_X1 U9386 ( .A(n8107), .ZN(n8059) );
  NOR3_X1 U9387 ( .A1(n8057), .A2(n8056), .A3(n8055), .ZN(n8058) );
  OAI21_X1 U9388 ( .B1(n8059), .B2(n8058), .A(n8706), .ZN(n8065) );
  INV_X1 U9389 ( .A(n8060), .ZN(n8099) );
  AOI21_X1 U9390 ( .B1(n8710), .B2(n8923), .A(n8061), .ZN(n8062) );
  OAI21_X1 U9391 ( .B1(n8820), .B2(n8712), .A(n8062), .ZN(n8063) );
  AOI21_X1 U9392 ( .B1(n8099), .B2(n8715), .A(n8063), .ZN(n8064) );
  OAI211_X1 U9393 ( .C1(n8101), .C2(n8719), .A(n8065), .B(n8064), .ZN(P2_U3176) );
  MUX2_X1 U9394 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9417), .Z(n8932) );
  XNOR2_X1 U9395 ( .A(n8932), .B(n8931), .ZN(n8933) );
  INV_X1 U9396 ( .A(n8066), .ZN(n8067) );
  XOR2_X1 U9397 ( .A(n8933), .B(n8934), .Z(n8089) );
  INV_X1 U9398 ( .A(n8070), .ZN(n8071) );
  MUX2_X1 U9399 ( .A(n8075), .B(P2_REG1_REG_12__SCAN_IN), .S(n8939), .Z(n8076)
         );
  OAI21_X1 U9400 ( .B1(n8077), .B2(n8076), .A(n8938), .ZN(n8087) );
  AOI22_X1 U9401 ( .A1(n8939), .A2(n6363), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n8931), .ZN(n8082) );
  NAND2_X1 U9402 ( .A1(n8078), .A2(n5391), .ZN(n8080) );
  OAI21_X1 U9403 ( .B1(n8082), .B2(n8081), .A(n8935), .ZN(n8083) );
  NAND2_X1 U9404 ( .A1(n8083), .A2(n10578), .ZN(n8085) );
  NOR2_X1 U9405 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9717), .ZN(n8112) );
  AOI21_X1 U9406 ( .B1(n10564), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8112), .ZN(
        n8084) );
  OAI211_X1 U9407 ( .C1(n9008), .C2(n8931), .A(n8085), .B(n8084), .ZN(n8086)
         );
  AOI21_X1 U9408 ( .B1(n10579), .B2(n8087), .A(n8086), .ZN(n8088) );
  OAI21_X1 U9409 ( .B1(n8089), .B2(n10536), .A(n8088), .ZN(P2_U3194) );
  NAND2_X1 U9410 ( .A1(n8090), .A2(n8804), .ZN(n8091) );
  XNOR2_X1 U9411 ( .A(n8091), .B(n8754), .ZN(n10742) );
  INV_X1 U9412 ( .A(n10742), .ZN(n8104) );
  INV_X1 U9413 ( .A(n8092), .ZN(n8095) );
  AOI21_X1 U9414 ( .B1(n8093), .B2(n8754), .A(n9323), .ZN(n8094) );
  OAI21_X1 U9415 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8098) );
  AOI22_X1 U9416 ( .A1(n9334), .A2(n8923), .B1(n8195), .B2(n9335), .ZN(n8097)
         );
  NAND2_X1 U9417 ( .A1(n8098), .A2(n8097), .ZN(n10744) );
  AOI22_X1 U9418 ( .A1(n9189), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n9188), .B2(
        n8099), .ZN(n8100) );
  OAI21_X1 U9419 ( .B1(n8101), .B2(n9265), .A(n8100), .ZN(n8102) );
  AOI21_X1 U9420 ( .B1(n10744), .B2(n9269), .A(n8102), .ZN(n8103) );
  OAI21_X1 U9421 ( .B1(n9274), .B2(n8104), .A(n8103), .ZN(P2_U3222) );
  INV_X1 U9422 ( .A(n8105), .ZN(n8106) );
  XOR2_X1 U9423 ( .A(n8574), .B(n10766), .Z(n8108) );
  MUX2_X1 U9424 ( .A(n8109), .B(n8821), .S(n8574), .Z(n8190) );
  NAND2_X1 U9425 ( .A1(n4997), .A2(n8190), .ZN(n8110) );
  XNOR2_X1 U9426 ( .A(n8191), .B(n8110), .ZN(n8116) );
  NOR2_X1 U9427 ( .A1(n8827), .A2(n8712), .ZN(n8111) );
  AOI211_X1 U9428 ( .C1(n8710), .C2(n8163), .A(n8112), .B(n8111), .ZN(n8113)
         );
  OAI21_X1 U9429 ( .B1(n8165), .B2(n8654), .A(n8113), .ZN(n8114) );
  AOI21_X1 U9430 ( .B1(n10766), .B2(n8689), .A(n8114), .ZN(n8115) );
  OAI21_X1 U9431 ( .B1(n8116), .B2(n8691), .A(n8115), .ZN(P2_U3164) );
  INV_X1 U9432 ( .A(n8117), .ZN(n8127) );
  OAI21_X1 U9433 ( .B1(n8120), .B2(n8119), .A(n8118), .ZN(n8121) );
  NAND2_X1 U9434 ( .A1(n8121), .A2(n9768), .ZN(n8126) );
  OAI22_X1 U9435 ( .A1(n9774), .A2(n8122), .B1(n9770), .B2(n9427), .ZN(n8123)
         );
  AOI211_X1 U9436 ( .C1(n9529), .C2(n9792), .A(n8124), .B(n8123), .ZN(n8125)
         );
  OAI211_X1 U9437 ( .C1(n8127), .C2(n9779), .A(n8126), .B(n8125), .ZN(P1_U3224) );
  INV_X1 U9438 ( .A(n8128), .ZN(n8146) );
  AOI22_X1 U9439 ( .A1(n8129), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10241), .ZN(n8130) );
  OAI21_X1 U9440 ( .B1(n8146), .B2(n7238), .A(n8130), .ZN(P1_U3330) );
  OAI21_X1 U9441 ( .B1(n8141), .B2(n8132), .A(n8131), .ZN(n8134) );
  AOI222_X1 U9442 ( .A1(n10659), .A2(n8134), .B1(n9787), .B2(n10089), .C1(
        n9789), .C2(n8133), .ZN(n10174) );
  AOI211_X1 U9443 ( .C1(n10171), .C2(n8136), .A(n10660), .B(n8135), .ZN(n10170) );
  INV_X1 U9444 ( .A(n10171), .ZN(n8138) );
  AOI22_X1 U9445 ( .A1(n10714), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9481), .B2(
        n10638), .ZN(n8137) );
  OAI21_X1 U9446 ( .B1(n8138), .B2(n10670), .A(n8137), .ZN(n8139) );
  AOI21_X1 U9447 ( .B1(n10170), .B2(n10674), .A(n8139), .ZN(n8144) );
  NAND2_X1 U9448 ( .A1(n8142), .A2(n8141), .ZN(n10172) );
  NAND3_X1 U9449 ( .A1(n8140), .A2(n10172), .A3(n10016), .ZN(n8143) );
  OAI211_X1 U9450 ( .C1(n10174), .C2(n10714), .A(n8144), .B(n8143), .ZN(
        P1_U3277) );
  OAI222_X1 U9451 ( .A1(n9415), .A2(n8147), .B1(n4925), .B2(n8146), .C1(n8145), 
        .C2(P2_U3151), .ZN(P2_U3270) );
  NAND2_X1 U9452 ( .A1(n8149), .A2(n8148), .ZN(n8752) );
  INV_X1 U9453 ( .A(n8752), .ZN(n8150) );
  XNOR2_X1 U9454 ( .A(n8151), .B(n8150), .ZN(n10734) );
  INV_X1 U9455 ( .A(n10735), .ZN(n8153) );
  OAI22_X1 U9456 ( .A1(n8153), .A2(n9265), .B1(n8152), .B2(n9267), .ZN(n8160)
         );
  XNOR2_X1 U9457 ( .A(n8154), .B(n8752), .ZN(n8158) );
  NAND2_X1 U9458 ( .A1(n10734), .A2(n8155), .ZN(n8157) );
  AOI22_X1 U9459 ( .A1(n9334), .A2(n8924), .B1(n8163), .B2(n9335), .ZN(n8156)
         );
  OAI211_X1 U9460 ( .C1(n8158), .C2(n9323), .A(n8157), .B(n8156), .ZN(n10739)
         );
  MUX2_X1 U9461 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10739), .S(n9269), .Z(n8159) );
  AOI211_X1 U9462 ( .C1(n10734), .C2(n8526), .A(n8160), .B(n8159), .ZN(n8161)
         );
  INV_X1 U9463 ( .A(n8161), .ZN(P2_U3223) );
  XNOR2_X1 U9464 ( .A(n8162), .B(n8819), .ZN(n8164) );
  AOI222_X1 U9465 ( .A1(n9340), .A2(n8164), .B1(n8163), .B2(n9334), .C1(n9262), 
        .C2(n9335), .ZN(n10763) );
  OAI22_X1 U9466 ( .A1(n9269), .A2(n6363), .B1(n8165), .B2(n9267), .ZN(n8168)
         );
  XNOR2_X1 U9467 ( .A(n8166), .B(n8819), .ZN(n10762) );
  NOR2_X1 U9468 ( .A1(n10762), .A2(n9274), .ZN(n8167) );
  AOI211_X1 U9469 ( .C1(n9253), .C2(n10766), .A(n8168), .B(n8167), .ZN(n8169)
         );
  OAI21_X1 U9470 ( .B1(n10763), .B2(n9194), .A(n8169), .ZN(P2_U3221) );
  OAI211_X1 U9471 ( .C1(n8171), .C2(n8756), .A(n8170), .B(n9340), .ZN(n8173)
         );
  AOI22_X1 U9472 ( .A1(n9334), .A2(n8195), .B1(n9246), .B2(n9335), .ZN(n8172)
         );
  NAND2_X1 U9473 ( .A1(n8173), .A2(n8172), .ZN(n10770) );
  INV_X1 U9474 ( .A(n8828), .ZN(n10769) );
  OAI22_X1 U9475 ( .A1(n10769), .A2(n8174), .B1(n8194), .B2(n9267), .ZN(n8175)
         );
  OAI21_X1 U9476 ( .B1(n10770), .B2(n8175), .A(n9269), .ZN(n8178) );
  XNOR2_X1 U9477 ( .A(n8176), .B(n8756), .ZN(n10772) );
  AOI22_X1 U9478 ( .A1(n10772), .A2(n9192), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9194), .ZN(n8177) );
  NAND2_X1 U9479 ( .A1(n8178), .A2(n8177), .ZN(P2_U3220) );
  INV_X1 U9480 ( .A(n8179), .ZN(n8183) );
  INV_X1 U9481 ( .A(n10665), .ZN(n8182) );
  AOI211_X1 U9482 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8186)
         );
  MUX2_X1 U9483 ( .A(n8184), .B(n8186), .S(n10757), .Z(n8185) );
  OAI21_X1 U9484 ( .B1(n8189), .B2(n10131), .A(n8185), .ZN(P1_U3536) );
  INV_X1 U9485 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8187) );
  MUX2_X1 U9486 ( .A(n8187), .B(n8186), .S(n10761), .Z(n8188) );
  OAI21_X1 U9487 ( .B1(n8189), .B2(n10220), .A(n8188), .ZN(P1_U3495) );
  XNOR2_X1 U9488 ( .A(n8828), .B(n8574), .ZN(n8530) );
  XNOR2_X1 U9489 ( .A(n8530), .B(n9262), .ZN(n8192) );
  OAI211_X1 U9490 ( .C1(n8193), .C2(n8192), .A(n8533), .B(n8706), .ZN(n8200)
         );
  INV_X1 U9491 ( .A(n8194), .ZN(n8198) );
  NOR2_X1 U9492 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6378), .ZN(n8937) );
  AOI21_X1 U9493 ( .B1(n8710), .B2(n8195), .A(n8937), .ZN(n8196) );
  OAI21_X1 U9494 ( .B1(n8833), .B2(n8712), .A(n8196), .ZN(n8197) );
  AOI21_X1 U9495 ( .B1(n8198), .B2(n8715), .A(n8197), .ZN(n8199) );
  OAI211_X1 U9496 ( .C1(n10769), .C2(n8719), .A(n8200), .B(n8199), .ZN(
        P2_U3174) );
  INV_X1 U9497 ( .A(n8201), .ZN(n8205) );
  AOI22_X1 U9498 ( .A1(n5542), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10241), .ZN(n8202) );
  OAI21_X1 U9499 ( .B1(n8205), .B2(n7238), .A(n8202), .ZN(P1_U3329) );
  OAI222_X1 U9500 ( .A1(n4925), .A2(n8205), .B1(P2_U3151), .B2(n8204), .C1(
        n8203), .C2(n9415), .ZN(P2_U3269) );
  XNOR2_X1 U9501 ( .A(n8206), .B(n8354), .ZN(n8207) );
  AOI22_X1 U9502 ( .A1(n8207), .A2(n10659), .B1(n10089), .B2(n9786), .ZN(
        n10168) );
  OAI21_X1 U9503 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n10169) );
  INV_X1 U9504 ( .A(n10169), .ZN(n8220) );
  INV_X1 U9505 ( .A(n10166), .ZN(n8218) );
  AOI21_X1 U9506 ( .B1(n10166), .B2(n8211), .A(n10660), .ZN(n8212) );
  AND2_X1 U9507 ( .A1(n8212), .A2(n10080), .ZN(n10164) );
  NAND2_X1 U9508 ( .A1(n10164), .A2(n10674), .ZN(n8217) );
  INV_X1 U9509 ( .A(n10085), .ZN(n8215) );
  OAI22_X1 U9510 ( .A1(n10707), .A2(n8213), .B1(n9490), .B2(n10718), .ZN(n8214) );
  AOI21_X1 U9511 ( .B1(n8215), .B2(n9788), .A(n8214), .ZN(n8216) );
  OAI211_X1 U9512 ( .C1(n8218), .C2(n10670), .A(n8217), .B(n8216), .ZN(n8219)
         );
  AOI21_X1 U9513 ( .B1(n8220), .B2(n10016), .A(n8219), .ZN(n8221) );
  OAI21_X1 U9514 ( .B1(n10714), .B2(n10168), .A(n8221), .ZN(P1_U3276) );
  INV_X1 U9515 ( .A(n8281), .ZN(n8265) );
  INV_X1 U9516 ( .A(SI_29_), .ZN(n9646) );
  INV_X1 U9517 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8226) );
  INV_X1 U9518 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8722) );
  MUX2_X1 U9519 ( .A(n8226), .B(n8722), .S(n5701), .Z(n8227) );
  INV_X1 U9520 ( .A(SI_30_), .ZN(n9645) );
  NAND2_X1 U9521 ( .A1(n8227), .A2(n9645), .ZN(n8266) );
  INV_X1 U9522 ( .A(n8227), .ZN(n8228) );
  NAND2_X1 U9523 ( .A1(n8228), .A2(SI_30_), .ZN(n8229) );
  NAND2_X1 U9524 ( .A1(n8266), .A2(n8229), .ZN(n8267) );
  NAND2_X1 U9525 ( .A1(n8230), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8231) );
  INV_X1 U9526 ( .A(n8434), .ZN(n8498) );
  NAND2_X1 U9527 ( .A1(n10159), .A2(n10074), .ZN(n8362) );
  AND2_X1 U9528 ( .A1(n8362), .A2(n8233), .ZN(n8356) );
  INV_X1 U9529 ( .A(n8356), .ZN(n8483) );
  INV_X1 U9530 ( .A(n8481), .ZN(n8254) );
  AND4_X1 U9531 ( .A1(n10652), .A2(n8235), .A3(n10604), .A4(n8234), .ZN(n8236)
         );
  NAND4_X1 U9532 ( .A1(n8237), .A2(n10696), .A3(n8236), .A4(n10187), .ZN(n8238) );
  NOR2_X1 U9533 ( .A1(n8239), .A2(n8238), .ZN(n8241) );
  NAND4_X1 U9534 ( .A1(n8292), .A2(n8242), .A3(n8241), .A4(n8240), .ZN(n8243)
         );
  NOR3_X1 U9535 ( .A1(n8248), .A2(n8247), .A3(n8246), .ZN(n8249) );
  NAND3_X1 U9536 ( .A1(n8251), .A2(n8250), .A3(n8249), .ZN(n8252) );
  OR4_X1 U9537 ( .A1(n8483), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n8257) );
  NAND2_X1 U9538 ( .A1(n8256), .A2(n8255), .ZN(n10071) );
  INV_X1 U9539 ( .A(n10071), .ZN(n10063) );
  NAND3_X1 U9540 ( .A1(n8482), .A2(n8359), .A3(n8352), .ZN(n8479) );
  OR4_X1 U9541 ( .A1(n8257), .A2(n10063), .A3(n10051), .A4(n8479), .ZN(n8258)
         );
  NOR2_X1 U9542 ( .A1(n10043), .A2(n8258), .ZN(n8259) );
  NAND4_X1 U9543 ( .A1(n9985), .A2(n10025), .A3(n10004), .A4(n8259), .ZN(n8260) );
  OR4_X1 U9544 ( .A1(n9936), .A2(n8283), .A3(n9972), .A4(n8260), .ZN(n8261) );
  NOR2_X1 U9545 ( .A1(n8387), .A2(n8261), .ZN(n8264) );
  INV_X1 U9546 ( .A(n8432), .ZN(n8263) );
  AND4_X1 U9547 ( .A1(n8265), .A2(n8498), .A3(n8264), .A4(n8263), .ZN(n8277)
         );
  MUX2_X1 U9548 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5701), .Z(n8270) );
  INV_X1 U9549 ( .A(SI_31_), .ZN(n8269) );
  XNOR2_X1 U9550 ( .A(n8270), .B(n8269), .ZN(n8271) );
  NAND2_X1 U9551 ( .A1(n9405), .A2(n8273), .ZN(n8276) );
  NAND2_X1 U9552 ( .A1(n8274), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8275) );
  INV_X1 U9553 ( .A(n10199), .ZN(n8403) );
  INV_X1 U9554 ( .A(n8433), .ZN(n9899) );
  INV_X1 U9555 ( .A(n8437), .ZN(n8499) );
  INV_X1 U9556 ( .A(n8439), .ZN(n8445) );
  INV_X1 U9557 ( .A(n8278), .ZN(n8428) );
  INV_X1 U9558 ( .A(n8421), .ZN(n8282) );
  NOR2_X1 U9559 ( .A1(n8283), .A2(n8282), .ZN(n8381) );
  NAND2_X1 U9560 ( .A1(n8374), .A2(n8284), .ZN(n8414) );
  NAND2_X1 U9561 ( .A1(n8481), .A2(n8288), .ZN(n8286) );
  NAND2_X1 U9562 ( .A1(n8352), .A2(n8476), .ZN(n8285) );
  MUX2_X1 U9563 ( .A(n8286), .B(n8285), .S(n8406), .Z(n8355) );
  NAND2_X1 U9564 ( .A1(n8476), .A2(n8472), .ZN(n8289) );
  NAND2_X1 U9565 ( .A1(n8288), .A2(n8287), .ZN(n8478) );
  MUX2_X1 U9566 ( .A(n8289), .B(n8478), .S(n8406), .Z(n8351) );
  INV_X1 U9567 ( .A(n8333), .ZN(n8291) );
  OAI211_X1 U9568 ( .C1(n8291), .C2(n8290), .A(n8341), .B(n8463), .ZN(n8294)
         );
  OAI211_X1 U9569 ( .C1(n8293), .C2(n8292), .A(n8334), .B(n8333), .ZN(n8467)
         );
  MUX2_X1 U9570 ( .A(n8294), .B(n8467), .S(n8400), .Z(n8344) );
  INV_X1 U9571 ( .A(n8298), .ZN(n8312) );
  MUX2_X1 U9572 ( .A(n8451), .B(n8304), .S(n8406), .Z(n8305) );
  INV_X1 U9573 ( .A(n8454), .ZN(n8295) );
  AOI21_X1 U9574 ( .B1(n8296), .B2(n8305), .A(n8295), .ZN(n8301) );
  INV_X1 U9575 ( .A(n8456), .ZN(n8299) );
  OAI21_X1 U9576 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8303) );
  INV_X1 U9577 ( .A(n8308), .ZN(n8302) );
  NAND2_X1 U9578 ( .A1(n8303), .A2(n8302), .ZN(n8311) );
  INV_X1 U9579 ( .A(n8304), .ZN(n8306) );
  OAI211_X1 U9580 ( .C1(n10631), .C2(n8306), .A(n8454), .B(n8305), .ZN(n8307)
         );
  NOR2_X1 U9581 ( .A1(n8307), .A2(n8456), .ZN(n8309) );
  NOR2_X1 U9582 ( .A1(n8309), .A2(n8308), .ZN(n8310) );
  OAI211_X1 U9583 ( .C1(n8312), .C2(n8457), .A(n8317), .B(n8318), .ZN(n8315)
         );
  AOI21_X1 U9584 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8325) );
  NAND2_X1 U9585 ( .A1(n8317), .A2(n8316), .ZN(n8323) );
  AND2_X1 U9586 ( .A1(n8319), .A2(n8318), .ZN(n8322) );
  INV_X1 U9587 ( .A(n8320), .ZN(n8321) );
  AOI21_X1 U9588 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8324) );
  MUX2_X1 U9589 ( .A(n8325), .B(n8324), .S(n8406), .Z(n8332) );
  MUX2_X1 U9590 ( .A(n8327), .B(n8326), .S(n8400), .Z(n8328) );
  OR2_X1 U9591 ( .A1(n8329), .A2(n8328), .ZN(n8330) );
  AOI21_X1 U9592 ( .B1(n8332), .B2(n8331), .A(n8330), .ZN(n8340) );
  OAI211_X1 U9593 ( .C1(n8344), .C2(n5505), .A(n8334), .B(n8338), .ZN(n8337)
         );
  AND2_X1 U9594 ( .A1(n8471), .A2(n8342), .ZN(n8336) );
  INV_X1 U9595 ( .A(n8339), .ZN(n8335) );
  AOI21_X1 U9596 ( .B1(n8337), .B2(n8336), .A(n8335), .ZN(n8348) );
  AND2_X1 U9597 ( .A1(n8339), .A2(n8338), .ZN(n8470) );
  AND2_X1 U9598 ( .A1(n8340), .A2(n8463), .ZN(n8343) );
  AND2_X1 U9599 ( .A1(n8342), .A2(n8341), .ZN(n8447) );
  OAI21_X1 U9600 ( .B1(n8344), .B2(n8343), .A(n8447), .ZN(n8346) );
  AOI21_X1 U9601 ( .B1(n8470), .B2(n8346), .A(n8345), .ZN(n8347) );
  MUX2_X1 U9602 ( .A(n8348), .B(n8347), .S(n8400), .Z(n8350) );
  MUX2_X1 U9603 ( .A(n8481), .B(n8352), .S(n8400), .Z(n8353) );
  NAND2_X1 U9604 ( .A1(n8356), .A2(n8360), .ZN(n8357) );
  NAND3_X1 U9605 ( .A1(n10071), .A2(n8482), .A3(n8357), .ZN(n8358) );
  NAND3_X1 U9606 ( .A1(n8487), .A2(n8362), .A3(n8361), .ZN(n8363) );
  MUX2_X1 U9607 ( .A(n8365), .B(n10042), .S(n8400), .Z(n8366) );
  MUX2_X1 U9608 ( .A(n8368), .B(n8367), .S(n8406), .Z(n8369) );
  NAND2_X1 U9609 ( .A1(n8370), .A2(n10025), .ZN(n8371) );
  NAND2_X1 U9610 ( .A1(n9986), .A2(n8406), .ZN(n8372) );
  NAND2_X1 U9611 ( .A1(n9986), .A2(n8373), .ZN(n8410) );
  NAND3_X1 U9612 ( .A1(n8410), .A2(n8374), .A3(n8400), .ZN(n8375) );
  INV_X1 U9613 ( .A(n9972), .ZN(n8376) );
  NAND3_X1 U9614 ( .A1(n8377), .A2(n8412), .A3(n8376), .ZN(n8380) );
  NAND2_X1 U9615 ( .A1(n8377), .A2(n8409), .ZN(n8378) );
  NAND2_X1 U9616 ( .A1(n8378), .A2(n8415), .ZN(n8379) );
  AOI21_X1 U9617 ( .B1(n8381), .B2(n8383), .A(n9936), .ZN(n8390) );
  INV_X1 U9618 ( .A(n8419), .ZN(n8386) );
  INV_X1 U9619 ( .A(n8426), .ZN(n8385) );
  MUX2_X1 U9620 ( .A(n8386), .B(n8385), .S(n8400), .Z(n8388) );
  AOI211_X1 U9621 ( .C1(n8390), .C2(n8389), .A(n8388), .B(n8387), .ZN(n8391)
         );
  INV_X1 U9622 ( .A(n8392), .ZN(n8431) );
  INV_X1 U9623 ( .A(n8393), .ZN(n8429) );
  AND2_X1 U9624 ( .A1(n9781), .A2(n8433), .ZN(n8396) );
  OAI22_X1 U9625 ( .A1(n8408), .A2(n8405), .B1(n6726), .B2(n7387), .ZN(n8444)
         );
  OAI211_X1 U9626 ( .C1(n4928), .C2(n7387), .A(n6726), .B(n6725), .ZN(n8443)
         );
  INV_X1 U9627 ( .A(n8409), .ZN(n8416) );
  NOR3_X1 U9628 ( .A1(n8416), .A2(n8411), .A3(n8410), .ZN(n8488) );
  INV_X1 U9629 ( .A(n8412), .ZN(n8413) );
  AOI21_X1 U9630 ( .B1(n9986), .B2(n8414), .A(n8413), .ZN(n8417) );
  OAI21_X1 U9631 ( .B1(n8417), .B2(n8416), .A(n8415), .ZN(n8489) );
  AOI21_X1 U9632 ( .B1(n8488), .B2(n8418), .A(n8489), .ZN(n8430) );
  NAND2_X1 U9633 ( .A1(n8420), .A2(n8419), .ZN(n8424) );
  INV_X1 U9634 ( .A(n8424), .ZN(n8423) );
  NAND3_X1 U9635 ( .A1(n8423), .A2(n8422), .A3(n8421), .ZN(n8446) );
  AOI21_X1 U9636 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8427) );
  NOR3_X1 U9637 ( .A1(n8429), .A2(n8428), .A3(n8427), .ZN(n8493) );
  OAI21_X1 U9638 ( .B1(n8430), .B2(n8446), .A(n8493), .ZN(n8435) );
  NOR3_X1 U9639 ( .A1(n8438), .A2(n8437), .A3(n8436), .ZN(n8440) );
  OAI21_X1 U9640 ( .B1(n8440), .B2(n8439), .A(n7387), .ZN(n8442) );
  INV_X1 U9641 ( .A(n8446), .ZN(n8496) );
  INV_X1 U9642 ( .A(n8447), .ZN(n8469) );
  INV_X1 U9643 ( .A(n8448), .ZN(n8460) );
  NAND2_X1 U9644 ( .A1(n6724), .A2(n10616), .ZN(n8449) );
  NAND4_X1 U9645 ( .A1(n8451), .A2(n8450), .A3(n6726), .A4(n8449), .ZN(n8453)
         );
  NAND2_X1 U9646 ( .A1(n8453), .A2(n8452), .ZN(n8455) );
  OAI21_X1 U9647 ( .B1(n10651), .B2(n8455), .A(n8454), .ZN(n8458) );
  AOI21_X1 U9648 ( .B1(n8458), .B2(n8457), .A(n8456), .ZN(n8459) );
  OR3_X1 U9649 ( .A1(n8461), .A2(n8460), .A3(n8459), .ZN(n8462) );
  NAND2_X1 U9650 ( .A1(n8463), .A2(n8462), .ZN(n8465) );
  NOR2_X1 U9651 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  NOR2_X1 U9652 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NOR2_X1 U9653 ( .A1(n8469), .A2(n8468), .ZN(n8474) );
  INV_X1 U9654 ( .A(n8470), .ZN(n8473) );
  OAI211_X1 U9655 ( .C1(n8474), .C2(n8473), .A(n8472), .B(n8471), .ZN(n8475)
         );
  INV_X1 U9656 ( .A(n8475), .ZN(n8477) );
  OAI21_X1 U9657 ( .B1(n8478), .B2(n8477), .A(n8476), .ZN(n8480) );
  AOI21_X1 U9658 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8484) );
  OAI21_X1 U9659 ( .B1(n8484), .B2(n8483), .A(n8482), .ZN(n8486) );
  AOI21_X1 U9660 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8492) );
  INV_X1 U9661 ( .A(n8488), .ZN(n8491) );
  INV_X1 U9662 ( .A(n8489), .ZN(n8490) );
  OAI21_X1 U9663 ( .B1(n8492), .B2(n8491), .A(n8490), .ZN(n8495) );
  INV_X1 U9664 ( .A(n8493), .ZN(n8494) );
  AOI21_X1 U9665 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8501) );
  INV_X1 U9666 ( .A(n8497), .ZN(n8500) );
  OAI211_X1 U9667 ( .C1(n8501), .C2(n8500), .A(n8499), .B(n8498), .ZN(n8502)
         );
  NAND2_X1 U9668 ( .A1(n8502), .A2(n4928), .ZN(n8504) );
  AOI21_X1 U9669 ( .B1(n8504), .B2(n10607), .A(n8509), .ZN(n8503) );
  OAI21_X1 U9670 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8512) );
  NOR3_X1 U9671 ( .A1(n10362), .A2(n8507), .A3(n8506), .ZN(n8511) );
  OAI21_X1 U9672 ( .B1(n8509), .B2(n8508), .A(P1_B_REG_SCAN_IN), .ZN(n8510) );
  OAI22_X1 U9673 ( .A1(n8513), .A2(n8512), .B1(n8511), .B2(n8510), .ZN(
        P1_U3242) );
  NAND2_X1 U9674 ( .A1(n8930), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8514) );
  OAI21_X1 U9675 ( .B1(n8515), .B2(n8930), .A(n8514), .ZN(P2_U3491) );
  OAI222_X1 U9676 ( .A1(n9415), .A2(n8518), .B1(n4925), .B2(n8517), .C1(n8516), 
        .C2(P2_U3151), .ZN(P2_U3271) );
  AOI22_X1 U9677 ( .A1(n10241), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9805), .ZN(n8519) );
  OAI21_X1 U9678 ( .B1(n8520), .B2(n7238), .A(n8519), .ZN(P1_U3354) );
  INV_X1 U9679 ( .A(n8726), .ZN(n8524) );
  NOR2_X1 U9680 ( .A1(n8522), .A2(n9267), .ZN(n9067) );
  AOI21_X1 U9681 ( .B1(n9194), .B2(P2_REG2_REG_29__SCAN_IN), .A(n9067), .ZN(
        n8523) );
  OAI21_X1 U9682 ( .B1(n8524), .B2(n9265), .A(n8523), .ZN(n8525) );
  AOI21_X1 U9683 ( .B1(n8527), .B2(n8526), .A(n8525), .ZN(n8528) );
  OAI21_X1 U9684 ( .B1(n8521), .B2(n9194), .A(n8528), .ZN(P2_U3204) );
  INV_X1 U9685 ( .A(n8529), .ZN(n10240) );
  OAI222_X1 U9686 ( .A1(n9415), .A2(n8722), .B1(n4925), .B2(n10240), .C1(
        P2_U3151), .C2(n6204), .ZN(P2_U3265) );
  XNOR2_X1 U9687 ( .A(n10778), .B(n8574), .ZN(n8534) );
  INV_X1 U9688 ( .A(n8530), .ZN(n8531) );
  XOR2_X1 U9689 ( .A(n9246), .B(n8534), .Z(n8598) );
  XNOR2_X1 U9690 ( .A(n9254), .B(n8574), .ZN(n8535) );
  XNOR2_X1 U9691 ( .A(n8535), .B(n9261), .ZN(n8708) );
  NAND2_X1 U9692 ( .A1(n8707), .A2(n8536), .ZN(n8642) );
  XNOR2_X1 U9693 ( .A(n8840), .B(n8574), .ZN(n8537) );
  XNOR2_X1 U9694 ( .A(n8537), .B(n9247), .ZN(n8643) );
  INV_X1 U9695 ( .A(n8537), .ZN(n8538) );
  XOR2_X1 U9696 ( .A(n8574), .B(n9355), .Z(n8649) );
  XNOR2_X1 U9697 ( .A(n9348), .B(n8574), .ZN(n8540) );
  XNOR2_X1 U9698 ( .A(n8540), .B(n9219), .ZN(n8683) );
  XNOR2_X1 U9699 ( .A(n8740), .B(n8574), .ZN(n8617) );
  INV_X1 U9700 ( .A(n8540), .ZN(n8541) );
  NAND2_X1 U9701 ( .A1(n8541), .A2(n9219), .ZN(n8610) );
  XNOR2_X1 U9702 ( .A(n9177), .B(n8542), .ZN(n8544) );
  NAND2_X1 U9703 ( .A1(n8544), .A2(n9325), .ZN(n8619) );
  INV_X1 U9704 ( .A(n8617), .ZN(n8543) );
  NAND3_X1 U9705 ( .A1(n8619), .A2(n8543), .A3(n9203), .ZN(n8546) );
  INV_X1 U9706 ( .A(n8544), .ZN(n8545) );
  NAND2_X1 U9707 ( .A1(n8545), .A2(n9182), .ZN(n8620) );
  XNOR2_X1 U9708 ( .A(n9385), .B(n8574), .ZN(n8550) );
  XNOR2_X1 U9709 ( .A(n8550), .B(n9336), .ZN(n8621) );
  XNOR2_X1 U9710 ( .A(n9320), .B(n8574), .ZN(n8552) );
  XOR2_X1 U9711 ( .A(n9326), .B(n8552), .Z(n8679) );
  NOR2_X1 U9712 ( .A1(n8552), .A2(n9134), .ZN(n8553) );
  XNOR2_X1 U9713 ( .A(n9137), .B(n8574), .ZN(n8556) );
  INV_X1 U9714 ( .A(n8556), .ZN(n8554) );
  NAND2_X1 U9715 ( .A1(n8555), .A2(n8554), .ZN(n8558) );
  NAND2_X1 U9716 ( .A1(n8557), .A2(n8556), .ZN(n8658) );
  XNOR2_X1 U9717 ( .A(n8873), .B(n8574), .ZN(n8560) );
  NAND2_X1 U9718 ( .A1(n8560), .A2(n9133), .ZN(n8632) );
  INV_X1 U9719 ( .A(n8560), .ZN(n8561) );
  NAND2_X1 U9720 ( .A1(n8561), .A2(n9300), .ZN(n8562) );
  XNOR2_X1 U9721 ( .A(n9301), .B(n8574), .ZN(n8564) );
  NAND2_X1 U9722 ( .A1(n8564), .A2(n9292), .ZN(n8693) );
  INV_X1 U9723 ( .A(n8564), .ZN(n8565) );
  NAND2_X1 U9724 ( .A1(n8565), .A2(n8922), .ZN(n8566) );
  XNOR2_X1 U9725 ( .A(n9295), .B(n8574), .ZN(n8569) );
  XNOR2_X1 U9726 ( .A(n8569), .B(n9103), .ZN(n8694) );
  AND2_X1 U9727 ( .A1(n8635), .A2(n8694), .ZN(n8568) );
  INV_X1 U9728 ( .A(n8694), .ZN(n8567) );
  NAND2_X1 U9729 ( .A1(n8569), .A2(n8570), .ZN(n8571) );
  XNOR2_X1 U9730 ( .A(n9287), .B(n8574), .ZN(n8572) );
  XOR2_X1 U9731 ( .A(n8921), .B(n8572), .Z(n8587) );
  XOR2_X1 U9732 ( .A(n8574), .B(n9073), .Z(n8575) );
  XNOR2_X1 U9733 ( .A(n8576), .B(n8575), .ZN(n8582) );
  INV_X1 U9734 ( .A(n9075), .ZN(n8578) );
  INV_X1 U9735 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8577) );
  OAI22_X1 U9736 ( .A1(n8578), .A2(n8654), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8577), .ZN(n8580) );
  OAI22_X1 U9737 ( .A1(n9279), .A2(n8712), .B1(n9293), .B2(n8700), .ZN(n8579)
         );
  AOI211_X1 U9738 ( .C1(n9281), .C2(n8689), .A(n8580), .B(n8579), .ZN(n8581)
         );
  OAI21_X1 U9739 ( .B1(n8582), .B2(n8691), .A(n8581), .ZN(P2_U3160) );
  INV_X1 U9740 ( .A(n8583), .ZN(n10247) );
  INV_X1 U9741 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8584) );
  OAI222_X1 U9742 ( .A1(n4925), .A2(n10247), .B1(n8585), .B2(P2_U3151), .C1(
        n8584), .C2(n9415), .ZN(P2_U3267) );
  INV_X1 U9743 ( .A(n9287), .ZN(n8595) );
  AOI21_X1 U9744 ( .B1(n8586), .B2(n8587), .A(n8691), .ZN(n8589) );
  NAND2_X1 U9745 ( .A1(n8589), .A2(n8588), .ZN(n8594) );
  INV_X1 U9746 ( .A(n9084), .ZN(n8591) );
  AOI22_X1 U9747 ( .A1(n9103), .A2(n8710), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8590) );
  OAI21_X1 U9748 ( .B1(n8591), .B2(n8654), .A(n8590), .ZN(n8592) );
  AOI21_X1 U9749 ( .B1(n8920), .B2(n8685), .A(n8592), .ZN(n8593) );
  OAI211_X1 U9750 ( .C1(n8595), .C2(n8719), .A(n8594), .B(n8593), .ZN(P2_U3154) );
  AOI21_X1 U9751 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8603) );
  INV_X1 U9752 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10583) );
  OAI22_X1 U9753 ( .A1(n8644), .A2(n8712), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10583), .ZN(n8599) );
  AOI21_X1 U9754 ( .B1(n8710), .B2(n9262), .A(n8599), .ZN(n8600) );
  OAI21_X1 U9755 ( .B1(n9268), .B2(n8654), .A(n8600), .ZN(n8601) );
  AOI21_X1 U9756 ( .B1(n10778), .B2(n8689), .A(n8601), .ZN(n8602) );
  OAI21_X1 U9757 ( .B1(n8603), .B2(n8691), .A(n8602), .ZN(P2_U3155) );
  AOI21_X1 U9758 ( .B1(n9146), .B2(n8604), .A(n4931), .ZN(n8609) );
  AOI22_X1 U9759 ( .A1(n9300), .A2(n8685), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8606) );
  NAND2_X1 U9760 ( .A1(n8715), .A2(n9138), .ZN(n8605) );
  OAI211_X1 U9761 ( .C1(n9134), .C2(n8700), .A(n8606), .B(n8605), .ZN(n8607)
         );
  AOI21_X1 U9762 ( .B1(n9137), .B2(n8689), .A(n8607), .ZN(n8608) );
  OAI21_X1 U9763 ( .B1(n8609), .B2(n8691), .A(n8608), .ZN(P2_U3156) );
  NAND2_X1 U9764 ( .A1(n8611), .A2(n8610), .ZN(n8618) );
  XNOR2_X1 U9765 ( .A(n8618), .B(n8617), .ZN(n8616) );
  NAND2_X1 U9766 ( .A1(n8715), .A2(n9187), .ZN(n8613) );
  NOR2_X1 U9767 ( .A1(n9708), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9055) );
  AOI21_X1 U9768 ( .B1(n8685), .B2(n9325), .A(n9055), .ZN(n8612) );
  OAI211_X1 U9769 ( .C1(n9183), .C2(n8700), .A(n8613), .B(n8612), .ZN(n8614)
         );
  AOI21_X1 U9770 ( .B1(n9186), .B2(n8689), .A(n8614), .ZN(n8615) );
  OAI21_X1 U9771 ( .B1(n8616), .B2(n8691), .A(n8615), .ZN(P2_U3159) );
  INV_X1 U9772 ( .A(n9385), .ZN(n8630) );
  MUX2_X1 U9773 ( .A(n9333), .B(n8618), .S(n8617), .Z(n8668) );
  NAND2_X1 U9774 ( .A1(n8619), .A2(n8620), .ZN(n8669) );
  NOR2_X1 U9775 ( .A1(n8668), .A2(n8669), .ZN(n8667) );
  INV_X1 U9776 ( .A(n8620), .ZN(n8622) );
  NOR3_X1 U9777 ( .A1(n8667), .A2(n8622), .A3(n8621), .ZN(n8625) );
  INV_X1 U9778 ( .A(n8623), .ZN(n8624) );
  OAI21_X1 U9779 ( .B1(n8625), .B2(n8624), .A(n8706), .ZN(n8629) );
  AOI22_X1 U9780 ( .A1(n9326), .A2(n8685), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8626) );
  OAI21_X1 U9781 ( .B1(n9182), .B2(n8700), .A(n8626), .ZN(n8627) );
  AOI21_X1 U9782 ( .B1(n9160), .B2(n8715), .A(n8627), .ZN(n8628) );
  OAI211_X1 U9783 ( .C1(n8630), .C2(n8719), .A(n8629), .B(n8628), .ZN(P2_U3163) );
  INV_X1 U9784 ( .A(n9301), .ZN(n8641) );
  INV_X1 U9785 ( .A(n8631), .ZN(n8661) );
  INV_X1 U9786 ( .A(n8632), .ZN(n8633) );
  NOR3_X1 U9787 ( .A1(n8661), .A2(n8633), .A3(n8635), .ZN(n8636) );
  OAI21_X1 U9788 ( .B1(n8636), .B2(n8696), .A(n8706), .ZN(n8640) );
  AOI22_X1 U9789 ( .A1(n9300), .A2(n8710), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8637) );
  OAI21_X1 U9790 ( .B1(n8570), .B2(n8712), .A(n8637), .ZN(n8638) );
  AOI21_X1 U9791 ( .B1(n9105), .B2(n8715), .A(n8638), .ZN(n8639) );
  OAI211_X1 U9792 ( .C1(n8641), .C2(n8719), .A(n8640), .B(n8639), .ZN(P2_U3165) );
  OAI211_X1 U9793 ( .C1(n8643), .C2(n8642), .A(n5016), .B(n8706), .ZN(n8648)
         );
  NAND2_X1 U9794 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8987) );
  OAI21_X1 U9795 ( .B1(n8644), .B2(n8700), .A(n8987), .ZN(n8646) );
  NOR2_X1 U9796 ( .A1(n8654), .A2(n9235), .ZN(n8645) );
  AOI211_X1 U9797 ( .C1(n8685), .C2(n9232), .A(n8646), .B(n8645), .ZN(n8647)
         );
  OAI211_X1 U9798 ( .C1(n9404), .C2(n8719), .A(n8648), .B(n8647), .ZN(P2_U3166) );
  XNOR2_X1 U9799 ( .A(n8649), .B(n9232), .ZN(n8650) );
  XNOR2_X1 U9800 ( .A(n8651), .B(n8650), .ZN(n8657) );
  AND2_X1 U9801 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9006) );
  NOR2_X1 U9802 ( .A1(n9183), .A2(n8712), .ZN(n8652) );
  AOI211_X1 U9803 ( .C1(n8710), .C2(n9247), .A(n9006), .B(n8652), .ZN(n8653)
         );
  OAI21_X1 U9804 ( .B1(n9223), .B2(n8654), .A(n8653), .ZN(n8655) );
  AOI21_X1 U9805 ( .B1(n9355), .B2(n8689), .A(n8655), .ZN(n8656) );
  OAI21_X1 U9806 ( .B1(n8657), .B2(n8691), .A(n8656), .ZN(P2_U3168) );
  INV_X1 U9807 ( .A(n8658), .ZN(n8660) );
  NOR3_X1 U9808 ( .A1(n4931), .A2(n8660), .A3(n8659), .ZN(n8662) );
  OAI21_X1 U9809 ( .B1(n8662), .B2(n8661), .A(n8706), .ZN(n8666) );
  AOI22_X1 U9810 ( .A1(n9146), .A2(n8710), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8663) );
  OAI21_X1 U9811 ( .B1(n9292), .B2(n8712), .A(n8663), .ZN(n8664) );
  AOI21_X1 U9812 ( .B1(n9122), .B2(n8715), .A(n8664), .ZN(n8665) );
  OAI211_X1 U9813 ( .C1(n9377), .C2(n8719), .A(n8666), .B(n8665), .ZN(P2_U3169) );
  AOI21_X1 U9814 ( .B1(n8669), .B2(n8668), .A(n8667), .ZN(n8674) );
  NAND2_X1 U9815 ( .A1(n8715), .A2(n9172), .ZN(n8671) );
  AOI22_X1 U9816 ( .A1(n9336), .A2(n8685), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8670) );
  OAI211_X1 U9817 ( .C1(n9203), .C2(n8700), .A(n8671), .B(n8670), .ZN(n8672)
         );
  AOI21_X1 U9818 ( .B1(n9177), .B2(n8689), .A(n8672), .ZN(n8673) );
  OAI21_X1 U9819 ( .B1(n8674), .B2(n8691), .A(n8673), .ZN(P2_U3173) );
  AOI22_X1 U9820 ( .A1(n9336), .A2(n8710), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8676) );
  NAND2_X1 U9821 ( .A1(n8715), .A2(n9147), .ZN(n8675) );
  OAI211_X1 U9822 ( .C1(n8559), .C2(n8712), .A(n8676), .B(n8675), .ZN(n8681)
         );
  AOI211_X1 U9823 ( .C1(n8679), .C2(n8678), .A(n8691), .B(n8677), .ZN(n8680)
         );
  AOI211_X1 U9824 ( .C1(n9320), .C2(n8689), .A(n8681), .B(n8680), .ZN(n8682)
         );
  INV_X1 U9825 ( .A(n8682), .ZN(P2_U3175) );
  XNOR2_X1 U9826 ( .A(n8684), .B(n8683), .ZN(n8692) );
  NAND2_X1 U9827 ( .A1(n8715), .A2(n9205), .ZN(n8687) );
  INV_X1 U9828 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9632) );
  NOR2_X1 U9829 ( .A1(n9632), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9036) );
  AOI21_X1 U9830 ( .B1(n8685), .B2(n9333), .A(n9036), .ZN(n8686) );
  OAI211_X1 U9831 ( .C1(n9204), .C2(n8700), .A(n8687), .B(n8686), .ZN(n8688)
         );
  AOI21_X1 U9832 ( .B1(n9348), .B2(n8689), .A(n8688), .ZN(n8690) );
  OAI21_X1 U9833 ( .B1(n8692), .B2(n8691), .A(n8690), .ZN(P2_U3178) );
  INV_X1 U9834 ( .A(n9295), .ZN(n8705) );
  INV_X1 U9835 ( .A(n8693), .ZN(n8695) );
  NOR3_X1 U9836 ( .A1(n8696), .A2(n8695), .A3(n8694), .ZN(n8699) );
  INV_X1 U9837 ( .A(n8697), .ZN(n8698) );
  OAI21_X1 U9838 ( .B1(n8699), .B2(n8698), .A(n8706), .ZN(n8704) );
  INV_X1 U9839 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9745) );
  OAI22_X1 U9840 ( .A1(n9292), .A2(n8700), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9745), .ZN(n8702) );
  NOR2_X1 U9841 ( .A1(n9293), .A2(n8712), .ZN(n8701) );
  AOI211_X1 U9842 ( .C1(n9094), .C2(n8715), .A(n8702), .B(n8701), .ZN(n8703)
         );
  OAI211_X1 U9843 ( .C1(n8705), .C2(n8719), .A(n8704), .B(n8703), .ZN(P2_U3180) );
  INV_X1 U9844 ( .A(n9254), .ZN(n10786) );
  OAI211_X1 U9845 ( .C1(n8709), .C2(n8708), .A(n8707), .B(n8706), .ZN(n8718)
         );
  INV_X1 U9846 ( .A(n9250), .ZN(n8716) );
  NOR2_X1 U9847 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9742), .ZN(n8961) );
  AOI21_X1 U9848 ( .B1(n8710), .B2(n9246), .A(n8961), .ZN(n8711) );
  OAI21_X1 U9849 ( .B1(n8713), .B2(n8712), .A(n8711), .ZN(n8714) );
  AOI21_X1 U9850 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8717) );
  OAI211_X1 U9851 ( .C1(n10786), .C2(n8719), .A(n8718), .B(n8717), .ZN(
        P2_U3181) );
  OR2_X1 U9852 ( .A1(n9279), .A2(n8726), .ZN(n8738) );
  NOR2_X1 U9853 ( .A1(n6274), .A2(n7062), .ZN(n8720) );
  INV_X1 U9854 ( .A(n9366), .ZN(n8733) );
  INV_X1 U9855 ( .A(n9066), .ZN(n8721) );
  INV_X1 U9856 ( .A(n9369), .ZN(n8725) );
  INV_X1 U9857 ( .A(n8919), .ZN(n8724) );
  NAND2_X1 U9858 ( .A1(n8725), .A2(n8724), .ZN(n8903) );
  NAND2_X1 U9859 ( .A1(n8726), .A2(n9279), .ZN(n8727) );
  NAND2_X1 U9860 ( .A1(n8903), .A2(n8727), .ZN(n8899) );
  NAND2_X1 U9861 ( .A1(n8764), .A2(n8729), .ZN(n8730) );
  AOI21_X1 U9862 ( .B1(n8731), .B2(n8738), .A(n8730), .ZN(n8732) );
  INV_X1 U9863 ( .A(n8732), .ZN(n8735) );
  AND2_X1 U9864 ( .A1(n9369), .A2(n8919), .ZN(n8737) );
  NOR2_X1 U9865 ( .A1(n9366), .A2(n9066), .ZN(n8908) );
  NAND2_X1 U9866 ( .A1(n8764), .A2(n8906), .ZN(n8736) );
  INV_X1 U9867 ( .A(n8737), .ZN(n8898) );
  INV_X1 U9868 ( .A(n8899), .ZN(n8763) );
  NAND2_X1 U9869 ( .A1(n8883), .A2(n8884), .ZN(n9089) );
  INV_X1 U9870 ( .A(n9118), .ZN(n9114) );
  INV_X1 U9871 ( .A(n8739), .ZN(n8877) );
  OR2_X1 U9872 ( .A1(n8878), .A2(n8877), .ZN(n8765) );
  INV_X1 U9873 ( .A(n8740), .ZN(n9184) );
  INV_X1 U9874 ( .A(n9244), .ZN(n9242) );
  INV_X1 U9875 ( .A(n8741), .ZN(n8743) );
  NAND4_X1 U9876 ( .A1(n8779), .A2(n8743), .A3(n8742), .A4(n8771), .ZN(n8749)
         );
  NAND2_X1 U9877 ( .A1(n8745), .A2(n8744), .ZN(n8748) );
  NAND2_X1 U9878 ( .A1(n8746), .A2(n8772), .ZN(n8747) );
  NOR3_X1 U9879 ( .A1(n8749), .A2(n8748), .A3(n8747), .ZN(n8750) );
  AND4_X1 U9880 ( .A1(n8752), .A2(n5329), .A3(n8751), .A4(n8750), .ZN(n8753)
         );
  NAND4_X1 U9881 ( .A1(n8819), .A2(n8754), .A3(n6621), .A4(n8753), .ZN(n8755)
         );
  NOR3_X1 U9882 ( .A1(n9259), .A2(n8756), .A3(n8755), .ZN(n8757) );
  NAND4_X1 U9883 ( .A1(n9200), .A2(n9242), .A3(n8757), .A4(n9212), .ZN(n8758)
         );
  INV_X1 U9884 ( .A(n9168), .ZN(n9166) );
  NAND2_X1 U9885 ( .A1(n9127), .A2(n9129), .ZN(n9150) );
  NAND4_X1 U9886 ( .A1(n9135), .A2(n5515), .A3(n9166), .A4(n9150), .ZN(n8759)
         );
  OR4_X1 U9887 ( .A1(n9098), .A2(n9114), .A3(n8765), .A4(n8759), .ZN(n8760) );
  OR2_X1 U9888 ( .A1(n9089), .A2(n8760), .ZN(n8761) );
  NOR2_X1 U9889 ( .A1(n9073), .A2(n8761), .ZN(n8762) );
  NAND4_X1 U9890 ( .A1(n8764), .A2(n8901), .A3(n8763), .A4(n8762), .ZN(n8907)
         );
  INV_X1 U9891 ( .A(n9159), .ZN(n8862) );
  NAND2_X1 U9892 ( .A1(n8767), .A2(n8772), .ZN(n8770) );
  AOI21_X1 U9893 ( .B1(n6617), .B2(n8768), .A(n5034), .ZN(n8769) );
  NAND3_X1 U9894 ( .A1(n8770), .A2(n8769), .A3(n8781), .ZN(n8780) );
  NAND2_X1 U9895 ( .A1(n7223), .A2(n8771), .ZN(n8773) );
  NAND4_X1 U9896 ( .A1(n8775), .A2(n8774), .A3(n8773), .A4(n8772), .ZN(n8776)
         );
  NAND4_X1 U9897 ( .A1(n8777), .A2(n5034), .A3(n8776), .A4(n8785), .ZN(n8778)
         );
  NAND3_X1 U9898 ( .A1(n8780), .A2(n8779), .A3(n8778), .ZN(n8789) );
  INV_X1 U9899 ( .A(n8781), .ZN(n8783) );
  OAI211_X1 U9900 ( .C1(n8789), .C2(n8783), .A(n8790), .B(n8782), .ZN(n8784)
         );
  NAND3_X1 U9901 ( .A1(n8784), .A2(n8794), .A3(n8787), .ZN(n8793) );
  INV_X1 U9902 ( .A(n8785), .ZN(n8788) );
  OAI211_X1 U9903 ( .C1(n8789), .C2(n8788), .A(n8787), .B(n8786), .ZN(n8791)
         );
  NAND3_X1 U9904 ( .A1(n8791), .A2(n8790), .A3(n8795), .ZN(n8792) );
  MUX2_X1 U9905 ( .A(n8795), .B(n8794), .S(n8887), .Z(n8796) );
  AND3_X1 U9906 ( .A1(n8811), .A2(n5329), .A3(n8796), .ZN(n8799) );
  NAND3_X1 U9907 ( .A1(n8800), .A2(n8799), .A3(n8801), .ZN(n8808) );
  INV_X1 U9908 ( .A(n8801), .ZN(n8815) );
  AND2_X1 U9909 ( .A1(n8803), .A2(n8802), .ZN(n8805) );
  NAND2_X1 U9910 ( .A1(n8806), .A2(n8887), .ZN(n8807) );
  INV_X1 U9911 ( .A(n8810), .ZN(n8812) );
  NAND2_X1 U9912 ( .A1(n8812), .A2(n8811), .ZN(n8814) );
  OAI211_X1 U9913 ( .C1(n8815), .C2(n8814), .A(n8813), .B(n5511), .ZN(n8817)
         );
  INV_X1 U9914 ( .A(n8819), .ZN(n8825) );
  NAND2_X1 U9915 ( .A1(n10766), .A2(n8820), .ZN(n8822) );
  MUX2_X1 U9916 ( .A(n8822), .B(n8821), .S(n8887), .Z(n8823) );
  NAND2_X1 U9917 ( .A1(n8828), .A2(n8827), .ZN(n8829) );
  MUX2_X1 U9918 ( .A(n8830), .B(n8829), .S(n8887), .Z(n8831) );
  NAND2_X1 U9919 ( .A1(n8832), .A2(n8831), .ZN(n8836) );
  NOR2_X1 U9920 ( .A1(n9244), .A2(n8834), .ZN(n8835) );
  NAND2_X1 U9921 ( .A1(n8836), .A2(n8835), .ZN(n8839) );
  MUX2_X1 U9922 ( .A(n9211), .B(n8837), .S(n8887), .Z(n8838) );
  NAND2_X1 U9923 ( .A1(n8840), .A2(n5034), .ZN(n8842) );
  OR2_X1 U9924 ( .A1(n8840), .A2(n5034), .ZN(n8841) );
  MUX2_X1 U9925 ( .A(n8842), .B(n8841), .S(n9247), .Z(n8843) );
  MUX2_X1 U9926 ( .A(n9232), .B(n9355), .S(n5034), .Z(n8844) );
  NAND3_X1 U9927 ( .A1(n8848), .A2(n9204), .A3(n8850), .ZN(n8846) );
  NAND3_X1 U9928 ( .A1(n9200), .A2(n8849), .A3(n9355), .ZN(n8845) );
  NAND3_X1 U9929 ( .A1(n8846), .A2(n8845), .A3(n8847), .ZN(n8854) );
  INV_X1 U9930 ( .A(n9355), .ZN(n9222) );
  NAND3_X1 U9931 ( .A1(n8848), .A2(n9222), .A3(n8847), .ZN(n8852) );
  NAND3_X1 U9932 ( .A1(n9200), .A2(n8849), .A3(n9232), .ZN(n8851) );
  NAND3_X1 U9933 ( .A1(n8852), .A2(n8851), .A3(n8850), .ZN(n8853) );
  NAND2_X1 U9934 ( .A1(n9186), .A2(n9203), .ZN(n8856) );
  MUX2_X1 U9935 ( .A(n8856), .B(n8855), .S(n5034), .Z(n8857) );
  NAND2_X1 U9936 ( .A1(n9325), .A2(n8887), .ZN(n8860) );
  NAND2_X1 U9937 ( .A1(n9182), .A2(n5034), .ZN(n8859) );
  MUX2_X1 U9938 ( .A(n8860), .B(n8859), .S(n9177), .Z(n8861) );
  MUX2_X1 U9939 ( .A(n8864), .B(n8863), .S(n5034), .Z(n8865) );
  MUX2_X1 U9940 ( .A(n9326), .B(n9320), .S(n8887), .Z(n8866) );
  OAI21_X1 U9941 ( .B1(n4952), .B2(n9127), .A(n8867), .ZN(n8868) );
  NOR2_X1 U9942 ( .A1(n9137), .A2(n8559), .ZN(n8870) );
  MUX2_X1 U9943 ( .A(n8870), .B(n8869), .S(n8887), .Z(n8871) );
  INV_X1 U9944 ( .A(n8871), .ZN(n8872) );
  NAND2_X1 U9945 ( .A1(n8873), .A2(n9133), .ZN(n8875) );
  MUX2_X1 U9946 ( .A(n8875), .B(n8874), .S(n8887), .Z(n8876) );
  MUX2_X1 U9947 ( .A(n8878), .B(n8877), .S(n8887), .Z(n8879) );
  INV_X1 U9948 ( .A(n8879), .ZN(n8880) );
  MUX2_X1 U9949 ( .A(n9081), .B(n5517), .S(n5034), .Z(n8882) );
  MUX2_X1 U9950 ( .A(n8884), .B(n8883), .S(n5034), .Z(n8885) );
  INV_X1 U9951 ( .A(n8890), .ZN(n8895) );
  NAND2_X1 U9952 ( .A1(n8891), .A2(n8890), .ZN(n8893) );
  MUX2_X1 U9953 ( .A(n8920), .B(n9281), .S(n5034), .Z(n8892) );
  AOI22_X1 U9954 ( .A1(n8895), .A2(n8894), .B1(n8893), .B2(n8892), .ZN(n8897)
         );
  INV_X1 U9955 ( .A(n8903), .ZN(n8904) );
  INV_X1 U9956 ( .A(n8908), .ZN(n8909) );
  XNOR2_X1 U9957 ( .A(n8911), .B(n9056), .ZN(n8918) );
  NAND3_X1 U9958 ( .A1(n8913), .A2(n8912), .A3(n9417), .ZN(n8914) );
  OAI211_X1 U9959 ( .C1(n8915), .C2(n8917), .A(n8914), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8916) );
  OAI21_X1 U9960 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(P2_U3296) );
  MUX2_X1 U9961 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8919), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9962 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8920), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8921), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9964 ( .A(n9103), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8930), .Z(
        P2_U3517) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8922), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9300), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9967 ( .A(n9146), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8930), .Z(
        P2_U3514) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9326), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9336), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9970 ( .A(n9325), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8930), .Z(
        P2_U3511) );
  MUX2_X1 U9971 ( .A(n9333), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8930), .Z(
        P2_U3510) );
  MUX2_X1 U9972 ( .A(n9219), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8930), .Z(
        P2_U3509) );
  MUX2_X1 U9973 ( .A(n9232), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8930), .Z(
        P2_U3508) );
  MUX2_X1 U9974 ( .A(n9247), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8930), .Z(
        P2_U3507) );
  MUX2_X1 U9975 ( .A(n9261), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8930), .Z(
        P2_U3506) );
  MUX2_X1 U9976 ( .A(n9246), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8930), .Z(
        P2_U3505) );
  MUX2_X1 U9977 ( .A(n9262), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8930), .Z(
        P2_U3504) );
  MUX2_X1 U9978 ( .A(n8923), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8930), .Z(
        P2_U3501) );
  MUX2_X1 U9979 ( .A(n8924), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8930), .Z(
        P2_U3500) );
  MUX2_X1 U9980 ( .A(n8925), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8930), .Z(
        P2_U3498) );
  MUX2_X1 U9981 ( .A(n8926), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8930), .Z(
        P2_U3497) );
  MUX2_X1 U9982 ( .A(n8927), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8930), .Z(
        P2_U3496) );
  MUX2_X1 U9983 ( .A(n8928), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8930), .Z(
        P2_U3495) );
  MUX2_X1 U9984 ( .A(n8929), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8930), .Z(
        P2_U3494) );
  MUX2_X1 U9985 ( .A(n6617), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8930), .Z(
        P2_U3493) );
  MUX2_X1 U9986 ( .A(n5475), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8930), .Z(
        P2_U3492) );
  MUX2_X1 U9987 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9417), .Z(n8950) );
  XNOR2_X1 U9988 ( .A(n8950), .B(n8952), .ZN(n8953) );
  XOR2_X1 U9989 ( .A(n8953), .B(n8954), .Z(n8948) );
  NAND2_X1 U9990 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n8936), .ZN(n8957) );
  OAI21_X1 U9991 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8936), .A(n8957), .ZN(
        n8946) );
  AOI21_X1 U9992 ( .B1(n10564), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n8937), .ZN(
        n8944) );
  INV_X1 U9993 ( .A(n8967), .ZN(n8940) );
  XNOR2_X1 U9994 ( .A(n8968), .B(n8940), .ZN(n8941) );
  NAND2_X1 U9995 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n8941), .ZN(n8969) );
  OAI21_X1 U9996 ( .B1(n8941), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8969), .ZN(
        n8942) );
  NAND2_X1 U9997 ( .A1(n10579), .A2(n8942), .ZN(n8943) );
  OAI211_X1 U9998 ( .C1(n9008), .C2(n8968), .A(n8944), .B(n8943), .ZN(n8945)
         );
  AOI21_X1 U9999 ( .B1(n8946), .B2(n10578), .A(n8945), .ZN(n8947) );
  OAI21_X1 U10000 ( .B1(n8948), .B2(n10536), .A(n8947), .ZN(P2_U3195) );
  MUX2_X1 U10001 ( .A(n9251), .B(n8949), .S(n9417), .Z(n8977) );
  XNOR2_X1 U10002 ( .A(n8977), .B(n8991), .ZN(n8979) );
  INV_X1 U10003 ( .A(n8950), .ZN(n8951) );
  MUX2_X1 U10004 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9417), .Z(n8955) );
  XNOR2_X1 U10005 ( .A(n8955), .B(n8965), .ZN(n10573) );
  XOR2_X1 U10006 ( .A(n8979), .B(n8980), .Z(n8976) );
  NAND2_X1 U10007 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8965), .ZN(n8959) );
  AOI22_X1 U10008 ( .A1(n10565), .A2(n6395), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n8965), .ZN(n10572) );
  NAND2_X1 U10009 ( .A1(n8968), .A2(n8956), .ZN(n8958) );
  NAND2_X1 U10010 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8960), .ZN(n8992) );
  OAI21_X1 U10011 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8960), .A(n8992), .ZN(
        n8964) );
  AOI21_X1 U10012 ( .B1(n10564), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8961), .ZN(
        n8962) );
  OAI21_X1 U10013 ( .B1(n9008), .B2(n8991), .A(n8962), .ZN(n8963) );
  AOI21_X1 U10014 ( .B1(n8964), .B2(n10578), .A(n8963), .ZN(n8975) );
  NAND2_X1 U10015 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8965), .ZN(n8971) );
  MUX2_X1 U10016 ( .A(n8966), .B(P2_REG1_REG_14__SCAN_IN), .S(n10565), .Z(
        n10568) );
  NAND2_X1 U10017 ( .A1(n8968), .A2(n8967), .ZN(n8970) );
  NAND2_X1 U10018 ( .A1(n8970), .A2(n8969), .ZN(n10569) );
  NAND2_X1 U10019 ( .A1(n10568), .A2(n10569), .ZN(n10567) );
  NAND2_X1 U10020 ( .A1(n8971), .A2(n10567), .ZN(n8981) );
  XNOR2_X1 U10021 ( .A(n8981), .B(n8978), .ZN(n8972) );
  NAND2_X1 U10022 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8972), .ZN(n8982) );
  OAI21_X1 U10023 ( .B1(n8972), .B2(P2_REG1_REG_15__SCAN_IN), .A(n8982), .ZN(
        n8973) );
  NAND2_X1 U10024 ( .A1(n8973), .A2(n10579), .ZN(n8974) );
  OAI211_X1 U10025 ( .C1(n8976), .C2(n10536), .A(n8975), .B(n8974), .ZN(
        P2_U3197) );
  MUX2_X1 U10026 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9417), .Z(n9001) );
  XNOR2_X1 U10027 ( .A(n9000), .B(n9001), .ZN(n9002) );
  AOI22_X1 U10028 ( .A1(n8980), .A2(n8979), .B1(n8978), .B2(n8977), .ZN(n9003)
         );
  XOR2_X1 U10029 ( .A(n9002), .B(n9003), .Z(n8999) );
  NAND2_X1 U10030 ( .A1(n8991), .A2(n8981), .ZN(n8983) );
  NAND2_X1 U10031 ( .A1(n8983), .A2(n8982), .ZN(n8985) );
  XNOR2_X1 U10032 ( .A(n9012), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U10033 ( .A1(n8984), .A2(n8985), .ZN(n9004) );
  OAI21_X1 U10034 ( .B1(n8985), .B2(n8984), .A(n9004), .ZN(n8989) );
  NAND2_X1 U10035 ( .A1(n10564), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8986) );
  OAI211_X1 U10036 ( .C1(n9008), .C2(n9000), .A(n8987), .B(n8986), .ZN(n8988)
         );
  AOI21_X1 U10037 ( .B1(n8989), .B2(n10579), .A(n8988), .ZN(n8998) );
  AOI22_X1 U10038 ( .A1(n9012), .A2(n9236), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n9000), .ZN(n8995) );
  NAND2_X1 U10039 ( .A1(n8991), .A2(n8990), .ZN(n8993) );
  NAND2_X1 U10040 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  NAND2_X1 U10041 ( .A1(n8995), .A2(n8994), .ZN(n9011) );
  OAI21_X1 U10042 ( .B1(n8995), .B2(n8994), .A(n9011), .ZN(n8996) );
  NAND2_X1 U10043 ( .A1(n8996), .A2(n10578), .ZN(n8997) );
  OAI211_X1 U10044 ( .C1(n8999), .C2(n10536), .A(n8998), .B(n8997), .ZN(
        P2_U3198) );
  MUX2_X1 U10045 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9417), .Z(n9026) );
  XNOR2_X1 U10046 ( .A(n9028), .B(n9026), .ZN(n9029) );
  XOR2_X1 U10047 ( .A(n9029), .B(n9030), .Z(n9017) );
  OAI21_X1 U10048 ( .B1(n9012), .B2(n9360), .A(n9004), .ZN(n9022) );
  XNOR2_X1 U10049 ( .A(n9028), .B(n9022), .ZN(n9005) );
  NAND2_X1 U10050 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n9005), .ZN(n9024) );
  OAI21_X1 U10051 ( .B1(n9005), .B2(P2_REG1_REG_17__SCAN_IN), .A(n9024), .ZN(
        n9010) );
  AOI21_X1 U10052 ( .B1(n10564), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9006), .ZN(
        n9007) );
  OAI21_X1 U10053 ( .B1(n9008), .B2(n9023), .A(n9007), .ZN(n9009) );
  AOI21_X1 U10054 ( .B1(n10579), .B2(n9010), .A(n9009), .ZN(n9016) );
  OAI21_X1 U10055 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9013), .A(n9019), .ZN(
        n9014) );
  NAND2_X1 U10056 ( .A1(n9014), .A2(n10578), .ZN(n9015) );
  OAI211_X1 U10057 ( .C1(n9017), .C2(n10536), .A(n9016), .B(n9015), .ZN(
        P2_U3199) );
  NAND2_X1 U10058 ( .A1(n9023), .A2(n9018), .ZN(n9020) );
  XNOR2_X1 U10059 ( .A(n9052), .B(n9207), .ZN(n9021) );
  XNOR2_X1 U10060 ( .A(n9042), .B(n9021), .ZN(n9039) );
  NAND2_X1 U10061 ( .A1(n9023), .A2(n9022), .ZN(n9025) );
  NAND2_X1 U10062 ( .A1(n9025), .A2(n9024), .ZN(n9046) );
  XNOR2_X1 U10063 ( .A(n9052), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9045) );
  XNOR2_X1 U10064 ( .A(n9046), .B(n9045), .ZN(n9038) );
  INV_X1 U10065 ( .A(n9026), .ZN(n9027) );
  AOI22_X1 U10066 ( .A1(n9030), .A2(n9029), .B1(n9028), .B2(n9027), .ZN(n9032)
         );
  MUX2_X1 U10067 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n9417), .Z(n9031) );
  NOR2_X1 U10068 ( .A1(n9032), .A2(n9031), .ZN(n9050) );
  NAND2_X1 U10069 ( .A1(n9032), .A2(n9031), .ZN(n9051) );
  INV_X1 U10070 ( .A(n9051), .ZN(n9033) );
  AOI21_X1 U10071 ( .B1(n9034), .B2(P2_U3893), .A(n10566), .ZN(n9037) );
  NOR3_X1 U10072 ( .A1(n9034), .A2(n9052), .A3(n10536), .ZN(n9035) );
  MUX2_X1 U10073 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n6461), .S(n9056), .Z(n9049) );
  INV_X1 U10074 ( .A(n9042), .ZN(n9040) );
  OAI21_X1 U10075 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9042), .A(n9041), .ZN(
        n9043) );
  XOR2_X1 U10076 ( .A(n9049), .B(n9043), .Z(n9063) );
  AOI22_X1 U10077 ( .A1(n9046), .A2(n9045), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9044), .ZN(n9047) );
  XNOR2_X1 U10078 ( .A(n9056), .B(n9346), .ZN(n9048) );
  XNOR2_X1 U10079 ( .A(n9047), .B(n9048), .ZN(n9061) );
  MUX2_X1 U10080 ( .A(n9049), .B(n9048), .S(n9417), .Z(n9054) );
  AOI21_X1 U10081 ( .B1(n9052), .B2(n9051), .A(n9050), .ZN(n9053) );
  XOR2_X1 U10082 ( .A(n9054), .B(n9053), .Z(n9059) );
  AOI21_X1 U10083 ( .B1(n10564), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9055), .ZN(
        n9058) );
  NAND2_X1 U10084 ( .A1(n10566), .A2(n9056), .ZN(n9057) );
  OAI211_X1 U10085 ( .C1(n9059), .C2(n10536), .A(n9058), .B(n9057), .ZN(n9060)
         );
  AOI21_X1 U10086 ( .B1(n10579), .B2(n9061), .A(n9060), .ZN(n9062) );
  OAI21_X1 U10087 ( .B1(n9064), .B2(n9063), .A(n9062), .ZN(P2_U3201) );
  NAND2_X1 U10088 ( .A1(n9066), .A2(n9065), .ZN(n9364) );
  INV_X1 U10089 ( .A(n9364), .ZN(n9068) );
  NOR3_X1 U10090 ( .A1(n9068), .A2(n9194), .A3(n9067), .ZN(n9071) );
  NOR2_X1 U10091 ( .A1(n9269), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9069) );
  OAI22_X1 U10092 ( .A1(n9366), .A2(n9265), .B1(n9071), .B2(n9069), .ZN(
        P2_U3202) );
  NOR2_X1 U10093 ( .A1(n9269), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9070) );
  OAI22_X1 U10094 ( .A1(n9369), .A2(n9265), .B1(n9071), .B2(n9070), .ZN(
        P2_U3203) );
  XNOR2_X1 U10095 ( .A(n9072), .B(n9073), .ZN(n9284) );
  XNOR2_X1 U10096 ( .A(n9074), .B(n9073), .ZN(n9278) );
  NAND2_X1 U10097 ( .A1(n9278), .A2(n9170), .ZN(n9080) );
  NOR2_X1 U10098 ( .A1(n9279), .A2(n9093), .ZN(n9078) );
  AOI22_X1 U10099 ( .A1(n9075), .A2(n9188), .B1(n9194), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n9076) );
  OAI21_X1 U10100 ( .B1(n9293), .B2(n9175), .A(n9076), .ZN(n9077) );
  AOI211_X1 U10101 ( .C1(n9281), .C2(n9253), .A(n9078), .B(n9077), .ZN(n9079)
         );
  OAI211_X1 U10102 ( .C1(n9284), .C2(n9274), .A(n9080), .B(n9079), .ZN(
        P2_U3205) );
  NAND2_X1 U10103 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  XOR2_X1 U10104 ( .A(n9083), .B(n9089), .Z(n9291) );
  NOR2_X1 U10105 ( .A1(n9285), .A2(n9093), .ZN(n9087) );
  AOI22_X1 U10106 ( .A1(n9084), .A2(n9188), .B1(n9194), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9085) );
  OAI21_X1 U10107 ( .B1(n8570), .B2(n9175), .A(n9085), .ZN(n9086) );
  AOI211_X1 U10108 ( .C1(n9287), .C2(n9253), .A(n9087), .B(n9086), .ZN(n9091)
         );
  XOR2_X1 U10109 ( .A(n9089), .B(n9088), .Z(n9288) );
  NAND2_X1 U10110 ( .A1(n9288), .A2(n9170), .ZN(n9090) );
  OAI211_X1 U10111 ( .C1(n9291), .C2(n9274), .A(n9091), .B(n9090), .ZN(
        P2_U3206) );
  XNOR2_X1 U10112 ( .A(n9092), .B(n9098), .ZN(n9299) );
  NOR2_X1 U10113 ( .A1(n9293), .A2(n9093), .ZN(n9097) );
  AOI22_X1 U10114 ( .A1(n9094), .A2(n9188), .B1(n9194), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9095) );
  OAI21_X1 U10115 ( .B1(n9292), .B2(n9175), .A(n9095), .ZN(n9096) );
  AOI211_X1 U10116 ( .C1(n9295), .C2(n9253), .A(n9097), .B(n9096), .ZN(n9101)
         );
  XNOR2_X1 U10117 ( .A(n9099), .B(n9098), .ZN(n9296) );
  NAND2_X1 U10118 ( .A1(n9296), .A2(n9170), .ZN(n9100) );
  OAI211_X1 U10119 ( .C1(n9299), .C2(n9274), .A(n9101), .B(n9100), .ZN(
        P2_U3207) );
  XNOR2_X1 U10120 ( .A(n9102), .B(n9107), .ZN(n9104) );
  AOI22_X1 U10121 ( .A1(n9104), .A2(n9340), .B1(n9335), .B2(n9103), .ZN(n9303)
         );
  AOI22_X1 U10122 ( .A1(n9105), .A2(n9188), .B1(n9189), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9106) );
  OAI21_X1 U10123 ( .B1(n9133), .B2(n9175), .A(n9106), .ZN(n9110) );
  XNOR2_X1 U10124 ( .A(n9108), .B(n9107), .ZN(n9304) );
  NOR2_X1 U10125 ( .A1(n9304), .A2(n9274), .ZN(n9109) );
  AOI211_X1 U10126 ( .C1(n9253), .C2(n9301), .A(n9110), .B(n9109), .ZN(n9111)
         );
  OAI21_X1 U10127 ( .B1(n9194), .B2(n9303), .A(n9111), .ZN(P2_U3208) );
  NAND2_X1 U10128 ( .A1(n9113), .A2(n9112), .ZN(n9115) );
  XNOR2_X1 U10129 ( .A(n9115), .B(n9114), .ZN(n9117) );
  OAI22_X1 U10130 ( .A1(n9292), .A2(n9316), .B1(n8559), .B2(n9314), .ZN(n9116)
         );
  AOI21_X1 U10131 ( .B1(n9117), .B2(n9340), .A(n9116), .ZN(n9307) );
  OR2_X1 U10132 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  AND2_X1 U10133 ( .A1(n9121), .A2(n9120), .ZN(n9305) );
  AOI22_X1 U10134 ( .A1(n9122), .A2(n9188), .B1(n9194), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n9123) );
  OAI21_X1 U10135 ( .B1(n9377), .B2(n9265), .A(n9123), .ZN(n9124) );
  AOI21_X1 U10136 ( .B1(n9305), .B2(n9192), .A(n9124), .ZN(n9125) );
  OAI21_X1 U10137 ( .B1(n9307), .B2(n9194), .A(n9125), .ZN(P2_U3209) );
  NAND2_X1 U10138 ( .A1(n9126), .A2(n9159), .ZN(n9144) );
  AND2_X1 U10139 ( .A1(n9143), .A2(n9127), .ZN(n9128) );
  NAND2_X1 U10140 ( .A1(n9144), .A2(n9128), .ZN(n9130) );
  AND2_X1 U10141 ( .A1(n9130), .A2(n9129), .ZN(n9131) );
  XNOR2_X1 U10142 ( .A(n9131), .B(n9135), .ZN(n9132) );
  OAI222_X1 U10143 ( .A1(n9314), .A2(n9134), .B1(n9316), .B2(n9133), .C1(n9132), .C2(n9323), .ZN(n9310) );
  INV_X1 U10144 ( .A(n9310), .ZN(n9142) );
  XNOR2_X1 U10145 ( .A(n9136), .B(n9135), .ZN(n9311) );
  INV_X1 U10146 ( .A(n9137), .ZN(n9381) );
  AOI22_X1 U10147 ( .A1(n9138), .A2(n9188), .B1(n9194), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n9139) );
  OAI21_X1 U10148 ( .B1(n9381), .B2(n9265), .A(n9139), .ZN(n9140) );
  AOI21_X1 U10149 ( .B1(n9311), .B2(n9192), .A(n9140), .ZN(n9141) );
  OAI21_X1 U10150 ( .B1(n9142), .B2(n9194), .A(n9141), .ZN(P2_U3210) );
  NAND2_X1 U10151 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  XNOR2_X1 U10152 ( .A(n9145), .B(n9150), .ZN(n9322) );
  NAND2_X1 U10153 ( .A1(n9146), .A2(n9171), .ZN(n9149) );
  AOI22_X1 U10154 ( .A1(n9189), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9147), .B2(
        n9188), .ZN(n9148) );
  OAI211_X1 U10155 ( .C1(n9315), .C2(n9175), .A(n9149), .B(n9148), .ZN(n9153)
         );
  XNOR2_X1 U10156 ( .A(n9151), .B(n9150), .ZN(n9317) );
  NOR2_X1 U10157 ( .A1(n9317), .A2(n9274), .ZN(n9152) );
  AOI211_X1 U10158 ( .C1(n9253), .C2(n9320), .A(n9153), .B(n9152), .ZN(n9154)
         );
  OAI21_X1 U10159 ( .B1(n9155), .B2(n9322), .A(n9154), .ZN(P2_U3211) );
  NAND2_X1 U10160 ( .A1(n9156), .A2(n9159), .ZN(n9157) );
  NAND2_X1 U10161 ( .A1(n9158), .A2(n9157), .ZN(n9329) );
  XNOR2_X1 U10162 ( .A(n9126), .B(n9159), .ZN(n9324) );
  NAND2_X1 U10163 ( .A1(n9324), .A2(n9170), .ZN(n9165) );
  NAND2_X1 U10164 ( .A1(n9171), .A2(n9326), .ZN(n9162) );
  AOI22_X1 U10165 ( .A1(n9189), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9188), .B2(
        n9160), .ZN(n9161) );
  OAI211_X1 U10166 ( .C1(n9182), .C2(n9175), .A(n9162), .B(n9161), .ZN(n9163)
         );
  AOI21_X1 U10167 ( .B1(n9385), .B2(n9253), .A(n9163), .ZN(n9164) );
  OAI211_X1 U10168 ( .C1(n9329), .C2(n9274), .A(n9165), .B(n9164), .ZN(
        P2_U3212) );
  XNOR2_X1 U10169 ( .A(n9167), .B(n9166), .ZN(n9338) );
  XNOR2_X1 U10170 ( .A(n9169), .B(n9168), .ZN(n9341) );
  NAND2_X1 U10171 ( .A1(n9341), .A2(n9170), .ZN(n9179) );
  NAND2_X1 U10172 ( .A1(n9171), .A2(n9336), .ZN(n9174) );
  AOI22_X1 U10173 ( .A1(n9189), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9188), .B2(
        n9172), .ZN(n9173) );
  OAI211_X1 U10174 ( .C1(n9203), .C2(n9175), .A(n9174), .B(n9173), .ZN(n9176)
         );
  AOI21_X1 U10175 ( .B1(n9177), .B2(n9253), .A(n9176), .ZN(n9178) );
  OAI211_X1 U10176 ( .C1(n9338), .C2(n9274), .A(n9179), .B(n9178), .ZN(
        P2_U3213) );
  XNOR2_X1 U10177 ( .A(n9180), .B(n9184), .ZN(n9181) );
  OAI222_X1 U10178 ( .A1(n9314), .A2(n9183), .B1(n9316), .B2(n9182), .C1(n9323), .C2(n9181), .ZN(n9344) );
  INV_X1 U10179 ( .A(n9344), .ZN(n9195) );
  XNOR2_X1 U10180 ( .A(n9185), .B(n9184), .ZN(n9345) );
  AOI22_X1 U10181 ( .A1(n9189), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9188), .B2(
        n9187), .ZN(n9190) );
  OAI21_X1 U10182 ( .B1(n5324), .B2(n9265), .A(n9190), .ZN(n9191) );
  AOI21_X1 U10183 ( .B1(n9345), .B2(n9192), .A(n9191), .ZN(n9193) );
  OAI21_X1 U10184 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(P2_U3214) );
  AND2_X1 U10185 ( .A1(n9197), .A2(n9196), .ZN(n9199) );
  OAI21_X1 U10186 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n9349) );
  XOR2_X1 U10187 ( .A(n9201), .B(n9200), .Z(n9202) );
  OAI222_X1 U10188 ( .A1(n9314), .A2(n9204), .B1(n9316), .B2(n9203), .C1(n9202), .C2(n9323), .ZN(n9350) );
  NAND2_X1 U10189 ( .A1(n9350), .A2(n9269), .ZN(n9210) );
  INV_X1 U10190 ( .A(n9205), .ZN(n9206) );
  OAI22_X1 U10191 ( .A1(n9269), .A2(n9207), .B1(n9206), .B2(n9267), .ZN(n9208)
         );
  AOI21_X1 U10192 ( .B1(n9348), .B2(n9253), .A(n9208), .ZN(n9209) );
  OAI211_X1 U10193 ( .C1(n9349), .C2(n9274), .A(n9210), .B(n9209), .ZN(
        P2_U3215) );
  NAND2_X1 U10194 ( .A1(n9241), .A2(n9211), .ZN(n9228) );
  NAND2_X1 U10195 ( .A1(n9228), .A2(n9212), .ZN(n9214) );
  NAND2_X1 U10196 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  XOR2_X1 U10197 ( .A(n9215), .B(n9217), .Z(n9357) );
  OAI211_X1 U10198 ( .C1(n9218), .C2(n9217), .A(n9216), .B(n9340), .ZN(n9221)
         );
  AOI22_X1 U10199 ( .A1(n9335), .A2(n9219), .B1(n9247), .B2(n9334), .ZN(n9220)
         );
  NAND2_X1 U10200 ( .A1(n9221), .A2(n9220), .ZN(n9354) );
  NOR2_X1 U10201 ( .A1(n9222), .A2(n9265), .ZN(n9226) );
  OAI22_X1 U10202 ( .A1(n9269), .A2(n9224), .B1(n9223), .B2(n9267), .ZN(n9225)
         );
  AOI211_X1 U10203 ( .C1(n9354), .C2(n9269), .A(n9226), .B(n9225), .ZN(n9227)
         );
  OAI21_X1 U10204 ( .B1(n9274), .B2(n9357), .A(n9227), .ZN(P2_U3216) );
  XNOR2_X1 U10205 ( .A(n9228), .B(n9230), .ZN(n9359) );
  INV_X1 U10206 ( .A(n9359), .ZN(n9240) );
  OAI211_X1 U10207 ( .C1(n9231), .C2(n9230), .A(n9229), .B(n9340), .ZN(n9234)
         );
  AOI22_X1 U10208 ( .A1(n9335), .A2(n9232), .B1(n9261), .B2(n9334), .ZN(n9233)
         );
  NAND2_X1 U10209 ( .A1(n9234), .A2(n9233), .ZN(n9358) );
  NOR2_X1 U10210 ( .A1(n9404), .A2(n9265), .ZN(n9238) );
  OAI22_X1 U10211 ( .A1(n9269), .A2(n9236), .B1(n9235), .B2(n9267), .ZN(n9237)
         );
  AOI211_X1 U10212 ( .C1(n9358), .C2(n9269), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10213 ( .B1(n9274), .B2(n9240), .A(n9239), .ZN(P2_U3217) );
  OAI21_X1 U10214 ( .B1(n4989), .B2(n9242), .A(n9241), .ZN(n10788) );
  OAI211_X1 U10215 ( .C1(n9245), .C2(n9244), .A(n9243), .B(n9340), .ZN(n9249)
         );
  AOI22_X1 U10216 ( .A1(n9335), .A2(n9247), .B1(n9246), .B2(n9334), .ZN(n9248)
         );
  NAND2_X1 U10217 ( .A1(n9249), .A2(n9248), .ZN(n10789) );
  NAND2_X1 U10218 ( .A1(n10789), .A2(n9269), .ZN(n9256) );
  OAI22_X1 U10219 ( .A1(n9269), .A2(n9251), .B1(n9250), .B2(n9267), .ZN(n9252)
         );
  AOI21_X1 U10220 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9255) );
  OAI211_X1 U10221 ( .C1(n9274), .C2(n10788), .A(n9256), .B(n9255), .ZN(
        P2_U3218) );
  XNOR2_X1 U10222 ( .A(n9257), .B(n9259), .ZN(n10776) );
  INV_X1 U10223 ( .A(n10776), .ZN(n9273) );
  OAI211_X1 U10224 ( .C1(n9260), .C2(n9259), .A(n9258), .B(n9340), .ZN(n9264)
         );
  AOI22_X1 U10225 ( .A1(n9334), .A2(n9262), .B1(n9261), .B2(n9335), .ZN(n9263)
         );
  NAND2_X1 U10226 ( .A1(n9264), .A2(n9263), .ZN(n10781) );
  NOR2_X1 U10227 ( .A1(n9266), .A2(n9265), .ZN(n9271) );
  OAI22_X1 U10228 ( .A1(n9269), .A2(n6395), .B1(n9268), .B2(n9267), .ZN(n9270)
         );
  AOI211_X1 U10229 ( .C1(n10781), .C2(n9269), .A(n9271), .B(n9270), .ZN(n9272)
         );
  OAI21_X1 U10230 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(P2_U3219) );
  NOR2_X1 U10231 ( .A1(n9364), .A2(n10782), .ZN(n9276) );
  AOI21_X1 U10232 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10782), .A(n9276), .ZN(
        n9275) );
  OAI21_X1 U10233 ( .B1(n9366), .B2(n9362), .A(n9275), .ZN(P2_U3490) );
  AOI21_X1 U10234 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10782), .A(n9276), .ZN(
        n9277) );
  OAI21_X1 U10235 ( .B1(n9369), .B2(n9362), .A(n9277), .ZN(P2_U3489) );
  NAND2_X1 U10236 ( .A1(n9278), .A2(n9340), .ZN(n9283) );
  OAI22_X1 U10237 ( .A1(n9279), .A2(n9316), .B1(n9293), .B2(n9314), .ZN(n9280)
         );
  AOI21_X1 U10238 ( .B1(n9281), .B2(n10777), .A(n9280), .ZN(n9282) );
  OAI211_X1 U10239 ( .C1(n10787), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9370)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9370), .S(n10791), .Z(
        P2_U3487) );
  OAI22_X1 U10241 ( .A1(n9285), .A2(n9316), .B1(n8570), .B2(n9314), .ZN(n9286)
         );
  AOI21_X1 U10242 ( .B1(n9287), .B2(n10777), .A(n9286), .ZN(n9290) );
  NAND2_X1 U10243 ( .A1(n9288), .A2(n9340), .ZN(n9289) );
  OAI211_X1 U10244 ( .C1(n9291), .C2(n10787), .A(n9290), .B(n9289), .ZN(n9371)
         );
  MUX2_X1 U10245 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9371), .S(n10791), .Z(
        P2_U3486) );
  OAI22_X1 U10246 ( .A1(n9293), .A2(n9316), .B1(n9292), .B2(n9314), .ZN(n9294)
         );
  AOI21_X1 U10247 ( .B1(n9295), .B2(n10777), .A(n9294), .ZN(n9298) );
  NAND2_X1 U10248 ( .A1(n9296), .A2(n9340), .ZN(n9297) );
  OAI211_X1 U10249 ( .C1(n9299), .C2(n10787), .A(n9298), .B(n9297), .ZN(n9372)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9372), .S(n10791), .Z(
        P2_U3485) );
  AOI22_X1 U10251 ( .A1(n9301), .A2(n10777), .B1(n9334), .B2(n9300), .ZN(n9302) );
  OAI211_X1 U10252 ( .C1(n10787), .C2(n9304), .A(n9303), .B(n9302), .ZN(n9373)
         );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9373), .S(n10791), .Z(
        P2_U3484) );
  NAND2_X1 U10254 ( .A1(n9305), .A2(n10775), .ZN(n9306) );
  AND2_X1 U10255 ( .A1(n9307), .A2(n9306), .ZN(n9375) );
  MUX2_X1 U10256 ( .A(n9375), .B(n9308), .S(n10782), .Z(n9309) );
  OAI21_X1 U10257 ( .B1(n9377), .B2(n9362), .A(n9309), .ZN(P2_U3483) );
  AOI21_X1 U10258 ( .B1(n10775), .B2(n9311), .A(n9310), .ZN(n9378) );
  MUX2_X1 U10259 ( .A(n9312), .B(n9378), .S(n10791), .Z(n9313) );
  OAI21_X1 U10260 ( .B1(n9381), .B2(n9362), .A(n9313), .ZN(P2_U3482) );
  OAI22_X1 U10261 ( .A1(n8559), .A2(n9316), .B1(n9315), .B2(n9314), .ZN(n9319)
         );
  NOR2_X1 U10262 ( .A1(n9317), .A2(n10787), .ZN(n9318) );
  AOI211_X1 U10263 ( .C1(n10777), .C2(n9320), .A(n9319), .B(n9318), .ZN(n9321)
         );
  OAI21_X1 U10264 ( .B1(n9323), .B2(n9322), .A(n9321), .ZN(n9382) );
  MUX2_X1 U10265 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9382), .S(n10791), .Z(
        P2_U3481) );
  NAND2_X1 U10266 ( .A1(n9324), .A2(n9340), .ZN(n9328) );
  AOI22_X1 U10267 ( .A1(n9326), .A2(n9335), .B1(n9334), .B2(n9325), .ZN(n9327)
         );
  OAI211_X1 U10268 ( .C1(n10787), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9383)
         );
  MUX2_X1 U10269 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9383), .S(n10791), .Z(
        n9330) );
  AOI21_X1 U10270 ( .B1(n9331), .B2(n9385), .A(n9330), .ZN(n9332) );
  INV_X1 U10271 ( .A(n9332), .ZN(P2_U3480) );
  INV_X1 U10272 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9342) );
  AOI22_X1 U10273 ( .A1(n9336), .A2(n9335), .B1(n9334), .B2(n9333), .ZN(n9337)
         );
  OAI21_X1 U10274 ( .B1(n9338), .B2(n10787), .A(n9337), .ZN(n9339) );
  AOI21_X1 U10275 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(n9388) );
  MUX2_X1 U10276 ( .A(n9342), .B(n9388), .S(n10791), .Z(n9343) );
  OAI21_X1 U10277 ( .B1(n9391), .B2(n9362), .A(n9343), .ZN(P2_U3479) );
  AOI21_X1 U10278 ( .B1(n9345), .B2(n10775), .A(n9344), .ZN(n9392) );
  MUX2_X1 U10279 ( .A(n9346), .B(n9392), .S(n10791), .Z(n9347) );
  OAI21_X1 U10280 ( .B1(n5324), .B2(n9362), .A(n9347), .ZN(P2_U3478) );
  INV_X1 U10281 ( .A(n9348), .ZN(n9398) );
  INV_X1 U10282 ( .A(n9349), .ZN(n9351) );
  AOI21_X1 U10283 ( .B1(n9351), .B2(n10775), .A(n9350), .ZN(n9395) );
  MUX2_X1 U10284 ( .A(n9352), .B(n9395), .S(n10791), .Z(n9353) );
  OAI21_X1 U10285 ( .B1(n9398), .B2(n9362), .A(n9353), .ZN(P2_U3477) );
  AOI21_X1 U10286 ( .B1(n10777), .B2(n9355), .A(n9354), .ZN(n9356) );
  OAI21_X1 U10287 ( .B1(n10787), .B2(n9357), .A(n9356), .ZN(n9399) );
  MUX2_X1 U10288 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9399), .S(n10791), .Z(
        P2_U3476) );
  AOI21_X1 U10289 ( .B1(n9359), .B2(n10775), .A(n9358), .ZN(n9400) );
  MUX2_X1 U10290 ( .A(n9360), .B(n9400), .S(n10791), .Z(n9361) );
  OAI21_X1 U10291 ( .B1(n9404), .B2(n9362), .A(n9361), .ZN(P2_U3475) );
  MUX2_X1 U10292 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9363), .S(n10791), .Z(
        P2_U3459) );
  NOR2_X1 U10293 ( .A1(n9364), .A2(n10792), .ZN(n9367) );
  AOI21_X1 U10294 ( .B1(n10792), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9367), .ZN(
        n9365) );
  OAI21_X1 U10295 ( .B1(n9366), .B2(n9403), .A(n9365), .ZN(P2_U3458) );
  AOI21_X1 U10296 ( .B1(n10792), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9367), .ZN(
        n9368) );
  OAI21_X1 U10297 ( .B1(n9369), .B2(n9403), .A(n9368), .ZN(P2_U3457) );
  MUX2_X1 U10298 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9370), .S(n6696), .Z(
        P2_U3455) );
  MUX2_X1 U10299 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9371), .S(n6696), .Z(
        P2_U3454) );
  MUX2_X1 U10300 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9372), .S(n6696), .Z(
        P2_U3453) );
  MUX2_X1 U10301 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9373), .S(n6696), .Z(
        P2_U3452) );
  INV_X1 U10302 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9374) );
  MUX2_X1 U10303 ( .A(n9375), .B(n9374), .S(n10792), .Z(n9376) );
  OAI21_X1 U10304 ( .B1(n9377), .B2(n9403), .A(n9376), .ZN(P2_U3451) );
  INV_X1 U10305 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9379) );
  MUX2_X1 U10306 ( .A(n9379), .B(n9378), .S(n6696), .Z(n9380) );
  OAI21_X1 U10307 ( .B1(n9381), .B2(n9403), .A(n9380), .ZN(P2_U3450) );
  MUX2_X1 U10308 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9382), .S(n6696), .Z(
        P2_U3449) );
  MUX2_X1 U10309 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9383), .S(n6696), .Z(n9384) );
  AOI21_X1 U10310 ( .B1(n9386), .B2(n9385), .A(n9384), .ZN(n9387) );
  INV_X1 U10311 ( .A(n9387), .ZN(P2_U3448) );
  INV_X1 U10312 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9389) );
  MUX2_X1 U10313 ( .A(n9389), .B(n9388), .S(n6696), .Z(n9390) );
  OAI21_X1 U10314 ( .B1(n9391), .B2(n9403), .A(n9390), .ZN(P2_U3447) );
  MUX2_X1 U10315 ( .A(n9393), .B(n9392), .S(n6696), .Z(n9394) );
  OAI21_X1 U10316 ( .B1(n5324), .B2(n9403), .A(n9394), .ZN(P2_U3446) );
  MUX2_X1 U10317 ( .A(n9396), .B(n9395), .S(n6696), .Z(n9397) );
  OAI21_X1 U10318 ( .B1(n9398), .B2(n9403), .A(n9397), .ZN(P2_U3444) );
  MUX2_X1 U10319 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9399), .S(n6696), .Z(
        P2_U3441) );
  INV_X1 U10320 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9401) );
  MUX2_X1 U10321 ( .A(n9401), .B(n9400), .S(n6696), .Z(n9402) );
  OAI21_X1 U10322 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(P2_U3438) );
  INV_X1 U10323 ( .A(n9405), .ZN(n10237) );
  NOR4_X1 U10324 ( .A1(n5049), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9406), .ZN(n9408) );
  AOI21_X1 U10325 ( .B1(n9409), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9408), .ZN(
        n9410) );
  OAI21_X1 U10326 ( .B1(n10237), .B2(n4925), .A(n9410), .ZN(P2_U3264) );
  INV_X1 U10327 ( .A(n9411), .ZN(n10244) );
  OAI222_X1 U10328 ( .A1(n4925), .A2(n10244), .B1(n6203), .B2(P2_U3151), .C1(
        n9412), .C2(n9415), .ZN(P2_U3266) );
  INV_X1 U10329 ( .A(n9414), .ZN(n10249) );
  OAI222_X1 U10330 ( .A1(n4925), .A2(n10249), .B1(n9417), .B2(P2_U3151), .C1(
        n9416), .C2(n9415), .ZN(P2_U3268) );
  MUX2_X1 U10331 ( .A(n9418), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10332 ( .A(n9419), .ZN(n9515) );
  NAND2_X1 U10333 ( .A1(n9420), .A2(n9515), .ZN(n9424) );
  XNOR2_X1 U10334 ( .A(n9422), .B(n9421), .ZN(n9423) );
  XNOR2_X1 U10335 ( .A(n9424), .B(n9423), .ZN(n9433) );
  OAI22_X1 U10336 ( .A1(n9770), .A2(n9426), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9425), .ZN(n9430) );
  OAI22_X1 U10337 ( .A1(n9774), .A2(n9428), .B1(n9772), .B2(n9427), .ZN(n9429)
         );
  AOI211_X1 U10338 ( .C1(n9431), .C2(n9546), .A(n9430), .B(n9429), .ZN(n9432)
         );
  OAI21_X1 U10339 ( .B1(n9433), .B2(n9541), .A(n9432), .ZN(P1_U3215) );
  INV_X1 U10340 ( .A(n9434), .ZN(n9437) );
  NOR3_X1 U10341 ( .A1(n9528), .A2(n9523), .A3(n9435), .ZN(n9436) );
  OAI21_X1 U10342 ( .B1(n9437), .B2(n9436), .A(n9768), .ZN(n9442) );
  NOR2_X1 U10343 ( .A1(n10126), .A2(n9772), .ZN(n9440) );
  OAI22_X1 U10344 ( .A1(n10007), .A2(n9774), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9438), .ZN(n9439) );
  AOI211_X1 U10345 ( .C1(n10005), .C2(n9762), .A(n9440), .B(n9439), .ZN(n9441)
         );
  OAI211_X1 U10346 ( .C1(n10221), .C2(n9779), .A(n9442), .B(n9441), .ZN(
        P1_U3216) );
  XOR2_X1 U10347 ( .A(n9444), .B(n9443), .Z(n9445) );
  XNOR2_X1 U10348 ( .A(n9446), .B(n9445), .ZN(n9450) );
  NAND2_X1 U10349 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9893) );
  OAI21_X1 U10350 ( .B1(n9772), .B2(n10074), .A(n9893), .ZN(n9448) );
  OAI22_X1 U10351 ( .A1(n10139), .A2(n9770), .B1(n9774), .B2(n10067), .ZN(
        n9447) );
  AOI211_X1 U10352 ( .C1(n10153), .C2(n9546), .A(n9448), .B(n9447), .ZN(n9449)
         );
  OAI21_X1 U10353 ( .B1(n9450), .B2(n9541), .A(n9449), .ZN(P1_U3219) );
  INV_X1 U10354 ( .A(n9451), .ZN(n9452) );
  NOR2_X1 U10355 ( .A1(n9453), .A2(n9452), .ZN(n9458) );
  INV_X1 U10356 ( .A(n9456), .ZN(n9457) );
  AOI21_X1 U10357 ( .B1(n9458), .B2(n9455), .A(n9457), .ZN(n9463) );
  OAI22_X1 U10358 ( .A1(n10139), .A2(n9772), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9459), .ZN(n9461) );
  OAI22_X1 U10359 ( .A1(n10126), .A2(n9770), .B1(n9774), .B2(n10035), .ZN(
        n9460) );
  AOI211_X1 U10360 ( .C1(n10142), .C2(n9546), .A(n9461), .B(n9460), .ZN(n9462)
         );
  OAI21_X1 U10361 ( .B1(n9463), .B2(n9541), .A(n9462), .ZN(P1_U3223) );
  AOI21_X1 U10362 ( .B1(n9464), .B2(n9466), .A(n9465), .ZN(n9473) );
  INV_X1 U10363 ( .A(n9467), .ZN(n9979) );
  AOI22_X1 U10364 ( .A1(n9979), .A2(n9759), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9469) );
  NAND2_X1 U10365 ( .A1(n10005), .A2(n9529), .ZN(n9468) );
  OAI211_X1 U10366 ( .C1(n10103), .C2(n9770), .A(n9469), .B(n9468), .ZN(n9470)
         );
  AOI21_X1 U10367 ( .B1(n9471), .B2(n9546), .A(n9470), .ZN(n9472) );
  OAI21_X1 U10368 ( .B1(n9473), .B2(n9541), .A(n9472), .ZN(P1_U3225) );
  INV_X1 U10369 ( .A(n9475), .ZN(n9476) );
  XNOR2_X1 U10370 ( .A(n9474), .B(n9475), .ZN(n9766) );
  NAND2_X1 U10371 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  OAI21_X1 U10372 ( .B1(n9476), .B2(n9474), .A(n9765), .ZN(n9480) );
  XNOR2_X1 U10373 ( .A(n9478), .B(n9477), .ZN(n9479) );
  XNOR2_X1 U10374 ( .A(n9480), .B(n9479), .ZN(n9485) );
  AOI22_X1 U10375 ( .A1(n9529), .A2(n9789), .B1(n9481), .B2(n9759), .ZN(n9482)
         );
  NAND2_X1 U10376 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9849) );
  OAI211_X1 U10377 ( .C1(n10156), .C2(n9770), .A(n9482), .B(n9849), .ZN(n9483)
         );
  AOI21_X1 U10378 ( .B1(n10171), .B2(n9546), .A(n9483), .ZN(n9484) );
  OAI21_X1 U10379 ( .B1(n9485), .B2(n9541), .A(n9484), .ZN(P1_U3226) );
  XNOR2_X1 U10380 ( .A(n9488), .B(n9487), .ZN(n9489) );
  XNOR2_X1 U10381 ( .A(n9486), .B(n9489), .ZN(n9494) );
  NAND2_X1 U10382 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9877) );
  OAI21_X1 U10383 ( .B1(n9772), .B2(n10163), .A(n9877), .ZN(n9492) );
  OAI22_X1 U10384 ( .A1(n9774), .A2(n9490), .B1(n9770), .B2(n10074), .ZN(n9491) );
  AOI211_X1 U10385 ( .C1(n10166), .C2(n9546), .A(n9492), .B(n9491), .ZN(n9493)
         );
  OAI21_X1 U10386 ( .B1(n9494), .B2(n9541), .A(n9493), .ZN(P1_U3228) );
  AND3_X1 U10387 ( .A1(n9434), .A2(n9496), .A3(n9495), .ZN(n9497) );
  OAI21_X1 U10388 ( .B1(n9498), .B2(n9497), .A(n9768), .ZN(n9503) );
  AOI22_X1 U10389 ( .A1(n9996), .A2(n9759), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9499) );
  OAI21_X1 U10390 ( .B1(n9991), .B2(n9772), .A(n9499), .ZN(n9500) );
  AOI21_X1 U10391 ( .B1(n9501), .B2(n9762), .A(n9500), .ZN(n9502) );
  OAI211_X1 U10392 ( .C1(n10216), .C2(n9779), .A(n9503), .B(n9502), .ZN(
        P1_U3229) );
  INV_X1 U10393 ( .A(n9455), .ZN(n9504) );
  AOI21_X1 U10394 ( .B1(n9506), .B2(n9505), .A(n9504), .ZN(n9512) );
  OAI22_X1 U10395 ( .A1(n10132), .A2(n9770), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9507), .ZN(n9510) );
  INV_X1 U10396 ( .A(n10057), .ZN(n9508) );
  OAI22_X1 U10397 ( .A1(n9774), .A2(n9508), .B1(n10054), .B2(n9772), .ZN(n9509) );
  AOI211_X1 U10398 ( .C1(n10148), .C2(n9546), .A(n9510), .B(n9509), .ZN(n9511)
         );
  OAI21_X1 U10399 ( .B1(n9512), .B2(n9541), .A(n9511), .ZN(P1_U3233) );
  NAND2_X1 U10400 ( .A1(n9515), .A2(n9514), .ZN(n9516) );
  XNOR2_X1 U10401 ( .A(n9513), .B(n9516), .ZN(n9522) );
  NAND2_X1 U10402 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10488)
         );
  OAI21_X1 U10403 ( .B1(n9770), .B2(n9771), .A(n10488), .ZN(n9520) );
  OAI22_X1 U10404 ( .A1(n9774), .A2(n9518), .B1(n9772), .B2(n9517), .ZN(n9519)
         );
  AOI211_X1 U10405 ( .C1(n10180), .C2(n9546), .A(n9520), .B(n9519), .ZN(n9521)
         );
  OAI21_X1 U10406 ( .B1(n9522), .B2(n9541), .A(n9521), .ZN(P1_U3234) );
  INV_X1 U10407 ( .A(n9523), .ZN(n9527) );
  AOI21_X1 U10408 ( .B1(n9527), .B2(n9525), .A(n9524), .ZN(n9526) );
  AOI21_X1 U10409 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9534) );
  NAND2_X1 U10410 ( .A1(n10027), .A2(n9762), .ZN(n9531) );
  AOI22_X1 U10411 ( .A1(n9784), .A2(n9529), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9530) );
  OAI211_X1 U10412 ( .C1(n9774), .C2(n10021), .A(n9531), .B(n9530), .ZN(n9532)
         );
  AOI21_X1 U10413 ( .B1(n10135), .B2(n9546), .A(n9532), .ZN(n9533) );
  OAI21_X1 U10414 ( .B1(n9534), .B2(n9541), .A(n9533), .ZN(P1_U3235) );
  AOI22_X1 U10415 ( .A1(n10088), .A2(n9762), .B1(n10082), .B2(n9759), .ZN(
        n9536) );
  AND2_X1 U10416 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10478) );
  INV_X1 U10417 ( .A(n10478), .ZN(n9535) );
  OAI211_X1 U10418 ( .C1(n10156), .C2(n9772), .A(n9536), .B(n9535), .ZN(n9545)
         );
  INV_X1 U10419 ( .A(n9537), .ZN(n9543) );
  AOI21_X1 U10420 ( .B1(n9539), .B2(n9542), .A(n9538), .ZN(n9540) );
  AOI211_X1 U10421 ( .C1(n9543), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9544)
         );
  AOI211_X1 U10422 ( .C1(n10159), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9753)
         );
  OAI22_X1 U10423 ( .A1(n9742), .A2(keyinput_127), .B1(keyinput_126), .B2(
        P2_REG3_REG_26__SCAN_IN), .ZN(n9547) );
  AOI221_X1 U10424 ( .B1(n9742), .B2(keyinput_127), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_126), .A(n9547), .ZN(n9635) );
  INV_X1 U10425 ( .A(keyinput_124), .ZN(n9633) );
  INV_X1 U10426 ( .A(keyinput_117), .ZN(n9622) );
  AOI22_X1 U10427 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_114), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .ZN(n9548) );
  OAI221_X1 U10428 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_115), .A(n9548), .ZN(n9618) );
  INV_X1 U10429 ( .A(keyinput_113), .ZN(n9616) );
  INV_X1 U10430 ( .A(keyinput_112), .ZN(n9614) );
  INV_X1 U10431 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9723) );
  INV_X1 U10432 ( .A(keyinput_111), .ZN(n9612) );
  INV_X1 U10433 ( .A(keyinput_110), .ZN(n9610) );
  OAI22_X1 U10434 ( .A1(n9708), .A2(keyinput_105), .B1(n9550), .B2(
        keyinput_104), .ZN(n9549) );
  AOI221_X1 U10435 ( .B1(n9708), .B2(keyinput_105), .C1(keyinput_104), .C2(
        n9550), .A(n9549), .ZN(n9608) );
  OAI22_X1 U10436 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_102), .B1(
        keyinput_101), .B2(P2_REG3_REG_14__SCAN_IN), .ZN(n9551) );
  AOI221_X1 U10437 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_101), .A(n9551), .ZN(n9601) );
  OAI22_X1 U10438 ( .A1(P2_U3151), .A2(keyinput_98), .B1(n6294), .B2(
        keyinput_99), .ZN(n9552) );
  AOI221_X1 U10439 ( .B1(P2_U3151), .B2(keyinput_98), .C1(keyinput_99), .C2(
        n6294), .A(n9552), .ZN(n9598) );
  OAI22_X1 U10440 ( .A1(SI_12_), .A2(keyinput_84), .B1(keyinput_86), .B2(
        SI_10_), .ZN(n9553) );
  AOI221_X1 U10441 ( .B1(SI_12_), .B2(keyinput_84), .C1(SI_10_), .C2(
        keyinput_86), .A(n9553), .ZN(n9583) );
  OAI22_X1 U10442 ( .A1(SI_16_), .A2(keyinput_80), .B1(SI_15_), .B2(
        keyinput_81), .ZN(n9554) );
  AOI221_X1 U10443 ( .B1(SI_16_), .B2(keyinput_80), .C1(keyinput_81), .C2(
        SI_15_), .A(n9554), .ZN(n9581) );
  INV_X1 U10444 ( .A(SI_21_), .ZN(n9655) );
  OAI22_X1 U10445 ( .A1(n9655), .A2(keyinput_75), .B1(SI_20_), .B2(keyinput_76), .ZN(n9555) );
  AOI221_X1 U10446 ( .B1(n9655), .B2(keyinput_75), .C1(keyinput_76), .C2(
        SI_20_), .A(n9555), .ZN(n9575) );
  INV_X1 U10447 ( .A(SI_27_), .ZN(n9654) );
  AOI22_X1 U10448 ( .A1(n9557), .A2(keyinput_77), .B1(keyinput_69), .B2(n9654), 
        .ZN(n9556) );
  OAI221_X1 U10449 ( .B1(n9557), .B2(keyinput_77), .C1(n9654), .C2(keyinput_69), .A(n9556), .ZN(n9565) );
  AOI22_X1 U10450 ( .A1(n9559), .A2(keyinput_73), .B1(n9657), .B2(keyinput_71), 
        .ZN(n9558) );
  OAI221_X1 U10451 ( .B1(n9559), .B2(keyinput_73), .C1(n9657), .C2(keyinput_71), .A(n9558), .ZN(n9564) );
  AOI22_X1 U10452 ( .A1(SI_17_), .A2(keyinput_79), .B1(SI_24_), .B2(
        keyinput_72), .ZN(n9560) );
  OAI221_X1 U10453 ( .B1(SI_17_), .B2(keyinput_79), .C1(SI_24_), .C2(
        keyinput_72), .A(n9560), .ZN(n9563) );
  AOI22_X1 U10454 ( .A1(SI_18_), .A2(keyinput_78), .B1(SI_26_), .B2(
        keyinput_70), .ZN(n9561) );
  OAI221_X1 U10455 ( .B1(SI_18_), .B2(keyinput_78), .C1(SI_26_), .C2(
        keyinput_70), .A(n9561), .ZN(n9562) );
  NOR4_X1 U10456 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n9574)
         );
  OAI22_X1 U10457 ( .A1(SI_29_), .A2(keyinput_67), .B1(SI_30_), .B2(
        keyinput_66), .ZN(n9566) );
  AOI221_X1 U10458 ( .B1(SI_29_), .B2(keyinput_67), .C1(keyinput_66), .C2(
        SI_30_), .A(n9566), .ZN(n9569) );
  AOI22_X1 U10459 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n9567) );
  OAI221_X1 U10460 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n9567), .ZN(n9568) );
  AOI22_X1 U10461 ( .A1(keyinput_68), .A2(n9571), .B1(n9569), .B2(n9568), .ZN(
        n9570) );
  OAI21_X1 U10462 ( .B1(n9571), .B2(keyinput_68), .A(n9570), .ZN(n9573) );
  XNOR2_X1 U10463 ( .A(SI_22_), .B(keyinput_74), .ZN(n9572) );
  NAND4_X1 U10464 ( .A1(n9575), .A2(n9574), .A3(n9573), .A4(n9572), .ZN(n9580)
         );
  AOI22_X1 U10465 ( .A1(SI_9_), .A2(keyinput_87), .B1(n9674), .B2(keyinput_83), 
        .ZN(n9576) );
  OAI221_X1 U10466 ( .B1(SI_9_), .B2(keyinput_87), .C1(n9674), .C2(keyinput_83), .A(n9576), .ZN(n9579) );
  AOI22_X1 U10467 ( .A1(SI_11_), .A2(keyinput_85), .B1(SI_14_), .B2(
        keyinput_82), .ZN(n9577) );
  OAI221_X1 U10468 ( .B1(SI_11_), .B2(keyinput_85), .C1(SI_14_), .C2(
        keyinput_82), .A(n9577), .ZN(n9578) );
  AOI211_X1 U10469 ( .C1(n9581), .C2(n9580), .A(n9579), .B(n9578), .ZN(n9582)
         );
  AOI22_X1 U10470 ( .A1(SI_8_), .A2(keyinput_88), .B1(n9583), .B2(n9582), .ZN(
        n9586) );
  AOI22_X1 U10471 ( .A1(SI_6_), .A2(keyinput_90), .B1(SI_7_), .B2(keyinput_89), 
        .ZN(n9584) );
  OAI221_X1 U10472 ( .B1(SI_6_), .B2(keyinput_90), .C1(SI_7_), .C2(keyinput_89), .A(n9584), .ZN(n9585) );
  AOI221_X1 U10473 ( .B1(SI_8_), .B2(n9586), .C1(keyinput_88), .C2(n9586), .A(
        n9585), .ZN(n9590) );
  AOI22_X1 U10474 ( .A1(SI_4_), .A2(keyinput_92), .B1(SI_5_), .B2(keyinput_91), 
        .ZN(n9587) );
  OAI221_X1 U10475 ( .B1(SI_4_), .B2(keyinput_92), .C1(SI_5_), .C2(keyinput_91), .A(n9587), .ZN(n9589) );
  XNOR2_X1 U10476 ( .A(SI_3_), .B(keyinput_93), .ZN(n9588) );
  OAI21_X1 U10477 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9593) );
  XNOR2_X1 U10478 ( .A(n9691), .B(keyinput_95), .ZN(n9592) );
  XNOR2_X1 U10479 ( .A(SI_2_), .B(keyinput_94), .ZN(n9591) );
  NAND3_X1 U10480 ( .A1(n9593), .A2(n9592), .A3(n9591), .ZN(n9596) );
  INV_X1 U10481 ( .A(SI_0_), .ZN(n9697) );
  OAI22_X1 U10482 ( .A1(n5223), .A2(keyinput_97), .B1(n9697), .B2(keyinput_96), 
        .ZN(n9594) );
  AOI221_X1 U10483 ( .B1(n5223), .B2(keyinput_97), .C1(keyinput_96), .C2(n9697), .A(n9594), .ZN(n9595) );
  NAND2_X1 U10484 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  AOI22_X1 U10485 ( .A1(n9598), .A2(n9597), .B1(keyinput_100), .B2(
        P2_REG3_REG_27__SCAN_IN), .ZN(n9599) );
  OAI21_X1 U10486 ( .B1(keyinput_100), .B2(P2_REG3_REG_27__SCAN_IN), .A(n9599), 
        .ZN(n9600) );
  AOI22_X1 U10487 ( .A1(n9601), .A2(n9600), .B1(keyinput_103), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9602) );
  OAI21_X1 U10488 ( .B1(keyinput_103), .B2(P2_REG3_REG_10__SCAN_IN), .A(n9602), 
        .ZN(n9607) );
  AOI22_X1 U10489 ( .A1(n8577), .A2(keyinput_106), .B1(keyinput_108), .B2(
        n7490), .ZN(n9603) );
  OAI221_X1 U10490 ( .B1(n8577), .B2(keyinput_106), .C1(n7490), .C2(
        keyinput_108), .A(n9603), .ZN(n9606) );
  AOI22_X1 U10491 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .ZN(n9604) );
  OAI221_X1 U10492 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_109), .A(n9604), .ZN(n9605) );
  AOI211_X1 U10493 ( .C1(n9608), .C2(n9607), .A(n9606), .B(n9605), .ZN(n9609)
         );
  AOI221_X1 U10494 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n9610), .C1(n9717), 
        .C2(keyinput_110), .A(n9609), .ZN(n9611) );
  AOI221_X1 U10495 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(
        n9720), .C2(n9612), .A(n9611), .ZN(n9613) );
  AOI221_X1 U10496 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(n9614), .C1(n9723), 
        .C2(keyinput_112), .A(n9613), .ZN(n9615) );
  AOI221_X1 U10497 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(n9616), .C1(n6262), .C2(
        keyinput_113), .A(n9615), .ZN(n9617) );
  OAI22_X1 U10498 ( .A1(keyinput_116), .A2(n9620), .B1(n9618), .B2(n9617), 
        .ZN(n9619) );
  AOI21_X1 U10499 ( .B1(keyinput_116), .B2(n9620), .A(n9619), .ZN(n9621) );
  AOI221_X1 U10500 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(n9622), .C1(n6329), .C2(
        keyinput_117), .A(n9621), .ZN(n9630) );
  AOI22_X1 U10501 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_118), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .ZN(n9623) );
  OAI221_X1 U10502 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_119), .A(n9623), .ZN(n9629) );
  OAI22_X1 U10503 ( .A1(n9625), .A2(keyinput_122), .B1(keyinput_120), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n9624) );
  AOI221_X1 U10504 ( .B1(n9625), .B2(keyinput_122), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_120), .A(n9624), .ZN(n9628) );
  OAI22_X1 U10505 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_121), .B1(
        keyinput_123), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n9626) );
  AOI221_X1 U10506 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_123), .A(n9626), .ZN(n9627) );
  OAI211_X1 U10507 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9631)
         );
  OAI221_X1 U10508 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n9633), .C1(n9632), 
        .C2(keyinput_124), .A(n9631), .ZN(n9634) );
  OAI211_X1 U10509 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_125), .A(n9635), 
        .B(n9634), .ZN(n9636) );
  AOI21_X1 U10510 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .A(n9636), 
        .ZN(n9751) );
  INV_X1 U10511 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9638) );
  OAI22_X1 U10512 ( .A1(n9638), .A2(keyinput_55), .B1(n10512), .B2(keyinput_54), .ZN(n9637) );
  AOI221_X1 U10513 ( .B1(n9638), .B2(keyinput_55), .C1(keyinput_54), .C2(
        n10512), .A(n9637), .ZN(n9738) );
  INV_X1 U10514 ( .A(keyinput_53), .ZN(n9731) );
  OAI22_X1 U10515 ( .A1(n9640), .A2(keyinput_51), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(keyinput_50), .ZN(n9639) );
  AOI221_X1 U10516 ( .B1(n9640), .B2(keyinput_51), .C1(keyinput_50), .C2(
        P2_REG3_REG_17__SCAN_IN), .A(n9639), .ZN(n9728) );
  INV_X1 U10517 ( .A(keyinput_49), .ZN(n9726) );
  INV_X1 U10518 ( .A(keyinput_48), .ZN(n9724) );
  INV_X1 U10519 ( .A(keyinput_47), .ZN(n9721) );
  INV_X1 U10520 ( .A(keyinput_46), .ZN(n9718) );
  INV_X1 U10521 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9642) );
  AOI22_X1 U10522 ( .A1(n9642), .A2(keyinput_38), .B1(keyinput_37), .B2(n10583), .ZN(n9641) );
  OAI221_X1 U10523 ( .B1(n9642), .B2(keyinput_38), .C1(n10583), .C2(
        keyinput_37), .A(n9641), .ZN(n9705) );
  AOI22_X1 U10524 ( .A1(P2_U3151), .A2(keyinput_34), .B1(keyinput_35), .B2(
        n6294), .ZN(n9643) );
  OAI221_X1 U10525 ( .B1(P2_U3151), .B2(keyinput_34), .C1(n6294), .C2(
        keyinput_35), .A(n9643), .ZN(n9701) );
  AOI22_X1 U10526 ( .A1(n9646), .A2(keyinput_3), .B1(keyinput_2), .B2(n9645), 
        .ZN(n9644) );
  OAI221_X1 U10527 ( .B1(n9646), .B2(keyinput_3), .C1(n9645), .C2(keyinput_2), 
        .A(n9644), .ZN(n9649) );
  OAI22_X1 U10528 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n9647) );
  AOI221_X1 U10529 ( .B1(SI_31_), .B2(keyinput_1), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n9647), .ZN(n9648) );
  OAI22_X1 U10530 ( .A1(n9649), .A2(n9648), .B1(keyinput_4), .B2(SI_28_), .ZN(
        n9650) );
  AOI21_X1 U10531 ( .B1(keyinput_4), .B2(SI_28_), .A(n9650), .ZN(n9668) );
  XNOR2_X1 U10532 ( .A(SI_23_), .B(keyinput_9), .ZN(n9667) );
  AOI22_X1 U10533 ( .A1(SI_19_), .A2(keyinput_13), .B1(n9652), .B2(keyinput_14), .ZN(n9651) );
  OAI221_X1 U10534 ( .B1(SI_19_), .B2(keyinput_13), .C1(n9652), .C2(
        keyinput_14), .A(n9651), .ZN(n9666) );
  OAI22_X1 U10535 ( .A1(n9655), .A2(keyinput_11), .B1(n9654), .B2(keyinput_5), 
        .ZN(n9653) );
  AOI221_X1 U10536 ( .B1(n9655), .B2(keyinput_11), .C1(keyinput_5), .C2(n9654), 
        .A(n9653), .ZN(n9664) );
  OAI22_X1 U10537 ( .A1(n9658), .A2(keyinput_6), .B1(n9657), .B2(keyinput_7), 
        .ZN(n9656) );
  AOI221_X1 U10538 ( .B1(n9658), .B2(keyinput_6), .C1(keyinput_7), .C2(n9657), 
        .A(n9656), .ZN(n9663) );
  OAI22_X1 U10539 ( .A1(SI_20_), .A2(keyinput_12), .B1(keyinput_15), .B2(
        SI_17_), .ZN(n9659) );
  AOI221_X1 U10540 ( .B1(SI_20_), .B2(keyinput_12), .C1(SI_17_), .C2(
        keyinput_15), .A(n9659), .ZN(n9662) );
  OAI22_X1 U10541 ( .A1(SI_24_), .A2(keyinput_8), .B1(keyinput_10), .B2(SI_22_), .ZN(n9660) );
  AOI221_X1 U10542 ( .B1(SI_24_), .B2(keyinput_8), .C1(SI_22_), .C2(
        keyinput_10), .A(n9660), .ZN(n9661) );
  NAND4_X1 U10543 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9665)
         );
  NOR4_X1 U10544 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n9678)
         );
  AOI22_X1 U10545 ( .A1(SI_15_), .A2(keyinput_17), .B1(SI_16_), .B2(
        keyinput_16), .ZN(n9669) );
  OAI221_X1 U10546 ( .B1(SI_15_), .B2(keyinput_17), .C1(SI_16_), .C2(
        keyinput_16), .A(n9669), .ZN(n9677) );
  OAI22_X1 U10547 ( .A1(n9671), .A2(keyinput_18), .B1(keyinput_22), .B2(SI_10_), .ZN(n9670) );
  AOI221_X1 U10548 ( .B1(n9671), .B2(keyinput_18), .C1(SI_10_), .C2(
        keyinput_22), .A(n9670), .ZN(n9676) );
  INV_X1 U10549 ( .A(SI_12_), .ZN(n9673) );
  OAI22_X1 U10550 ( .A1(n9674), .A2(keyinput_19), .B1(n9673), .B2(keyinput_20), 
        .ZN(n9672) );
  AOI221_X1 U10551 ( .B1(n9674), .B2(keyinput_19), .C1(keyinput_20), .C2(n9673), .A(n9672), .ZN(n9675) );
  OAI211_X1 U10552 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9681)
         );
  AOI22_X1 U10553 ( .A1(SI_9_), .A2(keyinput_23), .B1(SI_11_), .B2(keyinput_21), .ZN(n9679) );
  OAI221_X1 U10554 ( .B1(SI_9_), .B2(keyinput_23), .C1(SI_11_), .C2(
        keyinput_21), .A(n9679), .ZN(n9680) );
  OAI22_X1 U10555 ( .A1(keyinput_24), .A2(n9683), .B1(n9681), .B2(n9680), .ZN(
        n9682) );
  AOI21_X1 U10556 ( .B1(keyinput_24), .B2(n9683), .A(n9682), .ZN(n9689) );
  AOI22_X1 U10557 ( .A1(SI_7_), .A2(keyinput_25), .B1(n9685), .B2(keyinput_26), 
        .ZN(n9684) );
  OAI221_X1 U10558 ( .B1(SI_7_), .B2(keyinput_25), .C1(n9685), .C2(keyinput_26), .A(n9684), .ZN(n9688) );
  OAI22_X1 U10559 ( .A1(SI_5_), .A2(keyinput_27), .B1(SI_4_), .B2(keyinput_28), 
        .ZN(n9686) );
  AOI221_X1 U10560 ( .B1(SI_5_), .B2(keyinput_27), .C1(keyinput_28), .C2(SI_4_), .A(n9686), .ZN(n9687) );
  OAI21_X1 U10561 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9695) );
  INV_X1 U10562 ( .A(keyinput_29), .ZN(n9690) );
  MUX2_X1 U10563 ( .A(n9690), .B(keyinput_29), .S(SI_3_), .Z(n9694) );
  XNOR2_X1 U10564 ( .A(n9691), .B(keyinput_31), .ZN(n9693) );
  XNOR2_X1 U10565 ( .A(SI_2_), .B(keyinput_30), .ZN(n9692) );
  AOI211_X1 U10566 ( .C1(n9695), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9699)
         );
  AOI22_X1 U10567 ( .A1(n9697), .A2(keyinput_32), .B1(n5223), .B2(keyinput_33), 
        .ZN(n9696) );
  OAI221_X1 U10568 ( .B1(n9697), .B2(keyinput_32), .C1(n5223), .C2(keyinput_33), .A(n9696), .ZN(n9698) );
  NOR2_X1 U10569 ( .A1(n9699), .A2(n9698), .ZN(n9700) );
  OAI22_X1 U10570 ( .A1(keyinput_36), .A2(n9703), .B1(n9701), .B2(n9700), .ZN(
        n9702) );
  AOI21_X1 U10571 ( .B1(keyinput_36), .B2(n9703), .A(n9702), .ZN(n9704) );
  OAI22_X1 U10572 ( .A1(n9705), .A2(n9704), .B1(keyinput_39), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9706) );
  AOI21_X1 U10573 ( .B1(keyinput_39), .B2(P2_REG3_REG_10__SCAN_IN), .A(n9706), 
        .ZN(n9715) );
  AOI22_X1 U10574 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(n9708), 
        .B2(keyinput_41), .ZN(n9707) );
  OAI221_X1 U10575 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(n9708), 
        .C2(keyinput_41), .A(n9707), .ZN(n9714) );
  OAI22_X1 U10576 ( .A1(n9710), .A2(keyinput_45), .B1(keyinput_42), .B2(
        P2_REG3_REG_28__SCAN_IN), .ZN(n9709) );
  AOI221_X1 U10577 ( .B1(n9710), .B2(keyinput_45), .C1(P2_REG3_REG_28__SCAN_IN), .C2(keyinput_42), .A(n9709), .ZN(n9713) );
  OAI22_X1 U10578 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(
        keyinput_44), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n9711) );
  AOI221_X1 U10579 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_44), .A(n9711), .ZN(n9712) );
  OAI211_X1 U10580 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9716)
         );
  OAI221_X1 U10581 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n9718), .C1(n9717), 
        .C2(keyinput_46), .A(n9716), .ZN(n9719) );
  OAI221_X1 U10582 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n9721), .C1(n9720), 
        .C2(keyinput_47), .A(n9719), .ZN(n9722) );
  OAI221_X1 U10583 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(n9724), .C1(n9723), 
        .C2(keyinput_48), .A(n9722), .ZN(n9725) );
  OAI221_X1 U10584 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(n6262), 
        .C2(n9726), .A(n9725), .ZN(n9727) );
  AOI22_X1 U10585 ( .A1(n9728), .A2(n9727), .B1(keyinput_52), .B2(
        P2_REG3_REG_4__SCAN_IN), .ZN(n9729) );
  OAI21_X1 U10586 ( .B1(keyinput_52), .B2(P2_REG3_REG_4__SCAN_IN), .A(n9729), 
        .ZN(n9730) );
  OAI221_X1 U10587 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(n9731), .C1(n6329), .C2(
        keyinput_53), .A(n9730), .ZN(n9737) );
  INV_X1 U10588 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9733) );
  AOI22_X1 U10589 ( .A1(n6378), .A2(keyinput_56), .B1(n9733), .B2(keyinput_57), 
        .ZN(n9732) );
  OAI221_X1 U10590 ( .B1(n6378), .B2(keyinput_56), .C1(n9733), .C2(keyinput_57), .A(n9732), .ZN(n9736) );
  AOI22_X1 U10591 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n9734) );
  OAI221_X1 U10592 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n9734), .ZN(n9735) );
  AOI211_X1 U10593 ( .C1(n9738), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9740)
         );
  XNOR2_X1 U10594 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n9739)
         );
  OR2_X1 U10595 ( .A1(n9740), .A2(n9739), .ZN(n9749) );
  INV_X1 U10596 ( .A(keyinput_63), .ZN(n9741) );
  NAND2_X1 U10597 ( .A1(n9741), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9744) );
  AOI22_X1 U10598 ( .A1(n9745), .A2(keyinput_62), .B1(keyinput_63), .B2(n9742), 
        .ZN(n9743) );
  OAI211_X1 U10599 ( .C1(n9745), .C2(keyinput_62), .A(n9744), .B(n9743), .ZN(
        n9746) );
  INV_X1 U10600 ( .A(n9746), .ZN(n9748) );
  XNOR2_X1 U10601 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n9747) );
  NAND3_X1 U10602 ( .A1(n9749), .A2(n9748), .A3(n9747), .ZN(n9750) );
  NOR2_X1 U10603 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  XNOR2_X1 U10604 ( .A(n9753), .B(n9752), .ZN(P1_U3238) );
  OAI21_X1 U10605 ( .B1(n9465), .B2(n9755), .A(n9754), .ZN(n9756) );
  NAND3_X1 U10606 ( .A1(n9757), .A2(n9768), .A3(n9756), .ZN(n9764) );
  INV_X1 U10607 ( .A(n9758), .ZN(n9956) );
  AOI22_X1 U10608 ( .A1(n9956), .A2(n9759), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9760) );
  OAI21_X1 U10609 ( .B1(n10111), .B2(n9772), .A(n9760), .ZN(n9761) );
  AOI21_X1 U10610 ( .B1(n9954), .B2(n9762), .A(n9761), .ZN(n9763) );
  OAI211_X1 U10611 ( .C1(n10211), .C2(n9779), .A(n9764), .B(n9763), .ZN(
        P1_U3240) );
  OAI21_X1 U10612 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9769) );
  NAND2_X1 U10613 ( .A1(n9769), .A2(n9768), .ZN(n9778) );
  NOR2_X1 U10614 ( .A1(n9770), .A2(n10163), .ZN(n9776) );
  OAI22_X1 U10615 ( .A1(n9774), .A2(n9773), .B1(n9772), .B2(n9771), .ZN(n9775)
         );
  AOI211_X1 U10616 ( .C1(P1_REG3_REG_15__SCAN_IN), .C2(P1_U3086), .A(n9776), 
        .B(n9775), .ZN(n9777) );
  OAI211_X1 U10617 ( .C1(n9780), .C2(n9779), .A(n9778), .B(n9777), .ZN(
        P1_U3241) );
  MUX2_X1 U10618 ( .A(n9781), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9799), .Z(
        P1_U3584) );
  MUX2_X1 U10619 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9782), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9954), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10621 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9783), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10622 ( .A(n10005), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9799), .Z(
        P1_U3578) );
  MUX2_X1 U10623 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10045), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10624 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9784), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10625 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9785), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10626 ( .A(n10088), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9799), .Z(
        P1_U3573) );
  MUX2_X1 U10627 ( .A(n9786), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9799), .Z(
        P1_U3572) );
  MUX2_X1 U10628 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9787), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10629 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9788), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10630 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9789), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10631 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9790), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10632 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9791), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10633 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9792), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10634 ( .A(n9793), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9799), .Z(
        P1_U3564) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9794), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10636 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9795), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10637 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9796), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10638 ( .A(n9797), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9799), .Z(
        P1_U3558) );
  MUX2_X1 U10639 ( .A(n9798), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9799), .Z(
        P1_U3557) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5746), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10641 ( .A(n6724), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9799), .Z(
        P1_U3555) );
  MUX2_X1 U10642 ( .A(n6739), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9799), .Z(
        P1_U3554) );
  OAI211_X1 U10643 ( .C1(n9802), .C2(n9801), .A(n10591), .B(n9800), .ZN(n9809)
         );
  OAI211_X1 U10644 ( .C1(n9804), .C2(n9814), .A(n10587), .B(n9803), .ZN(n9808)
         );
  AOI22_X1 U10645 ( .A1(n10585), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9807) );
  NAND2_X1 U10646 ( .A1(n10595), .A2(n9805), .ZN(n9806) );
  NAND4_X1 U10647 ( .A1(n9809), .A2(n9808), .A3(n9807), .A4(n9806), .ZN(
        P1_U3244) );
  INV_X1 U10648 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9811) );
  AOI21_X1 U10649 ( .B1(n10364), .B2(n9811), .A(n9810), .ZN(n10363) );
  INV_X1 U10650 ( .A(n10364), .ZN(n9815) );
  NAND3_X1 U10651 ( .A1(n9812), .A2(n9815), .A3(n7090), .ZN(n9813) );
  OAI211_X1 U10652 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n10245), .ZN(n9816)
         );
  OAI211_X1 U10653 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10363), .A(n9816), .B(
        P1_U3973), .ZN(n10599) );
  INV_X1 U10654 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9818) );
  OAI22_X1 U10655 ( .A1(n10491), .A2(n9818), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9817), .ZN(n9819) );
  AOI21_X1 U10656 ( .B1(n9820), .B2(n10595), .A(n9819), .ZN(n9829) );
  OAI211_X1 U10657 ( .C1(n9823), .C2(n9822), .A(n10591), .B(n9821), .ZN(n9828)
         );
  OAI211_X1 U10658 ( .C1(n9826), .C2(n9825), .A(n10587), .B(n9824), .ZN(n9827)
         );
  NAND4_X1 U10659 ( .A1(n10599), .A2(n9829), .A3(n9828), .A4(n9827), .ZN(
        P1_U3245) );
  INV_X1 U10660 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9831) );
  OAI21_X1 U10661 ( .B1(n10491), .B2(n9831), .A(n9830), .ZN(n9832) );
  AOI21_X1 U10662 ( .B1(n9833), .B2(n10595), .A(n9832), .ZN(n9842) );
  OAI211_X1 U10663 ( .C1(n9836), .C2(n9835), .A(n10587), .B(n9834), .ZN(n9841)
         );
  OAI211_X1 U10664 ( .C1(n9839), .C2(n9838), .A(n10591), .B(n9837), .ZN(n9840)
         );
  NAND3_X1 U10665 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(P1_U3246) );
  INV_X1 U10666 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10667 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n9874), .B1(n9851), .B2(
        n9843), .ZN(n9848) );
  OAI21_X1 U10668 ( .B1(n9855), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9844), .ZN(
        n10481) );
  XNOR2_X1 U10669 ( .A(n10487), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10480) );
  NOR2_X1 U10670 ( .A1(n10481), .A2(n10480), .ZN(n10479) );
  AOI21_X1 U10671 ( .B1(n10487), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10479), 
        .ZN(n10445) );
  XNOR2_X1 U10672 ( .A(n10439), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10446) );
  NOR2_X1 U10673 ( .A1(n10445), .A2(n10446), .ZN(n10444) );
  AOI21_X1 U10674 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10439), .A(n10444), 
        .ZN(n9845) );
  NOR2_X1 U10675 ( .A1(n9845), .A2(n9857), .ZN(n9846) );
  XNOR2_X1 U10676 ( .A(n9857), .B(n9845), .ZN(n10458) );
  NOR2_X1 U10677 ( .A1(n10457), .A2(n10458), .ZN(n10456) );
  NOR2_X1 U10678 ( .A1(n9846), .A2(n10456), .ZN(n9847) );
  NAND2_X1 U10679 ( .A1(n9848), .A2(n9847), .ZN(n9873) );
  OAI21_X1 U10680 ( .B1(n9848), .B2(n9847), .A(n9873), .ZN(n9865) );
  NAND2_X1 U10681 ( .A1(n10585), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9850) );
  OAI211_X1 U10682 ( .C1(n10451), .C2(n9851), .A(n9850), .B(n9849), .ZN(n9864)
         );
  AOI22_X1 U10683 ( .A1(n10487), .A2(n9853), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9852), .ZN(n10483) );
  AOI21_X1 U10684 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10487), .A(n10482), 
        .ZN(n10441) );
  NAND2_X1 U10685 ( .A1(n10439), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9856) );
  OAI21_X1 U10686 ( .B1(n10439), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9856), .ZN(
        n10442) );
  NOR2_X1 U10687 ( .A1(n10441), .A2(n10442), .ZN(n10440) );
  NOR2_X1 U10688 ( .A1(n9858), .A2(n9857), .ZN(n9859) );
  INV_X1 U10689 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U10690 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9874), .ZN(n9860) );
  OAI21_X1 U10691 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9874), .A(n9860), .ZN(
        n9861) );
  NOR2_X1 U10692 ( .A1(n9862), .A2(n9861), .ZN(n9868) );
  AOI211_X1 U10693 ( .C1(n9862), .C2(n9861), .A(n9868), .B(n10496), .ZN(n9863)
         );
  AOI211_X1 U10694 ( .C1(n10591), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9866)
         );
  INV_X1 U10695 ( .A(n9866), .ZN(P1_U3259) );
  NOR2_X1 U10696 ( .A1(n9890), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9867) );
  AOI21_X1 U10697 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9890), .A(n9867), .ZN(
        n9870) );
  AOI21_X1 U10698 ( .B1(n9874), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9868), .ZN(
        n9869) );
  NAND2_X1 U10699 ( .A1(n9870), .A2(n9869), .ZN(n9884) );
  OAI21_X1 U10700 ( .B1(n9870), .B2(n9869), .A(n9884), .ZN(n9871) );
  INV_X1 U10701 ( .A(n9871), .ZN(n9883) );
  INV_X1 U10702 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U10703 ( .A1(n9890), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9872), .B2(
        n9879), .ZN(n9876) );
  OAI21_X1 U10704 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9874), .A(n9873), .ZN(
        n9875) );
  NAND2_X1 U10705 ( .A1(n9876), .A2(n9875), .ZN(n9889) );
  OAI21_X1 U10706 ( .B1(n9876), .B2(n9875), .A(n9889), .ZN(n9881) );
  NAND2_X1 U10707 ( .A1(n10585), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9878) );
  OAI211_X1 U10708 ( .C1(n10451), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9880)
         );
  AOI21_X1 U10709 ( .B1(n9881), .B2(n10591), .A(n9880), .ZN(n9882) );
  OAI21_X1 U10710 ( .B1(n9883), .B2(n10496), .A(n9882), .ZN(P1_U3260) );
  OAI21_X1 U10711 ( .B1(n9890), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9884), .ZN(
        n10474) );
  NAND2_X1 U10712 ( .A1(n10477), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9885) );
  OAI21_X1 U10713 ( .B1(n10477), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9885), .ZN(
        n10473) );
  OR2_X1 U10714 ( .A1(n10474), .A2(n10473), .ZN(n10471) );
  NAND2_X1 U10715 ( .A1(n10471), .A2(n9885), .ZN(n9888) );
  MUX2_X1 U10716 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10068), .S(n9886), .Z(
        n9887) );
  XNOR2_X1 U10717 ( .A(n9888), .B(n9887), .ZN(n9898) );
  OAI21_X1 U10718 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9890), .A(n9889), .ZN(
        n10470) );
  XNOR2_X1 U10719 ( .A(n10477), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10469) );
  NOR2_X1 U10720 ( .A1(n10470), .A2(n10469), .ZN(n10468) );
  AOI21_X1 U10721 ( .B1(n10477), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10468), 
        .ZN(n9892) );
  XNOR2_X1 U10722 ( .A(n7387), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9891) );
  XNOR2_X1 U10723 ( .A(n9892), .B(n9891), .ZN(n9896) );
  NAND2_X1 U10724 ( .A1(n10585), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9894) );
  OAI211_X1 U10725 ( .C1(n10451), .C2(n7387), .A(n9894), .B(n9893), .ZN(n9895)
         );
  AOI21_X1 U10726 ( .B1(n9896), .B2(n10591), .A(n9895), .ZN(n9897) );
  OAI21_X1 U10727 ( .B1(n9898), .B2(n10496), .A(n9897), .ZN(P1_U3262) );
  NAND2_X1 U10728 ( .A1(n10096), .A2(n10674), .ZN(n9902) );
  NOR2_X1 U10729 ( .A1(n9900), .A2(n9899), .ZN(n10095) );
  NOR2_X1 U10730 ( .A1(n10714), .A2(n5140), .ZN(n9909) );
  AOI21_X1 U10731 ( .B1(n10714), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9909), .ZN(
        n9901) );
  OAI211_X1 U10732 ( .C1(n10199), .C2(n10670), .A(n9902), .B(n9901), .ZN(
        P1_U3263) );
  NAND2_X1 U10733 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  NAND2_X1 U10734 ( .A1(n9905), .A2(n10192), .ZN(n9906) );
  NOR2_X1 U10735 ( .A1(n8399), .A2(n10670), .ZN(n9908) );
  AOI211_X1 U10736 ( .C1(n10714), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9909), .B(
        n9908), .ZN(n9910) );
  OAI21_X1 U10737 ( .B1(n10099), .B2(n10010), .A(n9910), .ZN(P1_U3264) );
  NAND2_X1 U10738 ( .A1(n9911), .A2(n10016), .ZN(n9921) );
  INV_X1 U10739 ( .A(n9912), .ZN(n9919) );
  INV_X1 U10740 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9913) );
  OAI22_X1 U10741 ( .A1(n9914), .A2(n10718), .B1(n9913), .B2(n10707), .ZN(
        n9918) );
  NOR2_X1 U10742 ( .A1(n9916), .A2(n9915), .ZN(n9917) );
  AOI211_X1 U10743 ( .C1(n9919), .C2(n10674), .A(n9918), .B(n9917), .ZN(n9920)
         );
  OAI211_X1 U10744 ( .C1(n9922), .C2(n10714), .A(n9921), .B(n9920), .ZN(
        P1_U3356) );
  INV_X1 U10745 ( .A(n9923), .ZN(n9932) );
  AOI22_X1 U10746 ( .A1(n9924), .A2(n10638), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10714), .ZN(n9925) );
  OAI21_X1 U10747 ( .B1(n9926), .B2(n10085), .A(n9925), .ZN(n9927) );
  AOI21_X1 U10748 ( .B1(n9928), .B2(n10081), .A(n9927), .ZN(n9929) );
  OAI21_X1 U10749 ( .B1(n9930), .B2(n10010), .A(n9929), .ZN(n9931) );
  AOI21_X1 U10750 ( .B1(n9932), .B2(n10016), .A(n9931), .ZN(n9933) );
  OAI21_X1 U10751 ( .B1(n10714), .B2(n9934), .A(n9933), .ZN(P1_U3265) );
  XNOR2_X1 U10752 ( .A(n9935), .B(n5310), .ZN(n10106) );
  INV_X1 U10753 ( .A(n10106), .ZN(n9951) );
  AOI21_X1 U10754 ( .B1(n9937), .B2(n9936), .A(n4961), .ZN(n9939) );
  OAI22_X1 U10755 ( .A1(n9939), .A2(n10698), .B1(n9938), .B2(n10703), .ZN(
        n10104) );
  AOI21_X1 U10756 ( .B1(n9947), .B2(n9958), .A(n10660), .ZN(n9942) );
  NAND2_X1 U10757 ( .A1(n9942), .A2(n9941), .ZN(n10102) );
  NAND2_X1 U10758 ( .A1(n10714), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9945) );
  NAND2_X1 U10759 ( .A1(n9943), .A2(n10638), .ZN(n9944) );
  OAI211_X1 U10760 ( .C1(n10103), .C2(n10085), .A(n9945), .B(n9944), .ZN(n9946) );
  AOI21_X1 U10761 ( .B1(n9947), .B2(n10081), .A(n9946), .ZN(n9948) );
  OAI21_X1 U10762 ( .B1(n10102), .B2(n10010), .A(n9948), .ZN(n9949) );
  AOI21_X1 U10763 ( .B1(n10104), .B2(n10707), .A(n9949), .ZN(n9950) );
  OAI21_X1 U10764 ( .B1(n10094), .B2(n9951), .A(n9950), .ZN(P1_U3266) );
  OAI21_X1 U10765 ( .B1(n9964), .B2(n9953), .A(n9952), .ZN(n9955) );
  AOI22_X1 U10766 ( .A1(n9955), .A2(n10659), .B1(n10089), .B2(n9954), .ZN(
        n10110) );
  AOI22_X1 U10767 ( .A1(n9956), .A2(n10638), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10714), .ZN(n9957) );
  OAI21_X1 U10768 ( .B1(n10111), .B2(n10085), .A(n9957), .ZN(n9961) );
  INV_X1 U10769 ( .A(n9968), .ZN(n9959) );
  OAI211_X1 U10770 ( .C1(n10211), .C2(n9959), .A(n10192), .B(n9958), .ZN(
        n10109) );
  NOR2_X1 U10771 ( .A1(n10109), .A2(n10010), .ZN(n9960) );
  AOI211_X1 U10772 ( .C1(n10081), .C2(n9962), .A(n9961), .B(n9960), .ZN(n9966)
         );
  XNOR2_X1 U10773 ( .A(n9963), .B(n9964), .ZN(n10113) );
  NAND2_X1 U10774 ( .A1(n10113), .A2(n10016), .ZN(n9965) );
  OAI211_X1 U10775 ( .C1(n10714), .C2(n10110), .A(n9966), .B(n9965), .ZN(
        P1_U3267) );
  XOR2_X1 U10776 ( .A(n9972), .B(n9967), .Z(n10118) );
  OAI211_X1 U10777 ( .C1(n5142), .C2(n4983), .A(n10192), .B(n9968), .ZN(n10116) );
  INV_X1 U10778 ( .A(n9969), .ZN(n9970) );
  AOI21_X1 U10779 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(n9973) );
  OAI22_X1 U10780 ( .A1(n9973), .A2(n10698), .B1(n10103), .B2(n10703), .ZN(
        n9977) );
  OAI22_X1 U10781 ( .A1(n5142), .A2(n10750), .B1(n9974), .B2(n10701), .ZN(
        n9975) );
  NOR2_X1 U10782 ( .A1(n9977), .A2(n9975), .ZN(n10117) );
  INV_X1 U10783 ( .A(n10117), .ZN(n9976) );
  OAI211_X1 U10784 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n10707), .ZN(n9981)
         );
  AOI22_X1 U10785 ( .A1(n9979), .A2(n10638), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10714), .ZN(n9980) );
  OAI211_X1 U10786 ( .C1(n10116), .C2(n10010), .A(n9981), .B(n9980), .ZN(n9982) );
  INV_X1 U10787 ( .A(n9982), .ZN(n9983) );
  OAI21_X1 U10788 ( .B1(n10118), .B2(n10094), .A(n9983), .ZN(P1_U3268) );
  XNOR2_X1 U10789 ( .A(n9984), .B(n9985), .ZN(n10121) );
  INV_X1 U10790 ( .A(n10121), .ZN(n10001) );
  INV_X1 U10791 ( .A(n9985), .ZN(n9988) );
  NAND2_X1 U10792 ( .A1(n10002), .A2(n9986), .ZN(n9987) );
  NAND2_X1 U10793 ( .A1(n9988), .A2(n9987), .ZN(n9990) );
  NAND3_X1 U10794 ( .A1(n9990), .A2(n10659), .A3(n9989), .ZN(n9994) );
  OAI22_X1 U10795 ( .A1(n10111), .A2(n10703), .B1(n9991), .B2(n10701), .ZN(
        n9992) );
  INV_X1 U10796 ( .A(n9992), .ZN(n9993) );
  NAND2_X1 U10797 ( .A1(n9994), .A2(n9993), .ZN(n10120) );
  AOI211_X1 U10798 ( .C1(n9995), .C2(n4930), .A(n10660), .B(n4983), .ZN(n10119) );
  NAND2_X1 U10799 ( .A1(n10119), .A2(n10674), .ZN(n9998) );
  AOI22_X1 U10800 ( .A1(n9996), .A2(n10638), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10714), .ZN(n9997) );
  OAI211_X1 U10801 ( .C1(n10216), .C2(n10670), .A(n9998), .B(n9997), .ZN(n9999) );
  AOI21_X1 U10802 ( .B1(n10707), .B2(n10120), .A(n9999), .ZN(n10000) );
  OAI21_X1 U10803 ( .B1(n10094), .B2(n10001), .A(n10000), .ZN(P1_U3269) );
  OAI21_X1 U10804 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(n10006) );
  AOI22_X1 U10805 ( .A1(n10006), .A2(n10659), .B1(n10089), .B2(n10005), .ZN(
        n10125) );
  INV_X1 U10806 ( .A(n10007), .ZN(n10008) );
  AOI22_X1 U10807 ( .A1(n10008), .A2(n10638), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10714), .ZN(n10009) );
  OAI21_X1 U10808 ( .B1(n10126), .B2(n10085), .A(n10009), .ZN(n10012) );
  OAI211_X1 U10809 ( .C1(n10221), .C2(n4984), .A(n4930), .B(n10192), .ZN(
        n10124) );
  NOR2_X1 U10810 ( .A1(n10124), .A2(n10010), .ZN(n10011) );
  AOI211_X1 U10811 ( .C1(n10081), .C2(n10013), .A(n10012), .B(n10011), .ZN(
        n10018) );
  XNOR2_X1 U10812 ( .A(n10014), .B(n10015), .ZN(n10128) );
  NAND2_X1 U10813 ( .A1(n10128), .A2(n10016), .ZN(n10017) );
  OAI211_X1 U10814 ( .C1(n10714), .C2(n10125), .A(n10018), .B(n10017), .ZN(
        P1_U3270) );
  XNOR2_X1 U10815 ( .A(n10019), .B(n10025), .ZN(n10138) );
  AOI211_X1 U10816 ( .C1(n10135), .C2(n10034), .A(n10660), .B(n4984), .ZN(
        n10133) );
  NAND2_X1 U10817 ( .A1(n10135), .A2(n10081), .ZN(n10024) );
  INV_X1 U10818 ( .A(n10021), .ZN(n10022) );
  AOI22_X1 U10819 ( .A1(n10022), .A2(n10638), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10714), .ZN(n10023) );
  OAI211_X1 U10820 ( .C1(n10132), .C2(n10085), .A(n10024), .B(n10023), .ZN(
        n10030) );
  XNOR2_X1 U10821 ( .A(n10026), .B(n10025), .ZN(n10028) );
  AOI22_X1 U10822 ( .A1(n10028), .A2(n10659), .B1(n10089), .B2(n10027), .ZN(
        n10136) );
  NOR2_X1 U10823 ( .A1(n10136), .A2(n10714), .ZN(n10029) );
  AOI211_X1 U10824 ( .C1(n10133), .C2(n10674), .A(n10030), .B(n10029), .ZN(
        n10031) );
  OAI21_X1 U10825 ( .B1(n10138), .B2(n10094), .A(n10031), .ZN(P1_U3271) );
  XNOR2_X1 U10826 ( .A(n10032), .B(n10033), .ZN(n10145) );
  AOI211_X1 U10827 ( .C1(n10142), .C2(n10055), .A(n10660), .B(n10020), .ZN(
        n10140) );
  NAND2_X1 U10828 ( .A1(n10142), .A2(n10081), .ZN(n10038) );
  INV_X1 U10829 ( .A(n10035), .ZN(n10036) );
  AOI22_X1 U10830 ( .A1(n10036), .A2(n10638), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10714), .ZN(n10037) );
  OAI211_X1 U10831 ( .C1(n10139), .C2(n10085), .A(n10038), .B(n10037), .ZN(
        n10048) );
  INV_X1 U10832 ( .A(n10039), .ZN(n10040) );
  NOR2_X1 U10833 ( .A1(n10041), .A2(n10040), .ZN(n10052) );
  OAI21_X1 U10834 ( .B1(n10052), .B2(n10051), .A(n10042), .ZN(n10044) );
  XNOR2_X1 U10835 ( .A(n10044), .B(n10043), .ZN(n10046) );
  AOI22_X1 U10836 ( .A1(n10046), .A2(n10659), .B1(n10089), .B2(n10045), .ZN(
        n10143) );
  NOR2_X1 U10837 ( .A1(n10143), .A2(n10714), .ZN(n10047) );
  AOI211_X1 U10838 ( .C1(n10140), .C2(n10674), .A(n10048), .B(n10047), .ZN(
        n10049) );
  OAI21_X1 U10839 ( .B1(n10145), .B2(n10094), .A(n10049), .ZN(P1_U3272) );
  XOR2_X1 U10840 ( .A(n10050), .B(n10051), .Z(n10150) );
  XNOR2_X1 U10841 ( .A(n10052), .B(n10051), .ZN(n10053) );
  OAI222_X1 U10842 ( .A1(n10703), .A2(n10132), .B1(n10701), .B2(n10054), .C1(
        n10698), .C2(n10053), .ZN(n10146) );
  INV_X1 U10843 ( .A(n10055), .ZN(n10056) );
  AOI211_X1 U10844 ( .C1(n10148), .C2(n5151), .A(n10660), .B(n10056), .ZN(
        n10147) );
  NAND2_X1 U10845 ( .A1(n10147), .A2(n10674), .ZN(n10059) );
  AOI22_X1 U10846 ( .A1(n10057), .A2(n10638), .B1(n10714), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n10058) );
  OAI211_X1 U10847 ( .C1(n10060), .C2(n10670), .A(n10059), .B(n10058), .ZN(
        n10061) );
  AOI21_X1 U10848 ( .B1(n10146), .B2(n10707), .A(n10061), .ZN(n10062) );
  OAI21_X1 U10849 ( .B1(n10150), .B2(n10094), .A(n10062), .ZN(P1_U3273) );
  XNOR2_X1 U10850 ( .A(n10064), .B(n10063), .ZN(n10155) );
  AOI211_X1 U10851 ( .C1(n10153), .C2(n10078), .A(n10660), .B(n10065), .ZN(
        n10152) );
  INV_X1 U10852 ( .A(n10153), .ZN(n10066) );
  NOR2_X1 U10853 ( .A1(n10066), .A2(n10670), .ZN(n10070) );
  OAI22_X1 U10854 ( .A1(n10068), .A2(n10707), .B1(n10067), .B2(n10718), .ZN(
        n10069) );
  AOI211_X1 U10855 ( .C1(n10152), .C2(n10674), .A(n10070), .B(n10069), .ZN(
        n10076) );
  XNOR2_X1 U10856 ( .A(n10072), .B(n10071), .ZN(n10073) );
  OAI222_X1 U10857 ( .A1(n10703), .A2(n10139), .B1(n10701), .B2(n10074), .C1(
        n10073), .C2(n10698), .ZN(n10151) );
  NAND2_X1 U10858 ( .A1(n10151), .A2(n10707), .ZN(n10075) );
  OAI211_X1 U10859 ( .C1(n10155), .C2(n10094), .A(n10076), .B(n10075), .ZN(
        P1_U3274) );
  XOR2_X1 U10860 ( .A(n10077), .B(n10086), .Z(n10162) );
  INV_X1 U10861 ( .A(n10078), .ZN(n10079) );
  AOI211_X1 U10862 ( .C1(n10159), .C2(n10080), .A(n10660), .B(n10079), .ZN(
        n10157) );
  NAND2_X1 U10863 ( .A1(n10159), .A2(n10081), .ZN(n10084) );
  AOI22_X1 U10864 ( .A1(n10714), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10082), 
        .B2(n10638), .ZN(n10083) );
  OAI211_X1 U10865 ( .C1(n10156), .C2(n10085), .A(n10084), .B(n10083), .ZN(
        n10092) );
  XOR2_X1 U10866 ( .A(n10087), .B(n10086), .Z(n10090) );
  AOI22_X1 U10867 ( .A1(n10090), .A2(n10659), .B1(n10089), .B2(n10088), .ZN(
        n10161) );
  NOR2_X1 U10868 ( .A1(n10161), .A2(n10714), .ZN(n10091) );
  AOI211_X1 U10869 ( .C1(n10157), .C2(n10674), .A(n10092), .B(n10091), .ZN(
        n10093) );
  OAI21_X1 U10870 ( .B1(n10162), .B2(n10094), .A(n10093), .ZN(P1_U3275) );
  MUX2_X1 U10871 ( .A(n10097), .B(n10196), .S(n10757), .Z(n10098) );
  OAI21_X1 U10872 ( .B1(n10199), .B2(n10131), .A(n10098), .ZN(P1_U3553) );
  NAND2_X1 U10873 ( .A1(n10099), .A2(n5140), .ZN(n10200) );
  MUX2_X1 U10874 ( .A(n10200), .B(P1_REG1_REG_30__SCAN_IN), .S(n10756), .Z(
        n10100) );
  INV_X1 U10875 ( .A(n10100), .ZN(n10101) );
  OAI21_X1 U10876 ( .B1(n8399), .B2(n10131), .A(n10101), .ZN(P1_U3552) );
  OAI21_X1 U10877 ( .B1(n10103), .B2(n10701), .A(n10102), .ZN(n10105) );
  AOI211_X1 U10878 ( .C1(n10106), .C2(n10754), .A(n10105), .B(n10104), .ZN(
        n10204) );
  MUX2_X1 U10879 ( .A(n10107), .B(n10204), .S(n10757), .Z(n10108) );
  OAI21_X1 U10880 ( .B1(n10207), .B2(n10131), .A(n10108), .ZN(P1_U3549) );
  OAI211_X1 U10881 ( .C1(n10111), .C2(n10701), .A(n10110), .B(n10109), .ZN(
        n10112) );
  AOI21_X1 U10882 ( .B1(n10113), .B2(n10754), .A(n10112), .ZN(n10208) );
  MUX2_X1 U10883 ( .A(n10114), .B(n10208), .S(n10757), .Z(n10115) );
  OAI21_X1 U10884 ( .B1(n10211), .B2(n10131), .A(n10115), .ZN(P1_U3548) );
  OAI211_X1 U10885 ( .C1(n10183), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        n10212) );
  MUX2_X1 U10886 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10212), .S(n10757), .Z(
        P1_U3547) );
  AOI211_X1 U10887 ( .C1(n10121), .C2(n10754), .A(n10120), .B(n10119), .ZN(
        n10213) );
  MUX2_X1 U10888 ( .A(n10122), .B(n10213), .S(n10757), .Z(n10123) );
  OAI21_X1 U10889 ( .B1(n10216), .B2(n10131), .A(n10123), .ZN(P1_U3546) );
  OAI211_X1 U10890 ( .C1(n10126), .C2(n10701), .A(n10125), .B(n10124), .ZN(
        n10127) );
  AOI21_X1 U10891 ( .B1(n10754), .B2(n10128), .A(n10127), .ZN(n10217) );
  MUX2_X1 U10892 ( .A(n10129), .B(n10217), .S(n10757), .Z(n10130) );
  OAI21_X1 U10893 ( .B1(n10221), .B2(n10131), .A(n10130), .ZN(P1_U3545) );
  NOR2_X1 U10894 ( .A1(n10132), .A2(n10701), .ZN(n10134) );
  AOI211_X1 U10895 ( .C1(n10663), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10137) );
  OAI211_X1 U10896 ( .C1(n10183), .C2(n10138), .A(n10137), .B(n10136), .ZN(
        n10222) );
  MUX2_X1 U10897 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10222), .S(n10757), .Z(
        P1_U3544) );
  NOR2_X1 U10898 ( .A1(n10139), .A2(n10701), .ZN(n10141) );
  AOI211_X1 U10899 ( .C1(n10663), .C2(n10142), .A(n10141), .B(n10140), .ZN(
        n10144) );
  OAI211_X1 U10900 ( .C1(n10183), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10223) );
  MUX2_X1 U10901 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10223), .S(n10757), .Z(
        P1_U3543) );
  AOI211_X1 U10902 ( .C1(n10663), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10149) );
  OAI21_X1 U10903 ( .B1(n10183), .B2(n10150), .A(n10149), .ZN(n10224) );
  MUX2_X1 U10904 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10224), .S(n10757), .Z(
        P1_U3542) );
  AOI211_X1 U10905 ( .C1(n10663), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10154) );
  OAI21_X1 U10906 ( .B1(n10183), .B2(n10155), .A(n10154), .ZN(n10225) );
  MUX2_X1 U10907 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10225), .S(n10757), .Z(
        P1_U3541) );
  NOR2_X1 U10908 ( .A1(n10156), .A2(n10701), .ZN(n10158) );
  AOI211_X1 U10909 ( .C1(n10663), .C2(n10159), .A(n10158), .B(n10157), .ZN(
        n10160) );
  OAI211_X1 U10910 ( .C1(n10162), .C2(n10183), .A(n10161), .B(n10160), .ZN(
        n10226) );
  MUX2_X1 U10911 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10226), .S(n10757), .Z(
        P1_U3540) );
  NOR2_X1 U10912 ( .A1(n10163), .A2(n10701), .ZN(n10165) );
  AOI211_X1 U10913 ( .C1(n10663), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        n10167) );
  OAI211_X1 U10914 ( .C1(n10169), .C2(n10183), .A(n10168), .B(n10167), .ZN(
        n10227) );
  MUX2_X1 U10915 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10227), .S(n10757), .Z(
        P1_U3539) );
  AOI21_X1 U10916 ( .B1(n10663), .B2(n10171), .A(n10170), .ZN(n10175) );
  NAND3_X1 U10917 ( .A1(n8140), .A2(n10754), .A3(n10172), .ZN(n10173) );
  NAND3_X1 U10918 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n10228) );
  MUX2_X1 U10919 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10228), .S(n10757), .Z(
        P1_U3538) );
  OAI211_X1 U10920 ( .C1(n10183), .C2(n10178), .A(n10177), .B(n10176), .ZN(
        n10229) );
  MUX2_X1 U10921 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10229), .S(n10757), .Z(
        P1_U3537) );
  AOI21_X1 U10922 ( .B1(n10663), .B2(n10180), .A(n10179), .ZN(n10181) );
  OAI211_X1 U10923 ( .C1(n10184), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        n10230) );
  MUX2_X1 U10924 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10230), .S(n10757), .Z(
        P1_U3535) );
  XOR2_X1 U10925 ( .A(n10187), .B(n10185), .Z(n10618) );
  XNOR2_X1 U10926 ( .A(n10187), .B(n10186), .ZN(n10191) );
  OAI22_X1 U10927 ( .A1(n10188), .A2(n10701), .B1(n10653), .B2(n10703), .ZN(
        n10190) );
  NOR2_X1 U10928 ( .A1(n10618), .A2(n10655), .ZN(n10189) );
  AOI211_X1 U10929 ( .C1(n10191), .C2(n10659), .A(n10190), .B(n10189), .ZN(
        n10624) );
  NAND2_X1 U10930 ( .A1(n10192), .A2(n10626), .ZN(n10627) );
  AND2_X1 U10931 ( .A1(n10193), .A2(n6731), .ZN(n10194) );
  NOR2_X1 U10932 ( .A1(n10627), .A2(n10194), .ZN(n10620) );
  AOI21_X1 U10933 ( .B1(n10663), .B2(n6731), .A(n10620), .ZN(n10195) );
  OAI211_X1 U10934 ( .C1(n10665), .C2(n10618), .A(n10624), .B(n10195), .ZN(
        n10613) );
  MUX2_X1 U10935 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10613), .S(n10757), .Z(
        P1_U3523) );
  INV_X1 U10936 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10197) );
  MUX2_X1 U10937 ( .A(n10197), .B(n10196), .S(n10761), .Z(n10198) );
  OAI21_X1 U10938 ( .B1(n10199), .B2(n10220), .A(n10198), .ZN(P1_U3521) );
  MUX2_X1 U10939 ( .A(n10200), .B(P1_REG0_REG_30__SCAN_IN), .S(n10758), .Z(
        n10201) );
  INV_X1 U10940 ( .A(n10201), .ZN(n10202) );
  OAI21_X1 U10941 ( .B1(n8399), .B2(n10220), .A(n10202), .ZN(P1_U3520) );
  MUX2_X1 U10942 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10203), .S(n10761), .Z(
        P1_U3519) );
  INV_X1 U10943 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10205) );
  MUX2_X1 U10944 ( .A(n10205), .B(n10204), .S(n10761), .Z(n10206) );
  OAI21_X1 U10945 ( .B1(n10207), .B2(n10220), .A(n10206), .ZN(P1_U3517) );
  INV_X1 U10946 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10209) );
  MUX2_X1 U10947 ( .A(n10209), .B(n10208), .S(n10761), .Z(n10210) );
  OAI21_X1 U10948 ( .B1(n10211), .B2(n10220), .A(n10210), .ZN(P1_U3516) );
  MUX2_X1 U10949 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10212), .S(n10761), .Z(
        P1_U3515) );
  INV_X1 U10950 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10214) );
  MUX2_X1 U10951 ( .A(n10214), .B(n10213), .S(n10761), .Z(n10215) );
  OAI21_X1 U10952 ( .B1(n10216), .B2(n10220), .A(n10215), .ZN(P1_U3514) );
  INV_X1 U10953 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10218) );
  MUX2_X1 U10954 ( .A(n10218), .B(n10217), .S(n10761), .Z(n10219) );
  OAI21_X1 U10955 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(P1_U3513) );
  MUX2_X1 U10956 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10222), .S(n10761), .Z(
        P1_U3512) );
  MUX2_X1 U10957 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10223), .S(n10761), .Z(
        P1_U3511) );
  MUX2_X1 U10958 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10224), .S(n10761), .Z(
        P1_U3510) );
  MUX2_X1 U10959 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10225), .S(n10761), .Z(
        P1_U3509) );
  MUX2_X1 U10960 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10226), .S(n10761), .Z(
        P1_U3507) );
  MUX2_X1 U10961 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10227), .S(n10761), .Z(
        P1_U3504) );
  MUX2_X1 U10962 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10228), .S(n10761), .Z(
        P1_U3501) );
  MUX2_X1 U10963 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10229), .S(n10761), .Z(
        P1_U3498) );
  MUX2_X1 U10964 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10230), .S(n10761), .Z(
        P1_U3492) );
  CLKBUF_X1 U10965 ( .A(n10269), .Z(n10283) );
  MUX2_X1 U10966 ( .A(P1_D_REG_0__SCAN_IN), .B(n10232), .S(n10283), .Z(
        P1_U3439) );
  NOR4_X1 U10967 ( .A1(n10234), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n10233), .ZN(n10235) );
  AOI21_X1 U10968 ( .B1(n10241), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10235), 
        .ZN(n10236) );
  OAI21_X1 U10969 ( .B1(n10237), .B2(n7238), .A(n10236), .ZN(P1_U3324) );
  AOI22_X1 U10970 ( .A1(n10238), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10241), .ZN(n10239) );
  OAI21_X1 U10971 ( .B1(n10240), .B2(n7238), .A(n10239), .ZN(P1_U3325) );
  AOI22_X1 U10972 ( .A1(n10242), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10241), .ZN(n10243) );
  OAI21_X1 U10973 ( .B1(n10244), .B2(n7238), .A(n10243), .ZN(P1_U3326) );
  AOI22_X1 U10974 ( .A1(n10245), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10241), .ZN(n10246) );
  OAI21_X1 U10975 ( .B1(n10247), .B2(n7238), .A(n10246), .ZN(P1_U3327) );
  AOI22_X1 U10976 ( .A1(n10364), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10241), .ZN(n10248) );
  OAI21_X1 U10977 ( .B1(n10249), .B2(n7238), .A(n10248), .ZN(P1_U3328) );
  INV_X1 U10978 ( .A(n10250), .ZN(n10251) );
  MUX2_X1 U10979 ( .A(n10251), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10980 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U10981 ( .A1(n10269), .A2(n10252), .ZN(P1_U3323) );
  INV_X1 U10982 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10253) );
  NOR2_X1 U10983 ( .A1(n10269), .A2(n10253), .ZN(P1_U3322) );
  INV_X1 U10984 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10254) );
  NOR2_X1 U10985 ( .A1(n10283), .A2(n10254), .ZN(P1_U3321) );
  INV_X1 U10986 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U10987 ( .A1(n10283), .A2(n10255), .ZN(P1_U3320) );
  INV_X1 U10988 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10256) );
  NOR2_X1 U10989 ( .A1(n10283), .A2(n10256), .ZN(P1_U3319) );
  INV_X1 U10990 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10257) );
  NOR2_X1 U10991 ( .A1(n10283), .A2(n10257), .ZN(P1_U3318) );
  INV_X1 U10992 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U10993 ( .A1(n10283), .A2(n10258), .ZN(P1_U3317) );
  INV_X1 U10994 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U10995 ( .A1(n10283), .A2(n10259), .ZN(P1_U3316) );
  INV_X1 U10996 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10260) );
  NOR2_X1 U10997 ( .A1(n10283), .A2(n10260), .ZN(P1_U3315) );
  INV_X1 U10998 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U10999 ( .A1(n10269), .A2(n10261), .ZN(P1_U3314) );
  INV_X1 U11000 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10262) );
  NOR2_X1 U11001 ( .A1(n10269), .A2(n10262), .ZN(P1_U3313) );
  INV_X1 U11002 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10263) );
  NOR2_X1 U11003 ( .A1(n10269), .A2(n10263), .ZN(P1_U3312) );
  INV_X1 U11004 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U11005 ( .A1(n10269), .A2(n10264), .ZN(P1_U3311) );
  INV_X1 U11006 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10265) );
  NOR2_X1 U11007 ( .A1(n10269), .A2(n10265), .ZN(P1_U3310) );
  INV_X1 U11008 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10266) );
  NOR2_X1 U11009 ( .A1(n10269), .A2(n10266), .ZN(P1_U3309) );
  INV_X1 U11010 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U11011 ( .A1(n10269), .A2(n10267), .ZN(P1_U3308) );
  INV_X1 U11012 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10268) );
  NOR2_X1 U11013 ( .A1(n10269), .A2(n10268), .ZN(P1_U3307) );
  INV_X1 U11014 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U11015 ( .A1(n10283), .A2(n10270), .ZN(P1_U3306) );
  INV_X1 U11016 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U11017 ( .A1(n10283), .A2(n10271), .ZN(P1_U3305) );
  INV_X1 U11018 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10272) );
  NOR2_X1 U11019 ( .A1(n10283), .A2(n10272), .ZN(P1_U3304) );
  INV_X1 U11020 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U11021 ( .A1(n10283), .A2(n10273), .ZN(P1_U3303) );
  INV_X1 U11022 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U11023 ( .A1(n10283), .A2(n10274), .ZN(P1_U3302) );
  INV_X1 U11024 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U11025 ( .A1(n10283), .A2(n10275), .ZN(P1_U3301) );
  INV_X1 U11026 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10276) );
  NOR2_X1 U11027 ( .A1(n10283), .A2(n10276), .ZN(P1_U3300) );
  INV_X1 U11028 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10277) );
  NOR2_X1 U11029 ( .A1(n10283), .A2(n10277), .ZN(P1_U3299) );
  INV_X1 U11030 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U11031 ( .A1(n10283), .A2(n10278), .ZN(P1_U3298) );
  INV_X1 U11032 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10279) );
  NOR2_X1 U11033 ( .A1(n10283), .A2(n10279), .ZN(P1_U3297) );
  INV_X1 U11034 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10280) );
  NOR2_X1 U11035 ( .A1(n10283), .A2(n10280), .ZN(P1_U3296) );
  INV_X1 U11036 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10281) );
  NOR2_X1 U11037 ( .A1(n10283), .A2(n10281), .ZN(P1_U3295) );
  INV_X1 U11038 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10282) );
  NOR2_X1 U11039 ( .A1(n10283), .A2(n10282), .ZN(P1_U3294) );
  NAND2_X1 U11040 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10287) );
  OAI21_X1 U11041 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10287), .ZN(n10284) );
  INV_X1 U11042 ( .A(n10284), .ZN(ADD_1068_U46) );
  INV_X1 U11043 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U11044 ( .A1(n10285), .A2(n10287), .ZN(n10288) );
  OAI21_X1 U11045 ( .B1(n10285), .B2(n10287), .A(n10288), .ZN(n10286) );
  XNOR2_X1 U11046 ( .A(n10286), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  INV_X1 U11047 ( .A(n10287), .ZN(n10289) );
  AOI22_X1 U11048 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10289), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10288), .ZN(n10292) );
  NAND2_X1 U11049 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10290) );
  OAI21_X1 U11050 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10290), .ZN(n10291) );
  NOR2_X1 U11051 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  AOI21_X1 U11052 ( .B1(n10292), .B2(n10291), .A(n10293), .ZN(ADD_1068_U54) );
  AOI21_X1 U11053 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10293), .ZN(n10296) );
  NAND2_X1 U11054 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10294) );
  OAI21_X1 U11055 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10294), .ZN(n10295) );
  NOR2_X1 U11056 ( .A1(n10296), .A2(n10295), .ZN(n10297) );
  AOI21_X1 U11057 ( .B1(n10296), .B2(n10295), .A(n10297), .ZN(ADD_1068_U53) );
  AOI21_X1 U11058 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10297), .ZN(n10300) );
  NOR2_X1 U11059 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10298) );
  AOI21_X1 U11060 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10298), .ZN(n10299) );
  NAND2_X1 U11061 ( .A1(n10300), .A2(n10299), .ZN(n10302) );
  OAI21_X1 U11062 ( .B1(n10300), .B2(n10299), .A(n10302), .ZN(ADD_1068_U52) );
  NOR2_X1 U11063 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10301) );
  AOI21_X1 U11064 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10301), .ZN(n10304) );
  OAI21_X1 U11065 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10302), .ZN(n10303) );
  NAND2_X1 U11066 ( .A1(n10304), .A2(n10303), .ZN(n10306) );
  OAI21_X1 U11067 ( .B1(n10304), .B2(n10303), .A(n10306), .ZN(ADD_1068_U51) );
  NOR2_X1 U11068 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10305) );
  AOI21_X1 U11069 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10305), .ZN(n10308) );
  OAI21_X1 U11070 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10306), .ZN(n10307) );
  NAND2_X1 U11071 ( .A1(n10308), .A2(n10307), .ZN(n10310) );
  OAI21_X1 U11072 ( .B1(n10308), .B2(n10307), .A(n10310), .ZN(ADD_1068_U50) );
  NOR2_X1 U11073 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10309) );
  AOI21_X1 U11074 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10309), .ZN(n10312) );
  OAI21_X1 U11075 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10310), .ZN(n10311) );
  NAND2_X1 U11076 ( .A1(n10312), .A2(n10311), .ZN(n10314) );
  OAI21_X1 U11077 ( .B1(n10312), .B2(n10311), .A(n10314), .ZN(ADD_1068_U49) );
  NOR2_X1 U11078 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10313) );
  AOI21_X1 U11079 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10313), .ZN(n10316) );
  OAI21_X1 U11080 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10314), .ZN(n10315) );
  NAND2_X1 U11081 ( .A1(n10316), .A2(n10315), .ZN(n10318) );
  OAI21_X1 U11082 ( .B1(n10316), .B2(n10315), .A(n10318), .ZN(ADD_1068_U48) );
  NOR2_X1 U11083 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10317) );
  AOI21_X1 U11084 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10317), .ZN(n10320) );
  OAI21_X1 U11085 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10318), .ZN(n10319) );
  NAND2_X1 U11086 ( .A1(n10320), .A2(n10319), .ZN(n10322) );
  OAI21_X1 U11087 ( .B1(n10320), .B2(n10319), .A(n10322), .ZN(ADD_1068_U47) );
  NOR2_X1 U11088 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10321) );
  AOI21_X1 U11089 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10321), .ZN(n10324) );
  OAI21_X1 U11090 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10322), .ZN(n10323) );
  NAND2_X1 U11091 ( .A1(n10324), .A2(n10323), .ZN(n10326) );
  OAI21_X1 U11092 ( .B1(n10324), .B2(n10323), .A(n10326), .ZN(ADD_1068_U63) );
  NOR2_X1 U11093 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10325) );
  AOI21_X1 U11094 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10325), .ZN(n10328) );
  OAI21_X1 U11095 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10326), .ZN(n10327) );
  NAND2_X1 U11096 ( .A1(n10328), .A2(n10327), .ZN(n10330) );
  OAI21_X1 U11097 ( .B1(n10328), .B2(n10327), .A(n10330), .ZN(ADD_1068_U62) );
  NOR2_X1 U11098 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10329) );
  AOI21_X1 U11099 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10329), .ZN(n10332) );
  OAI21_X1 U11100 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10330), .ZN(n10331) );
  NAND2_X1 U11101 ( .A1(n10332), .A2(n10331), .ZN(n10334) );
  OAI21_X1 U11102 ( .B1(n10332), .B2(n10331), .A(n10334), .ZN(ADD_1068_U61) );
  NOR2_X1 U11103 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10333) );
  AOI21_X1 U11104 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10333), .ZN(n10336) );
  OAI21_X1 U11105 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10334), .ZN(n10335) );
  NAND2_X1 U11106 ( .A1(n10336), .A2(n10335), .ZN(n10338) );
  OAI21_X1 U11107 ( .B1(n10336), .B2(n10335), .A(n10338), .ZN(ADD_1068_U60) );
  NOR2_X1 U11108 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10337) );
  AOI21_X1 U11109 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10337), .ZN(n10340) );
  OAI21_X1 U11110 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10338), .ZN(n10339) );
  NAND2_X1 U11111 ( .A1(n10340), .A2(n10339), .ZN(n10342) );
  OAI21_X1 U11112 ( .B1(n10340), .B2(n10339), .A(n10342), .ZN(ADD_1068_U59) );
  NOR2_X1 U11113 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10341) );
  AOI21_X1 U11114 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10341), .ZN(n10344) );
  OAI21_X1 U11115 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10342), .ZN(n10343) );
  NAND2_X1 U11116 ( .A1(n10344), .A2(n10343), .ZN(n10346) );
  OAI21_X1 U11117 ( .B1(n10344), .B2(n10343), .A(n10346), .ZN(ADD_1068_U58) );
  NOR2_X1 U11118 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10345) );
  AOI21_X1 U11119 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10345), .ZN(n10348) );
  OAI21_X1 U11120 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10346), .ZN(n10347) );
  NAND2_X1 U11121 ( .A1(n10348), .A2(n10347), .ZN(n10350) );
  OAI21_X1 U11122 ( .B1(n10348), .B2(n10347), .A(n10350), .ZN(ADD_1068_U57) );
  NOR2_X1 U11123 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10349) );
  AOI21_X1 U11124 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10349), .ZN(n10352) );
  OAI21_X1 U11125 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10350), .ZN(n10351) );
  NAND2_X1 U11126 ( .A1(n10352), .A2(n10351), .ZN(n10354) );
  OAI21_X1 U11127 ( .B1(n10352), .B2(n10351), .A(n10354), .ZN(ADD_1068_U56) );
  NOR2_X1 U11128 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n10353) );
  AOI21_X1 U11129 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n10353), .ZN(n10356) );
  OAI21_X1 U11130 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10354), .ZN(n10355) );
  NAND2_X1 U11131 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  OAI21_X1 U11132 ( .B1(n10356), .B2(n10355), .A(n10357), .ZN(ADD_1068_U55) );
  OAI21_X1 U11133 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10357), .ZN(n10359) );
  XOR2_X1 U11134 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10358) );
  XNOR2_X1 U11135 ( .A(n10359), .B(n10358), .ZN(ADD_1068_U4) );
  INV_X1 U11136 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10361) );
  AOI21_X1 U11137 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(P1_U3440) );
  OAI21_X1 U11138 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n10364), .A(n10363), .ZN(
        n10366) );
  XNOR2_X1 U11139 ( .A(n10366), .B(n10365), .ZN(n10368) );
  AOI22_X1 U11140 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10585), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10367) );
  OAI21_X1 U11141 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(P1_U3243) );
  INV_X1 U11142 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10384) );
  INV_X1 U11143 ( .A(n10370), .ZN(n10371) );
  OAI211_X1 U11144 ( .C1(n10373), .C2(n10372), .A(n10591), .B(n10371), .ZN(
        n10381) );
  AOI21_X1 U11145 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(n10377) );
  NAND2_X1 U11146 ( .A1(n10587), .A2(n10377), .ZN(n10380) );
  NAND2_X1 U11147 ( .A1(n10595), .A2(n10378), .ZN(n10379) );
  AND3_X1 U11148 ( .A1(n10381), .A2(n10380), .A3(n10379), .ZN(n10383) );
  OAI211_X1 U11149 ( .C1(n10491), .C2(n10384), .A(n10383), .B(n10382), .ZN(
        P1_U3248) );
  AOI211_X1 U11150 ( .C1(n10387), .C2(n10386), .A(n10385), .B(n10496), .ZN(
        n10392) );
  AOI211_X1 U11151 ( .C1(n10390), .C2(n10389), .A(n10388), .B(n10492), .ZN(
        n10391) );
  AOI211_X1 U11152 ( .C1(n10595), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        n10394) );
  INV_X1 U11153 ( .A(n10394), .ZN(n10396) );
  AOI211_X1 U11154 ( .C1(n10585), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10396), .B(
        n10395), .ZN(n10397) );
  INV_X1 U11155 ( .A(n10397), .ZN(P1_U3249) );
  INV_X1 U11156 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10409) );
  AOI211_X1 U11157 ( .C1(n10400), .C2(n10399), .A(n10398), .B(n10496), .ZN(
        n10405) );
  AOI211_X1 U11158 ( .C1(n10403), .C2(n10402), .A(n10492), .B(n10401), .ZN(
        n10404) );
  AOI211_X1 U11159 ( .C1(n10595), .C2(n10406), .A(n10405), .B(n10404), .ZN(
        n10408) );
  OAI211_X1 U11160 ( .C1(n10491), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        P1_U3250) );
  OAI211_X1 U11161 ( .C1(n10412), .C2(n10411), .A(n10410), .B(n10591), .ZN(
        n10419) );
  INV_X1 U11162 ( .A(n10413), .ZN(n10417) );
  INV_X1 U11163 ( .A(n10414), .ZN(n10416) );
  OAI211_X1 U11164 ( .C1(n10417), .C2(n10416), .A(n10587), .B(n10415), .ZN(
        n10418) );
  OAI211_X1 U11165 ( .C1(n10451), .C2(n10420), .A(n10419), .B(n10418), .ZN(
        n10422) );
  AOI211_X1 U11166 ( .C1(n10585), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10422), .B(
        n10421), .ZN(n10423) );
  INV_X1 U11167 ( .A(n10423), .ZN(P1_U3251) );
  INV_X1 U11168 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10438) );
  AOI21_X1 U11169 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(n10427) );
  NAND2_X1 U11170 ( .A1(n10591), .A2(n10427), .ZN(n10433) );
  AOI21_X1 U11171 ( .B1(n10430), .B2(n10429), .A(n10428), .ZN(n10431) );
  NAND2_X1 U11172 ( .A1(n10587), .A2(n10431), .ZN(n10432) );
  OAI211_X1 U11173 ( .C1(n10451), .C2(n10434), .A(n10433), .B(n10432), .ZN(
        n10435) );
  INV_X1 U11174 ( .A(n10435), .ZN(n10437) );
  OAI211_X1 U11175 ( .C1(n10491), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        P1_U3254) );
  INV_X1 U11176 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10455) );
  INV_X1 U11177 ( .A(n10439), .ZN(n10450) );
  AOI21_X1 U11178 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(n10443) );
  NAND2_X1 U11179 ( .A1(n10587), .A2(n10443), .ZN(n10449) );
  AOI21_X1 U11180 ( .B1(n10446), .B2(n10445), .A(n10444), .ZN(n10447) );
  NAND2_X1 U11181 ( .A1(n10591), .A2(n10447), .ZN(n10448) );
  OAI211_X1 U11182 ( .C1(n10451), .C2(n10450), .A(n10449), .B(n10448), .ZN(
        n10452) );
  INV_X1 U11183 ( .A(n10452), .ZN(n10454) );
  NAND2_X1 U11184 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10453)
         );
  OAI211_X1 U11185 ( .C1(n10491), .C2(n10455), .A(n10454), .B(n10453), .ZN(
        P1_U3257) );
  INV_X1 U11186 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10467) );
  AOI211_X1 U11187 ( .C1(n10458), .C2(n10457), .A(n10456), .B(n10492), .ZN(
        n10463) );
  AOI211_X1 U11188 ( .C1(n10461), .C2(n10460), .A(n10459), .B(n10496), .ZN(
        n10462) );
  AOI211_X1 U11189 ( .C1(n10595), .C2(n10464), .A(n10463), .B(n10462), .ZN(
        n10466) );
  NAND2_X1 U11190 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n10465)
         );
  OAI211_X1 U11191 ( .C1(n10491), .C2(n10467), .A(n10466), .B(n10465), .ZN(
        P1_U3258) );
  AOI211_X1 U11192 ( .C1(n10470), .C2(n10469), .A(n10492), .B(n10468), .ZN(
        n10476) );
  INV_X1 U11193 ( .A(n10471), .ZN(n10472) );
  AOI211_X1 U11194 ( .C1(n10474), .C2(n10473), .A(n10496), .B(n10472), .ZN(
        n10475) );
  INV_X1 U11195 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10490) );
  AOI211_X1 U11196 ( .C1(n10481), .C2(n10480), .A(n10479), .B(n10492), .ZN(
        n10486) );
  AOI211_X1 U11197 ( .C1(n10484), .C2(n10483), .A(n10482), .B(n10496), .ZN(
        n10485) );
  AOI211_X1 U11198 ( .C1(n10595), .C2(n10487), .A(n10486), .B(n10485), .ZN(
        n10489) );
  OAI211_X1 U11199 ( .C1(n10491), .C2(n10490), .A(n10489), .B(n10488), .ZN(
        P1_U3256) );
  AOI211_X1 U11200 ( .C1(n10495), .C2(n10494), .A(n10493), .B(n10492), .ZN(
        n10501) );
  AOI211_X1 U11201 ( .C1(n10499), .C2(n10498), .A(n10497), .B(n10496), .ZN(
        n10500) );
  AOI211_X1 U11202 ( .C1(n10595), .C2(n10502), .A(n10501), .B(n10500), .ZN(
        n10503) );
  INV_X1 U11203 ( .A(n10503), .ZN(n10505) );
  AOI211_X1 U11204 ( .C1(n10585), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n10505), 
        .B(n10504), .ZN(n10506) );
  INV_X1 U11205 ( .A(n10506), .ZN(P1_U3253) );
  AOI22_X1 U11206 ( .A1(n10566), .A2(P2_IR_REG_0__SCAN_IN), .B1(n10564), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10511) );
  INV_X1 U11207 ( .A(n10536), .ZN(n10575) );
  XOR2_X1 U11208 ( .A(n10507), .B(P2_IR_REG_0__SCAN_IN), .Z(n10508) );
  OAI21_X1 U11209 ( .B1(n10509), .B2(n10575), .A(n10508), .ZN(n10510) );
  OAI211_X1 U11210 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10512), .A(n10511), .B(
        n10510), .ZN(P2_U3182) );
  INV_X1 U11211 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10528) );
  OAI21_X1 U11212 ( .B1(n10514), .B2(P2_REG2_REG_3__SCAN_IN), .A(n10513), .ZN(
        n10515) );
  AOI22_X1 U11213 ( .A1(n10566), .A2(n10516), .B1(n10578), .B2(n10515), .ZN(
        n10527) );
  OAI21_X1 U11214 ( .B1(n10519), .B2(n10518), .A(n10517), .ZN(n10525) );
  OAI21_X1 U11215 ( .B1(n10521), .B2(P2_REG1_REG_3__SCAN_IN), .A(n10520), .ZN(
        n10522) );
  AND2_X1 U11216 ( .A1(n10579), .A2(n10522), .ZN(n10523) );
  AOI211_X1 U11217 ( .C1(n10525), .C2(n10575), .A(n10524), .B(n10523), .ZN(
        n10526) );
  OAI211_X1 U11218 ( .C1(n10563), .C2(n10528), .A(n10527), .B(n10526), .ZN(
        P2_U3185) );
  INV_X1 U11219 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10544) );
  OAI21_X1 U11220 ( .B1(n10531), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10530), .ZN(
        n10532) );
  AOI22_X1 U11221 ( .A1(n10566), .A2(n5220), .B1(n10578), .B2(n10532), .ZN(
        n10543) );
  OAI21_X1 U11222 ( .B1(n10534), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10533), .ZN(
        n10541) );
  AOI211_X1 U11223 ( .C1(n10538), .C2(n10537), .A(n10536), .B(n10535), .ZN(
        n10539) );
  AOI211_X1 U11224 ( .C1(n10579), .C2(n10541), .A(n10540), .B(n10539), .ZN(
        n10542) );
  OAI211_X1 U11225 ( .C1(n10563), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        P2_U3187) );
  INV_X1 U11226 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10562) );
  OAI21_X1 U11227 ( .B1(n10547), .B2(n10546), .A(n10545), .ZN(n10548) );
  AOI22_X1 U11228 ( .A1(n10549), .A2(n10566), .B1(n10548), .B2(n10578), .ZN(
        n10561) );
  OAI21_X1 U11229 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(n10559) );
  OAI21_X1 U11230 ( .B1(n10555), .B2(n10554), .A(n10553), .ZN(n10556) );
  AND2_X1 U11231 ( .A1(n10556), .A2(n10579), .ZN(n10557) );
  AOI211_X1 U11232 ( .C1(n10559), .C2(n10575), .A(n10558), .B(n10557), .ZN(
        n10560) );
  OAI211_X1 U11233 ( .C1(n10563), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        P2_U3188) );
  AOI22_X1 U11234 ( .A1(n10566), .A2(n10565), .B1(n10564), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10582) );
  OAI21_X1 U11235 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(n10580) );
  OAI21_X1 U11236 ( .B1(n10572), .B2(n10571), .A(n10570), .ZN(n10577) );
  XNOR2_X1 U11237 ( .A(n10574), .B(n10573), .ZN(n10576) );
  AOI222_X1 U11238 ( .A1(n10580), .A2(n10579), .B1(n10578), .B2(n10577), .C1(
        n10576), .C2(n10575), .ZN(n10581) );
  OAI211_X1 U11239 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10583), .A(n10582), .B(
        n10581), .ZN(P2_U3196) );
  XNOR2_X1 U11240 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11241 ( .B1(n10585), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10584), .ZN(
        n10601) );
  OAI211_X1 U11242 ( .C1(n10589), .C2(n10588), .A(n10587), .B(n10586), .ZN(
        n10598) );
  OAI211_X1 U11243 ( .C1(n10593), .C2(n10592), .A(n10591), .B(n10590), .ZN(
        n10597) );
  NAND2_X1 U11244 ( .A1(n10595), .A2(n10594), .ZN(n10596) );
  AND3_X1 U11245 ( .A1(n10598), .A2(n10597), .A3(n10596), .ZN(n10600) );
  NAND3_X1 U11246 ( .A1(n10601), .A2(n10600), .A3(n10599), .ZN(P1_U3247) );
  NOR3_X1 U11247 ( .A1(n10604), .A2(n10603), .A3(n10602), .ZN(n10611) );
  NOR2_X1 U11248 ( .A1(n10718), .A2(n10605), .ZN(n10609) );
  NOR3_X1 U11249 ( .A1(n10688), .A2(n10607), .A3(n10606), .ZN(n10608) );
  NOR4_X1 U11250 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  AOI22_X1 U11251 ( .A1(n10714), .A2(n9811), .B1(n10612), .B2(n10707), .ZN(
        P1_U3293) );
  INV_X1 U11252 ( .A(n10613), .ZN(n10615) );
  INV_X1 U11253 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U11254 ( .A1(n10761), .A2(n10615), .B1(n10614), .B2(n10758), .ZN(
        P1_U3456) );
  OAI22_X1 U11255 ( .A1(n10670), .A2(n10616), .B1(n7158), .B2(n10718), .ZN(
        n10617) );
  AOI21_X1 U11256 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n10714), .A(n10617), .ZN(
        n10623) );
  INV_X1 U11257 ( .A(n10618), .ZN(n10621) );
  INV_X1 U11258 ( .A(n10619), .ZN(n10675) );
  AOI22_X1 U11259 ( .A1(n10621), .A2(n10675), .B1(n10674), .B2(n10620), .ZN(
        n10622) );
  OAI211_X1 U11260 ( .C1(n10714), .C2(n10624), .A(n10623), .B(n10622), .ZN(
        P1_U3292) );
  XNOR2_X1 U11261 ( .A(n10625), .B(n10632), .ZN(n10637) );
  OAI21_X1 U11262 ( .B1(n10660), .B2(n10626), .A(n10750), .ZN(n10630) );
  INV_X1 U11263 ( .A(n10627), .ZN(n10629) );
  MUX2_X1 U11264 ( .A(n10630), .B(n10629), .S(n10628), .Z(n10639) );
  XNOR2_X1 U11265 ( .A(n10632), .B(n10631), .ZN(n10633) );
  OAI222_X1 U11266 ( .A1(n10701), .A2(n10634), .B1(n10703), .B2(n10700), .C1(
        n10633), .C2(n10698), .ZN(n10636) );
  AOI211_X1 U11267 ( .C1(n10754), .C2(n10637), .A(n10639), .B(n10636), .ZN(
        n10635) );
  AOI22_X1 U11268 ( .A1(n10757), .A2(n10635), .B1(n5732), .B2(n10756), .ZN(
        P1_U3524) );
  AOI22_X1 U11269 ( .A1(n10761), .A2(n10635), .B1(n5731), .B2(n10758), .ZN(
        P1_U3459) );
  AOI21_X1 U11270 ( .B1(n10713), .B2(n10637), .A(n10636), .ZN(n10642) );
  INV_X1 U11271 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U11272 ( .A1(n10639), .A2(n10709), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10638), .ZN(n10640) );
  OAI221_X1 U11273 ( .B1(n10714), .B2(n10642), .C1(n10707), .C2(n10641), .A(
        n10640), .ZN(P1_U3291) );
  INV_X1 U11274 ( .A(n10643), .ZN(n10644) );
  AOI211_X1 U11275 ( .C1(n10733), .C2(n10646), .A(n10645), .B(n10644), .ZN(
        n10648) );
  AOI22_X1 U11276 ( .A1(n10791), .A2(n10648), .B1(n6226), .B2(n10782), .ZN(
        P2_U3461) );
  INV_X1 U11277 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U11278 ( .A1(n6696), .A2(n10648), .B1(n10647), .B2(n10792), .ZN(
        P2_U3396) );
  XNOR2_X1 U11279 ( .A(n10649), .B(n10652), .ZN(n10672) );
  OAI21_X1 U11280 ( .B1(n10652), .B2(n10651), .A(n10650), .ZN(n10658) );
  OAI22_X1 U11281 ( .A1(n10654), .A2(n10703), .B1(n10653), .B2(n10701), .ZN(
        n10657) );
  NOR2_X1 U11282 ( .A1(n10672), .A2(n10655), .ZN(n10656) );
  AOI211_X1 U11283 ( .C1(n10659), .C2(n10658), .A(n10657), .B(n10656), .ZN(
        n10679) );
  OR2_X1 U11284 ( .A1(n10690), .A2(n10660), .ZN(n10687) );
  AOI21_X1 U11285 ( .B1(n10662), .B2(n10661), .A(n10687), .ZN(n10673) );
  AOI21_X1 U11286 ( .B1(n10663), .B2(n10662), .A(n10673), .ZN(n10664) );
  OAI211_X1 U11287 ( .C1(n10672), .C2(n10665), .A(n10679), .B(n10664), .ZN(
        n10666) );
  INV_X1 U11288 ( .A(n10666), .ZN(n10668) );
  AOI22_X1 U11289 ( .A1(n10757), .A2(n10668), .B1(n7099), .B2(n10756), .ZN(
        P1_U3525) );
  INV_X1 U11290 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U11291 ( .A1(n10761), .A2(n10668), .B1(n10667), .B2(n10758), .ZN(
        P1_U3462) );
  OAI22_X1 U11292 ( .A1(n10670), .A2(n10669), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n10718), .ZN(n10671) );
  AOI21_X1 U11293 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n10714), .A(n10671), .ZN(
        n10678) );
  INV_X1 U11294 ( .A(n10672), .ZN(n10676) );
  AOI22_X1 U11295 ( .A1(n10676), .A2(n10675), .B1(n10674), .B2(n10673), .ZN(
        n10677) );
  OAI211_X1 U11296 ( .C1(n10714), .C2(n10679), .A(n10678), .B(n10677), .ZN(
        P1_U3290) );
  NOR2_X1 U11297 ( .A1(n10680), .A2(n10785), .ZN(n10682) );
  AOI211_X1 U11298 ( .C1(n10775), .C2(n10683), .A(n10682), .B(n10681), .ZN(
        n10685) );
  AOI22_X1 U11299 ( .A1(n10791), .A2(n10685), .B1(n7340), .B2(n10782), .ZN(
        P2_U3463) );
  INV_X1 U11300 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U11301 ( .A1(n6696), .A2(n10685), .B1(n10684), .B2(n10792), .ZN(
        P2_U3402) );
  XOR2_X1 U11302 ( .A(n10696), .B(n10686), .Z(n10712) );
  OAI21_X1 U11303 ( .B1(n10689), .B2(n10688), .A(n10687), .ZN(n10695) );
  INV_X1 U11304 ( .A(n10690), .ZN(n10693) );
  NAND3_X1 U11305 ( .A1(n10693), .A2(n10692), .A3(n10691), .ZN(n10694) );
  AND2_X1 U11306 ( .A1(n10695), .A2(n10694), .ZN(n10710) );
  XOR2_X1 U11307 ( .A(n10697), .B(n10696), .Z(n10699) );
  OAI222_X1 U11308 ( .A1(n10703), .A2(n10702), .B1(n10701), .B2(n10700), .C1(
        n10699), .C2(n10698), .ZN(n10711) );
  AOI211_X1 U11309 ( .C1(n10754), .C2(n10712), .A(n10710), .B(n10711), .ZN(
        n10705) );
  AOI22_X1 U11310 ( .A1(n10757), .A2(n10705), .B1(n7101), .B2(n10756), .ZN(
        P1_U3526) );
  INV_X1 U11311 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U11312 ( .A1(n10761), .A2(n10705), .B1(n10704), .B2(n10758), .ZN(
        P1_U3465) );
  NOR2_X1 U11313 ( .A1(n10707), .A2(n10706), .ZN(n10708) );
  AOI21_X1 U11314 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(n10717) );
  AOI21_X1 U11315 ( .B1(n10713), .B2(n10712), .A(n10711), .ZN(n10715) );
  OR2_X1 U11316 ( .A1(n10715), .A2(n10714), .ZN(n10716) );
  OAI211_X1 U11317 ( .C1(n10719), .C2(n10718), .A(n10717), .B(n10716), .ZN(
        P1_U3289) );
  NOR2_X1 U11318 ( .A1(n10720), .A2(n10785), .ZN(n10722) );
  AOI211_X1 U11319 ( .C1(n10733), .C2(n10723), .A(n10722), .B(n10721), .ZN(
        n10725) );
  AOI22_X1 U11320 ( .A1(n10791), .A2(n10725), .B1(n6266), .B2(n10782), .ZN(
        P2_U3464) );
  INV_X1 U11321 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U11322 ( .A1(n6696), .A2(n10725), .B1(n10724), .B2(n10792), .ZN(
        P2_U3405) );
  INV_X1 U11323 ( .A(n10726), .ZN(n10730) );
  OAI22_X1 U11324 ( .A1(n10728), .A2(n10787), .B1(n10727), .B2(n10785), .ZN(
        n10729) );
  NOR2_X1 U11325 ( .A1(n10730), .A2(n10729), .ZN(n10732) );
  AOI22_X1 U11326 ( .A1(n10791), .A2(n10732), .B1(n6281), .B2(n10782), .ZN(
        P2_U3465) );
  INV_X1 U11327 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U11328 ( .A1(n6696), .A2(n10732), .B1(n10731), .B2(n10792), .ZN(
        P2_U3408) );
  NAND2_X1 U11329 ( .A1(n10734), .A2(n10733), .ZN(n10737) );
  NAND2_X1 U11330 ( .A1(n10735), .A2(n10777), .ZN(n10736) );
  NAND2_X1 U11331 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  NOR2_X1 U11332 ( .A1(n10739), .A2(n10738), .ZN(n10741) );
  AOI22_X1 U11333 ( .A1(n10791), .A2(n10741), .B1(n7923), .B2(n10782), .ZN(
        P2_U3469) );
  INV_X1 U11334 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U11335 ( .A1(n6696), .A2(n10741), .B1(n10740), .B2(n10792), .ZN(
        P2_U3420) );
  AND2_X1 U11336 ( .A1(n10742), .A2(n10775), .ZN(n10746) );
  AND2_X1 U11337 ( .A1(n10743), .A2(n10777), .ZN(n10745) );
  NOR3_X1 U11338 ( .A1(n10746), .A2(n10745), .A3(n10744), .ZN(n10748) );
  AOI22_X1 U11339 ( .A1(n10791), .A2(n10748), .B1(n8073), .B2(n10782), .ZN(
        P2_U3470) );
  INV_X1 U11340 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U11341 ( .A1(n6696), .A2(n10748), .B1(n10747), .B2(n10792), .ZN(
        P2_U3423) );
  OAI21_X1 U11342 ( .B1(n10751), .B2(n10750), .A(n10749), .ZN(n10752) );
  AOI211_X1 U11343 ( .C1(n10755), .C2(n10754), .A(n10753), .B(n10752), .ZN(
        n10760) );
  AOI22_X1 U11344 ( .A1(n10757), .A2(n10760), .B1(n7272), .B2(n10756), .ZN(
        P1_U3533) );
  INV_X1 U11345 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U11346 ( .A1(n10761), .A2(n10760), .B1(n10759), .B2(n10758), .ZN(
        P1_U3486) );
  NOR2_X1 U11347 ( .A1(n10762), .A2(n10787), .ZN(n10765) );
  INV_X1 U11348 ( .A(n10763), .ZN(n10764) );
  AOI211_X1 U11349 ( .C1(n10777), .C2(n10766), .A(n10765), .B(n10764), .ZN(
        n10768) );
  AOI22_X1 U11350 ( .A1(n10791), .A2(n10768), .B1(n8075), .B2(n10782), .ZN(
        P2_U3471) );
  INV_X1 U11351 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U11352 ( .A1(n6696), .A2(n10768), .B1(n10767), .B2(n10792), .ZN(
        P2_U3426) );
  NOR2_X1 U11353 ( .A1(n10769), .A2(n10785), .ZN(n10771) );
  AOI211_X1 U11354 ( .C1(n10772), .C2(n10775), .A(n10771), .B(n10770), .ZN(
        n10774) );
  AOI22_X1 U11355 ( .A1(n10791), .A2(n10774), .B1(n6382), .B2(n10782), .ZN(
        P2_U3472) );
  INV_X1 U11356 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U11357 ( .A1(n6696), .A2(n10774), .B1(n10773), .B2(n10792), .ZN(
        P2_U3429) );
  AND2_X1 U11358 ( .A1(n10776), .A2(n10775), .ZN(n10780) );
  AND2_X1 U11359 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  NOR3_X1 U11360 ( .A1(n10781), .A2(n10780), .A3(n10779), .ZN(n10784) );
  AOI22_X1 U11361 ( .A1(n10791), .A2(n10784), .B1(n8966), .B2(n10782), .ZN(
        P2_U3473) );
  INV_X1 U11362 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U11363 ( .A1(n6696), .A2(n10784), .B1(n10783), .B2(n10792), .ZN(
        P2_U3432) );
  OAI22_X1 U11364 ( .A1(n10788), .A2(n10787), .B1(n10786), .B2(n10785), .ZN(
        n10790) );
  NOR2_X1 U11365 ( .A1(n10790), .A2(n10789), .ZN(n10794) );
  AOI22_X1 U11366 ( .A1(n10791), .A2(n10794), .B1(n8949), .B2(n10782), .ZN(
        P2_U3474) );
  INV_X1 U11367 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U11368 ( .A1(n6696), .A2(n10794), .B1(n10793), .B2(n10792), .ZN(
        P2_U3435) );
  XNOR2_X1 U11369 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND2_X2 U5007 ( .A1(n5224), .A2(n5222), .ZN(n5701) );
  CLKBUF_X2 U4989 ( .A(n5013), .Z(n8574) );
  CLKBUF_X1 U4992 ( .A(n6244), .Z(n6401) );
  CLKBUF_X1 U5003 ( .A(n5759), .Z(n7060) );
  AND2_X1 U5008 ( .A1(n5701), .A2(P2_U3151), .ZN(n10798) );
endmodule

