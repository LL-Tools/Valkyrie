

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
         n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
         n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
         n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
         n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
         n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
         n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22789;

  NOR2_X1 U11260 ( .A1(n21745), .A2(n21673), .ZN(n21967) );
  INV_X2 U11261 ( .A(n16956), .ZN(n16955) );
  XNOR2_X1 U11262 ( .A(n13321), .B(n22179), .ZN(n15171) );
  OR2_X1 U11263 ( .A1(n11858), .A2(n11842), .ZN(n11931) );
  INV_X2 U11264 ( .A(n12113), .ZN(n11961) );
  NAND2_X1 U11265 ( .A1(n14249), .A2(n15025), .ZN(n14345) );
  OR2_X1 U11266 ( .A1(n13252), .A2(n13251), .ZN(n13258) );
  NAND2_X1 U11267 ( .A1(n11945), .A2(n11946), .ZN(n12115) );
  INV_X2 U11268 ( .A(n14125), .ZN(n18713) );
  CLKBUF_X2 U11269 ( .A(n11752), .Z(n20269) );
  INV_X1 U11271 ( .A(n18547), .ZN(n18366) );
  BUF_X1 U11272 ( .A(n18424), .Z(n18409) );
  BUF_X1 U11274 ( .A(n14064), .Z(n18522) );
  AND2_X1 U11275 ( .A1(n11169), .A2(n11739), .ZN(n11807) );
  CLKBUF_X2 U11276 ( .A(n13325), .Z(n13816) );
  NAND2_X1 U11277 ( .A1(n12572), .A2(n11737), .ZN(n15276) );
  NAND2_X1 U11278 ( .A1(n12351), .A2(n14565), .ZN(n11761) );
  CLKBUF_X1 U11279 ( .A(n11304), .Z(n19249) );
  AND2_X2 U11280 ( .A1(n11213), .A2(n11713), .ZN(n11567) );
  INV_X1 U11281 ( .A(n15025), .ZN(n15130) );
  BUF_X2 U11282 ( .A(n11589), .Z(n12788) );
  NAND2_X2 U11283 ( .A1(n11304), .A2(n12954), .ZN(n12132) );
  AND4_X1 U11284 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        n13149) );
  NAND2_X2 U11285 ( .A1(n11524), .A2(n11523), .ZN(n20528) );
  NAND3_X1 U11286 ( .A1(n13042), .A2(n13035), .A3(n11508), .ZN(n13167) );
  AND2_X2 U11287 ( .A1(n13038), .A2(n13037), .ZN(n11225) );
  AND2_X1 U11288 ( .A1(n13038), .A2(n17222), .ZN(n13325) );
  AND2_X1 U11289 ( .A1(n17222), .A2(n14712), .ZN(n13126) );
  CLKBUF_X3 U11290 ( .A(n13191), .Z(n11161) );
  AND2_X2 U11291 ( .A1(n17222), .A2(n14713), .ZN(n11227) );
  AND2_X1 U11292 ( .A1(n11390), .A2(n13036), .ZN(n13191) );
  INV_X4 U11293 ( .A(n18693), .ZN(n18689) );
  INV_X1 U11295 ( .A(n22789), .ZN(n11154) );
  AND3_X1 U11296 ( .A1(n13162), .A2(n11273), .A3(n13169), .ZN(n11245) );
  INV_X1 U11298 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11512) );
  AND2_X1 U11299 ( .A1(n13038), .A2(n14897), .ZN(n11228) );
  AND2_X1 U11300 ( .A1(n12970), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12129) );
  AND2_X2 U11301 ( .A1(n13038), .A2(n13037), .ZN(n13116) );
  OAI21_X2 U11302 ( .B1(n14705), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13234), 
        .ZN(n13252) );
  NAND3_X1 U11303 ( .A1(n13061), .A2(n11510), .A3(n13060), .ZN(n13092) );
  INV_X1 U11304 ( .A(n14107), .ZN(n14125) );
  NAND2_X1 U11305 ( .A1(n13274), .A2(n13273), .ZN(n13481) );
  AND2_X1 U11306 ( .A1(n11170), .A2(n11171), .ZN(n20851) );
  AND2_X1 U11307 ( .A1(n11390), .A2(n14713), .ZN(n13136) );
  NOR2_X1 U11308 ( .A1(n11770), .A2(n12132), .ZN(n11737) );
  NAND2_X1 U11309 ( .A1(n11847), .A2(n11846), .ZN(n11924) );
  INV_X1 U11310 ( .A(n18547), .ZN(n18455) );
  NOR3_X2 U11311 ( .A1(n18760), .A2(n18820), .A3(n11347), .ZN(n18856) );
  NAND2_X1 U11312 ( .A1(n13167), .A2(n13156), .ZN(n14256) );
  NAND2_X1 U11313 ( .A1(n11179), .A2(n16645), .ZN(n16592) );
  INV_X2 U11314 ( .A(n13412), .ZN(n16956) );
  XNOR2_X1 U11315 ( .A(n13241), .B(n13242), .ZN(n14870) );
  INV_X1 U11316 ( .A(n13156), .ZN(n15026) );
  AND2_X1 U11317 ( .A1(n11736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12312) );
  INV_X2 U11318 ( .A(n12415), .ZN(n11163) );
  XNOR2_X1 U11319 ( .A(n11343), .B(n14459), .ZN(n14471) );
  NOR2_X1 U11320 ( .A1(n14497), .A2(n19313), .ZN(n14496) );
  NOR2_X1 U11321 ( .A1(n14207), .A2(n14185), .ZN(n13013) );
  NAND2_X1 U11322 ( .A1(n11441), .A2(n11444), .ZN(n17598) );
  NAND2_X1 U11323 ( .A1(n12565), .A2(n12575), .ZN(n11773) );
  INV_X2 U11324 ( .A(n12345), .ZN(n11727) );
  NAND2_X1 U11325 ( .A1(n14028), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14029) );
  INV_X2 U11326 ( .A(n21214), .ZN(n21199) );
  OR2_X1 U11327 ( .A1(n11352), .A2(n11351), .ZN(n11350) );
  OR3_X1 U11328 ( .A1(n21206), .A2(n21221), .A3(n21201), .ZN(n18983) );
  AND2_X1 U11329 ( .A1(n18794), .A2(n11353), .ZN(n18992) );
  INV_X1 U11330 ( .A(n22119), .ZN(n21745) );
  AND2_X1 U11331 ( .A1(n16263), .A2(n16300), .ZN(n16299) );
  AND3_X1 U11332 ( .A1(n11276), .A2(n16796), .A3(n11275), .ZN(n11249) );
  NAND2_X1 U11333 ( .A1(n14870), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14871) );
  NAND2_X1 U11334 ( .A1(n17521), .A2(n17520), .ZN(n17503) );
  NAND2_X1 U11335 ( .A1(n14907), .A2(n14906), .ZN(n14905) );
  INV_X1 U11336 ( .A(n13007), .ZN(n15513) );
  AND3_X1 U11337 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14489) );
  OAI21_X2 U11338 ( .B1(n18016), .B2(n11445), .A(n11442), .ZN(n17578) );
  AND2_X1 U11339 ( .A1(n11826), .A2(n11831), .ZN(n19505) );
  INV_X1 U11340 ( .A(n21375), .ZN(n21399) );
  NAND2_X1 U11341 ( .A1(n21522), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21526) );
  INV_X1 U11342 ( .A(n20937), .ZN(n19855) );
  INV_X1 U11343 ( .A(n22357), .ZN(n22384) );
  INV_X1 U11345 ( .A(n18589), .ZN(n18602) );
  INV_X1 U11346 ( .A(n19137), .ZN(n19128) );
  INV_X2 U11347 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21656) );
  OR2_X1 U11348 ( .A1(n12577), .A2(n11730), .ZN(n11155) );
  NOR4_X1 U11349 ( .A1(n19905), .A2(n19855), .A3(n21425), .A4(n22088), .ZN(
        n18691) );
  NOR2_X1 U11350 ( .A1(n14029), .A2(n18897), .ZN(n14034) );
  OAI221_X1 U11351 ( .B1(n18589), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18689), 
        .C2(n21557), .A(n18588), .ZN(P3_U2676) );
  OR2_X1 U11352 ( .A1(n11858), .A2(n11856), .ZN(n20194) );
  OR2_X2 U11353 ( .A1(n15274), .A2(n12677), .ZN(n11858) );
  AND2_X1 U11354 ( .A1(n11736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11156) );
  AND2_X1 U11355 ( .A1(n11736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11157) );
  AND2_X1 U11356 ( .A1(n11736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11203) );
  NOR3_X4 U11357 ( .A1(n12031), .A2(n12029), .A3(n12013), .ZN(n12039) );
  NAND2_X2 U11358 ( .A1(n12016), .A2(n12017), .ZN(n12031) );
  NAND2_X2 U11359 ( .A1(n15312), .A2(n11512), .ZN(n11536) );
  NAND2_X2 U11360 ( .A1(n15485), .A2(n15484), .ZN(n15486) );
  NAND2_X2 U11361 ( .A1(n11416), .A2(n12161), .ZN(n12167) );
  NAND2_X4 U11362 ( .A1(n12378), .A2(n12377), .ZN(n12529) );
  AND2_X2 U11363 ( .A1(n12039), .A2(n12040), .ZN(n12033) );
  NOR2_X2 U11364 ( .A1(n14905), .A2(n11468), .ZN(n15092) );
  INV_X1 U11365 ( .A(n14024), .ZN(n21214) );
  INV_X4 U11366 ( .A(n15311), .ZN(n12937) );
  NAND3_X2 U11367 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15311) );
  INV_X1 U11368 ( .A(n21628), .ZN(n21015) );
  XNOR2_X2 U11369 ( .A(n13367), .B(n13368), .ZN(n13558) );
  AND2_X2 U11370 ( .A1(n13027), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11390) );
  BUF_X4 U11371 ( .A(n18408), .Z(n11158) );
  OAI21_X2 U11374 ( .B1(n15565), .B2(n12114), .A(n16450), .ZN(n11979) );
  AND2_X4 U11375 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14713) );
  NOR2_X2 U11376 ( .A1(n15035), .A2(n15029), .ZN(n22333) );
  XNOR2_X2 U11377 ( .A(n11993), .B(n18068), .ZN(n17703) );
  NAND2_X2 U11378 ( .A1(n11950), .A2(n19287), .ZN(n11993) );
  AND2_X4 U11379 ( .A1(n13217), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13038) );
  AOI21_X2 U11380 ( .B1(n18730), .B2(n18729), .A(n18728), .ZN(n18769) );
  XNOR2_X2 U11381 ( .A(n12158), .B(n12159), .ZN(n16272) );
  AOI21_X1 U11382 ( .B1(n16477), .B2(n20860), .A(n14021), .ZN(n14022) );
  NAND2_X1 U11383 ( .A1(n12987), .A2(n12986), .ZN(n19476) );
  CLKBUF_X1 U11384 ( .A(n16517), .Z(n16518) );
  CLKBUF_X1 U11385 ( .A(n16543), .Z(n16544) );
  OR2_X1 U11386 ( .A1(n12982), .A2(n14181), .ZN(n19458) );
  CLKBUF_X1 U11387 ( .A(n16593), .Z(n16594) );
  AND2_X1 U11388 ( .A1(n17267), .A2(n16403), .ZN(n14180) );
  NAND2_X1 U11389 ( .A1(n12553), .A2(n12552), .ZN(n17484) );
  NAND2_X1 U11390 ( .A1(n15092), .A2(n12698), .ZN(n15192) );
  CLKBUF_X1 U11391 ( .A(n12168), .Z(n12179) );
  INV_X1 U11392 ( .A(n18935), .ZN(n18898) );
  INV_X4 U11393 ( .A(n19141), .ZN(n19097) );
  AND2_X2 U11394 ( .A1(n17951), .A2(n17950), .ZN(n17326) );
  OAI22_X1 U11395 ( .A1(n12866), .A2(n20194), .B1(n11931), .B2(n11896), .ZN(
        n11897) );
  NAND2_X1 U11396 ( .A1(n14914), .A2(n14924), .ZN(n14923) );
  OR2_X2 U11397 ( .A1(n11858), .A2(n11860), .ZN(n11918) );
  OR2_X1 U11398 ( .A1(n11859), .A2(n11851), .ZN(n11236) );
  INV_X1 U11399 ( .A(n15274), .ZN(n11162) );
  INV_X1 U11400 ( .A(n22333), .ZN(n22373) );
  BUF_X1 U11401 ( .A(n14903), .Z(n11223) );
  AND2_X1 U11402 ( .A1(n11296), .A2(n11251), .ZN(n19020) );
  OR2_X1 U11404 ( .A1(n14961), .A2(n13222), .ZN(n13263) );
  AND2_X1 U11405 ( .A1(n13158), .A2(n13157), .ZN(n13169) );
  NAND2_X1 U11406 ( .A1(n11187), .A2(n15026), .ZN(n14710) );
  NOR2_X1 U11407 ( .A1(n21467), .A2(n16239), .ZN(n21934) );
  INV_X2 U11408 ( .A(n12529), .ZN(n12379) );
  INV_X4 U11409 ( .A(n11961), .ZN(n12114) );
  CLKBUF_X2 U11410 ( .A(n12403), .Z(n12563) );
  AOI211_X1 U11412 ( .C1(n18712), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n14098), .B(n14097), .ZN(n14099) );
  NOR2_X2 U11413 ( .A1(n15025), .A2(n11221), .ZN(n13166) );
  CLKBUF_X1 U11414 ( .A(n13170), .Z(n14977) );
  NAND2_X2 U11415 ( .A1(n13091), .A2(n11240), .ZN(n13153) );
  BUF_X2 U11417 ( .A(n13093), .Z(n14411) );
  AND3_X1 U11418 ( .A1(n13090), .A2(n13089), .A3(n11509), .ZN(n11240) );
  CLKBUF_X2 U11419 ( .A(n14102), .Z(n18708) );
  AND4_X1 U11420 ( .A1(n13069), .A2(n13068), .A3(n13067), .A4(n13066), .ZN(
        n13070) );
  CLKBUF_X2 U11421 ( .A(n16155), .Z(n18712) );
  BUF_X2 U11422 ( .A(n14067), .Z(n18707) );
  BUF_X2 U11423 ( .A(n13136), .Z(n13985) );
  BUF_X2 U11424 ( .A(n16134), .Z(n18524) );
  CLKBUF_X2 U11425 ( .A(n13126), .Z(n13993) );
  BUF_X2 U11426 ( .A(n14079), .Z(n18711) );
  CLKBUF_X2 U11427 ( .A(n13081), .Z(n13963) );
  CLKBUF_X2 U11428 ( .A(n13179), .Z(n13988) );
  CLKBUF_X2 U11429 ( .A(n20708), .Z(n22130) );
  CLKBUF_X2 U11430 ( .A(n13137), .Z(n13986) );
  CLKBUF_X2 U11431 ( .A(n13117), .Z(n13987) );
  NAND2_X2 U11432 ( .A1(n11541), .A2(n15277), .ZN(n12934) );
  INV_X4 U11433 ( .A(n11536), .ZN(n12938) );
  AND2_X2 U11434 ( .A1(n12968), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11566) );
  AND2_X2 U11435 ( .A1(n12130), .A2(n11512), .ZN(n11213) );
  INV_X4 U11436 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21609) );
  NAND2_X4 U11437 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21638) );
  AOI21_X1 U11438 ( .B1(n12634), .B2(n18200), .A(n12633), .ZN(n12641) );
  AOI211_X1 U11439 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17890), .A(
        n17889), .B(n17888), .ZN(n17891) );
  OR2_X1 U11440 ( .A1(n17852), .A2(n18184), .ZN(n12665) );
  OAI211_X1 U11441 ( .C1(n12626), .C2(n12629), .A(n12627), .B(n13021), .ZN(
        n12118) );
  XNOR2_X1 U11442 ( .A(n14198), .B(n12097), .ZN(n17555) );
  OR2_X1 U11443 ( .A1(n17608), .A2(n17607), .ZN(n17825) );
  NAND2_X1 U11444 ( .A1(n12196), .A2(n12195), .ZN(n14207) );
  OAI21_X1 U11445 ( .B1(n16956), .B2(n11500), .A(n14216), .ZN(n14217) );
  AND2_X1 U11446 ( .A1(n11449), .A2(n11451), .ZN(n17363) );
  OAI21_X1 U11447 ( .B1(n17655), .B2(n17652), .A(n17651), .ZN(n17638) );
  NAND2_X1 U11448 ( .A1(n12194), .A2(n11272), .ZN(n17565) );
  AOI21_X1 U11449 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14440), .A(
        n14439), .ZN(n14441) );
  NAND2_X1 U11450 ( .A1(n17661), .A2(n12649), .ZN(n17655) );
  NAND2_X1 U11451 ( .A1(n17591), .A2(n17590), .ZN(n17589) );
  NAND2_X1 U11452 ( .A1(n18016), .A2(n11230), .ZN(n11441) );
  OAI21_X1 U11453 ( .B1(n14209), .B2(n14211), .A(n14210), .ZN(n16506) );
  NAND2_X1 U11454 ( .A1(n12639), .A2(n12638), .ZN(n19478) );
  CLKBUF_X1 U11455 ( .A(n14468), .Z(n14469) );
  OAI21_X1 U11456 ( .B1(n16830), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16956), .ZN(n13430) );
  NAND2_X1 U11457 ( .A1(n18053), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18054) );
  AND2_X1 U11458 ( .A1(n11329), .A2(n12185), .ZN(n11194) );
  NAND2_X1 U11459 ( .A1(n11447), .A2(n12177), .ZN(n18053) );
  OAI21_X1 U11460 ( .B1(n17395), .B2(n11268), .A(n11458), .ZN(n12885) );
  INV_X1 U11461 ( .A(n11180), .ZN(n16606) );
  CLKBUF_X1 U11462 ( .A(n12178), .Z(n11190) );
  NAND2_X1 U11463 ( .A1(n11277), .A2(n13424), .ZN(n16869) );
  AND2_X2 U11464 ( .A1(n11229), .A2(n16646), .ZN(n16645) );
  INV_X1 U11465 ( .A(n17482), .ZN(n12553) );
  NOR2_X1 U11466 ( .A1(n21923), .A2(n21922), .ZN(n21933) );
  AND2_X2 U11467 ( .A1(n16299), .A2(n11475), .ZN(n11229) );
  XNOR2_X1 U11468 ( .A(n14356), .B(n14355), .ZN(n16677) );
  NAND2_X1 U11469 ( .A1(n11302), .A2(n11988), .ZN(n11301) );
  NAND2_X1 U11470 ( .A1(n20849), .A2(n13402), .ZN(n16343) );
  AND2_X2 U11471 ( .A1(n16253), .A2(n12699), .ZN(n16367) );
  OR2_X1 U11472 ( .A1(n18914), .A2(n19044), .ZN(n11297) );
  NOR2_X1 U11473 ( .A1(n12658), .A2(n12659), .ZN(n11389) );
  NAND2_X1 U11474 ( .A1(n15563), .A2(n12157), .ZN(n12158) );
  NAND2_X1 U11475 ( .A1(n17311), .A2(n17312), .ZN(n12658) );
  NAND2_X1 U11476 ( .A1(n12155), .A2(n12154), .ZN(n15563) );
  INV_X1 U11477 ( .A(n17548), .ZN(n12538) );
  NAND3_X1 U11478 ( .A1(n12142), .A2(n12143), .A3(n11448), .ZN(n12162) );
  OAI21_X1 U11479 ( .B1(n15495), .B2(n15497), .A(n15496), .ZN(n20262) );
  OR2_X1 U11480 ( .A1(n16379), .A2(n11237), .ZN(n11278) );
  NAND2_X1 U11481 ( .A1(n21322), .A2(n21323), .ZN(n21321) );
  XNOR2_X1 U11482 ( .A(n16955), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16379) );
  NAND2_X1 U11483 ( .A1(n15664), .A2(n11379), .ZN(n11382) );
  AND2_X1 U11484 ( .A1(n16920), .A2(n13420), .ZN(n16899) );
  OR2_X1 U11485 ( .A1(n17310), .A2(n11961), .ZN(n12046) );
  AND2_X1 U11486 ( .A1(n11944), .A2(n11943), .ZN(n12181) );
  AND2_X1 U11487 ( .A1(n12068), .A2(n12067), .ZN(n12075) );
  NAND2_X1 U11488 ( .A1(n21313), .A2(n21314), .ZN(n21312) );
  OAI21_X1 U11489 ( .B1(n21012), .B2(n18980), .A(n19653), .ZN(n18935) );
  NAND2_X1 U11490 ( .A1(n15640), .A2(n15639), .ZN(n15666) );
  OR3_X1 U11491 ( .A1(n12048), .A2(n11961), .A3(n17866), .ZN(n17639) );
  NAND2_X1 U11492 ( .A1(n14933), .A2(n13527), .ZN(n15172) );
  AND2_X1 U11493 ( .A1(n14928), .A2(n11254), .ZN(n15640) );
  NAND2_X1 U11494 ( .A1(n19142), .A2(n19097), .ZN(n18980) );
  AND2_X1 U11495 ( .A1(n17669), .A2(n12026), .ZN(n12644) );
  NAND2_X1 U11496 ( .A1(n13364), .A2(n13363), .ZN(n13365) );
  NOR2_X2 U11497 ( .A1(n14923), .A2(n14929), .ZN(n14928) );
  NAND2_X1 U11498 ( .A1(n13380), .A2(n13379), .ZN(n13394) );
  NAND2_X1 U11499 ( .A1(n11861), .A2(n11828), .ZN(n20065) );
  NAND2_X1 U11500 ( .A1(n11241), .A2(n12694), .ZN(n15497) );
  OAI22_X1 U11501 ( .A1(n11853), .A2(n15509), .B1(n11236), .B2(n11852), .ZN(
        n11854) );
  NAND2_X1 U11502 ( .A1(n21287), .A2(n21288), .ZN(n21286) );
  OR2_X1 U11503 ( .A1(n11857), .A2(n11856), .ZN(n11926) );
  NAND2_X1 U11504 ( .A1(n19082), .A2(n21459), .ZN(n18965) );
  NOR2_X1 U11505 ( .A1(n14915), .A2(n14916), .ZN(n14914) );
  NAND2_X1 U11506 ( .A1(n17989), .A2(n17990), .ZN(n17991) );
  NAND2_X1 U11507 ( .A1(n11280), .A2(n11279), .ZN(n13382) );
  INV_X1 U11508 ( .A(n11162), .ZN(n11196) );
  AND2_X2 U11509 ( .A1(n18733), .A2(n22115), .ZN(n22124) );
  OR2_X1 U11510 ( .A1(n11859), .A2(n11856), .ZN(n11927) );
  AND2_X1 U11511 ( .A1(n11239), .A2(n11828), .ZN(n15716) );
  NAND2_X1 U11512 ( .A1(n11495), .A2(n11263), .ZN(n17098) );
  NAND2_X1 U11513 ( .A1(n11239), .A2(n11846), .ZN(n15509) );
  NAND2_X1 U11514 ( .A1(n13538), .A2(n13537), .ZN(n15173) );
  NAND2_X1 U11515 ( .A1(n14910), .A2(n14909), .ZN(n14915) );
  NAND2_X1 U11516 ( .A1(n13515), .A2(n13514), .ZN(n14885) );
  OR2_X1 U11517 ( .A1(n18752), .A2(n22012), .ZN(n18751) );
  AOI22_X1 U11518 ( .A1(n14471), .A2(n19251), .B1(n14472), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14531) );
  OR2_X1 U11519 ( .A1(n19505), .A2(n17360), .ZN(n11856) );
  NOR2_X2 U11520 ( .A1(n15199), .A2(n15198), .ZN(n15197) );
  NAND2_X1 U11521 ( .A1(n16584), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15035) );
  AND2_X1 U11522 ( .A1(n16705), .A2(n16698), .ZN(n16699) );
  NOR2_X2 U11523 ( .A1(n16707), .A2(n16706), .ZN(n16705) );
  OR2_X1 U11524 ( .A1(n19046), .A2(n18748), .ZN(n11296) );
  NOR2_X1 U11525 ( .A1(n15141), .A2(n15140), .ZN(n22773) );
  NAND2_X2 U11526 ( .A1(n16791), .A2(n14882), .ZN(n16782) );
  NAND2_X1 U11527 ( .A1(n14415), .A2(n14414), .ZN(n16791) );
  INV_X1 U11528 ( .A(n19505), .ZN(n15304) );
  OR2_X1 U11529 ( .A1(n16303), .A2(n16350), .ZN(n16707) );
  NOR2_X1 U11530 ( .A1(n11235), .A2(n13017), .ZN(n13016) );
  NAND2_X1 U11531 ( .A1(n13257), .A2(n13404), .ZN(n13509) );
  AND2_X1 U11532 ( .A1(n14943), .A2(n16463), .ZN(n14623) );
  OR2_X1 U11533 ( .A1(n18127), .A2(n14621), .ZN(n14943) );
  NOR2_X2 U11534 ( .A1(n20213), .A2(n20525), .ZN(n20214) );
  NOR2_X2 U11535 ( .A1(n20269), .A2(n20527), .ZN(n20270) );
  OR2_X2 U11536 ( .A1(n16463), .A2(n11221), .ZN(n14808) );
  NAND2_X1 U11537 ( .A1(n13272), .A2(n13271), .ZN(n14740) );
  AND2_X1 U11538 ( .A1(n12200), .A2(n11816), .ZN(n12201) );
  OR2_X1 U11539 ( .A1(n13272), .A2(n13271), .ZN(n11484) );
  NOR2_X2 U11540 ( .A1(n20037), .A2(n20525), .ZN(n15512) );
  NOR2_X2 U11541 ( .A1(n20817), .A2(n20816), .ZN(n20819) );
  NAND2_X1 U11542 ( .A1(n11824), .A2(n11823), .ZN(n11826) );
  INV_X2 U11543 ( .A(n17411), .ZN(n17432) );
  OR2_X1 U11544 ( .A1(n20825), .A2(n15661), .ZN(n20817) );
  NAND2_X1 U11545 ( .A1(n13207), .A2(n13206), .ZN(n13255) );
  NAND2_X1 U11546 ( .A1(n18204), .A2(n12315), .ZN(n18190) );
  NAND2_X1 U11547 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  NAND2_X1 U11548 ( .A1(n13302), .A2(n13301), .ZN(n15211) );
  NOR2_X1 U11549 ( .A1(n20990), .A2(n20951), .ZN(n21001) );
  NAND3_X1 U11550 ( .A1(n11790), .A2(n11789), .A3(n11788), .ZN(n11821) );
  CLKBUF_X1 U11551 ( .A(n13518), .Z(n11176) );
  OR2_X1 U11552 ( .A1(n13296), .A2(n13030), .ZN(n13270) );
  OR2_X2 U11553 ( .A1(n14514), .A2(n14473), .ZN(n14475) );
  INV_X2 U11554 ( .A(n20951), .ZN(n21004) );
  AOI21_X1 U11555 ( .B1(n11157), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11795), .ZN(n11798) );
  OR2_X1 U11556 ( .A1(n13296), .A2(n13027), .ZN(n13302) );
  OR2_X1 U11557 ( .A1(n11787), .A2(n19251), .ZN(n11788) );
  CLKBUF_X1 U11558 ( .A(n18691), .Z(n11217) );
  AOI22_X1 U11559 ( .A1(n12371), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12317), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11763) );
  OAI211_X1 U11560 ( .C1(n13177), .C2(n13176), .A(n13175), .B(n13174), .ZN(
        n13215) );
  NOR2_X2 U11561 ( .A1(n14036), .A2(n18903), .ZN(n14035) );
  NAND2_X1 U11562 ( .A1(n14950), .A2(n14949), .ZN(n15373) );
  AND4_X1 U11563 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n15558) );
  OAI211_X1 U11564 ( .C1(n14836), .C2(n11794), .A(n11741), .B(n11740), .ZN(
        n11742) );
  NAND2_X1 U11565 ( .A1(n13220), .A2(n11245), .ZN(n11396) );
  BUF_X4 U11566 ( .A(n11807), .Z(n12306) );
  MUX2_X1 U11567 ( .A(n12134), .B(P2_EBX_REG_2__SCAN_IN), .S(n20269), .Z(
        n11974) );
  MUX2_X1 U11568 ( .A(n11747), .B(n12582), .S(n12584), .Z(n11785) );
  NAND3_X2 U11569 ( .A1(n21934), .A2(n21932), .A3(n21673), .ZN(n19044) );
  AND3_X1 U11570 ( .A1(n12573), .A2(n11429), .A3(n11252), .ZN(n12565) );
  AND2_X1 U11571 ( .A1(n12149), .A2(n11738), .ZN(n11346) );
  MUX2_X1 U11572 ( .A(n12358), .B(n12352), .S(n12357), .Z(n11745) );
  NOR2_X1 U11573 ( .A1(n19692), .A2(n21487), .ZN(n16123) );
  AND2_X1 U11574 ( .A1(n14706), .A2(n14363), .ZN(n13157) );
  INV_X1 U11575 ( .A(n11770), .ZN(n12575) );
  INV_X2 U11576 ( .A(n12132), .ZN(n11738) );
  INV_X1 U11577 ( .A(n12333), .ZN(n19490) );
  OR2_X1 U11578 ( .A1(n14707), .A2(n14428), .ZN(n14359) );
  OR2_X1 U11579 ( .A1(n13476), .A2(n14256), .ZN(n14706) );
  NOR2_X1 U11580 ( .A1(n13447), .A2(n14409), .ZN(n13160) );
  AND2_X1 U11581 ( .A1(n11752), .A2(n13007), .ZN(n12998) );
  AND3_X1 U11582 ( .A1(n14426), .A2(n14364), .A3(n13151), .ZN(n14357) );
  NAND2_X1 U11583 ( .A1(n18743), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18760) );
  OR2_X1 U11584 ( .A1(n21598), .A2(n21482), .ZN(n16227) );
  CLKBUF_X3 U11585 ( .A(n11743), .Z(n12377) );
  CLKBUF_X1 U11586 ( .A(n11744), .Z(n12357) );
  INV_X1 U11587 ( .A(n12954), .ZN(n12819) );
  NAND3_X1 U11588 ( .A1(n14101), .A2(n14100), .A3(n14099), .ZN(n19652) );
  OR2_X1 U11589 ( .A1(n11613), .A2(n11612), .ZN(n12416) );
  NAND3_X1 U11590 ( .A1(n14052), .A2(n14051), .A3(n14050), .ZN(n20937) );
  OR2_X1 U11591 ( .A1(n11550), .A2(n11549), .ZN(n12149) );
  AND2_X1 U11592 ( .A1(n13167), .A2(n14966), .ZN(n14364) );
  OR2_X1 U11593 ( .A1(n11598), .A2(n11597), .ZN(n11909) );
  OR2_X1 U11594 ( .A1(n11884), .A2(n11883), .ZN(n12375) );
  NAND2_X1 U11595 ( .A1(n12376), .A2(n20165), .ZN(n12382) );
  NOR2_X1 U11596 ( .A1(n12376), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12402) );
  NAND2_X2 U11597 ( .A1(n11694), .A2(n11693), .ZN(n13007) );
  AND4_X1 U11598 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11653) );
  INV_X2 U11599 ( .A(U212), .ZN(n11164) );
  MUX2_X1 U11600 ( .A(n11681), .B(n11680), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12584) );
  NAND2_X1 U11601 ( .A1(n11517), .A2(n11713), .ZN(n11524) );
  NAND2_X1 U11602 ( .A1(n18992), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n21201) );
  NAND4_X2 U11603 ( .A1(n13149), .A2(n13148), .A3(n13147), .A4(n13146), .ZN(
        n11221) );
  AND4_X1 U11604 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11517) );
  NAND4_X1 U11605 ( .A1(n13052), .A2(n13051), .A3(n13050), .A4(n13049), .ZN(
        n13150) );
  BUF_X4 U11606 ( .A(n12129), .Z(n11206) );
  AND4_X1 U11607 ( .A1(n13085), .A2(n13084), .A3(n13083), .A4(n13082), .ZN(
        n13091) );
  NAND2_X2 U11608 ( .A1(U214), .A2(n20869), .ZN(n20933) );
  AND4_X1 U11609 ( .A1(n13109), .A2(n13108), .A3(n13107), .A4(n13106), .ZN(
        n13124) );
  AND4_X1 U11610 ( .A1(n13103), .A2(n13102), .A3(n13101), .A4(n13100), .ZN(
        n13125) );
  NAND2_X1 U11611 ( .A1(n11511), .A2(n13070), .ZN(n13093) );
  AND4_X1 U11612 ( .A1(n13034), .A2(n13033), .A3(n13032), .A4(n13031), .ZN(
        n13042) );
  AND4_X1 U11613 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11652) );
  AND4_X1 U11614 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n13148) );
  AND4_X1 U11615 ( .A1(n13141), .A2(n13140), .A3(n13139), .A4(n13138), .ZN(
        n13147) );
  AND4_X1 U11616 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13142), .ZN(
        n13146) );
  BUF_X2 U11617 ( .A(n18424), .Z(n21637) );
  AND4_X1 U11618 ( .A1(n13121), .A2(n13120), .A3(n13119), .A4(n13118), .ZN(
        n13122) );
  AND4_X1 U11619 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13051) );
  AND4_X1 U11620 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        n13123) );
  AND4_X1 U11621 ( .A1(n13056), .A2(n13055), .A3(n13054), .A4(n13053), .ZN(
        n13061) );
  AND2_X1 U11622 ( .A1(n11525), .A2(n11713), .ZN(n11529) );
  AND2_X2 U11623 ( .A1(n12969), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11871) );
  INV_X1 U11624 ( .A(n11620), .ZN(n11211) );
  INV_X1 U11625 ( .A(n11620), .ZN(n11210) );
  INV_X2 U11626 ( .A(n19227), .ZN(n19233) );
  AND2_X1 U11627 ( .A1(n11518), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11521) );
  BUF_X2 U11628 ( .A(n16134), .Z(n18705) );
  NAND2_X1 U11629 ( .A1(n19060), .A2(n14023), .ZN(n21115) );
  INV_X2 U11630 ( .A(n22435), .ZN(n18306) );
  BUF_X2 U11631 ( .A(n11201), .Z(n12969) );
  AND2_X1 U11632 ( .A1(n11315), .A2(n11314), .ZN(n11533) );
  BUF_X2 U11633 ( .A(n14092), .Z(n18660) );
  BUF_X2 U11634 ( .A(n14079), .Z(n21034) );
  CLKBUF_X3 U11635 ( .A(n11715), .Z(n12970) );
  BUF_X2 U11636 ( .A(n16155), .Z(n18397) );
  NAND2_X2 U11637 ( .A1(n22113), .A2(n18696), .ZN(n18767) );
  BUF_X2 U11638 ( .A(n14068), .Z(n18714) );
  NAND2_X2 U11639 ( .A1(n22787), .A2(n20720), .ZN(n20776) );
  NAND2_X2 U11640 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22787), .ZN(n20772) );
  INV_X2 U11641 ( .A(n20643), .ZN(n20693) );
  AND2_X1 U11642 ( .A1(n19006), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19060) );
  AND2_X2 U11643 ( .A1(n12796), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11878) );
  NAND2_X1 U11644 ( .A1(n12937), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11620) );
  AND2_X2 U11645 ( .A1(n13036), .A2(n13037), .ZN(n13104) );
  AND2_X2 U11646 ( .A1(n11543), .A2(n12797), .ZN(n11591) );
  NOR2_X1 U11647 ( .A1(n14042), .A2(n14040), .ZN(n18408) );
  BUF_X4 U11648 ( .A(n14090), .Z(n11165) );
  OR2_X2 U11649 ( .A1(n14019), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16939) );
  INV_X1 U11650 ( .A(n12944), .ZN(n11218) );
  AND2_X2 U11651 ( .A1(n12968), .A2(n11713), .ZN(n11607) );
  AND2_X2 U11652 ( .A1(n13036), .A2(n17222), .ZN(n13131) );
  NOR2_X1 U11653 ( .A1(n19086), .A2(n19085), .ZN(n19006) );
  INV_X1 U11654 ( .A(n21639), .ZN(n14040) );
  AND2_X1 U11655 ( .A1(n13029), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13036) );
  AND2_X2 U11656 ( .A1(n12130), .A2(n11512), .ZN(n12796) );
  AND2_X2 U11657 ( .A1(n14712), .A2(n14897), .ZN(n13110) );
  AND2_X2 U11658 ( .A1(n13030), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17222) );
  INV_X1 U11659 ( .A(n11213), .ZN(n11166) );
  AND2_X2 U11660 ( .A1(n12797), .A2(n11542), .ZN(n11590) );
  AND2_X2 U11661 ( .A1(n12797), .A2(n11544), .ZN(n11592) );
  NOR2_X2 U11662 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11544) );
  NOR2_X1 U11663 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12797) );
  INV_X1 U11664 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13217) );
  CLKBUF_X1 U11665 ( .A(n17610), .Z(n11167) );
  INV_X1 U11666 ( .A(n15300), .ZN(n11168) );
  NAND2_X1 U11667 ( .A1(n11762), .A2(n11155), .ZN(n12371) );
  NAND2_X1 U11668 ( .A1(n17609), .A2(n17611), .ZN(n17610) );
  AND2_X1 U11669 ( .A1(n11726), .A2(n12998), .ZN(n11169) );
  AND2_X2 U11670 ( .A1(n11726), .A2(n12998), .ZN(n11756) );
  AND2_X1 U11671 ( .A1(n11755), .A2(n11732), .ZN(n11726) );
  NOR2_X2 U11672 ( .A1(n21256), .A2(n18667), .ZN(n18584) );
  BUF_X4 U11673 ( .A(n18424), .Z(n14127) );
  NAND2_X1 U11674 ( .A1(n20837), .A2(n11173), .ZN(n11170) );
  OR2_X1 U11675 ( .A1(n11172), .A2(n20844), .ZN(n11171) );
  INV_X1 U11676 ( .A(n13390), .ZN(n11172) );
  AND2_X1 U11677 ( .A1(n13366), .A2(n13390), .ZN(n11173) );
  NAND2_X1 U11678 ( .A1(n15171), .A2(n15170), .ZN(n11174) );
  NOR2_X1 U11679 ( .A1(n16806), .A2(n11492), .ZN(n11175) );
  NAND2_X1 U11680 ( .A1(n15171), .A2(n15170), .ZN(n15169) );
  NOR2_X1 U11681 ( .A1(n16806), .A2(n11492), .ZN(n13439) );
  XNOR2_X1 U11682 ( .A(n13216), .B(n13178), .ZN(n13518) );
  INV_X1 U11683 ( .A(n11817), .ZN(n11177) );
  INV_X1 U11684 ( .A(n11177), .ZN(n11178) );
  NAND2_X1 U11685 ( .A1(n11768), .A2(n11767), .ZN(n11817) );
  NAND2_X1 U11686 ( .A1(n13240), .A2(n13239), .ZN(n13242) );
  AND2_X1 U11687 ( .A1(n13776), .A2(n16777), .ZN(n11179) );
  NAND2_X1 U11688 ( .A1(n16645), .A2(n16777), .ZN(n11180) );
  CLKBUF_X1 U11689 ( .A(n15349), .Z(n11181) );
  NAND3_X2 U11690 ( .A1(n11735), .A2(n11155), .A3(n11773), .ZN(n11736) );
  NAND2_X1 U11691 ( .A1(n11305), .A2(n11885), .ZN(n11965) );
  INV_X1 U11692 ( .A(n11804), .ZN(n11322) );
  INV_X1 U11693 ( .A(n15140), .ZN(n11182) );
  INV_X1 U11694 ( .A(n14999), .ZN(n11183) );
  OR2_X2 U11695 ( .A1(n11188), .A2(n11189), .ZN(n14410) );
  AND2_X2 U11696 ( .A1(n18856), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14028) );
  AND2_X2 U11697 ( .A1(n14712), .A2(n13037), .ZN(n13137) );
  OR3_X4 U11698 ( .A1(n16105), .A2(n16127), .A3(n21620), .ZN(n18086) );
  INV_X1 U11699 ( .A(n14531), .ZN(n11184) );
  INV_X1 U11700 ( .A(n11184), .ZN(n11185) );
  INV_X1 U11701 ( .A(n11184), .ZN(n11186) );
  INV_X1 U11702 ( .A(n11187), .ZN(n14238) );
  OR4_X1 U11703 ( .A1(n21486), .A2(n16105), .A3(n14141), .A4(n19905), .ZN(
        n14139) );
  NOR3_X2 U11704 ( .A1(n21587), .A2(n21433), .A3(n21432), .ZN(n21575) );
  NOR2_X2 U11705 ( .A1(n11999), .A2(n11998), .ZN(n11997) );
  AND2_X2 U11706 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12130) );
  XNOR2_X2 U11707 ( .A(n12086), .B(n12087), .ZN(n12100) );
  AND2_X2 U11708 ( .A1(n14372), .A2(n15130), .ZN(n11187) );
  OR2_X2 U11709 ( .A1(n12636), .A2(n12637), .ZN(n12639) );
  NOR2_X2 U11710 ( .A1(n11382), .A2(n11257), .ZN(n17438) );
  NOR2_X2 U11711 ( .A1(n17270), .A2(n17271), .ZN(n14201) );
  NAND4_X1 U11712 ( .A1(n13074), .A2(n13073), .A3(n13072), .A4(n13071), .ZN(
        n11188) );
  NAND4_X1 U11713 ( .A1(n13078), .A2(n13077), .A3(n13076), .A4(n13075), .ZN(
        n11189) );
  NOR2_X4 U11714 ( .A1(n21616), .A2(n21621), .ZN(n21884) );
  AND2_X2 U11715 ( .A1(n17297), .A2(n17298), .ZN(n17283) );
  NOR2_X2 U11716 ( .A1(n17991), .A2(n17343), .ZN(n17951) );
  NOR2_X2 U11717 ( .A1(n17503), .A2(n12546), .ZN(n17297) );
  NAND2_X1 U11718 ( .A1(n18054), .A2(n11194), .ZN(n11191) );
  AND2_X2 U11719 ( .A1(n11191), .A2(n11192), .ZN(n18016) );
  OR2_X1 U11720 ( .A1(n11193), .A2(n17738), .ZN(n11192) );
  INV_X1 U11721 ( .A(n12185), .ZN(n11193) );
  NOR2_X2 U11722 ( .A1(n17878), .A2(n12654), .ZN(n11195) );
  OAI21_X1 U11723 ( .B1(n11760), .B2(n11771), .A(n11759), .ZN(n11197) );
  NOR2_X1 U11724 ( .A1(n17878), .A2(n12654), .ZN(n17645) );
  OAI21_X1 U11725 ( .B1(n11760), .B2(n11771), .A(n11759), .ZN(n11806) );
  NAND2_X1 U11726 ( .A1(n11306), .A2(n11910), .ZN(n11966) );
  AOI21_X2 U11727 ( .B1(n12642), .B2(n12061), .A(n12060), .ZN(n17609) );
  INV_X2 U11728 ( .A(n16861), .ZN(n13431) );
  AND2_X2 U11729 ( .A1(n16857), .A2(n16858), .ZN(n16861) );
  AND2_X2 U11730 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n18611), .ZN(n18605) );
  NOR2_X2 U11731 ( .A1(n21326), .A2(n18606), .ZN(n18611) );
  NOR4_X4 U11732 ( .A1(n21571), .A2(n21520), .A3(n21519), .A4(n21518), .ZN(
        n21565) );
  NAND2_X2 U11733 ( .A1(n21579), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21571) );
  NAND2_X1 U11734 ( .A1(n14710), .A2(n13152), .ZN(n14222) );
  INV_X1 U11735 ( .A(n11965), .ZN(n12142) );
  OAI21_X1 U11736 ( .B1(n16606), .B2(n16636), .A(n16635), .ZN(n16911) );
  NAND2_X1 U11737 ( .A1(n11825), .A2(n11834), .ZN(n17360) );
  OR2_X1 U11738 ( .A1(n11825), .A2(n11827), .ZN(n11860) );
  AOI21_X2 U11739 ( .B1(n11156), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11742), .ZN(n11768) );
  AND2_X1 U11740 ( .A1(n14897), .A2(n14713), .ZN(n11198) );
  AND2_X1 U11741 ( .A1(n14897), .A2(n14713), .ZN(n11199) );
  OAI211_X1 U11743 ( .C1(n14871), .C2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11392), .B(n11391), .ZN(n14940) );
  INV_X2 U11744 ( .A(n11743), .ZN(n11752) );
  AND2_X2 U11745 ( .A1(n13203), .A2(n14410), .ZN(n13448) );
  INV_X1 U11746 ( .A(n12944), .ZN(n11200) );
  BUF_X4 U11747 ( .A(n11682), .Z(n11201) );
  AOI21_X2 U11748 ( .B1(n11784), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11779), 
        .ZN(n11759) );
  AND2_X1 U11749 ( .A1(n11736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11202) );
  NOR2_X2 U11750 ( .A1(n21152), .A2(n18448), .ZN(n18420) );
  INV_X1 U11751 ( .A(n12934), .ZN(n11204) );
  INV_X1 U11752 ( .A(n12934), .ZN(n11205) );
  NAND2_X2 U11753 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21609), .ZN(
        n14042) );
  NAND2_X2 U11754 ( .A1(n13079), .A2(n14239), .ZN(n13161) );
  INV_X2 U11755 ( .A(n11536), .ZN(n11207) );
  NAND2_X2 U11756 ( .A1(n11732), .A2(n11743), .ZN(n11746) );
  NAND2_X1 U11757 ( .A1(n11397), .A2(n13164), .ZN(n13216) );
  NOR2_X2 U11758 ( .A1(n22116), .A2(n18086), .ZN(n18319) );
  NAND2_X1 U11759 ( .A1(n16272), .A2(n16325), .ZN(n11416) );
  AND2_X1 U11760 ( .A1(n14897), .A2(n14713), .ZN(n11208) );
  AND2_X1 U11761 ( .A1(n14897), .A2(n14713), .ZN(n11209) );
  OR2_X2 U11762 ( .A1(n11857), .A2(n11851), .ZN(n11912) );
  AND2_X1 U11763 ( .A1(n13150), .A2(n13092), .ZN(n13079) );
  NAND2_X1 U11764 ( .A1(n14411), .A2(n13150), .ZN(n14428) );
  NOR3_X4 U11765 ( .A1(n14475), .A2(n17583), .A3(n17574), .ZN(n14518) );
  XNOR2_X1 U11766 ( .A(n13255), .B(n13254), .ZN(n13516) );
  NOR2_X4 U11767 ( .A1(n17930), .A2(n17908), .ZN(n17896) );
  NOR2_X2 U11768 ( .A1(n14505), .A2(n19358), .ZN(n14507) );
  AND2_X1 U11769 ( .A1(n12130), .A2(n11512), .ZN(n11214) );
  INV_X2 U11770 ( .A(n12934), .ZN(n11216) );
  NAND2_X1 U11771 ( .A1(n13263), .A2(n15434), .ZN(n14705) );
  INV_X1 U11773 ( .A(n12944), .ZN(n11219) );
  NAND2_X2 U11774 ( .A1(n11542), .A2(n15277), .ZN(n12944) );
  NOR2_X2 U11775 ( .A1(n15673), .A2(n16262), .ZN(n16263) );
  NOR2_X2 U11776 ( .A1(n15251), .A2(n15653), .ZN(n15652) );
  AND2_X2 U11777 ( .A1(n12969), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11220) );
  NOR2_X2 U11778 ( .A1(n16543), .A2(n16545), .ZN(n16529) );
  NAND4_X1 U11779 ( .A1(n13149), .A2(n13148), .A3(n13147), .A4(n13146), .ZN(
        n13156) );
  NOR2_X1 U11780 ( .A1(n13220), .A2(n22396), .ZN(n13260) );
  XNOR2_X1 U11781 ( .A(n13510), .B(n13509), .ZN(n14903) );
  AND2_X1 U11782 ( .A1(n13038), .A2(n13037), .ZN(n11224) );
  AND2_X1 U11783 ( .A1(n17222), .A2(n14713), .ZN(n11226) );
  AND2_X2 U11784 ( .A1(n17222), .A2(n14713), .ZN(n13086) );
  OAI21_X1 U11785 ( .B1(n16465), .B2(n14551), .A(n14359), .ZN(n11274) );
  INV_X1 U11786 ( .A(n13345), .ZN(n11280) );
  NAND2_X1 U11787 ( .A1(n11396), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13264) );
  NOR2_X1 U11788 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13773) );
  OR2_X1 U11789 ( .A1(n14411), .A2(n22489), .ZN(n13701) );
  OR2_X1 U11790 ( .A1(n11182), .A2(n22489), .ZN(n13519) );
  INV_X1 U11791 ( .A(n13322), .ZN(n11410) );
  OR2_X1 U11792 ( .A1(n13202), .A2(n13201), .ZN(n13237) );
  NAND2_X1 U11793 ( .A1(n13263), .A2(n13262), .ZN(n13272) );
  OAI21_X1 U11794 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13261), .A(
        n13260), .ZN(n13262) );
  INV_X1 U11795 ( .A(n13773), .ZN(n13982) );
  NAND2_X1 U11796 ( .A1(n11951), .A2(n11962), .ZN(n11960) );
  NAND2_X1 U11797 ( .A1(n11728), .A2(n11727), .ZN(n11770) );
  NAND2_X1 U11798 ( .A1(n17684), .A2(n17683), .ZN(n17668) );
  OR2_X1 U11799 ( .A1(n11995), .A2(n11996), .ZN(n11439) );
  NAND2_X1 U11800 ( .A1(n19020), .A2(n11295), .ZN(n18791) );
  AND2_X1 U11801 ( .A1(n19022), .A2(n22024), .ZN(n11295) );
  INV_X1 U11802 ( .A(n13519), .ZN(n14010) );
  AND2_X1 U11803 ( .A1(n22489), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14009) );
  NAND2_X1 U11804 ( .A1(n14345), .A2(n14256), .ZN(n14814) );
  AND2_X1 U11805 ( .A1(n16850), .A2(n16994), .ZN(n11411) );
  NAND2_X1 U11806 ( .A1(n11453), .A2(n11452), .ZN(n11451) );
  AND2_X1 U11807 ( .A1(n12696), .A2(n12695), .ZN(n12697) );
  NOR2_X1 U11808 ( .A1(n12098), .A2(n12105), .ZN(n12106) );
  NAND2_X1 U11809 ( .A1(n13014), .A2(n13015), .ZN(n12636) );
  INV_X1 U11810 ( .A(n17565), .ZN(n12196) );
  NAND2_X1 U11811 ( .A1(n11438), .A2(n11437), .ZN(n11436) );
  INV_X1 U11812 ( .A(n17712), .ZN(n11437) );
  INV_X1 U11813 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20165) );
  AND2_X1 U11814 ( .A1(n20199), .A2(n20167), .ZN(n20195) );
  NAND2_X1 U11815 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20199), .ZN(n20527) );
  INV_X1 U11816 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20146) );
  AND2_X1 U11817 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11355) );
  AOI21_X1 U11818 ( .B1(n13223), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n11361), .ZN(n13333) );
  AND2_X1 U11819 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11361) );
  NAND2_X1 U11820 ( .A1(n15716), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11428) );
  NOR2_X1 U11821 ( .A1(n12566), .A2(n12342), .ZN(n11779) );
  AND2_X1 U11822 ( .A1(n13346), .A2(n13368), .ZN(n11279) );
  AOI21_X1 U11823 ( .B1(n13223), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11360), .ZN(n13182) );
  AND2_X1 U11824 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11360) );
  AOI21_X1 U11825 ( .B1(n13086), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n11357), .ZN(n13277) );
  AND2_X1 U11826 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11357) );
  OR3_X1 U11827 ( .A1(n12122), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n18108), .ZN(n12120) );
  INV_X1 U11828 ( .A(n17390), .ZN(n11461) );
  AND2_X1 U11829 ( .A1(n12861), .A2(n17390), .ZN(n11459) );
  NAND4_X1 U11830 ( .A1(n11752), .A2(n15513), .A3(n11725), .A4(n11729), .ZN(
        n11747) );
  NAND2_X1 U11831 ( .A1(n12182), .A2(n12181), .ZN(n12186) );
  AND2_X1 U11832 ( .A1(n19813), .A2(n14138), .ZN(n16115) );
  NAND2_X1 U11833 ( .A1(n14211), .A2(n11481), .ZN(n11480) );
  INV_X1 U11834 ( .A(n16519), .ZN(n11481) );
  AND2_X1 U11835 ( .A1(n11259), .A2(n16556), .ZN(n11472) );
  OR2_X1 U11836 ( .A1(n16625), .A2(n16634), .ZN(n16607) );
  AND2_X1 U11837 ( .A1(n13637), .A2(n16349), .ZN(n11477) );
  AND2_X1 U11838 ( .A1(n11479), .A2(n16349), .ZN(n11478) );
  INV_X1 U11839 ( .A(n16704), .ZN(n11479) );
  XNOR2_X1 U11840 ( .A(n13394), .B(n13393), .ZN(n13572) );
  NAND2_X1 U11841 ( .A1(n11280), .A2(n13346), .ZN(n13367) );
  AND2_X1 U11842 ( .A1(n13450), .A2(n13449), .ZN(n14362) );
  INV_X1 U11843 ( .A(n13411), .ZN(n11402) );
  NAND2_X1 U11844 ( .A1(n14625), .A2(n15033), .ZN(n14347) );
  INV_X1 U11845 ( .A(n13163), .ZN(n11273) );
  NOR2_X1 U11846 ( .A1(n13167), .A2(n13153), .ZN(n17198) );
  NAND2_X1 U11847 ( .A1(n13216), .A2(n13215), .ZN(n13222) );
  AOI22_X1 U11848 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13075) );
  INV_X1 U11849 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22475) );
  NAND2_X1 U11850 ( .A1(n11955), .A2(n11342), .ZN(n11341) );
  INV_X1 U11851 ( .A(n11952), .ZN(n11342) );
  NAND2_X1 U11852 ( .A1(n11333), .A2(n11615), .ZN(n11984) );
  INV_X1 U11853 ( .A(n11981), .ZN(n11333) );
  NAND2_X1 U11854 ( .A1(n17381), .A2(n12888), .ZN(n12909) );
  NAND3_X1 U11855 ( .A1(n11732), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12954), 
        .ZN(n12905) );
  NAND2_X1 U11856 ( .A1(n19249), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12342) );
  AND2_X1 U11857 ( .A1(n15194), .A2(n15087), .ZN(n11378) );
  NOR2_X2 U11858 ( .A1(n11984), .A2(n11628), .ZN(n11945) );
  INV_X1 U11859 ( .A(n11983), .ZN(n11628) );
  AND2_X1 U11860 ( .A1(n12167), .A2(n12179), .ZN(n12169) );
  AOI21_X1 U11861 ( .B1(n11202), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11811), .ZN(n11813) );
  NAND2_X1 U11862 ( .A1(n11430), .A2(n11728), .ZN(n11429) );
  NAND2_X1 U11863 ( .A1(n11801), .A2(n11802), .ZN(n11384) );
  NAND2_X1 U11864 ( .A1(n11457), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U11865 ( .A1(n11196), .A2(n15498), .ZN(n11457) );
  AND2_X1 U11866 ( .A1(n12124), .A2(n12123), .ZN(n12343) );
  OR2_X1 U11867 ( .A1(n12122), .A2(n12121), .ZN(n12124) );
  NAND2_X1 U11868 ( .A1(n11162), .A2(n12677), .ZN(n11857) );
  NAND2_X1 U11869 ( .A1(n11714), .A2(n11713), .ZN(n11722) );
  NOR2_X1 U11870 ( .A1(n14041), .A2(n14040), .ZN(n14068) );
  NOR2_X1 U11871 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21015), .ZN(
        n14102) );
  NOR2_X1 U11872 ( .A1(n21177), .A2(n21165), .ZN(n11353) );
  INV_X1 U11873 ( .A(n21939), .ZN(n11299) );
  NAND2_X1 U11874 ( .A1(n19100), .A2(n16232), .ZN(n16236) );
  NAND2_X1 U11875 ( .A1(n16227), .A2(n16223), .ZN(n16224) );
  AND3_X1 U11876 ( .A1(n19905), .A2(n19773), .A3(n21521), .ZN(n14148) );
  NAND2_X1 U11877 ( .A1(n14408), .A2(n14407), .ZN(n14720) );
  OR2_X1 U11878 ( .A1(n14620), .A2(n22389), .ZN(n14408) );
  AND2_X1 U11879 ( .A1(n14008), .A2(n14007), .ZN(n14402) );
  OR2_X1 U11880 ( .A1(n13922), .A2(n13921), .ZN(n13958) );
  AND2_X1 U11881 ( .A1(n13722), .A2(n13721), .ZN(n16750) );
  NAND2_X1 U11882 ( .A1(n13772), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13751) );
  AOI21_X1 U11883 ( .B1(n13548), .B2(n13632), .A(n13547), .ZN(n15253) );
  OAI21_X1 U11884 ( .B1(n14902), .B2(n13701), .A(n13507), .ZN(n13508) );
  NAND2_X1 U11885 ( .A1(n13432), .A2(n13433), .ZN(n13434) );
  AND2_X1 U11886 ( .A1(n16831), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13432) );
  NAND2_X1 U11887 ( .A1(n13430), .A2(n16850), .ZN(n16819) );
  INV_X1 U11888 ( .A(n16612), .ZN(n11371) );
  INV_X1 U11889 ( .A(n17081), .ZN(n17161) );
  NAND2_X1 U11890 ( .A1(n11406), .A2(n15169), .ZN(n11405) );
  AND2_X1 U11891 ( .A1(n14376), .A2(n14864), .ZN(n22182) );
  NAND2_X1 U11892 ( .A1(n13518), .A2(n22396), .ZN(n13207) );
  NAND2_X1 U11893 ( .A1(n13253), .A2(n11485), .ZN(n11482) );
  INV_X1 U11894 ( .A(n13509), .ZN(n11485) );
  NAND2_X1 U11895 ( .A1(n11483), .A2(n13285), .ZN(n13286) );
  NAND2_X1 U11896 ( .A1(n15432), .A2(n15427), .ZN(n15429) );
  OR2_X1 U11897 ( .A1(n13528), .A2(n15426), .ZN(n22483) );
  INV_X1 U11898 ( .A(n11212), .ZN(n15428) );
  NOR2_X1 U11899 ( .A1(n22540), .A2(n15602), .ZN(n22529) );
  NAND2_X1 U11900 ( .A1(n13528), .A2(n14902), .ZN(n15058) );
  INV_X1 U11901 ( .A(n15098), .ZN(n15431) );
  NOR2_X1 U11902 ( .A1(n11223), .A2(n15428), .ZN(n15102) );
  NOR2_X1 U11903 ( .A1(n22521), .A2(n15602), .ZN(n22548) );
  OR2_X1 U11904 ( .A1(n14902), .A2(n14957), .ZN(n15081) );
  AOI21_X1 U11905 ( .B1(n22524), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n15602), 
        .ZN(n22492) );
  AND2_X1 U11906 ( .A1(n11223), .A2(n11212), .ZN(n22470) );
  INV_X1 U11907 ( .A(n15081), .ZN(n15103) );
  AND2_X1 U11908 ( .A1(n11761), .A2(n14564), .ZN(n15331) );
  AND2_X1 U11909 ( .A1(n19251), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15498) );
  AND2_X1 U11910 ( .A1(n12537), .A2(n11320), .ZN(n11319) );
  INV_X1 U11911 ( .A(n17314), .ZN(n11320) );
  NAND2_X1 U11912 ( .A1(n11997), .A2(n12006), .ZN(n12024) );
  NOR2_X1 U11913 ( .A1(n11724), .A2(n11304), .ZN(n11325) );
  NAND2_X1 U11914 ( .A1(n11467), .A2(n15638), .ZN(n11466) );
  INV_X1 U11915 ( .A(n15593), .ZN(n11467) );
  NOR2_X1 U11916 ( .A1(n11466), .A2(n12490), .ZN(n11465) );
  AND2_X1 U11917 ( .A1(n12955), .A2(n11450), .ZN(n11449) );
  INV_X1 U11918 ( .A(n17364), .ZN(n11450) );
  AND3_X1 U11919 ( .A1(n12515), .A2(n12514), .A3(n12513), .ZN(n17922) );
  INV_X1 U11920 ( .A(n12342), .ZN(n14682) );
  NAND2_X1 U11921 ( .A1(n13016), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11343) );
  AND2_X1 U11922 ( .A1(n11253), .A2(n12085), .ZN(n11334) );
  AND2_X1 U11923 ( .A1(n11381), .A2(n11380), .ZN(n11379) );
  INV_X1 U11924 ( .A(n14535), .ZN(n11380) );
  OR2_X1 U11925 ( .A1(n11436), .A2(n11435), .ZN(n11432) );
  NOR2_X1 U11926 ( .A1(n12005), .A2(n11435), .ZN(n11434) );
  NAND2_X1 U11927 ( .A1(n18054), .A2(n11329), .ZN(n17739) );
  NAND2_X1 U11928 ( .A1(n12180), .A2(n12179), .ZN(n11329) );
  AND2_X1 U11929 ( .A1(n12114), .A2(n12379), .ZN(n12425) );
  INV_X1 U11930 ( .A(n11822), .ZN(n11823) );
  INV_X1 U11931 ( .A(n11821), .ZN(n11824) );
  NAND2_X1 U11932 ( .A1(n12376), .A2(n20528), .ZN(n12333) );
  NAND2_X1 U11933 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20195), .ZN(n20164) );
  NOR2_X1 U11934 ( .A1(n20076), .A2(n20192), .ZN(n20079) );
  INV_X1 U11935 ( .A(n11856), .ZN(n11848) );
  INV_X1 U11936 ( .A(n15710), .ZN(n15720) );
  NAND2_X1 U11937 ( .A1(n15502), .A2(n15501), .ZN(n20199) );
  NAND2_X1 U11938 ( .A1(n19529), .A2(n19251), .ZN(n15502) );
  OR2_X1 U11939 ( .A1(n20262), .A2(n20409), .ZN(n15710) );
  INV_X1 U11940 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20103) );
  NAND2_X1 U11941 ( .A1(n21312), .A2(n21199), .ZN(n21322) );
  AOI22_X1 U11942 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U11943 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18712), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14051) );
  AOI211_X1 U11944 ( .C1(n11165), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n14049), .B(n14048), .ZN(n14050) );
  NOR2_X1 U11945 ( .A1(n19692), .A2(n19652), .ZN(n21607) );
  NOR2_X1 U11946 ( .A1(n19855), .A2(n14139), .ZN(n20948) );
  NAND2_X1 U11947 ( .A1(n14035), .A2(n11348), .ZN(n11352) );
  NOR2_X1 U11948 ( .A1(n18961), .A2(n11349), .ZN(n11348) );
  NAND3_X1 U11949 ( .A1(n18726), .A2(n18725), .A3(n18724), .ZN(n21673) );
  NOR2_X1 U11950 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18894), .ZN(
        n21939) );
  NAND2_X1 U11951 ( .A1(n11299), .A2(n11298), .ZN(n18914) );
  INV_X1 U11952 ( .A(n18945), .ZN(n11298) );
  NAND2_X1 U11953 ( .A1(n18754), .A2(n11246), .ZN(n11293) );
  AND2_X1 U11954 ( .A1(n18749), .A2(n21752), .ZN(n18748) );
  NAND2_X2 U11955 ( .A1(n21888), .A2(n22035), .ZN(n21911) );
  NOR2_X1 U11956 ( .A1(n21599), .A2(n21767), .ZN(n11300) );
  AND2_X1 U11957 ( .A1(n11187), .A2(n16471), .ZN(n16474) );
  NAND2_X1 U11958 ( .A1(n14353), .A2(n14352), .ZN(n14356) );
  AND2_X1 U11959 ( .A1(n14378), .A2(n14360), .ZN(n22231) );
  OR2_X1 U11960 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n22534) );
  NAND2_X1 U11961 ( .A1(n11484), .A2(n14740), .ZN(n17208) );
  INV_X1 U11962 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15681) );
  NAND2_X1 U11963 ( .A1(n19482), .A2(n19483), .ZN(n19480) );
  NAND2_X1 U11964 ( .A1(n15094), .A2(n11469), .ZN(n11468) );
  INV_X1 U11965 ( .A(n11471), .ZN(n11469) );
  NAND2_X1 U11966 ( .A1(n11503), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11471) );
  AND2_X1 U11967 ( .A1(n20008), .A2(n15508), .ZN(n20005) );
  INV_X1 U11968 ( .A(n17462), .ZN(n20003) );
  AND2_X1 U11969 ( .A1(n20513), .A2(n12352), .ZN(n20461) );
  INV_X1 U11970 ( .A(n20515), .ZN(n20459) );
  INV_X1 U11971 ( .A(n12313), .ZN(n11383) );
  INV_X1 U11972 ( .A(n18185), .ZN(n18198) );
  XNOR2_X1 U11973 ( .A(n12197), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12619) );
  OAI21_X1 U11974 ( .B1(n13014), .B2(n13015), .A(n12636), .ZN(n19457) );
  OAI21_X1 U11975 ( .B1(n17556), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14207), .ZN(n16409) );
  NAND2_X1 U11976 ( .A1(n11313), .A2(n11310), .ZN(n11309) );
  NOR2_X1 U11977 ( .A1(n11312), .A2(n11311), .ZN(n11310) );
  NAND2_X1 U11978 ( .A1(n19445), .A2(n19504), .ZN(n11313) );
  NAND2_X1 U11979 ( .A1(n11427), .A2(n14200), .ZN(n11422) );
  NAND2_X1 U11980 ( .A1(n11421), .A2(n11417), .ZN(n11419) );
  XNOR2_X1 U11981 ( .A(n11195), .B(n17853), .ZN(n17863) );
  INV_X1 U11982 ( .A(n19508), .ZN(n18055) );
  INV_X1 U11983 ( .A(n18066), .ZN(n19500) );
  INV_X1 U11984 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20122) );
  INV_X1 U11985 ( .A(n20192), .ZN(n20167) );
  NOR2_X1 U11986 ( .A1(n14743), .A2(n14747), .ZN(n19269) );
  XNOR2_X1 U11987 ( .A(n14835), .B(n14834), .ZN(n20255) );
  INV_X1 U11988 ( .A(n11724), .ZN(n11324) );
  INV_X1 U11989 ( .A(n20640), .ZN(n20533) );
  OR3_X1 U11990 ( .A1(n15357), .A2(n15356), .A3(n15355), .ZN(n19520) );
  NAND2_X1 U11991 ( .A1(n22115), .A2(n22063), .ZN(n20949) );
  OAI211_X1 U11992 ( .C1(n16121), .C2(n16111), .A(n16110), .B(n16122), .ZN(
        n22116) );
  NAND2_X1 U11993 ( .A1(n21390), .A2(n14024), .ZN(n21406) );
  NAND2_X1 U11994 ( .A1(n21294), .A2(n21199), .ZN(n21313) );
  NAND2_X1 U11995 ( .A1(n21270), .A2(n21199), .ZN(n21287) );
  CLKBUF_X2 U11996 ( .A(n21002), .Z(n20990) );
  NAND2_X1 U11997 ( .A1(n11289), .A2(n21925), .ZN(n11288) );
  NAND2_X1 U11998 ( .A1(n11290), .A2(n22027), .ZN(n11289) );
  NAND2_X1 U11999 ( .A1(n11291), .A2(n11498), .ZN(n11290) );
  NAND2_X1 U12000 ( .A1(n11287), .A2(n11285), .ZN(n11284) );
  NOR2_X1 U12001 ( .A1(n21937), .A2(n11286), .ZN(n11285) );
  OAI21_X1 U12002 ( .B1(n21933), .B2(n21925), .A(n21924), .ZN(n11287) );
  AOI21_X1 U12003 ( .B1(n11228), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n11365), .ZN(n13997) );
  AND2_X1 U12004 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11365) );
  AOI21_X1 U12005 ( .B1(n11227), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n11359), .ZN(n13932) );
  AND2_X1 U12006 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11359) );
  AOI21_X1 U12007 ( .B1(n13223), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n11363), .ZN(n13887) );
  AND2_X1 U12008 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11363) );
  AOI21_X1 U12009 ( .B1(n13993), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11366), .ZN(n13726) );
  AND2_X1 U12010 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11366) );
  AOI22_X1 U12011 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13086), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U12012 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11560) );
  INV_X1 U12013 ( .A(n13474), .ZN(n13473) );
  AOI21_X1 U12014 ( .B1(n13105), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n11355), .ZN(n13822) );
  AOI21_X1 U12015 ( .B1(n13105), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n11356), .ZN(n13707) );
  AND2_X1 U12016 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11356) );
  AOI21_X1 U12017 ( .B1(n11228), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n11364), .ZN(n13743) );
  AND2_X1 U12018 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11364) );
  AOI21_X1 U12019 ( .B1(n13985), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n11368), .ZN(n13766) );
  AND2_X1 U12020 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11368) );
  AOI21_X1 U12021 ( .B1(n13110), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11367), .ZN(n13673) );
  AND2_X1 U12022 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11367) );
  AOI21_X1 U12023 ( .B1(n13223), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n11362), .ZN(n13641) );
  AND2_X1 U12024 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11362) );
  CLKBUF_X1 U12025 ( .A(n13115), .Z(n13994) );
  AOI21_X1 U12026 ( .B1(n13963), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n11369), .ZN(n13609) );
  AND2_X1 U12027 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11369) );
  AOI21_X1 U12028 ( .B1(n13086), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n11358), .ZN(n13583) );
  AND2_X1 U12029 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11358) );
  NAND2_X1 U12030 ( .A1(n13324), .A2(n15079), .ZN(n13345) );
  NAND2_X1 U12031 ( .A1(n13154), .A2(n11182), .ZN(n13447) );
  OR2_X1 U12032 ( .A1(n13335), .A2(n13334), .ZN(n13359) );
  INV_X1 U12033 ( .A(n14364), .ZN(n14377) );
  NAND2_X1 U12034 ( .A1(n13204), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13274) );
  OR2_X1 U12035 ( .A1(n15025), .A2(n22396), .ZN(n13273) );
  AOI22_X1 U12036 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13088) );
  AND2_X1 U12037 ( .A1(n13116), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13028) );
  AOI22_X1 U12038 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13078) );
  AND2_X1 U12039 ( .A1(n11911), .A2(n12416), .ZN(n11448) );
  OAI22_X1 U12040 ( .A1(n11850), .A2(n11924), .B1(n20060), .B2(n11849), .ZN(
        n11855) );
  OAI22_X1 U12041 ( .A1(n11900), .A2(n11924), .B1(n20117), .B2(n11899), .ZN(
        n11904) );
  OAI21_X1 U12042 ( .B1(n11892), .B2(n11919), .A(n11428), .ZN(n11893) );
  XNOR2_X1 U12043 ( .A(n11729), .B(n11743), .ZN(n12358) );
  AND2_X1 U12044 ( .A1(n11746), .A2(n12376), .ZN(n12574) );
  OAI211_X1 U12045 ( .C1(n14894), .C2(n11794), .A(n11793), .B(n11792), .ZN(
        n11795) );
  NAND2_X1 U12046 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11314) );
  AOI21_X1 U12047 ( .B1(n11214), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n11713), .ZN(n11315) );
  AOI22_X1 U12048 ( .A1(n11205), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U12049 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20122), .ZN(
        n12125) );
  NOR2_X1 U12050 ( .A1(n21640), .A2(n21005), .ZN(n14126) );
  NAND2_X1 U12051 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21033), .ZN(
        n14043) );
  NOR2_X1 U12052 ( .A1(n16227), .A2(n21477), .ZN(n16233) );
  INV_X1 U12053 ( .A(n16113), .ZN(n16105) );
  AND2_X1 U12054 ( .A1(n13467), .A2(n13466), .ZN(n14232) );
  NAND2_X1 U12055 ( .A1(n11370), .A2(n14248), .ZN(n14254) );
  INV_X1 U12056 ( .A(n14347), .ZN(n11370) );
  NAND2_X1 U12057 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13114) );
  INV_X1 U12058 ( .A(n16568), .ZN(n11473) );
  AND2_X1 U12059 ( .A1(n16579), .A2(n13815), .ZN(n11474) );
  AND2_X1 U12060 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13529), .ZN(
        n13539) );
  AND2_X1 U12061 ( .A1(n13503), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13536) );
  NAND2_X1 U12062 ( .A1(n11374), .A2(n16505), .ZN(n11373) );
  INV_X1 U12063 ( .A(n16520), .ZN(n11374) );
  NOR2_X1 U12064 ( .A1(n16599), .A2(n17069), .ZN(n11376) );
  NOR2_X1 U12065 ( .A1(n11237), .A2(n11402), .ZN(n11401) );
  INV_X1 U12066 ( .A(n13381), .ZN(n13379) );
  INV_X1 U12067 ( .A(n13382), .ZN(n13380) );
  NOR2_X1 U12068 ( .A1(n14411), .A2(n13092), .ZN(n13151) );
  OR2_X1 U12069 ( .A1(n13189), .A2(n13188), .ZN(n13406) );
  NOR2_X1 U12070 ( .A1(n13173), .A2(n13172), .ZN(n13174) );
  OR2_X1 U12071 ( .A1(n13284), .A2(n13283), .ZN(n13290) );
  AND2_X1 U12072 ( .A1(n18166), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13458) );
  OAI21_X1 U12073 ( .B1(n13264), .B2(n13217), .A(n13219), .ZN(n13221) );
  AND2_X1 U12074 ( .A1(n15005), .A2(n13298), .ZN(n15604) );
  AOI21_X1 U12075 ( .B1(n18159), .B2(n22395), .A(n22400), .ZN(n14965) );
  AND2_X2 U12076 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14897) );
  NAND2_X1 U12077 ( .A1(n12094), .A2(n12095), .ZN(n12091) );
  NAND2_X1 U12078 ( .A1(n12088), .A2(n12089), .ZN(n12109) );
  INV_X1 U12079 ( .A(n12091), .ZN(n12088) );
  INV_X1 U12080 ( .A(n17535), .ZN(n12537) );
  NAND2_X1 U12081 ( .A1(n12909), .A2(n12910), .ZN(n17368) );
  OR2_X1 U12082 ( .A1(n12861), .A2(n11461), .ZN(n11460) );
  INV_X1 U12083 ( .A(n12905), .ZN(n12881) );
  NAND2_X1 U12084 ( .A1(n12097), .A2(n17557), .ZN(n11335) );
  NAND2_X1 U12085 ( .A1(n14508), .A2(n11266), .ZN(n11337) );
  NAND2_X1 U12086 ( .A1(n17283), .A2(n17284), .ZN(n17482) );
  NAND2_X1 U12087 ( .A1(n12538), .A2(n12537), .ZN(n17537) );
  AND2_X1 U12088 ( .A1(n16364), .A2(n12236), .ZN(n11381) );
  INV_X1 U12089 ( .A(n16256), .ZN(n12236) );
  AND2_X1 U12090 ( .A1(n17339), .A2(n12054), .ZN(n12643) );
  INV_X1 U12091 ( .A(n17694), .ZN(n11435) );
  XNOR2_X1 U12092 ( .A(n12186), .B(n11961), .ZN(n12183) );
  NAND2_X1 U12093 ( .A1(n12141), .A2(n12146), .ZN(n12159) );
  NAND2_X1 U12094 ( .A1(n12676), .A2(n12678), .ZN(n12694) );
  AOI21_X1 U12095 ( .B1(n22069), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14150), .ZN(n14156) );
  NOR2_X1 U12096 ( .A1(n14157), .A2(n16107), .ZN(n14150) );
  NOR2_X1 U12097 ( .A1(n21005), .A2(n14043), .ZN(n14064) );
  INV_X1 U12098 ( .A(n22089), .ZN(n20947) );
  NAND2_X1 U12099 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11347) );
  INV_X1 U12100 ( .A(n19060), .ZN(n21074) );
  NOR2_X1 U12101 ( .A1(n16112), .A2(n21619), .ZN(n18321) );
  AND2_X1 U12102 ( .A1(n18727), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18728) );
  INV_X1 U12103 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21033) );
  NOR2_X2 U12104 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21639) );
  AND2_X1 U12105 ( .A1(n13589), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13605) );
  AND2_X1 U12106 ( .A1(n16569), .A2(n16562), .ZN(n16560) );
  AND2_X1 U12107 ( .A1(n14255), .A2(n11372), .ZN(n14950) );
  NAND2_X1 U12108 ( .A1(n14816), .A2(n15033), .ZN(n11372) );
  XNOR2_X1 U12109 ( .A(n14255), .B(n14816), .ZN(n15463) );
  AND2_X1 U12110 ( .A1(n14999), .A2(n13150), .ZN(n14426) );
  AND2_X1 U12111 ( .A1(n14945), .A2(n14944), .ZN(n20697) );
  OR2_X1 U12112 ( .A1(n13961), .A2(n13960), .ZN(n14014) );
  AOI21_X1 U12113 ( .B1(n15010), .B2(n16514), .A(n13957), .ZN(n14211) );
  OAI21_X1 U12114 ( .B1(n13982), .B2(n16815), .A(n13939), .ZN(n16519) );
  NAND2_X1 U12115 ( .A1(n13897), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13920) );
  NAND2_X1 U12116 ( .A1(n13834), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13836) );
  OR2_X1 U12117 ( .A1(n13836), .A2(n13835), .ZN(n13896) );
  OR2_X1 U12118 ( .A1(n22385), .A2(n13982), .ZN(n13813) );
  AND2_X1 U12119 ( .A1(n16750), .A2(n16608), .ZN(n13776) );
  NOR2_X1 U12120 ( .A1(n13751), .A2(n13752), .ZN(n13738) );
  INV_X1 U12121 ( .A(n13717), .ZN(n13718) );
  NAND2_X1 U12122 ( .A1(n13697), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13717) );
  AND2_X1 U12123 ( .A1(n13670), .A2(n13669), .ZN(n13697) );
  AND2_X1 U12124 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13669) );
  INV_X1 U12125 ( .A(n11476), .ZN(n11475) );
  OAI21_X1 U12126 ( .B1(n11477), .B2(n11478), .A(n11267), .ZN(n11476) );
  NAND2_X1 U12127 ( .A1(n13605), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13633) );
  INV_X1 U12128 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13566) );
  NOR2_X1 U12129 ( .A1(n13567), .A2(n13566), .ZN(n13589) );
  AND2_X1 U12130 ( .A1(n13551), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13560) );
  AOI21_X1 U12131 ( .B1(n13558), .B2(n13632), .A(n13557), .ZN(n15653) );
  INV_X1 U12132 ( .A(n15253), .ZN(n13549) );
  NAND2_X1 U12133 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13530) );
  AND3_X1 U12134 ( .A1(n14362), .A2(n13451), .A3(n14242), .ZN(n18145) );
  OR2_X1 U12135 ( .A1(n16497), .A2(n14625), .ZN(n14353) );
  NOR2_X1 U12136 ( .A1(n16531), .A2(n16520), .ZN(n16522) );
  NOR2_X1 U12137 ( .A1(n16580), .A2(n16570), .ZN(n16569) );
  NAND2_X1 U12138 ( .A1(n11376), .A2(n11375), .ZN(n16580) );
  INV_X1 U12139 ( .A(n16582), .ZN(n11375) );
  NAND2_X1 U12140 ( .A1(n13426), .A2(n16955), .ZN(n16860) );
  NAND2_X1 U12141 ( .A1(n13429), .A2(n11414), .ZN(n11413) );
  AND2_X1 U12142 ( .A1(n11489), .A2(n11415), .ZN(n11414) );
  INV_X1 U12143 ( .A(n11376), .ZN(n17071) );
  NOR2_X2 U12144 ( .A1(n17098), .A2(n17097), .ZN(n17100) );
  AND2_X1 U12145 ( .A1(n14314), .A2(n14313), .ZN(n16612) );
  INV_X1 U12146 ( .A(n17149), .ZN(n14303) );
  NAND2_X1 U12147 ( .A1(n16699), .A2(n16663), .ZN(n16665) );
  AOI21_X1 U12148 ( .B1(n16379), .B2(n11402), .A(n11237), .ZN(n11399) );
  INV_X1 U12149 ( .A(n16379), .ZN(n11400) );
  INV_X1 U12150 ( .A(n16304), .ZN(n14282) );
  NAND2_X1 U12151 ( .A1(n16341), .A2(n13411), .ZN(n16380) );
  NAND2_X1 U12152 ( .A1(n20819), .A2(n16265), .ZN(n16305) );
  INV_X1 U12153 ( .A(n15256), .ZN(n14270) );
  NOR2_X1 U12154 ( .A1(n15373), .A2(n15374), .ZN(n15258) );
  AND2_X1 U12155 ( .A1(n17161), .A2(n17157), .ZN(n22221) );
  AND2_X1 U12156 ( .A1(n14378), .A2(n14371), .ZN(n17081) );
  AND2_X1 U12157 ( .A1(n17157), .A2(n14389), .ZN(n14865) );
  OAI21_X1 U12158 ( .B1(n13516), .B2(n13403), .A(n13214), .ZN(n14812) );
  NAND2_X1 U12159 ( .A1(n11396), .A2(n11395), .ZN(n11397) );
  NOR2_X1 U12160 ( .A1(n18128), .A2(n22396), .ZN(n11395) );
  NAND2_X1 U12161 ( .A1(n14961), .A2(n13222), .ZN(n15434) );
  NOR2_X1 U12162 ( .A1(n15377), .A2(n11223), .ZN(n15386) );
  OR2_X1 U12163 ( .A1(n11223), .A2(n11212), .ZN(n15098) );
  INV_X1 U12164 ( .A(n13153), .ZN(n14966) );
  CLKBUF_X1 U12165 ( .A(n13203), .Z(n13204) );
  INV_X1 U12166 ( .A(n14410), .ZN(n14999) );
  NOR2_X1 U12167 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14965), .ZN(n15139) );
  OR2_X1 U12168 ( .A1(n14954), .A2(n16972), .ZN(n15138) );
  OR3_X1 U12169 ( .A1(n15600), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14965), 
        .ZN(n15141) );
  INV_X1 U12170 ( .A(n14357), .ZN(n18156) );
  AND2_X1 U12171 ( .A1(n12140), .A2(n12139), .ZN(n15339) );
  AND2_X1 U12172 ( .A1(n12571), .A2(n12570), .ZN(n15341) );
  NAND2_X1 U12173 ( .A1(n14518), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14520) );
  NOR2_X1 U12174 ( .A1(n12086), .A2(n11339), .ZN(n12094) );
  INV_X1 U12175 ( .A(n12087), .ZN(n11339) );
  NAND2_X1 U12176 ( .A1(n12081), .A2(n12082), .ZN(n12086) );
  NAND2_X1 U12177 ( .A1(n17293), .A2(n11186), .ZN(n17286) );
  NAND2_X1 U12178 ( .A1(n17286), .A2(n17593), .ZN(n17285) );
  NAND2_X1 U12179 ( .A1(n12033), .A2(n12034), .ZN(n12038) );
  NAND2_X1 U12180 ( .A1(n11655), .A2(n11959), .ZN(n11999) );
  NAND2_X1 U12181 ( .A1(n11340), .A2(n11955), .ZN(n11953) );
  INV_X1 U12182 ( .A(n12115), .ZN(n11340) );
  NAND2_X1 U12183 ( .A1(n11967), .A2(n11968), .ZN(n11981) );
  NAND2_X1 U12184 ( .A1(n11465), .A2(n11464), .ZN(n11463) );
  INV_X1 U12185 ( .A(n12909), .ZN(n12912) );
  XNOR2_X1 U12186 ( .A(n12885), .B(n12886), .ZN(n17383) );
  NAND2_X1 U12187 ( .A1(n17383), .A2(n17382), .ZN(n17381) );
  AND2_X1 U12188 ( .A1(n17446), .A2(n17422), .ZN(n17428) );
  OR2_X1 U12189 ( .A1(n17427), .A2(n17443), .ZN(n17444) );
  AND2_X1 U12190 ( .A1(n16367), .A2(n16374), .ZN(n17416) );
  AND3_X1 U12191 ( .A1(n12477), .A2(n12476), .A3(n12475), .ZN(n17343) );
  AND3_X1 U12192 ( .A1(n12451), .A2(n12450), .A3(n12449), .ZN(n15266) );
  NOR2_X2 U12193 ( .A1(n15265), .A2(n15266), .ZN(n17989) );
  CLKBUF_X1 U12194 ( .A(n15265), .Z(n18032) );
  AND2_X1 U12195 ( .A1(n14681), .A2(n19252), .ZN(n18238) );
  INV_X1 U12196 ( .A(n14661), .ZN(n15508) );
  INV_X1 U12197 ( .A(n12312), .ZN(n12299) );
  OR2_X1 U12198 ( .A1(n11337), .A2(n11336), .ZN(n14514) );
  NAND2_X1 U12199 ( .A1(n14508), .A2(n11232), .ZN(n14479) );
  AND2_X1 U12200 ( .A1(n14508), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14480) );
  NAND2_X1 U12201 ( .A1(n17668), .A2(n12644), .ZN(n12647) );
  NAND2_X1 U12202 ( .A1(n14506), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14505) );
  AND2_X1 U12203 ( .A1(n14503), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14506) );
  NAND2_X1 U12204 ( .A1(n14500), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14504) );
  NOR2_X1 U12205 ( .A1(n14504), .A2(n11338), .ZN(n14503) );
  INV_X1 U12206 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14498) );
  NOR2_X1 U12207 ( .A1(n14499), .A2(n14498), .ZN(n14500) );
  INV_X1 U12208 ( .A(n15590), .ZN(n11377) );
  NAND2_X1 U12209 ( .A1(n14492), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14497) );
  AND2_X1 U12210 ( .A1(n14494), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14492) );
  NOR2_X1 U12211 ( .A1(n14490), .A2(n17741), .ZN(n14494) );
  NOR2_X1 U12212 ( .A1(n14488), .A2(n16332), .ZN(n14491) );
  NAND2_X1 U12213 ( .A1(n14489), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14488) );
  NAND2_X1 U12214 ( .A1(n11323), .A2(n11322), .ZN(n11385) );
  AND2_X1 U12215 ( .A1(n12201), .A2(n11386), .ZN(n11323) );
  NOR2_X1 U12216 ( .A1(n16408), .A2(n16407), .ZN(n11311) );
  OR2_X1 U12217 ( .A1(n16405), .A2(n16406), .ZN(n11312) );
  NAND2_X1 U12218 ( .A1(n11250), .A2(n11427), .ZN(n11417) );
  NOR2_X1 U12219 ( .A1(n11426), .A2(n12097), .ZN(n11420) );
  INV_X1 U12220 ( .A(n17385), .ZN(n11387) );
  AND2_X1 U12221 ( .A1(n19421), .A2(n12102), .ZN(n17580) );
  NAND2_X1 U12222 ( .A1(n17599), .A2(n12073), .ZN(n17591) );
  INV_X1 U12223 ( .A(n11443), .ZN(n11442) );
  OAI21_X1 U12224 ( .B1(n11230), .B2(n11445), .A(n12193), .ZN(n11443) );
  AND2_X1 U12225 ( .A1(n17964), .A2(n12607), .ZN(n17819) );
  NAND2_X1 U12226 ( .A1(n11389), .A2(n11388), .ZN(n17408) );
  INV_X1 U12227 ( .A(n17413), .ZN(n11388) );
  AND2_X1 U12228 ( .A1(n17514), .A2(n17513), .ZN(n19396) );
  AOI21_X1 U12229 ( .B1(n17638), .B2(n12652), .A(n12651), .ZN(n17617) );
  INV_X1 U12230 ( .A(n11389), .ZN(n17414) );
  XNOR2_X1 U12231 ( .A(n17617), .B(n17616), .ZN(n17619) );
  NAND2_X1 U12232 ( .A1(n11321), .A2(n11260), .ZN(n17546) );
  AND2_X1 U12233 ( .A1(n17722), .A2(n18020), .ZN(n17723) );
  XNOR2_X1 U12234 ( .A(n12187), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18015) );
  INV_X1 U12235 ( .A(n11988), .ZN(n11303) );
  AND2_X1 U12236 ( .A1(n12379), .A2(n12423), .ZN(n12424) );
  NAND2_X1 U12237 ( .A1(n16319), .A2(n12169), .ZN(n11447) );
  OAI21_X1 U12238 ( .B1(n12167), .B2(n12175), .A(n12174), .ZN(n12176) );
  AND2_X1 U12239 ( .A1(n12409), .A2(n11317), .ZN(n11316) );
  INV_X1 U12240 ( .A(n15558), .ZN(n11317) );
  NAND2_X1 U12241 ( .A1(n15554), .A2(n15553), .ZN(n16269) );
  INV_X1 U12242 ( .A(n11761), .ZN(n11762) );
  NAND2_X1 U12243 ( .A1(n15486), .A2(n12409), .ZN(n11318) );
  NAND2_X1 U12244 ( .A1(n19505), .A2(n15498), .ZN(n12686) );
  XNOR2_X1 U12245 ( .A(n14743), .B(n12690), .ZN(n14835) );
  AOI21_X1 U12246 ( .B1(n17360), .B2(n15498), .A(n12689), .ZN(n14834) );
  INV_X1 U12247 ( .A(n11384), .ZN(n11818) );
  NAND2_X1 U12248 ( .A1(n12346), .A2(n12344), .ZN(n15472) );
  AND2_X1 U12249 ( .A1(n11743), .A2(n12345), .ZN(n11723) );
  NAND2_X1 U12250 ( .A1(n20262), .A2(n20409), .ZN(n20184) );
  NAND2_X1 U12251 ( .A1(n20262), .A2(n18220), .ZN(n20133) );
  OR2_X1 U12252 ( .A1(n20255), .A2(n20519), .ZN(n20163) );
  NAND3_X1 U12253 ( .A1(n11522), .A2(n11521), .A3(n11496), .ZN(n11523) );
  NAND2_X1 U12254 ( .A1(n20255), .A2(n20519), .ZN(n20144) );
  NOR2_X2 U12255 ( .A1(n15508), .A2(n20164), .ZN(n20531) );
  INV_X1 U12256 ( .A(n15716), .ZN(n15713) );
  AOI21_X1 U12257 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n22080), .A(
        n14160), .ZN(n16110) );
  NAND2_X1 U12258 ( .A1(n21243), .A2(n21199), .ZN(n21258) );
  NAND2_X1 U12259 ( .A1(n14024), .A2(n11505), .ZN(n21234) );
  NAND2_X1 U12260 ( .A1(n21234), .A2(n21235), .ZN(n21233) );
  INV_X1 U12261 ( .A(n19007), .ZN(n14023) );
  OAI211_X1 U12262 ( .C1(n11234), .C2(n14074), .A(n14073), .B(n11493), .ZN(
        n14075) );
  NOR2_X1 U12263 ( .A1(n21616), .A2(n20948), .ZN(n21427) );
  NOR2_X1 U12264 ( .A1(n20949), .A2(n18097), .ZN(n19197) );
  NOR2_X1 U12265 ( .A1(n20947), .A2(n20949), .ZN(n20951) );
  NAND2_X1 U12266 ( .A1(n14035), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18937) );
  AND2_X1 U12267 ( .A1(n11297), .A2(n11299), .ZN(n18895) );
  NOR2_X1 U12268 ( .A1(n18895), .A2(n21938), .ZN(n21923) );
  NAND2_X1 U12269 ( .A1(n14034), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14036) );
  INV_X1 U12270 ( .A(n18794), .ZN(n21147) );
  AND2_X1 U12271 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19099) );
  NAND2_X1 U12272 ( .A1(n21933), .A2(n11292), .ZN(n11291) );
  AND2_X1 U12273 ( .A1(n21934), .A2(n21932), .ZN(n11292) );
  NOR2_X1 U12274 ( .A1(n18874), .A2(n18875), .ZN(n18882) );
  AND2_X1 U12275 ( .A1(n11293), .A2(n19044), .ZN(n18875) );
  NOR2_X1 U12276 ( .A1(n18875), .A2(n18758), .ZN(n18816) );
  AND2_X1 U12277 ( .A1(n21884), .A2(n16106), .ZN(n22035) );
  NOR2_X1 U12278 ( .A1(n18742), .A2(n19048), .ZN(n21990) );
  NOR2_X1 U12279 ( .A1(n19049), .A2(n21752), .ZN(n19048) );
  XNOR2_X1 U12280 ( .A(n16236), .B(n16235), .ZN(n19084) );
  NAND2_X1 U12281 ( .A1(n19110), .A2(n16230), .ZN(n19101) );
  XNOR2_X1 U12282 ( .A(n11294), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19102) );
  INV_X1 U12283 ( .A(n16231), .ZN(n11294) );
  NAND2_X1 U12284 ( .A1(n19101), .A2(n19102), .ZN(n19100) );
  INV_X2 U12285 ( .A(n19196), .ZN(n19905) );
  NOR2_X2 U12286 ( .A1(n14113), .A2(n14112), .ZN(n19813) );
  NOR2_X1 U12287 ( .A1(n14123), .A2(n14122), .ZN(n19773) );
  BUF_X1 U12288 ( .A(n14138), .Z(n19733) );
  INV_X1 U12289 ( .A(n19854), .ZN(n19902) );
  CLKBUF_X1 U12290 ( .A(n14661), .Z(n15507) );
  OR2_X1 U12291 ( .A1(n14620), .A2(n22406), .ZN(n14624) );
  OR2_X1 U12292 ( .A1(n16559), .A2(n20761), .ZN(n16549) );
  OR2_X1 U12293 ( .A1(n22333), .A2(n22279), .ZN(n22339) );
  NOR2_X2 U12294 ( .A1(n15035), .A2(n15034), .ZN(n22359) );
  INV_X1 U12295 ( .A(n22370), .ZN(n22355) );
  INV_X1 U12296 ( .A(n16666), .ZN(n22353) );
  AND2_X1 U12297 ( .A1(n15023), .A2(n15022), .ZN(n22357) );
  AND2_X1 U12298 ( .A1(n20830), .A2(n15140), .ZN(n20826) );
  NAND2_X1 U12299 ( .A1(n14843), .A2(n14842), .ZN(n20830) );
  INV_X1 U12300 ( .A(n20826), .ZN(n20820) );
  INV_X1 U12301 ( .A(n16791), .ZN(n16770) );
  INV_X1 U12302 ( .A(n16763), .ZN(n16771) );
  OR2_X1 U12303 ( .A1(n16770), .A2(n14882), .ZN(n16794) );
  NOR2_X1 U12304 ( .A1(n16463), .A2(n14749), .ZN(n14752) );
  XNOR2_X1 U12305 ( .A(n14015), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15022) );
  NOR2_X1 U12306 ( .A1(n14014), .A2(n16801), .ZN(n14015) );
  XNOR2_X1 U12307 ( .A(n16495), .B(n14403), .ZN(n16803) );
  INV_X1 U12308 ( .A(n20856), .ZN(n20859) );
  AND2_X2 U12309 ( .A1(n22386), .A2(n14016), .ZN(n20857) );
  INV_X1 U12310 ( .A(n16805), .ZN(n11275) );
  NAND2_X1 U12311 ( .A1(n16798), .A2(n16797), .ZN(n11276) );
  XNOR2_X1 U12312 ( .A(n14217), .B(n16991), .ZN(n17000) );
  NAND2_X1 U12313 ( .A1(n14215), .A2(n16956), .ZN(n14216) );
  INV_X1 U12314 ( .A(n13434), .ZN(n11412) );
  OAI211_X1 U12315 ( .C1(n11174), .C2(n11404), .A(n11403), .B(n13344), .ZN(
        n20839) );
  NAND2_X1 U12316 ( .A1(n11174), .A2(n13322), .ZN(n20833) );
  NOR2_X1 U12317 ( .A1(n22221), .A2(n14865), .ZN(n22160) );
  INV_X1 U12318 ( .A(n22226), .ZN(n22239) );
  INV_X1 U12319 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18135) );
  NAND2_X1 U12320 ( .A1(n13258), .A2(n11482), .ZN(n13287) );
  INV_X1 U12321 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18166) );
  INV_X1 U12322 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18128) );
  NOR2_X1 U12323 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20865) );
  NOR2_X1 U12324 ( .A1(n15429), .A2(n15428), .ZN(n22715) );
  OAI21_X1 U12325 ( .B1(n15430), .B2(n15435), .A(n22492), .ZN(n22677) );
  INV_X1 U12326 ( .A(n22715), .ZN(n15462) );
  OAI211_X1 U12327 ( .C1(n22479), .C2(n22478), .A(n22529), .B(n22477), .ZN(
        n22723) );
  INV_X1 U12328 ( .A(n22498), .ZN(n22730) );
  OAI211_X1 U12329 ( .C1(n15600), .C2(n22690), .A(n15520), .B(n22529), .ZN(
        n22694) );
  NOR2_X2 U12330 ( .A1(n15058), .A2(n15098), .ZN(n22750) );
  INV_X1 U12331 ( .A(n15126), .ZN(n15167) );
  NAND2_X1 U12332 ( .A1(n15103), .A2(n15102), .ZN(n22772) );
  OAI211_X1 U12333 ( .C1(n15683), .C2(n15688), .A(n22525), .B(n22548), .ZN(
        n22710) );
  INV_X1 U12334 ( .A(n17236), .ZN(n22605) );
  INV_X1 U12335 ( .A(n17244), .ZN(n22627) );
  INV_X1 U12336 ( .A(n22697), .ZN(n22705) );
  NOR2_X2 U12337 ( .A1(n15081), .A2(n15597), .ZN(n22778) );
  INV_X1 U12338 ( .A(n17230), .ZN(n22400) );
  AND2_X1 U12339 ( .A1(n18164), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22390) );
  INV_X1 U12340 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22489) );
  OR2_X1 U12341 ( .A1(n14565), .A2(n14566), .ZN(n14578) );
  NAND2_X1 U12342 ( .A1(n19450), .A2(n11186), .ZN(n19464) );
  NAND2_X1 U12343 ( .A1(n19464), .A2(n19465), .ZN(n19463) );
  NAND2_X1 U12344 ( .A1(n17265), .A2(n11185), .ZN(n19451) );
  NAND2_X1 U12345 ( .A1(n19451), .A2(n19452), .ZN(n19450) );
  NAND2_X1 U12346 ( .A1(n17266), .A2(n17558), .ZN(n17265) );
  NAND2_X1 U12347 ( .A1(n19435), .A2(n19436), .ZN(n19434) );
  NAND2_X1 U12348 ( .A1(n17285), .A2(n11185), .ZN(n19426) );
  NAND2_X1 U12349 ( .A1(n19426), .A2(n19427), .ZN(n19425) );
  NAND2_X1 U12350 ( .A1(n17294), .A2(n17603), .ZN(n17293) );
  NAND2_X1 U12351 ( .A1(n19371), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19443) );
  INV_X1 U12352 ( .A(n19441), .ZN(n19473) );
  AND2_X1 U12353 ( .A1(n18168), .A2(n14458), .ZN(n19470) );
  INV_X1 U12354 ( .A(n19443), .ZN(n19472) );
  INV_X1 U12355 ( .A(n15192), .ZN(n11462) );
  INV_X1 U12356 ( .A(n14905), .ZN(n11470) );
  INV_X1 U12357 ( .A(n17419), .ZN(n17452) );
  NAND2_X1 U12358 ( .A1(n11451), .A2(n12955), .ZN(n17365) );
  NAND2_X1 U12359 ( .A1(n17391), .A2(n17390), .ZN(n17389) );
  XNOR2_X1 U12360 ( .A(n17395), .B(n12861), .ZN(n17391) );
  AND2_X1 U12361 ( .A1(n20517), .A2(n20515), .ZN(n20209) );
  XNOR2_X1 U12362 ( .A(n14893), .B(n14892), .ZN(n20409) );
  CLKBUF_X1 U12364 ( .A(n18257), .Z(n18266) );
  NOR2_X1 U12365 ( .A1(n18238), .A2(n18266), .ZN(n18251) );
  INV_X1 U12366 ( .A(n14602), .ZN(n14636) );
  INV_X1 U12367 ( .A(n14636), .ZN(n14704) );
  INV_X1 U12368 ( .A(n18204), .ZN(n18174) );
  NOR2_X1 U12369 ( .A1(n12657), .A2(n17624), .ZN(n17850) );
  AND2_X1 U12370 ( .A1(n17448), .A2(n16399), .ZN(n19346) );
  INV_X1 U12371 ( .A(n12642), .ZN(n17697) );
  NAND2_X1 U12372 ( .A1(n11431), .A2(n11436), .ZN(n17693) );
  INV_X1 U12373 ( .A(n15564), .ZN(n12154) );
  INV_X1 U12374 ( .A(n12201), .ZN(n11455) );
  INV_X1 U12375 ( .A(n12677), .ZN(n16440) );
  INV_X1 U12376 ( .A(n17838), .ZN(n19502) );
  INV_X1 U12377 ( .A(n18061), .ZN(n19504) );
  INV_X1 U12378 ( .A(n19269), .ZN(n20519) );
  INV_X1 U12379 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20150) );
  INV_X1 U12380 ( .A(n20409), .ZN(n18220) );
  AND2_X1 U12381 ( .A1(n15472), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19529) );
  OAI21_X1 U12382 ( .B1(n20631), .B2(n20200), .A(n20199), .ZN(n20637) );
  AOI211_X2 U12383 ( .C1(n20195), .C2(n20171), .A(n20170), .B(n20169), .ZN(
        n20619) );
  OAI21_X1 U12384 ( .B1(n20174), .B2(n20162), .A(n20161), .ZN(n20617) );
  INV_X1 U12385 ( .A(n20615), .ZN(n20603) );
  OAI21_X1 U12386 ( .B1(n16293), .B2(n16292), .A(n16291), .ZN(n20604) );
  OR2_X1 U12387 ( .A1(n20133), .A2(n20183), .ZN(n20495) );
  NOR2_X1 U12388 ( .A1(n20133), .A2(n20163), .ZN(n20590) );
  OR2_X1 U12389 ( .A1(n20133), .A2(n20100), .ZN(n20581) );
  OAI21_X1 U12390 ( .B1(n20575), .B2(n20105), .A(n20199), .ZN(n20578) );
  NAND2_X1 U12391 ( .A1(n20109), .A2(n20108), .ZN(n20577) );
  OAI22_X1 U12392 ( .A1(n20085), .A2(n20084), .B1(n20195), .B2(n20083), .ZN(
        n20564) );
  INV_X1 U12393 ( .A(n20300), .ZN(n20305) );
  NAND2_X1 U12394 ( .A1(n20062), .A2(n20061), .ZN(n20553) );
  INV_X1 U12395 ( .A(n20450), .ZN(n20452) );
  NOR2_X2 U12396 ( .A1(n20183), .A2(n15710), .ZN(n20552) );
  INV_X1 U12397 ( .A(n20641), .ZN(n20618) );
  INV_X1 U12398 ( .A(n20185), .ZN(n20207) );
  AOI21_X1 U12399 ( .B1(n20537), .B2(n20199), .A(n20043), .ZN(n20540) );
  NAND2_X1 U12400 ( .A1(n20047), .A2(n20046), .ZN(n20539) );
  INV_X1 U12401 ( .A(n20188), .ZN(n20191) );
  INV_X1 U12402 ( .A(n20623), .ZN(n20634) );
  INV_X1 U12403 ( .A(n20512), .ZN(n20503) );
  INV_X1 U12404 ( .A(n20506), .ZN(n20508) );
  INV_X1 U12405 ( .A(n20456), .ZN(n20447) );
  INV_X1 U12406 ( .A(n20357), .ZN(n20348) );
  INV_X1 U12407 ( .A(n20309), .ZN(n20297) );
  NAND2_X1 U12408 ( .A1(n15720), .A2(n15718), .ZN(n20640) );
  INV_X1 U12409 ( .A(n20543), .ZN(n20471) );
  INV_X1 U12410 ( .A(n20252), .ZN(n20242) );
  INV_X1 U12411 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19251) );
  AND2_X1 U12412 ( .A1(n15362), .A2(n15361), .ZN(n19527) );
  CLKBUF_X1 U12413 ( .A(n18313), .Z(n18308) );
  INV_X1 U12414 ( .A(n22059), .ZN(n18697) );
  INV_X1 U12415 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n22091) );
  AND2_X1 U12416 ( .A1(n21339), .A2(n14170), .ZN(n21364) );
  NAND2_X1 U12417 ( .A1(n22090), .A2(n14168), .ZN(n21349) );
  NAND2_X1 U12418 ( .A1(n21271), .A2(n21272), .ZN(n21270) );
  NAND2_X1 U12419 ( .A1(n21257), .A2(n21199), .ZN(n21271) );
  NAND2_X1 U12420 ( .A1(n21244), .A2(n21245), .ZN(n21243) );
  NAND2_X1 U12421 ( .A1(n21233), .A2(n14024), .ZN(n21244) );
  NOR2_X1 U12422 ( .A1(n21242), .A2(n21241), .ZN(n21279) );
  INV_X1 U12423 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n21165) );
  NOR3_X1 U12424 ( .A1(n21349), .A2(n21126), .A3(n21125), .ZN(n21157) );
  INV_X1 U12425 ( .A(n22096), .ZN(n21391) );
  INV_X1 U12426 ( .A(n21349), .ZN(n21339) );
  INV_X1 U12427 ( .A(n21416), .ZN(n21306) );
  INV_X1 U12428 ( .A(n21385), .ZN(n21419) );
  NAND2_X1 U12429 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18605), .ZN(n18589) );
  NOR2_X1 U12430 ( .A1(n21297), .A2(n18630), .ZN(n18612) );
  NOR2_X1 U12431 ( .A1(n21273), .A2(n18641), .ZN(n18586) );
  NAND2_X1 U12432 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18686), .ZN(n18667) );
  NAND2_X1 U12433 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18464), .ZN(n18670) );
  NOR2_X2 U12434 ( .A1(n21237), .A2(n18670), .ZN(n18686) );
  BUF_X1 U12435 ( .A(n14137), .Z(n18687) );
  AND4_X1 U12436 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_7__SCAN_IN), .A4(n18364), .ZN(n18463) );
  AND2_X1 U12437 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18353), .ZN(n18364) );
  AND2_X1 U12438 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18351), .ZN(n18353) );
  AND4_X1 U12439 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18691), .A4(n18322), .ZN(n18351) );
  INV_X1 U12440 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18690) );
  NOR2_X1 U12441 ( .A1(n18692), .A2(n18687), .ZN(n18693) );
  NOR2_X1 U12442 ( .A1(n21553), .A2(n21548), .ZN(n21547) );
  NAND2_X1 U12443 ( .A1(n21554), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21553) );
  INV_X1 U12444 ( .A(n21559), .ZN(n21522) );
  NOR2_X1 U12445 ( .A1(n21521), .A2(n21564), .ZN(n21558) );
  INV_X1 U12446 ( .A(n21492), .ZN(n21488) );
  INV_X1 U12447 ( .A(n21513), .ZN(n21509) );
  NAND2_X1 U12448 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n21509), .ZN(n21508) );
  NAND4_X1 U12449 ( .A1(n21472), .A2(n21457), .A3(P3_EAX_REG_6__SCAN_IN), .A4(
        P3_EAX_REG_7__SCAN_IN), .ZN(n21587) );
  NOR2_X1 U12450 ( .A1(n16154), .A2(n16153), .ZN(n21467) );
  NOR2_X1 U12451 ( .A1(n21592), .A2(n21456), .ZN(n21472) );
  INV_X1 U12452 ( .A(n16228), .ZN(n21477) );
  NOR2_X1 U12453 ( .A1(n16196), .A2(n16195), .ZN(n21482) );
  INV_X1 U12454 ( .A(n21601), .ZN(n21593) );
  INV_X1 U12455 ( .A(n21592), .ZN(n21604) );
  INV_X1 U12456 ( .A(n21595), .ZN(n21606) );
  NOR2_X1 U12457 ( .A1(n22057), .A2(n19197), .ZN(n19208) );
  CLKBUF_X1 U12458 ( .A(n19206), .Z(n22057) );
  CLKBUF_X1 U12459 ( .A(n19208), .Z(n19214) );
  NOR3_X1 U12461 ( .A1(n22453), .A2(n20950), .A3(n20949), .ZN(n21002) );
  NOR2_X1 U12462 ( .A1(n21850), .A2(n18932), .ZN(n18919) );
  OR2_X1 U12463 ( .A1(n21857), .A2(n18891), .ZN(n18932) );
  NOR2_X1 U12464 ( .A1(n18760), .A2(n21255), .ZN(n18839) );
  INV_X1 U12465 ( .A(n18965), .ZN(n19047) );
  AND2_X1 U12466 ( .A1(n18733), .A2(n18704), .ZN(n19082) );
  INV_X1 U12467 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19085) );
  INV_X1 U12468 ( .A(n19082), .ZN(n19135) );
  AOI21_X2 U12469 ( .B1(n20944), .B2(n22113), .A(n22124), .ZN(n19141) );
  INV_X1 U12470 ( .A(n11297), .ZN(n18913) );
  NAND2_X1 U12471 ( .A1(n18754), .A2(n11497), .ZN(n18978) );
  INV_X1 U12472 ( .A(n11293), .ZN(n18977) );
  NOR2_X1 U12473 ( .A1(n21818), .A2(n18998), .ZN(n21820) );
  INV_X1 U12474 ( .A(n11296), .ZN(n18792) );
  INV_X1 U12475 ( .A(n22039), .ZN(n22055) );
  INV_X1 U12476 ( .A(n21884), .ZN(n22022) );
  AOI21_X1 U12477 ( .B1(n21767), .B2(n21599), .A(n11300), .ZN(n19143) );
  INV_X1 U12478 ( .A(n21950), .ZN(n21941) );
  INV_X1 U12479 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22076) );
  INV_X1 U12480 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n22080) );
  NOR2_X1 U12481 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n22100), .ZN(
        n22105) );
  CLKBUF_X1 U12482 ( .A(n19565), .Z(n19897) );
  AOI21_X1 U12483 ( .B1(n16677), .B2(n22231), .A(n14399), .ZN(n14400) );
  OAI211_X1 U12484 ( .C1(n14469), .C2(n19475), .A(n11231), .B(n11344), .ZN(
        P2_U2824) );
  INV_X1 U12485 ( .A(n14522), .ZN(n11344) );
  INV_X1 U12486 ( .A(n13010), .ZN(n13011) );
  OAI21_X1 U12487 ( .B1(n19478), .B2(n17432), .A(n13009), .ZN(n13010) );
  NOR2_X1 U12488 ( .A1(n14905), .A2(n11471), .ZN(n15095) );
  INV_X1 U12489 ( .A(n14469), .ZN(n20004) );
  OAI21_X1 U12490 ( .B1(n19476), .B2(n20515), .A(n13002), .ZN(n13003) );
  OR2_X1 U12491 ( .A1(n16442), .A2(n18190), .ZN(n11504) );
  NAND2_X1 U12492 ( .A1(n14434), .A2(n18198), .ZN(n12640) );
  NAND2_X1 U12493 ( .A1(n13024), .A2(n18200), .ZN(n13025) );
  INV_X1 U12494 ( .A(n11424), .ZN(n11423) );
  OAI21_X1 U12495 ( .B1(n16409), .B2(n18185), .A(n11425), .ZN(n11424) );
  AOI21_X1 U12496 ( .B1(n19445), .B2(n18199), .A(n14208), .ZN(n11425) );
  NOR2_X1 U12497 ( .A1(n17636), .A2(n17635), .ZN(n11331) );
  AOI21_X1 U12498 ( .B1(n17873), .B2(n18198), .A(n17649), .ZN(n17650) );
  INV_X1 U12499 ( .A(n14193), .ZN(n14194) );
  OAI21_X1 U12500 ( .B1(n16411), .B2(n19495), .A(n11247), .ZN(P2_U3018) );
  INV_X1 U12501 ( .A(n11308), .ZN(n11307) );
  NAND2_X1 U12502 ( .A1(n19493), .A2(n11327), .ZN(n19491) );
  NAND2_X1 U12503 ( .A1(n19490), .A2(n19489), .ZN(n11328) );
  NAND2_X1 U12504 ( .A1(n11283), .A2(n11281), .ZN(P3_U2834) );
  NOR2_X1 U12505 ( .A1(n11242), .A2(n11282), .ZN(n11281) );
  NOR2_X1 U12506 ( .A1(n18767), .A2(n21940), .ZN(n11282) );
  OR2_X1 U12507 ( .A1(n20869), .A2(n20920), .ZN(U212) );
  INV_X1 U12508 ( .A(n11870), .ZN(n12733) );
  NAND2_X1 U12509 ( .A1(n16593), .A2(n11474), .ZN(n16567) );
  INV_X1 U12510 ( .A(n13448), .ZN(n13476) );
  INV_X2 U12511 ( .A(n14625), .ZN(n14351) );
  AND2_X1 U12512 ( .A1(n16593), .A2(n11259), .ZN(n16555) );
  NAND2_X1 U12513 ( .A1(n16299), .A2(n16349), .ZN(n16348) );
  NAND2_X1 U12514 ( .A1(n17278), .A2(n17392), .ZN(n17384) );
  NAND2_X1 U12515 ( .A1(n12194), .A2(n11271), .ZN(n17563) );
  AND2_X1 U12516 ( .A1(n18015), .A2(n17925), .ZN(n11230) );
  NAND2_X1 U12517 ( .A1(n16380), .A2(n16379), .ZN(n16378) );
  XNOR2_X1 U12518 ( .A(n13323), .B(n15079), .ZN(n13528) );
  INV_X1 U12519 ( .A(n14200), .ZN(n11426) );
  NAND2_X1 U12520 ( .A1(n17278), .A2(n11264), .ZN(n17270) );
  OR2_X1 U12521 ( .A1(n14528), .A2(n19480), .ZN(n11231) );
  NAND2_X1 U12522 ( .A1(n12078), .A2(n17794), .ZN(n12079) );
  NAND2_X1 U12523 ( .A1(n11470), .A2(n11503), .ZN(n14921) );
  AND2_X1 U12524 ( .A1(n14928), .A2(n15087), .ZN(n15086) );
  NAND2_X1 U12525 ( .A1(n11462), .A2(n11465), .ZN(n15668) );
  AND2_X1 U12526 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11232) );
  OR2_X1 U12527 ( .A1(n17474), .A2(n17268), .ZN(n11233) );
  AND2_X2 U12528 ( .A1(n15026), .A2(n15025), .ZN(n13211) );
  INV_X1 U12529 ( .A(n15033), .ZN(n14866) );
  OR3_X2 U12530 ( .A1(n21640), .A2(n21622), .A3(n21609), .ZN(n11234) );
  INV_X2 U12531 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11713) );
  OR2_X1 U12532 ( .A1(n14520), .A2(n14204), .ZN(n11235) );
  AND2_X1 U12533 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11237) );
  NAND2_X1 U12534 ( .A1(n17739), .A2(n17738), .ZN(n17740) );
  NAND2_X1 U12535 ( .A1(n18014), .A2(n12189), .ZN(n17679) );
  NAND2_X1 U12536 ( .A1(n16299), .A2(n11477), .ZN(n16657) );
  NOR2_X1 U12537 ( .A1(n14222), .A2(n11274), .ZN(n13220) );
  OR2_X1 U12538 ( .A1(n17484), .A2(n17474), .ZN(n11238) );
  AND2_X1 U12539 ( .A1(n15274), .A2(n12677), .ZN(n11239) );
  INV_X1 U12540 ( .A(n11445), .ZN(n11444) );
  NOR2_X1 U12541 ( .A1(n12189), .A2(n11446), .ZN(n11445) );
  AND2_X1 U12542 ( .A1(n17279), .A2(n17280), .ZN(n17278) );
  AND2_X1 U12543 ( .A1(n16593), .A2(n13815), .ZN(n16578) );
  OR2_X1 U12544 ( .A1(n14893), .A2(n14892), .ZN(n11241) );
  AND3_X1 U12545 ( .A1(n21939), .A2(n22039), .A3(n21938), .ZN(n11242) );
  OR2_X1 U12546 ( .A1(n16531), .A2(n11373), .ZN(n11243) );
  OAI21_X1 U12547 ( .B1(n16341), .B2(n11400), .A(n11399), .ZN(n16898) );
  NOR2_X1 U12548 ( .A1(n11412), .A2(n16819), .ZN(n16812) );
  NAND2_X1 U12549 ( .A1(n14812), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13241) );
  NOR2_X1 U12550 ( .A1(n12098), .A2(n12093), .ZN(n11244) );
  AND2_X1 U12551 ( .A1(n14201), .A2(n14202), .ZN(n13014) );
  NAND2_X1 U12552 ( .A1(n17589), .A2(n12079), .ZN(n17566) );
  AND2_X1 U12553 ( .A1(n11497), .A2(n22004), .ZN(n11246) );
  AND2_X1 U12554 ( .A1(n17264), .A2(n12113), .ZN(n14199) );
  INV_X1 U12555 ( .A(n12005), .ZN(n11438) );
  NOR2_X1 U12556 ( .A1(n16410), .A2(n11307), .ZN(n11247) );
  AND2_X1 U12557 ( .A1(n14180), .A2(n14179), .ZN(n12982) );
  OR2_X1 U12558 ( .A1(n12031), .A2(n12029), .ZN(n11248) );
  AND2_X1 U12559 ( .A1(n17406), .A2(n17296), .ZN(n17279) );
  NAND2_X1 U12560 ( .A1(n14200), .A2(n17557), .ZN(n11250) );
  OR2_X1 U12561 ( .A1(n18749), .A2(n21752), .ZN(n11251) );
  OR2_X1 U12562 ( .A1(n16517), .A2(n11480), .ZN(n14210) );
  AND2_X1 U12563 ( .A1(n11734), .A2(n11733), .ZN(n11252) );
  AND2_X1 U12564 ( .A1(n12084), .A2(n12079), .ZN(n11253) );
  AND2_X1 U12565 ( .A1(n11378), .A2(n11377), .ZN(n11254) );
  AND2_X1 U12566 ( .A1(n11426), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11255) );
  INV_X1 U12567 ( .A(n11386), .ZN(n11803) );
  NAND2_X1 U12568 ( .A1(n11384), .A2(n11802), .ZN(n11386) );
  NAND4_X1 U12569 ( .A1(n11653), .A2(n11652), .A3(n11487), .A4(n11651), .ZN(
        n12113) );
  NAND2_X1 U12570 ( .A1(n11326), .A2(n11325), .ZN(n12351) );
  AND2_X1 U12571 ( .A1(n14897), .A2(n13036), .ZN(n13179) );
  NOR2_X1 U12572 ( .A1(n15192), .A2(n11466), .ZN(n15636) );
  NAND2_X1 U12573 ( .A1(n17326), .A2(n17328), .ZN(n17327) );
  NOR2_X1 U12574 ( .A1(n15192), .A2(n15593), .ZN(n15592) );
  NAND2_X1 U12575 ( .A1(n11495), .A2(n16637), .ZN(n11256) );
  OR2_X1 U12576 ( .A1(n17447), .A2(n16398), .ZN(n11257) );
  AND2_X1 U12577 ( .A1(n14310), .A2(n16637), .ZN(n11258) );
  AND2_X1 U12578 ( .A1(n17438), .A2(n17440), .ZN(n17311) );
  NAND2_X1 U12579 ( .A1(n15664), .A2(n11381), .ZN(n14534) );
  NAND2_X1 U12580 ( .A1(n12686), .A2(n12685), .ZN(n14743) );
  AND2_X1 U12581 ( .A1(n15664), .A2(n12236), .ZN(n16255) );
  NAND2_X1 U12582 ( .A1(n12132), .A2(n12333), .ZN(n12573) );
  AND2_X1 U12583 ( .A1(n12673), .A2(n12696), .ZN(n15495) );
  INV_X1 U12584 ( .A(n11321), .ZN(n14537) );
  AND2_X1 U12585 ( .A1(n11473), .A2(n11474), .ZN(n11259) );
  NOR2_X1 U12586 ( .A1(n12532), .A2(n16389), .ZN(n11260) );
  AND4_X1 U12587 ( .A1(n13099), .A2(n13098), .A3(n13097), .A4(n13448), .ZN(
        n14372) );
  OR2_X1 U12588 ( .A1(n16496), .A2(n11480), .ZN(n11261) );
  AND2_X1 U12589 ( .A1(n14282), .A2(n16265), .ZN(n11262) );
  AND2_X1 U12590 ( .A1(n11258), .A2(n11371), .ZN(n11263) );
  INV_X1 U12591 ( .A(n11345), .ZN(n14515) );
  NOR2_X1 U12592 ( .A1(n14475), .A2(n17583), .ZN(n11345) );
  INV_X1 U12593 ( .A(n13344), .ZN(n11409) );
  NOR2_X1 U12594 ( .A1(n15192), .A2(n11463), .ZN(n16253) );
  INV_X1 U12595 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U12596 ( .A1(n14928), .A2(n11378), .ZN(n15193) );
  NAND2_X1 U12597 ( .A1(n20819), .A2(n11262), .ZN(n16303) );
  AND2_X1 U12598 ( .A1(n15486), .A2(n11316), .ZN(n16276) );
  INV_X1 U12599 ( .A(n22027), .ZN(n22044) );
  AND2_X1 U12600 ( .A1(n16133), .A2(n22115), .ZN(n22027) );
  XNOR2_X1 U12601 ( .A(n13221), .B(n13260), .ZN(n14961) );
  NAND2_X1 U12602 ( .A1(n11495), .A2(n11258), .ZN(n16610) );
  INV_X1 U12603 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13030) );
  AND2_X1 U12604 ( .A1(n17392), .A2(n11387), .ZN(n11264) );
  OR2_X1 U12605 ( .A1(n12487), .A2(n12486), .ZN(n15669) );
  OR2_X1 U12606 ( .A1(n11627), .A2(n11626), .ZN(n11911) );
  AND2_X1 U12607 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11265) );
  AND2_X1 U12608 ( .A1(n11232), .A2(n11265), .ZN(n11266) );
  AND2_X1 U12609 ( .A1(n16661), .A2(n16696), .ZN(n11267) );
  AND2_X1 U12610 ( .A1(n11460), .A2(n12863), .ZN(n11268) );
  INV_X1 U12611 ( .A(n18184), .ZN(n18200) );
  OR2_X1 U12612 ( .A1(n19539), .A2(n12819), .ZN(n18184) );
  OR2_X1 U12613 ( .A1(n18760), .A2(n11347), .ZN(n11269) );
  AND2_X1 U12614 ( .A1(n18168), .A2(n15360), .ZN(n19459) );
  AND2_X1 U12615 ( .A1(n12953), .A2(n12928), .ZN(n11270) );
  AND2_X1 U12616 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11271) );
  INV_X1 U12617 ( .A(n16252), .ZN(n11464) );
  NAND2_X1 U12618 ( .A1(n11326), .A2(n11324), .ZN(n15349) );
  AND2_X1 U12619 ( .A1(n11271), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11272) );
  INV_X1 U12620 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11349) );
  INV_X1 U12621 ( .A(n17925), .ZN(n11446) );
  INV_X1 U12622 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11336) );
  INV_X1 U12623 ( .A(n22376), .ZN(n22342) );
  OAI21_X2 U12624 ( .B1(n15138), .B2(n16722), .A(n15003), .ZN(n22582) );
  OAI21_X2 U12625 ( .B1(n15138), .B2(n14956), .A(n14955), .ZN(n22602) );
  OAI21_X2 U12626 ( .B1(n15138), .B2(n14982), .A(n14981), .ZN(n22624) );
  NOR3_X2 U12627 ( .A1(n20132), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20601) );
  OAI21_X2 U12628 ( .B1(n13434), .B2(n16982), .A(n16955), .ZN(n16796) );
  NAND3_X1 U12629 ( .A1(n11398), .A2(n13419), .A3(n11278), .ZN(n11277) );
  NAND2_X1 U12630 ( .A1(n17229), .A2(n22396), .ZN(n13314) );
  XNOR2_X2 U12631 ( .A(n14740), .B(n15211), .ZN(n17229) );
  NAND2_X2 U12632 ( .A1(n13394), .A2(n13405), .ZN(n13412) );
  NAND3_X1 U12633 ( .A1(n13394), .A2(n13559), .A3(n13235), .ZN(n13388) );
  NAND3_X1 U12634 ( .A1(n11288), .A2(n18767), .A3(n11284), .ZN(n11283) );
  NAND3_X1 U12635 ( .A1(n21927), .A2(n21926), .A3(n21950), .ZN(n11286) );
  NOR2_X2 U12636 ( .A1(n19058), .A2(n18732), .ZN(n19046) );
  OAI21_X1 U12637 ( .B1(n11300), .B2(n19134), .A(n19133), .ZN(n21688) );
  NAND2_X1 U12638 ( .A1(n19134), .A2(n11300), .ZN(n19133) );
  NAND2_X2 U12639 ( .A1(n21622), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14041) );
  INV_X4 U12640 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21622) );
  NAND2_X1 U12641 ( .A1(n16269), .A2(n11982), .ZN(n16315) );
  OAI211_X2 U12642 ( .C1(n16269), .C2(n11303), .A(n11301), .B(n11989), .ZN(
        n17702) );
  INV_X1 U12643 ( .A(n11982), .ZN(n11302) );
  INV_X4 U12644 ( .A(n12376), .ZN(n12954) );
  NAND2_X1 U12645 ( .A1(n12642), .A2(n17696), .ZN(n17684) );
  XNOR2_X2 U12646 ( .A(n11966), .B(n11965), .ZN(n15565) );
  NAND4_X1 U12647 ( .A1(n11866), .A2(n11869), .A3(n11867), .A4(n11868), .ZN(
        n11305) );
  NAND4_X1 U12648 ( .A1(n11906), .A2(n11905), .A3(n11908), .A4(n11907), .ZN(
        n11306) );
  AOI21_X1 U12649 ( .B1(n17465), .B2(n19500), .A(n11309), .ZN(n11308) );
  XNOR2_X1 U12650 ( .A(n11318), .B(n15558), .ZN(n20263) );
  NOR2_X2 U12651 ( .A1(n17484), .A2(n11233), .ZN(n17267) );
  XNOR2_X1 U12652 ( .A(n17267), .B(n16403), .ZN(n19455) );
  AND2_X2 U12653 ( .A1(n12538), .A2(n11319), .ZN(n17521) );
  NOR2_X2 U12654 ( .A1(n17327), .A2(n17922), .ZN(n11321) );
  NAND2_X1 U12655 ( .A1(n15197), .A2(n18033), .ZN(n15265) );
  NOR2_X1 U12656 ( .A1(n18057), .A2(n12425), .ZN(n15199) );
  NAND2_X2 U12657 ( .A1(n11535), .A2(n11534), .ZN(n12376) );
  AND2_X2 U12658 ( .A1(n11825), .A2(n11796), .ZN(n11804) );
  INV_X1 U12659 ( .A(n11750), .ZN(n11326) );
  NOR2_X1 U12660 ( .A1(n11181), .A2(n11328), .ZN(n11327) );
  INV_X1 U12661 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11330) );
  NOR2_X2 U12662 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15312) );
  AND3_X2 U12663 ( .A1(n15277), .A2(n11330), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11682) );
  OAI211_X1 U12664 ( .C1(n17865), .C2(n18184), .A(n11332), .B(n11331), .ZN(
        P2_U2995) );
  NAND2_X1 U12665 ( .A1(n17863), .A2(n18198), .ZN(n11332) );
  NAND2_X2 U12666 ( .A1(n17598), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17930) );
  NAND3_X1 U12667 ( .A1(n11244), .A2(n17570), .A3(n11335), .ZN(n12107) );
  AND2_X2 U12668 ( .A1(n17589), .A2(n11334), .ZN(n17570) );
  INV_X1 U12669 ( .A(n11337), .ZN(n14512) );
  AND2_X2 U12670 ( .A1(n12075), .A2(n12074), .ZN(n12081) );
  NOR2_X2 U12671 ( .A1(n12115), .A2(n11341), .ZN(n11951) );
  NOR2_X1 U12672 ( .A1(n12337), .A2(n11346), .ZN(n12134) );
  INV_X1 U12673 ( .A(n11352), .ZN(n14025) );
  XNOR2_X2 U12674 ( .A(n11350), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14024) );
  INV_X1 U12675 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11351) );
  INV_X1 U12676 ( .A(n14034), .ZN(n14026) );
  NAND2_X1 U12677 ( .A1(n21406), .A2(n21407), .ZN(n14038) );
  NAND2_X1 U12678 ( .A1(n21392), .A2(n21393), .ZN(n21390) );
  NAND2_X1 U12679 ( .A1(n21380), .A2(n21199), .ZN(n21392) );
  NOR2_X2 U12680 ( .A1(n21115), .A2(n18795), .ZN(n18794) );
  NAND3_X1 U12681 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19086) );
  CLKBUF_X1 U12682 ( .A(n13131), .Z(n11354) );
  AND2_X4 U12683 ( .A1(n11221), .A2(n15025), .ZN(n15033) );
  OAI22_X1 U12684 ( .A1(n11243), .A2(n16487), .B1(n16497), .B2(n14351), .ZN(
        n16489) );
  NOR3_X2 U12685 ( .A1(n16531), .A2(n11373), .A3(n16498), .ZN(n16497) );
  XNOR2_X2 U12686 ( .A(n12639), .B(n11383), .ZN(n16442) );
  NAND2_X2 U12687 ( .A1(n11820), .A2(n11831), .ZN(n11825) );
  AND2_X2 U12688 ( .A1(n11385), .A2(n12200), .ZN(n14910) );
  NOR2_X2 U12689 ( .A1(n17408), .A2(n17407), .ZN(n17406) );
  AND2_X4 U12690 ( .A1(n11390), .A2(n14712), .ZN(n13115) );
  AND2_X2 U12691 ( .A1(n13038), .A2(n11390), .ZN(n13081) );
  NAND3_X1 U12692 ( .A1(n14871), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n13244), .ZN(n11391) );
  NAND2_X1 U12693 ( .A1(n14871), .A2(n13244), .ZN(n11394) );
  NAND2_X1 U12694 ( .A1(n11393), .A2(n22158), .ZN(n11392) );
  INV_X1 U12695 ( .A(n13244), .ZN(n11393) );
  NAND2_X1 U12696 ( .A1(n11394), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13295) );
  NAND2_X1 U12697 ( .A1(n16341), .A2(n11401), .ZN(n11398) );
  NAND2_X1 U12698 ( .A1(n11410), .A2(n20832), .ZN(n11403) );
  INV_X1 U12699 ( .A(n20832), .ZN(n11404) );
  NAND2_X1 U12700 ( .A1(n11407), .A2(n11405), .ZN(n20837) );
  NOR2_X1 U12701 ( .A1(n11410), .A2(n11409), .ZN(n11406) );
  INV_X1 U12702 ( .A(n11408), .ZN(n11407) );
  OAI21_X1 U12703 ( .B1(n11409), .B2(n20832), .A(n20838), .ZN(n11408) );
  NAND2_X1 U12704 ( .A1(n20833), .A2(n20832), .ZN(n20831) );
  NAND3_X1 U12705 ( .A1(n13434), .A2(n13430), .A3(n11411), .ZN(n16798) );
  NAND2_X1 U12706 ( .A1(n16798), .A2(n16796), .ZN(n16806) );
  NAND2_X1 U12707 ( .A1(n11413), .A2(n16956), .ZN(n16858) );
  NAND3_X1 U12708 ( .A1(n16857), .A2(n14330), .A3(n16858), .ZN(n16830) );
  NAND2_X2 U12709 ( .A1(n16860), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16857) );
  AND2_X1 U12710 ( .A1(n13428), .A2(n13427), .ZN(n11415) );
  NAND2_X1 U12711 ( .A1(n14198), .A2(n14199), .ZN(n11427) );
  OAI211_X1 U12712 ( .C1(n11422), .C2(n17555), .A(n11419), .B(n11418), .ZN(
        n16411) );
  NAND2_X1 U12713 ( .A1(n17555), .A2(n11255), .ZN(n11418) );
  OAI21_X1 U12714 ( .B1(n16411), .B2(n18184), .A(n11423), .ZN(P2_U2986) );
  NAND2_X1 U12715 ( .A1(n14198), .A2(n11420), .ZN(n11421) );
  NAND3_X1 U12716 ( .A1(n11752), .A2(n20528), .A3(n11732), .ZN(n11430) );
  NAND3_X1 U12717 ( .A1(n11322), .A2(n11386), .A3(n12201), .ZN(n11456) );
  NAND3_X1 U12718 ( .A1(n11440), .A2(n11439), .A3(n11438), .ZN(n11431) );
  AND2_X2 U12719 ( .A1(n11433), .A2(n11432), .ZN(n12642) );
  NAND3_X1 U12720 ( .A1(n11440), .A2(n11439), .A3(n11434), .ZN(n11433) );
  NAND2_X1 U12721 ( .A1(n11990), .A2(n17702), .ZN(n11440) );
  NAND2_X1 U12722 ( .A1(n18016), .A2(n18015), .ZN(n18014) );
  NAND3_X2 U12723 ( .A1(n12178), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n12166), .ZN(n16319) );
  AND2_X1 U12724 ( .A1(n11190), .A2(n12166), .ZN(n16318) );
  XNOR2_X1 U12725 ( .A(n12162), .B(n12181), .ZN(n12168) );
  NAND3_X1 U12726 ( .A1(n12142), .A2(n12143), .A3(n12416), .ZN(n12141) );
  INV_X2 U12727 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15277) );
  NAND3_X1 U12728 ( .A1(n12929), .A2(n12928), .A3(n17374), .ZN(n11453) );
  NAND3_X1 U12729 ( .A1(n12929), .A2(n11270), .A3(n17374), .ZN(n12955) );
  NOR2_X2 U12730 ( .A1(n17363), .A2(n12956), .ZN(n12977) );
  INV_X1 U12731 ( .A(n12953), .ZN(n11452) );
  NAND2_X2 U12732 ( .A1(n11456), .A2(n11454), .ZN(n15274) );
  OAI21_X2 U12733 ( .B1(n11804), .B2(n11803), .A(n11455), .ZN(n11454) );
  NAND2_X1 U12734 ( .A1(n17395), .A2(n11459), .ZN(n11458) );
  NAND3_X1 U12735 ( .A1(n13099), .A2(n13098), .A3(n13097), .ZN(n13165) );
  NAND2_X1 U12736 ( .A1(n16593), .A2(n11472), .ZN(n16543) );
  NOR2_X1 U12737 ( .A1(n16517), .A2(n16519), .ZN(n14209) );
  NOR2_X2 U12738 ( .A1(n16517), .A2(n11261), .ZN(n16495) );
  NAND2_X1 U12739 ( .A1(n13258), .A2(n13253), .ZN(n13510) );
  NAND3_X1 U12740 ( .A1(n13258), .A2(n13286), .A3(n11482), .ZN(n13323) );
  NAND3_X1 U12741 ( .A1(n11484), .A2(n14740), .A3(n22396), .ZN(n11483) );
  INV_X1 U12742 ( .A(n11731), .ZN(n11733) );
  AND2_X1 U12743 ( .A1(n17411), .A2(n13007), .ZN(n17419) );
  NAND2_X1 U12744 ( .A1(n11825), .A2(n11178), .ZN(n11819) );
  AOI22_X1 U12745 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13055) );
  OR2_X1 U12746 ( .A1(n12672), .A2(n12671), .ZN(n12673) );
  NAND2_X1 U12747 ( .A1(n17397), .A2(n17396), .ZN(n17395) );
  OAI21_X2 U12748 ( .B1(n17400), .B2(n17401), .A(n12821), .ZN(n17397) );
  OR2_X2 U12749 ( .A1(n11857), .A2(n11860), .ZN(n20117) );
  NAND2_X1 U12750 ( .A1(n11239), .A2(n11848), .ZN(n20060) );
  OAI22_X1 U12751 ( .A1(n11927), .A2(n12830), .B1(n11843), .B2(n20040), .ZN(
        n11844) );
  NAND2_X1 U12752 ( .A1(n11239), .A2(n11839), .ZN(n20040) );
  INV_X1 U12753 ( .A(n13093), .ZN(n13170) );
  NAND2_X1 U12754 ( .A1(n11731), .A2(n11707), .ZN(n11708) );
  CLKBUF_X1 U12755 ( .A(n13264), .Z(n13296) );
  NAND2_X1 U12756 ( .A1(n14357), .A2(n15025), .ZN(n16465) );
  INV_X1 U12757 ( .A(n13167), .ZN(n14249) );
  AOI22_X1 U12758 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13081), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13056) );
  AND2_X1 U12759 ( .A1(n12976), .A2(n12975), .ZN(n11486) );
  AND4_X1 U12760 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11487) );
  AND3_X1 U12761 ( .A1(n18145), .A2(n14840), .A3(n16472), .ZN(n20853) );
  INV_X1 U12762 ( .A(n19495), .ZN(n14175) );
  OR2_X1 U12763 ( .A1(n19478), .A2(n18190), .ZN(n11488) );
  AND2_X1 U12764 ( .A1(n17095), .A2(n16870), .ZN(n11489) );
  OR2_X1 U12765 ( .A1(n13443), .A2(n13442), .ZN(n11490) );
  OR4_X1 U12766 ( .A1(n18156), .A2(n22132), .A3(n18155), .A4(n18154), .ZN(
        n11491) );
  AND2_X1 U12767 ( .A1(n16955), .A2(n16797), .ZN(n11492) );
  AND4_X1 U12768 ( .A1(n14072), .A2(n14071), .A3(n14070), .A4(n14069), .ZN(
        n11493) );
  INV_X1 U12769 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22396) );
  OR2_X2 U12770 ( .A1(n11857), .A2(n11842), .ZN(n11919) );
  INV_X1 U12771 ( .A(n12838), .ZN(n12820) );
  AND2_X1 U12772 ( .A1(n17620), .A2(n17623), .ZN(n11494) );
  AND2_X2 U12773 ( .A1(n16648), .A2(n14303), .ZN(n11495) );
  INV_X1 U12774 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12635) );
  OR2_X1 U12775 ( .A1(n19596), .A2(n19902), .ZN(n19653) );
  AND2_X1 U12776 ( .A1(n11520), .A2(n11519), .ZN(n11496) );
  AND2_X1 U12777 ( .A1(n18751), .A2(n11506), .ZN(n11497) );
  OR2_X1 U12778 ( .A1(n21936), .A2(n21935), .ZN(n11498) );
  AND2_X1 U12779 ( .A1(n13022), .A2(n13021), .ZN(n11499) );
  INV_X1 U12780 ( .A(n11851), .ZN(n11846) );
  AND3_X1 U12781 ( .A1(n14212), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11500) );
  OR2_X1 U12782 ( .A1(n17710), .A2(n17709), .ZN(n11501) );
  INV_X1 U12783 ( .A(n11860), .ZN(n11828) );
  INV_X1 U12784 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18108) );
  AND2_X1 U12785 ( .A1(n11807), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11502) );
  AND2_X1 U12786 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U12787 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13035) );
  OR2_X1 U12788 ( .A1(n22419), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19239) );
  OR2_X1 U12789 ( .A1(n18983), .A2(n21200), .ZN(n11505) );
  NOR2_X2 U12790 ( .A1(n20939), .A2(n18086), .ZN(n21893) );
  INV_X1 U12791 ( .A(n21893), .ZN(n16106) );
  NAND2_X1 U12792 ( .A1(n11706), .A2(n11705), .ZN(n11744) );
  INV_X1 U12793 ( .A(n15191), .ZN(n12698) );
  OR2_X1 U12794 ( .A1(n19044), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11506) );
  INV_X1 U12795 ( .A(n19044), .ZN(n18749) );
  OR2_X1 U12796 ( .A1(n16506), .A2(n16972), .ZN(n11507) );
  AND3_X1 U12797 ( .A1(n13041), .A2(n13040), .A3(n13039), .ZN(n11508) );
  INV_X1 U12798 ( .A(n13110), .ZN(n13863) );
  AND2_X1 U12799 ( .A1(n13088), .A2(n13087), .ZN(n11509) );
  AND3_X1 U12800 ( .A1(n13059), .A2(n13058), .A3(n13057), .ZN(n11510) );
  AND4_X1 U12801 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n11511) );
  AND2_X1 U12802 ( .A1(n13168), .A2(n14361), .ZN(n13162) );
  INV_X1 U12803 ( .A(n14199), .ZN(n12097) );
  OR2_X1 U12804 ( .A1(n13356), .A2(n13355), .ZN(n13384) );
  OAI22_X1 U12805 ( .A1(n11891), .A2(n11918), .B1(n15509), .B2(n12729), .ZN(
        n11894) );
  INV_X1 U12806 ( .A(n13086), .ZN(n13190) );
  INV_X1 U12807 ( .A(n13323), .ZN(n13324) );
  OR2_X1 U12808 ( .A1(n13233), .A2(n13232), .ZN(n13246) );
  INV_X1 U12809 ( .A(n12023), .ZN(n11656) );
  NOR2_X1 U12810 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  INV_X1 U12811 ( .A(n11777), .ZN(n11794) );
  INV_X1 U12812 ( .A(n12394), .ZN(n12396) );
  OR2_X1 U12813 ( .A1(n14155), .A2(n14156), .ZN(n14151) );
  INV_X1 U12814 ( .A(n13489), .ZN(n13468) );
  AOI21_X1 U12815 ( .B1(n13115), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n13028), .ZN(n13034) );
  INV_X1 U12816 ( .A(n13833), .ZN(n13834) );
  OR2_X1 U12817 ( .A1(n13378), .A2(n13377), .ZN(n13396) );
  OR2_X1 U12818 ( .A1(n13312), .A2(n13311), .ZN(n13338) );
  INV_X1 U12819 ( .A(n13274), .ZN(n13256) );
  AOI22_X1 U12820 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13081), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13085) );
  AND2_X1 U12821 ( .A1(n12132), .A2(n12324), .ZN(n12337) );
  INV_X1 U12822 ( .A(n12584), .ZN(n11728) );
  INV_X1 U12823 ( .A(n12910), .ZN(n12911) );
  NAND2_X1 U12824 ( .A1(n12885), .A2(n12887), .ZN(n12888) );
  NAND2_X1 U12825 ( .A1(n12104), .A2(n14196), .ZN(n12105) );
  NAND2_X1 U12826 ( .A1(n12057), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12058) );
  NAND2_X1 U12827 ( .A1(n12666), .A2(n20165), .ZN(n12687) );
  AOI22_X1 U12828 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11218), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11673) );
  OAI21_X1 U12829 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21033), .A(
        n14151), .ZN(n14152) );
  NAND2_X1 U12830 ( .A1(n13468), .A2(n13235), .ZN(n13494) );
  INV_X1 U12831 ( .A(n16740), .ZN(n13815) );
  NOR2_X1 U12832 ( .A1(n13896), .A2(n13895), .ZN(n13897) );
  NAND2_X1 U12833 ( .A1(n14735), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13979) );
  NOR2_X1 U12834 ( .A1(n17126), .A2(n13423), .ZN(n13424) );
  NAND3_X1 U12835 ( .A1(n14409), .A2(n15025), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13489) );
  NAND2_X1 U12836 ( .A1(n13314), .A2(n13313), .ZN(n15079) );
  INV_X1 U12837 ( .A(n17370), .ZN(n12928) );
  NAND2_X1 U12838 ( .A1(n12375), .A2(n12379), .ZN(n12380) );
  AOI21_X1 U12839 ( .B1(n14189), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14188), .ZN(n14190) );
  INV_X1 U12840 ( .A(n19442), .ZN(n12099) );
  OR2_X1 U12841 ( .A1(n17737), .A2(n17734), .ZN(n18018) );
  INV_X1 U12842 ( .A(n12171), .ZN(n12164) );
  NAND2_X1 U12843 ( .A1(n11203), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11790) );
  INV_X1 U12844 ( .A(n11842), .ZN(n11839) );
  NOR2_X1 U12845 ( .A1(n21005), .A2(n21651), .ZN(n14090) );
  NOR2_X1 U12846 ( .A1(n14041), .A2(n14043), .ZN(n14092) );
  INV_X1 U12847 ( .A(n21475), .ZN(n16234) );
  INV_X1 U12848 ( .A(n21617), .ZN(n16241) );
  OR2_X1 U12849 ( .A1(n13494), .A2(n14233), .ZN(n13500) );
  OR2_X1 U12850 ( .A1(n13462), .A2(n13458), .ZN(n13459) );
  NAND2_X1 U12851 ( .A1(n15130), .A2(n11221), .ZN(n14363) );
  AND2_X1 U12852 ( .A1(n13048), .A2(n13047), .ZN(n13050) );
  OR2_X1 U12853 ( .A1(n13920), .A2(n13919), .ZN(n13922) );
  AND2_X1 U12854 ( .A1(n13738), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13719) );
  INV_X1 U12855 ( .A(n13979), .ZN(n14003) );
  NAND2_X1 U12856 ( .A1(n13565), .A2(n13564), .ZN(n15659) );
  INV_X1 U12857 ( .A(n13701), .ZN(n13632) );
  AND2_X1 U12858 ( .A1(n14296), .A2(n14295), .ZN(n16663) );
  NAND2_X1 U12859 ( .A1(n15033), .A2(n14351), .ZN(n14344) );
  INV_X1 U12860 ( .A(n20823), .ZN(n14269) );
  INV_X1 U12861 ( .A(n11223), .ZN(n15427) );
  INV_X1 U12862 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18150) );
  AND2_X1 U12863 ( .A1(n12540), .A2(n12539), .ZN(n17314) );
  INV_X1 U12864 ( .A(n11960), .ZN(n11655) );
  INV_X1 U12865 ( .A(n16369), .ZN(n12699) );
  NAND2_X1 U12866 ( .A1(n12677), .A2(n15498), .ZN(n12682) );
  INV_X1 U12867 ( .A(n17374), .ZN(n17376) );
  INV_X1 U12868 ( .A(n12401), .ZN(n12415) );
  INV_X1 U12869 ( .A(n11746), .ZN(n12352) );
  OAI21_X1 U12870 ( .B1(n19458), .B2(n18066), .A(n14190), .ZN(n14191) );
  NAND2_X1 U12871 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12654) );
  AND2_X1 U12872 ( .A1(n19343), .A2(n12053), .ZN(n12648) );
  OR2_X1 U12873 ( .A1(n12593), .A2(n12592), .ZN(n17964) );
  NAND2_X1 U12874 ( .A1(n12389), .A2(n12388), .ZN(n12394) );
  INV_X1 U12875 ( .A(n11873), .ZN(n15285) );
  NAND2_X1 U12876 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18897) );
  AND2_X1 U12877 ( .A1(n18873), .A2(n21665), .ZN(n18758) );
  INV_X1 U12878 ( .A(n19010), .ZN(n18771) );
  OAI211_X1 U12879 ( .C1(n14148), .C2(n14147), .A(n14146), .B(n14145), .ZN(
        n21642) );
  INV_X1 U12880 ( .A(n18318), .ZN(n14138) );
  CLKBUF_X2 U12881 ( .A(n14064), .Z(n18717) );
  NAND2_X1 U12882 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  NAND2_X1 U12883 ( .A1(n13459), .A2(n13461), .ZN(n14233) );
  AND2_X1 U12884 ( .A1(n16537), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16523) );
  NAND2_X1 U12885 ( .A1(n13809), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13811) );
  NOR2_X1 U12886 ( .A1(n13633), .A2(n16965), .ZN(n13634) );
  OR2_X1 U12887 ( .A1(n22127), .A2(n15015), .ZN(n16584) );
  INV_X1 U12888 ( .A(n16472), .ZN(n16466) );
  INV_X1 U12889 ( .A(n14402), .ZN(n14403) );
  OAI21_X1 U12890 ( .B1(n13982), .B2(n16853), .A(n13861), .ZN(n16568) );
  AND2_X1 U12891 ( .A1(n13719), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13809) );
  AND2_X1 U12892 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n13718), .ZN(
        n13772) );
  INV_X1 U12893 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16965) );
  AND2_X1 U12894 ( .A1(n13539), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13551) );
  INV_X1 U12895 ( .A(n20857), .ZN(n16966) );
  AND2_X1 U12896 ( .A1(n16935), .A2(n16932), .ZN(n16918) );
  AND2_X1 U12897 ( .A1(n14301), .A2(n14300), .ZN(n16649) );
  AND2_X1 U12898 ( .A1(n14286), .A2(n14285), .ZN(n16350) );
  AND2_X1 U12899 ( .A1(n14274), .A2(n14273), .ZN(n15661) );
  INV_X1 U12900 ( .A(n22406), .ZN(n14840) );
  INV_X1 U12901 ( .A(n22470), .ZN(n22471) );
  INV_X1 U12902 ( .A(n17252), .ZN(n15632) );
  NAND2_X1 U12903 ( .A1(n15217), .A2(n11212), .ZN(n22735) );
  NOR2_X1 U12904 ( .A1(n15377), .A2(n15427), .ZN(n15217) );
  INV_X1 U12905 ( .A(n15139), .ZN(n15602) );
  OR2_X1 U12906 ( .A1(n15058), .A2(n15597), .ZN(n22551) );
  INV_X1 U12907 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22524) );
  INV_X1 U12908 ( .A(n22639), .ZN(n22643) );
  NAND2_X1 U12909 ( .A1(n11223), .A2(n15428), .ZN(n15597) );
  INV_X1 U12910 ( .A(n13982), .ZN(n15010) );
  INV_X1 U12911 ( .A(n12361), .ZN(n15332) );
  OR2_X1 U12912 ( .A1(n12109), .A2(n12108), .ZN(n14464) );
  INV_X1 U12913 ( .A(n17330), .ZN(n17354) );
  NAND2_X1 U12914 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n14496), .ZN(
        n14499) );
  NOR2_X1 U12915 ( .A1(n12343), .A2(n12127), .ZN(n14564) );
  NAND2_X1 U12916 ( .A1(n15496), .A2(n12697), .ZN(n14907) );
  NAND2_X1 U12917 ( .A1(n12820), .A2(n12819), .ZN(n12821) );
  AND2_X1 U12918 ( .A1(n19356), .A2(n12049), .ZN(n17652) );
  AND3_X1 U12919 ( .A1(n12606), .A2(n12605), .A3(n19497), .ZN(n18003) );
  OR2_X1 U12920 ( .A1(n12186), .A2(n11961), .ZN(n12187) );
  AND3_X1 U12921 ( .A1(n12422), .A2(n12421), .A3(n12420), .ZN(n15182) );
  OR2_X1 U12922 ( .A1(n20262), .A2(n18220), .ZN(n20092) );
  NAND2_X1 U12923 ( .A1(n20165), .A2(n20103), .ZN(n20192) );
  INV_X1 U12924 ( .A(n16129), .ZN(n22063) );
  NOR2_X1 U12925 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n21232), .ZN(n21247) );
  NOR2_X1 U12926 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n21205), .ZN(n21219) );
  NOR2_X1 U12927 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n21146), .ZN(n21163) );
  INV_X1 U12928 ( .A(n21521), .ZN(n14137) );
  AND2_X1 U12929 ( .A1(n21604), .A2(n21521), .ZN(n21546) );
  NOR2_X1 U12930 ( .A1(n16185), .A2(n16184), .ZN(n21599) );
  INV_X1 U12931 ( .A(n14028), .ZN(n18854) );
  INV_X1 U12932 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n21177) );
  NOR2_X1 U12933 ( .A1(n21752), .A2(n18771), .ZN(n21769) );
  INV_X1 U12934 ( .A(n19099), .ZN(n19113) );
  INV_X1 U12935 ( .A(n21463), .ZN(n21932) );
  NOR2_X1 U12936 ( .A1(n16242), .A2(n21646), .ZN(n21998) );
  AND2_X1 U12937 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21820), .ZN(
        n21810) );
  INV_X1 U12938 ( .A(n21967), .ZN(n21928) );
  NAND2_X2 U12939 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21656), .ZN(
        n21651) );
  INV_X1 U12940 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22069) );
  CLKBUF_X3 U12941 ( .A(n18475), .Z(n18548) );
  AND2_X1 U12942 ( .A1(n13502), .A2(n13501), .ZN(n16472) );
  OR2_X1 U12943 ( .A1(n13811), .A2(n13810), .ZN(n13833) );
  AND2_X1 U12944 ( .A1(n13634), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13670) );
  NOR2_X1 U12945 ( .A1(n15021), .A2(n15022), .ZN(n22360) );
  INV_X1 U12946 ( .A(n20830), .ZN(n16708) );
  INV_X1 U12947 ( .A(n14447), .ZN(n14449) );
  AND2_X1 U12948 ( .A1(n16791), .A2(n14426), .ZN(n16773) );
  NAND2_X1 U12949 ( .A1(n14720), .A2(n14840), .ZN(n14415) );
  INV_X2 U12950 ( .A(n14752), .ZN(n14809) );
  NAND2_X1 U12951 ( .A1(n13560), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13567) );
  INV_X1 U12952 ( .A(n14398), .ZN(n14399) );
  INV_X1 U12953 ( .A(n16648), .ZN(n17148) );
  INV_X1 U12954 ( .A(n22151), .ZN(n22225) );
  INV_X1 U12955 ( .A(n22182), .ZN(n22163) );
  AND2_X1 U12956 ( .A1(n14246), .A2(n14840), .ZN(n14378) );
  NAND2_X1 U12957 ( .A1(n16472), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17230) );
  INV_X1 U12958 ( .A(n22483), .ZN(n15432) );
  INV_X1 U12959 ( .A(n22681), .ZN(n22722) );
  NOR2_X2 U12960 ( .A1(n22483), .A2(n22471), .ZN(n22729) );
  NOR2_X2 U12961 ( .A1(n22483), .A2(n15597), .ZN(n22728) );
  AND2_X1 U12962 ( .A1(n15386), .A2(n11212), .ZN(n17252) );
  AND2_X1 U12963 ( .A1(n15386), .A2(n15428), .ZN(n22737) );
  AND2_X1 U12964 ( .A1(n15217), .A2(n15428), .ZN(n22693) );
  INV_X1 U12965 ( .A(n15058), .ZN(n15083) );
  NOR2_X1 U12966 ( .A1(n15141), .A2(n14977), .ZN(n22697) );
  AND2_X1 U12967 ( .A1(n15083), .A2(n22470), .ZN(n22749) );
  INV_X1 U12968 ( .A(n22551), .ZN(n22759) );
  INV_X1 U12969 ( .A(n22772), .ZN(n22535) );
  INV_X1 U12970 ( .A(n15684), .ZN(n22768) );
  OR2_X1 U12971 ( .A1(n18153), .A2(n18152), .ZN(n22398) );
  INV_X1 U12972 ( .A(n11997), .ZN(n12008) );
  OR2_X1 U12973 ( .A1(n18168), .A2(n14454), .ZN(n19371) );
  INV_X1 U12974 ( .A(n19477), .ZN(n19461) );
  OR2_X1 U12975 ( .A1(n12435), .A2(n12434), .ZN(n15094) );
  OR2_X1 U12976 ( .A1(n17444), .A2(n17434), .ZN(n17435) );
  NAND2_X1 U12977 ( .A1(n17416), .A2(n16388), .ZN(n17427) );
  OAI21_X1 U12978 ( .B1(n12997), .B2(n12996), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14661) );
  INV_X1 U12979 ( .A(n14701), .ZN(n14687) );
  AND2_X1 U12980 ( .A1(n18204), .A2(n14633), .ZN(n18196) );
  OAI211_X1 U12981 ( .C1(n16442), .C2(n18061), .A(n12617), .B(n12616), .ZN(
        n12618) );
  OR2_X1 U12982 ( .A1(n17723), .A2(n17724), .ZN(n17981) );
  AND2_X1 U12983 ( .A1(n12370), .A2(n19511), .ZN(n12621) );
  INV_X1 U12984 ( .A(n20199), .ZN(n20525) );
  NAND2_X1 U12985 ( .A1(n20204), .A2(n20203), .ZN(n20636) );
  INV_X1 U12986 ( .A(n20630), .ZN(n20633) );
  NOR2_X1 U12987 ( .A1(n20184), .A2(n20144), .ZN(n20610) );
  OR2_X1 U12988 ( .A1(n20255), .A2(n19269), .ZN(n20183) );
  INV_X1 U12989 ( .A(n20495), .ZN(n20602) );
  NOR2_X1 U12990 ( .A1(n20133), .A2(n20144), .ZN(n20488) );
  INV_X1 U12991 ( .A(n20581), .ZN(n20584) );
  NOR2_X2 U12992 ( .A1(n20092), .A2(n20183), .ZN(n20576) );
  NOR2_X2 U12993 ( .A1(n20092), .A2(n20163), .ZN(n20569) );
  NOR2_X2 U12994 ( .A1(n20092), .A2(n20144), .ZN(n20563) );
  NOR2_X1 U12995 ( .A1(n20100), .A2(n20092), .ZN(n20055) );
  INV_X1 U12996 ( .A(n20549), .ZN(n20538) );
  OAI22_X1 U12997 ( .A1(n20932), .A2(n20212), .B1(n19569), .B2(n20211), .ZN(
        n20185) );
  INV_X1 U12998 ( .A(n20401), .ZN(n20403) );
  NOR2_X2 U12999 ( .A1(n15507), .A2(n20164), .ZN(n20532) );
  AND3_X1 U13000 ( .A1(n18105), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n19511) );
  NOR2_X1 U13001 ( .A1(n21616), .A2(n14149), .ZN(n22062) );
  NAND2_X1 U13002 ( .A1(n21366), .A2(n21367), .ZN(n21365) );
  INV_X1 U13003 ( .A(n14164), .ZN(n14168) );
  INV_X1 U13004 ( .A(n21420), .ZN(n21377) );
  NOR2_X1 U13005 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n21173), .ZN(n21193) );
  NOR2_X1 U13006 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n21117), .ZN(n21141) );
  NAND2_X1 U13007 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18463), .ZN(n18448) );
  AOI21_X1 U13008 ( .B1(n18321), .B2(n18320), .A(n18319), .ZN(n21425) );
  NOR2_X1 U13009 ( .A1(n21503), .A2(n21508), .ZN(n21502) );
  INV_X2 U13010 ( .A(n21546), .ZN(n21588) );
  OR2_X1 U13011 ( .A1(n18871), .A2(n21658), .ZN(n21946) );
  INV_X1 U13012 ( .A(n18822), .ZN(n18986) );
  INV_X1 U13013 ( .A(n19057), .ZN(n19040) );
  INV_X1 U13014 ( .A(n19140), .ZN(n19074) );
  XOR2_X1 U13015 ( .A(n21698), .B(n16224), .Z(n19123) );
  NAND2_X1 U13016 ( .A1(n18980), .A2(n18979), .ZN(n19137) );
  AOI21_X1 U13017 ( .B1(n21763), .B2(n21817), .A(n22044), .ZN(n22050) );
  NOR2_X2 U13018 ( .A1(n22044), .A2(n21922), .ZN(n22039) );
  AND2_X1 U13019 ( .A1(n22117), .A2(n22027), .ZN(n21853) );
  NOR2_X1 U13020 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19568), .ZN(n19854) );
  INV_X1 U13021 ( .A(n19925), .ZN(n19933) );
  INV_X1 U13022 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19617) );
  INV_X1 U13023 ( .A(n22088), .ZN(n22115) );
  AND2_X1 U13024 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22421), .ZN(n19229) );
  NAND2_X1 U13025 ( .A1(n14622), .A2(n16472), .ZN(n16463) );
  NAND2_X1 U13026 ( .A1(n14624), .A2(n14623), .ZN(n22127) );
  OR2_X1 U13027 ( .A1(n14552), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22784) );
  INV_X1 U13028 ( .A(n22359), .ZN(n22377) );
  INV_X1 U13029 ( .A(n22360), .ZN(n22379) );
  INV_X1 U13030 ( .A(n20697), .ZN(n20718) );
  INV_X1 U13031 ( .A(n20853), .ZN(n22386) );
  OR2_X1 U13032 ( .A1(n20857), .A2(n14877), .ZN(n20856) );
  OR2_X1 U13033 ( .A1(n22393), .A2(n22534), .ZN(n16972) );
  INV_X1 U13034 ( .A(n22231), .ZN(n22245) );
  NAND2_X1 U13035 ( .A1(n14247), .A2(n14378), .ZN(n22226) );
  AOI22_X1 U13036 ( .A1(n22461), .A2(n22466), .B1(n22460), .B2(n22521), .ZN(
        n22719) );
  NAND2_X1 U13037 ( .A1(n15432), .A2(n15431), .ZN(n22681) );
  AOI22_X1 U13038 ( .A1(n22474), .A2(n22478), .B1(n22521), .B2(n22503), .ZN(
        n22726) );
  INV_X1 U13039 ( .A(n22490), .ZN(n22733) );
  NOR2_X1 U13040 ( .A1(n15603), .A2(n22507), .ZN(n17235) );
  AOI22_X1 U13041 ( .A1(n22504), .A2(n22510), .B1(n22540), .B2(n22503), .ZN(
        n22741) );
  NAND2_X1 U13042 ( .A1(n15083), .A2(n15102), .ZN(n22747) );
  AOI22_X1 U13043 ( .A1(n22522), .A2(n22530), .B1(n22521), .B2(n22520), .ZN(
        n22754) );
  INV_X1 U13044 ( .A(n15622), .ZN(n22585) );
  AOI22_X1 U13045 ( .A1(n22541), .A2(n22549), .B1(n22540), .B2(n22539), .ZN(
        n22765) );
  NAND2_X1 U13046 ( .A1(n15103), .A2(n15431), .ZN(n15684) );
  NAND2_X1 U13047 ( .A1(n15103), .A2(n22470), .ZN(n22782) );
  INV_X1 U13048 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n18164) );
  AND2_X1 U13049 ( .A1(n15331), .A2(n19511), .ZN(n18168) );
  AND4_X1 U13050 ( .A1(n19449), .A2(n19448), .A3(n19447), .A4(n19446), .ZN(
        n19454) );
  OR2_X1 U13051 ( .A1(n14463), .A2(n14460), .ZN(n19477) );
  OR3_X1 U13052 ( .A1(n14463), .A2(n14462), .A3(n14461), .ZN(n19441) );
  INV_X1 U13053 ( .A(n19459), .ZN(n19475) );
  AND2_X1 U13054 ( .A1(n13006), .A2(n19511), .ZN(n17411) );
  INV_X1 U13055 ( .A(n13003), .ZN(n13004) );
  INV_X1 U13056 ( .A(n20461), .ZN(n20517) );
  NAND2_X2 U13057 ( .A1(n12981), .A2(n12980), .ZN(n20513) );
  AND2_X1 U13058 ( .A1(n20010), .A2(n20009), .ZN(n20465) );
  INV_X1 U13059 ( .A(n18238), .ZN(n18268) );
  NAND2_X1 U13060 ( .A1(n14580), .A2(n12819), .ZN(n14701) );
  NAND2_X1 U13061 ( .A1(n19539), .A2(n12314), .ZN(n18204) );
  INV_X1 U13062 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19313) );
  INV_X1 U13063 ( .A(n18196), .ZN(n18181) );
  INV_X1 U13064 ( .A(n12618), .ZN(n12625) );
  NAND2_X1 U13065 ( .A1(n12621), .A2(n15342), .ZN(n19495) );
  NAND2_X1 U13066 ( .A1(n12621), .A2(n12373), .ZN(n18061) );
  INV_X1 U13067 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20145) );
  OR2_X1 U13068 ( .A1(n20184), .A2(n20183), .ZN(n20630) );
  OR2_X1 U13069 ( .A1(n20184), .A2(n20100), .ZN(n20615) );
  INV_X1 U13070 ( .A(n20610), .ZN(n20622) );
  AOI21_X1 U13071 ( .B1(n16286), .B2(n16292), .A(n16285), .ZN(n20608) );
  INV_X1 U13072 ( .A(n20590), .ZN(n20600) );
  INV_X1 U13073 ( .A(n20488), .ZN(n20594) );
  INV_X1 U13074 ( .A(n20576), .ZN(n20487) );
  AND2_X1 U13075 ( .A1(n20091), .A2(n20090), .ZN(n20574) );
  AOI21_X1 U13076 ( .B1(n20079), .B2(n20084), .A(n20078), .ZN(n20567) );
  INV_X1 U13077 ( .A(n20055), .ZN(n20561) );
  NAND2_X1 U13078 ( .A1(n15720), .A2(n15506), .ZN(n20549) );
  NAND2_X1 U13079 ( .A1(n15720), .A2(n15719), .ZN(n20543) );
  INV_X1 U13080 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n18105) );
  INV_X1 U13081 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18270) );
  NOR2_X1 U13082 ( .A1(n22062), .A2(n20949), .ZN(n20942) );
  AND2_X1 U13083 ( .A1(n14171), .A2(n21402), .ZN(n14172) );
  NAND4_X1 U13084 ( .A1(n14168), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n20937), 
        .A4(n14162), .ZN(n21385) );
  OR2_X1 U13085 ( .A1(n21231), .A2(n21230), .ZN(n21241) );
  NAND2_X1 U13086 ( .A1(n21306), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21375) );
  NAND2_X1 U13087 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18586), .ZN(n18630) );
  NOR2_X1 U13088 ( .A1(n16144), .A2(n16143), .ZN(n21463) );
  NOR2_X1 U13089 ( .A1(n16206), .A2(n16205), .ZN(n21475) );
  INV_X1 U13090 ( .A(n19197), .ZN(n19195) );
  NAND3_X1 U13091 ( .A1(n22415), .A2(n19097), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18979) );
  NAND2_X1 U13092 ( .A1(n21673), .A2(n19082), .ZN(n19057) );
  INV_X1 U13093 ( .A(n21853), .ZN(n21805) );
  OR2_X1 U13094 ( .A1(n22027), .A2(n22043), .ZN(n21950) );
  INV_X1 U13095 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22079) );
  INV_X1 U13096 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n22113) );
  INV_X1 U13097 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n22100) );
  INV_X1 U13098 ( .A(n19239), .ZN(n22421) );
  NOR2_X2 U13099 ( .A1(n11330), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11541) );
  AOI22_X1 U13100 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11516) );
  AND2_X2 U13101 ( .A1(n11330), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11543) );
  AND2_X4 U13102 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11543), .ZN(
        n11715) );
  AND2_X2 U13103 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U13104 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11515) );
  AND2_X4 U13105 ( .A1(n11544), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12968) );
  AOI22_X1 U13106 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U13107 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U13108 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U13109 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U13110 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U13111 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U13112 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U13113 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U13114 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11218), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U13115 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U13116 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11535) );
  AOI22_X1 U13117 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U13118 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U13119 ( .A1(n11205), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U13120 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  AND2_X2 U13121 ( .A1(n11216), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12726) );
  AOI22_X1 U13122 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11540) );
  AND2_X1 U13123 ( .A1(n11715), .A2(n11713), .ZN(n11870) );
  INV_X2 U13124 ( .A(n12944), .ZN(n12795) );
  AND2_X2 U13125 ( .A1(n12795), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12730) );
  AOI22_X1 U13126 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11539) );
  AND2_X2 U13127 ( .A1(n12938), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11872) );
  AOI22_X1 U13128 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11872), .B1(
        n11871), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11538) );
  AND2_X2 U13129 ( .A1(n12937), .A2(n11713), .ZN(n11873) );
  AOI22_X1 U13130 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11537) );
  NAND4_X1 U13131 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11550) );
  AOI22_X1 U13132 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U13133 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11211), .B1(
        n11878), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11547) );
  AND2_X1 U13134 ( .A1(n11541), .A2(n12797), .ZN(n11589) );
  AOI22_X1 U13135 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U13136 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U13137 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11549) );
  XNOR2_X1 U13138 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12327) );
  INV_X1 U13139 ( .A(n12125), .ZN(n11551) );
  NAND2_X1 U13140 ( .A1(n12327), .A2(n11551), .ZN(n11553) );
  NAND2_X1 U13141 ( .A1(n20150), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11552) );
  NAND2_X1 U13142 ( .A1(n11553), .A2(n11552), .ZN(n11581) );
  XNOR2_X1 U13143 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11580) );
  XNOR2_X1 U13144 ( .A(n11581), .B(n11580), .ZN(n12332) );
  INV_X1 U13145 ( .A(n12332), .ZN(n12324) );
  AOI22_X1 U13146 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U13147 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U13148 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11218), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U13149 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11554) );
  NAND4_X1 U13150 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11558) );
  NAND2_X1 U13151 ( .A1(n11558), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11565) );
  AOI22_X1 U13152 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U13153 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U13154 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11559) );
  NAND4_X1 U13155 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11563) );
  NAND2_X1 U13156 ( .A1(n11563), .A2(n11713), .ZN(n11564) );
  NAND2_X2 U13157 ( .A1(n11565), .A2(n11564), .ZN(n11743) );
  AOI22_X1 U13158 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U13159 ( .A1(n11206), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U13160 ( .A1(n11607), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U13161 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11878), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U13162 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11577) );
  AOI22_X1 U13163 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13164 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11574) );
  INV_X2 U13165 ( .A(n12733), .ZN(n12783) );
  AOI22_X1 U13166 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12783), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U13167 ( .A1(n11871), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U13168 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  NOR2_X1 U13169 ( .A1(n11577), .A2(n11576), .ZN(n12390) );
  INV_X1 U13170 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11578) );
  INV_X1 U13171 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14836) );
  NAND2_X1 U13172 ( .A1(n11578), .A2(n14836), .ZN(n11579) );
  MUX2_X1 U13173 ( .A(n12390), .B(n11579), .S(n20269), .Z(n11975) );
  NOR2_X2 U13174 ( .A1(n11974), .A2(n11975), .ZN(n11967) );
  NAND2_X1 U13175 ( .A1(n11581), .A2(n11580), .ZN(n11583) );
  NAND2_X1 U13176 ( .A1(n20146), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U13177 ( .A1(n11583), .A2(n11582), .ZN(n11600) );
  XNOR2_X1 U13178 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11599) );
  INV_X1 U13179 ( .A(n11599), .ZN(n11584) );
  XNOR2_X1 U13180 ( .A(n11600), .B(n11584), .ZN(n12119) );
  AOI22_X1 U13181 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n11206), .B1(
        n11871), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U13182 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U13183 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13184 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U13185 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11598) );
  AOI22_X1 U13186 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U13187 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11211), .B1(
        n11878), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13188 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U13189 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11593) );
  NAND4_X1 U13190 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11597) );
  MUX2_X1 U13191 ( .A(n12119), .B(n11909), .S(n11738), .Z(n12137) );
  INV_X1 U13192 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11810) );
  MUX2_X1 U13193 ( .A(n12137), .B(n11810), .S(n20269), .Z(n11968) );
  NAND2_X1 U13194 ( .A1(n11600), .A2(n11599), .ZN(n11602) );
  NAND2_X1 U13195 ( .A1(n20145), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U13196 ( .A1(n11602), .A2(n11601), .ZN(n12122) );
  AOI22_X1 U13197 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13198 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U13199 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11872), .B1(
        n11871), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U13200 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U13201 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11613) );
  AOI22_X1 U13202 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U13203 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11211), .B1(
        n11878), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U13204 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U13205 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11608) );
  NAND4_X1 U13206 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11612) );
  MUX2_X1 U13207 ( .A(n12120), .B(n12416), .S(n11738), .Z(n12136) );
  INV_X1 U13208 ( .A(n12136), .ZN(n11614) );
  MUX2_X1 U13209 ( .A(n11614), .B(P2_EBX_REG_4__SCAN_IN), .S(n20269), .Z(
        n11980) );
  INV_X1 U13210 ( .A(n11980), .ZN(n11615) );
  AOI22_X1 U13211 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U13212 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U13213 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n11872), .B1(
        n11871), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U13214 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11616) );
  NAND4_X1 U13215 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11627) );
  AOI22_X1 U13216 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11625) );
  INV_X1 U13217 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U13218 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U13219 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U13220 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11622) );
  NAND4_X1 U13221 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11626) );
  INV_X1 U13222 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14918) );
  MUX2_X1 U13223 ( .A(n11911), .B(n14918), .S(n20269), .Z(n11983) );
  AOI22_X1 U13224 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U13225 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U13226 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11872), .B1(
        n11871), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U13227 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11567), .B1(
        n11878), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U13228 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11638) );
  AOI22_X1 U13229 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U13230 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11210), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U13231 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U13232 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11633) );
  NAND4_X1 U13233 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11637) );
  NOR2_X1 U13234 ( .A1(n11638), .A2(n11637), .ZN(n11942) );
  INV_X1 U13235 ( .A(n11942), .ZN(n12423) );
  INV_X1 U13236 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12209) );
  MUX2_X1 U13237 ( .A(n12423), .B(n12209), .S(n20269), .Z(n11946) );
  NAND2_X1 U13238 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11642) );
  NAND2_X1 U13239 ( .A1(n11206), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U13240 ( .A1(n11871), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U13241 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11639) );
  AOI22_X1 U13242 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U13243 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11645) );
  NAND2_X1 U13244 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U13245 ( .A1(n11607), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U13246 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U13247 ( .A1(n12730), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11649) );
  NAND2_X1 U13248 ( .A1(n11878), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U13249 ( .A1(n11873), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11647) );
  AOI22_X1 U13250 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11210), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11651) );
  NAND2_X1 U13251 ( .A1(n12113), .A2(n12377), .ZN(n11654) );
  OAI21_X1 U13252 ( .B1(n12377), .B2(P2_EBX_REG_7__SCAN_IN), .A(n11654), .ZN(
        n11955) );
  INV_X1 U13253 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n19298) );
  NOR2_X1 U13254 ( .A1(n12377), .A2(n19298), .ZN(n11952) );
  NAND2_X1 U13255 ( .A1(n20269), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U13256 ( .A1(n20269), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11959) );
  INV_X1 U13257 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12227) );
  NOR2_X1 U13258 ( .A1(n12377), .A2(n12227), .ZN(n11998) );
  NAND2_X1 U13259 ( .A1(n20269), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12006) );
  NAND2_X1 U13260 ( .A1(n20269), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12023) );
  NOR2_X2 U13261 ( .A1(n12024), .A2(n11656), .ZN(n12019) );
  NAND2_X1 U13262 ( .A1(n20269), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12020) );
  AND2_X2 U13263 ( .A1(n12019), .A2(n12020), .ZN(n12016) );
  NAND2_X1 U13264 ( .A1(n20269), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12017) );
  INV_X1 U13265 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12251) );
  NOR2_X1 U13266 ( .A1(n12377), .A2(n12251), .ZN(n12029) );
  INV_X1 U13267 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12247) );
  NOR2_X1 U13268 ( .A1(n12377), .A2(n12247), .ZN(n12013) );
  NAND2_X1 U13269 ( .A1(n20269), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12040) );
  NAND2_X1 U13270 ( .A1(n20269), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12034) );
  INV_X1 U13271 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12263) );
  NOR2_X1 U13272 ( .A1(n12377), .A2(n12263), .ZN(n12011) );
  OR2_X2 U13273 ( .A1(n12038), .A2(n12011), .ZN(n12066) );
  INV_X1 U13274 ( .A(n12066), .ZN(n11657) );
  NAND2_X1 U13275 ( .A1(n20269), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U13276 ( .A1(n11657), .A2(n12044), .ZN(n11659) );
  NAND2_X1 U13277 ( .A1(n20269), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11658) );
  XNOR2_X1 U13278 ( .A(n11659), .B(n11658), .ZN(n19414) );
  NAND2_X1 U13279 ( .A1(n19414), .A2(n12114), .ZN(n12062) );
  INV_X1 U13280 ( .A(n12062), .ZN(n12063) );
  AOI22_X1 U13281 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11218), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U13282 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U13283 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U13284 ( .A1(n11205), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U13285 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11664) );
  NAND2_X1 U13286 ( .A1(n11664), .A2(n11713), .ZN(n11671) );
  AOI22_X1 U13287 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U13288 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U13289 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U13290 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11669) );
  NAND2_X1 U13291 ( .A1(n11669), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11670) );
  NAND2_X2 U13292 ( .A1(n11671), .A2(n11670), .ZN(n11729) );
  INV_X2 U13293 ( .A(n11729), .ZN(n11732) );
  AOI22_X1 U13294 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U13295 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U13296 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11672) );
  NAND4_X1 U13297 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(
        n11681) );
  AOI22_X1 U13298 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U13299 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U13300 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U13301 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U13302 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11680) );
  NAND2_X1 U13303 ( .A1(n11746), .A2(n12584), .ZN(n11734) );
  AOI22_X1 U13304 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11715), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U13305 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U13306 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11218), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U13307 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11683) );
  NAND4_X1 U13308 ( .A1(n11686), .A2(n11685), .A3(n11684), .A4(n11683), .ZN(
        n11687) );
  NAND2_X1 U13309 ( .A1(n11687), .A2(n11713), .ZN(n11694) );
  AOI22_X1 U13310 ( .A1(n11201), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U13311 ( .A1(n11205), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11715), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U13312 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U13313 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11688) );
  NAND4_X1 U13314 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11692) );
  NAND2_X1 U13315 ( .A1(n11692), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11693) );
  AOI22_X1 U13316 ( .A1(n11205), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U13317 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U13318 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U13319 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U13320 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  NAND2_X1 U13321 ( .A1(n11699), .A2(n11713), .ZN(n11706) );
  AOI22_X1 U13322 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U13323 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U13324 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U13325 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11700) );
  NAND4_X1 U13326 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11704) );
  NAND2_X1 U13327 ( .A1(n11704), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U13328 ( .A1(n13007), .A2(n11744), .ZN(n11731) );
  NAND2_X1 U13329 ( .A1(n11725), .A2(n11729), .ZN(n11707) );
  NAND2_X1 U13330 ( .A1(n11734), .A2(n11708), .ZN(n11750) );
  INV_X2 U13331 ( .A(n11744), .ZN(n11725) );
  AOI22_X1 U13332 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U13333 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U13334 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U13335 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12796), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U13336 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11714) );
  AOI22_X1 U13337 ( .A1(n11216), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11201), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U13338 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12968), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U13339 ( .A1(n11715), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U13340 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11716) );
  NAND4_X1 U13341 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11720) );
  NAND2_X1 U13342 ( .A1(n11720), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11721) );
  NAND2_X2 U13343 ( .A1(n11722), .A2(n11721), .ZN(n12345) );
  NAND3_X1 U13344 ( .A1(n11725), .A2(n13007), .A3(n11723), .ZN(n11724) );
  AND3_X2 U13345 ( .A1(n11725), .A2(n11727), .A3(n12584), .ZN(n11755) );
  NAND2_X1 U13346 ( .A1(n11756), .A2(n19249), .ZN(n14565) );
  NAND2_X1 U13347 ( .A1(n11761), .A2(n12132), .ZN(n11735) );
  NAND2_X1 U13348 ( .A1(n12575), .A2(n19490), .ZN(n12577) );
  NAND2_X1 U13349 ( .A1(n13007), .A2(n11729), .ZN(n11753) );
  INV_X1 U13350 ( .A(n11753), .ZN(n12988) );
  NAND2_X1 U13351 ( .A1(n12988), .A2(n11752), .ZN(n11730) );
  INV_X1 U13352 ( .A(n11747), .ZN(n12572) );
  NOR2_X4 U13353 ( .A1(n15276), .A2(n19251), .ZN(n11777) );
  NAND2_X2 U13354 ( .A1(n11738), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11771) );
  INV_X1 U13355 ( .A(n11771), .ZN(n11739) );
  NAND2_X1 U13356 ( .A1(n11807), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11741) );
  NAND2_X1 U13357 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11740) );
  INV_X1 U13358 ( .A(n11768), .ZN(n11766) );
  NAND2_X1 U13359 ( .A1(n11745), .A2(n13007), .ZN(n12582) );
  INV_X1 U13360 ( .A(n11785), .ZN(n11760) );
  NAND2_X1 U13361 ( .A1(n12574), .A2(n11747), .ZN(n11786) );
  NAND2_X1 U13362 ( .A1(n11786), .A2(n20528), .ZN(n11751) );
  NAND2_X1 U13363 ( .A1(n12377), .A2(n11729), .ZN(n11748) );
  NAND2_X1 U13364 ( .A1(n11748), .A2(n11727), .ZN(n11749) );
  OAI211_X1 U13365 ( .C1(n11750), .C2(n11749), .A(n15349), .B(n20528), .ZN(
        n12588) );
  NAND2_X1 U13366 ( .A1(n11751), .A2(n12588), .ZN(n11784) );
  NOR2_X1 U13367 ( .A1(n11753), .A2(n11752), .ZN(n11754) );
  NAND2_X1 U13368 ( .A1(n11755), .A2(n11754), .ZN(n12323) );
  NAND3_X1 U13369 ( .A1(n12323), .A2(n11727), .A3(n12954), .ZN(n11758) );
  INV_X1 U13370 ( .A(n11756), .ZN(n11757) );
  NAND2_X1 U13371 ( .A1(n11758), .A2(n11757), .ZN(n12566) );
  NAND2_X1 U13372 ( .A1(n11806), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11764) );
  NOR2_X1 U13373 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12317) );
  AND2_X2 U13374 ( .A1(n11764), .A2(n11763), .ZN(n11767) );
  INV_X1 U13375 ( .A(n11767), .ZN(n11765) );
  NAND2_X1 U13376 ( .A1(n11766), .A2(n11765), .ZN(n11769) );
  AND2_X2 U13377 ( .A1(n11769), .A2(n11817), .ZN(n11820) );
  NOR2_X1 U13378 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  OAI22_X1 U13379 ( .A1(n11197), .A2(n11772), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11777), .ZN(n11776) );
  INV_X1 U13380 ( .A(n11773), .ZN(n11774) );
  AOI22_X1 U13381 ( .A1(n11774), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12317), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U13382 ( .A1(n11776), .A2(n11775), .ZN(n11822) );
  NAND2_X1 U13383 ( .A1(n11777), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11782) );
  INV_X1 U13384 ( .A(n12317), .ZN(n19510) );
  NAND2_X1 U13385 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11778) );
  AND2_X1 U13386 ( .A1(n19510), .A2(n11778), .ZN(n11781) );
  INV_X1 U13387 ( .A(n11779), .ZN(n11780) );
  NAND3_X1 U13388 ( .A1(n11782), .A2(n11781), .A3(n11780), .ZN(n11783) );
  NOR2_X1 U13389 ( .A1(n11502), .A2(n11783), .ZN(n11789) );
  AOI21_X1 U13390 ( .B1(n11786), .B2(n11785), .A(n11784), .ZN(n11787) );
  NAND2_X2 U13391 ( .A1(n11822), .A2(n11821), .ZN(n11831) );
  OAI21_X1 U13392 ( .B1(n20146), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n18105), 
        .ZN(n11791) );
  AOI21_X1 U13393 ( .B1(n11197), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11791), .ZN(n11797) );
  INV_X1 U13394 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14894) );
  NAND2_X1 U13395 ( .A1(n11807), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U13396 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11792) );
  NAND2_X1 U13397 ( .A1(n11797), .A2(n11798), .ZN(n11802) );
  AND2_X1 U13398 ( .A1(n11178), .A2(n11802), .ZN(n11796) );
  INV_X1 U13399 ( .A(n11797), .ZN(n11800) );
  INV_X1 U13400 ( .A(n11798), .ZN(n11799) );
  NAND2_X1 U13401 ( .A1(n11800), .A2(n11799), .ZN(n11801) );
  NOR2_X1 U13402 ( .A1(n19510), .A2(n20145), .ZN(n11805) );
  AOI21_X1 U13403 ( .B1(n11197), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11805), .ZN(n11812) );
  INV_X4 U13404 ( .A(n11777), .ZN(n12309) );
  NAND2_X1 U13405 ( .A1(n12306), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11809) );
  NAND2_X1 U13406 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11808) );
  OAI211_X1 U13407 ( .C1(n12309), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        n11811) );
  NAND2_X1 U13408 ( .A1(n11812), .A2(n11813), .ZN(n12200) );
  INV_X1 U13409 ( .A(n11812), .ZN(n11815) );
  INV_X1 U13410 ( .A(n11813), .ZN(n11814) );
  NAND2_X1 U13411 ( .A1(n11815), .A2(n11814), .ZN(n11816) );
  XNOR2_X2 U13412 ( .A(n11819), .B(n11818), .ZN(n12677) );
  INV_X1 U13413 ( .A(n11820), .ZN(n11832) );
  NAND2_X1 U13414 ( .A1(n11832), .A2(n19505), .ZN(n11851) );
  INV_X1 U13415 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11830) );
  INV_X1 U13416 ( .A(n11826), .ZN(n11827) );
  NAND2_X1 U13417 ( .A1(n15716), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11829) );
  OAI211_X1 U13418 ( .C1(n11912), .C2(n11830), .A(n11829), .B(n12954), .ZN(
        n11838) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11836) );
  INV_X1 U13420 ( .A(n11831), .ZN(n11833) );
  NAND2_X1 U13421 ( .A1(n11833), .A2(n11832), .ZN(n11834) );
  NAND2_X1 U13422 ( .A1(n17360), .A2(n15304), .ZN(n11842) );
  INV_X1 U13423 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11835) );
  OAI22_X1 U13424 ( .A1(n11836), .A2(n11931), .B1(n11919), .B2(n11835), .ZN(
        n11837) );
  NOR2_X1 U13425 ( .A1(n11838), .A2(n11837), .ZN(n11869) );
  INV_X1 U13426 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U13427 ( .A1(n15274), .A2(n16440), .ZN(n11859) );
  NAND2_X2 U13428 ( .A1(n11861), .A2(n11839), .ZN(n11915) );
  INV_X1 U13429 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11840) );
  OAI22_X1 U13430 ( .A1(n11841), .A2(n20117), .B1(n11915), .B2(n11840), .ZN(
        n11845) );
  INV_X1 U13431 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12830) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11843) );
  NOR2_X1 U13433 ( .A1(n11845), .A2(n11844), .ZN(n11868) );
  INV_X1 U13434 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11850) );
  INV_X1 U13435 ( .A(n11858), .ZN(n11847) );
  INV_X1 U13436 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11849) );
  INV_X1 U13437 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11853) );
  INV_X1 U13438 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11852) );
  NOR2_X1 U13439 ( .A1(n11855), .A2(n11854), .ZN(n11867) );
  INV_X1 U13440 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12823) );
  INV_X1 U13441 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20498) );
  OAI22_X1 U13442 ( .A1(n12823), .A2(n20194), .B1(n11926), .B2(n20498), .ZN(
        n11865) );
  INV_X1 U13443 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11863) );
  INV_X1 U13444 ( .A(n11859), .ZN(n11861) );
  INV_X1 U13445 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11862) );
  OAI22_X1 U13446 ( .A1(n11863), .A2(n11918), .B1(n20065), .B2(n11862), .ZN(
        n11864) );
  NOR2_X1 U13447 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  AOI22_X1 U13448 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12726), .B1(
        n12129), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U13449 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U13450 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11872), .B1(
        n11220), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U13451 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11874) );
  NAND4_X1 U13452 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11884) );
  AOI22_X1 U13453 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11882) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14745) );
  AOI22_X1 U13455 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11878), .B1(
        n11211), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U13456 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U13457 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U13458 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11883) );
  NAND2_X1 U13459 ( .A1(n12819), .A2(n12375), .ZN(n14630) );
  OR2_X1 U13460 ( .A1(n12390), .A2(n14630), .ZN(n12147) );
  INV_X1 U13461 ( .A(n12149), .ZN(n12398) );
  NAND2_X1 U13462 ( .A1(n12147), .A2(n12398), .ZN(n11885) );
  INV_X1 U13463 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12873) );
  INV_X1 U13464 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11886) );
  OAI22_X1 U13465 ( .A1(n12873), .A2(n11927), .B1(n11236), .B2(n11886), .ZN(
        n11890) );
  INV_X1 U13466 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11888) );
  INV_X1 U13467 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11887) );
  OAI22_X1 U13468 ( .A1(n11888), .A2(n20065), .B1(n11915), .B2(n11887), .ZN(
        n11889) );
  NOR2_X1 U13469 ( .A1(n11890), .A2(n11889), .ZN(n11908) );
  INV_X1 U13470 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11891) );
  INV_X1 U13471 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12729) );
  INV_X1 U13472 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11892) );
  NOR2_X1 U13473 ( .A1(n11894), .A2(n11893), .ZN(n11907) );
  INV_X1 U13474 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11895) );
  INV_X1 U13475 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12731) );
  OAI22_X1 U13476 ( .A1(n11895), .A2(n20060), .B1(n20040), .B2(n12731), .ZN(
        n11898) );
  INV_X1 U13477 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12866) );
  INV_X1 U13478 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11896) );
  NOR2_X1 U13479 ( .A1(n11898), .A2(n11897), .ZN(n11906) );
  INV_X1 U13480 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11900) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11899) );
  INV_X1 U13482 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11902) );
  INV_X1 U13483 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11901) );
  OAI22_X1 U13484 ( .A1(n11902), .A2(n11926), .B1(n11912), .B2(n11901), .ZN(
        n11903) );
  INV_X1 U13485 ( .A(n11909), .ZN(n12410) );
  NAND2_X1 U13486 ( .A1(n12410), .A2(n12819), .ZN(n11910) );
  INV_X1 U13487 ( .A(n11966), .ZN(n12143) );
  INV_X1 U13488 ( .A(n11911), .ZN(n12419) );
  INV_X1 U13489 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11914) );
  INV_X1 U13490 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11913) );
  OAI22_X1 U13491 ( .A1(n11914), .A2(n11912), .B1(n11236), .B2(n11913), .ZN(
        n11917) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12932) );
  INV_X1 U13493 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12933) );
  OAI22_X1 U13494 ( .A1(n12932), .A2(n11915), .B1(n20040), .B2(n12933), .ZN(
        n11916) );
  NOR2_X1 U13495 ( .A1(n11917), .A2(n11916), .ZN(n11941) );
  INV_X1 U13496 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12945) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11920) );
  OAI22_X1 U13498 ( .A1(n12945), .A2(n11918), .B1(n11919), .B2(n11920), .ZN(
        n11923) );
  INV_X1 U13499 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12942) );
  INV_X1 U13500 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11921) );
  OAI22_X1 U13501 ( .A1(n12942), .A2(n20194), .B1(n20060), .B2(n11921), .ZN(
        n11922) );
  NOR2_X1 U13502 ( .A1(n11923), .A2(n11922), .ZN(n11940) );
  INV_X1 U13503 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11925) );
  INV_X1 U13504 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12943) );
  OAI22_X1 U13505 ( .A1(n11925), .A2(n11924), .B1(n20117), .B2(n12943), .ZN(
        n11930) );
  INV_X1 U13506 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11928) );
  INV_X1 U13507 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12931) );
  OAI22_X1 U13508 ( .A1(n11928), .A2(n11926), .B1(n11927), .B2(n12931), .ZN(
        n11929) );
  NOR2_X1 U13509 ( .A1(n11930), .A2(n11929), .ZN(n11939) );
  INV_X1 U13510 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11933) );
  INV_X1 U13511 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11932) );
  OAI22_X1 U13512 ( .A1(n11933), .A2(n11931), .B1(n20065), .B2(n11932), .ZN(
        n11937) );
  INV_X1 U13513 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11935) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11934) );
  OAI22_X1 U13515 ( .A1(n11935), .A2(n15509), .B1(n15713), .B2(n11934), .ZN(
        n11936) );
  NOR2_X1 U13516 ( .A1(n11937), .A2(n11936), .ZN(n11938) );
  NAND4_X1 U13517 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11944) );
  NAND2_X1 U13518 ( .A1(n11942), .A2(n12819), .ZN(n11943) );
  NAND2_X1 U13519 ( .A1(n12168), .A2(n11961), .ZN(n11950) );
  INV_X1 U13520 ( .A(n11945), .ZN(n11948) );
  INV_X1 U13521 ( .A(n11946), .ZN(n11947) );
  NAND2_X1 U13522 ( .A1(n11948), .A2(n11947), .ZN(n11949) );
  NAND2_X1 U13523 ( .A1(n12115), .A2(n11949), .ZN(n19287) );
  INV_X1 U13524 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18068) );
  INV_X1 U13525 ( .A(n11951), .ZN(n11963) );
  NAND2_X1 U13526 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  NAND2_X1 U13527 ( .A1(n11963), .A2(n11954), .ZN(n19299) );
  NOR2_X1 U13528 ( .A1(n19299), .A2(n11961), .ZN(n11957) );
  NAND2_X1 U13529 ( .A1(n11957), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18020) );
  INV_X1 U13530 ( .A(n18020), .ZN(n11992) );
  XNOR2_X1 U13531 ( .A(n12115), .B(n11955), .ZN(n15207) );
  INV_X1 U13532 ( .A(n15207), .ZN(n11956) );
  INV_X1 U13533 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18046) );
  NAND2_X1 U13534 ( .A1(n11956), .A2(n18046), .ZN(n18017) );
  INV_X1 U13535 ( .A(n11957), .ZN(n11958) );
  INV_X1 U13536 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18037) );
  NAND2_X1 U13537 ( .A1(n11958), .A2(n18037), .ZN(n18019) );
  AND2_X1 U13538 ( .A1(n18017), .A2(n18019), .ZN(n17721) );
  OR2_X1 U13539 ( .A1(n11992), .A2(n17721), .ZN(n17707) );
  XNOR2_X1 U13540 ( .A(n11960), .B(n11959), .ZN(n19311) );
  AOI21_X1 U13541 ( .B1(n19311), .B2(n12114), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17983) );
  XNOR2_X1 U13542 ( .A(n11963), .B(n11962), .ZN(n15261) );
  AOI21_X1 U13543 ( .B1(n15261), .B2(n12113), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17724) );
  OR2_X1 U13544 ( .A1(n17983), .A2(n17724), .ZN(n17709) );
  INV_X1 U13545 ( .A(n17709), .ZN(n11964) );
  AND2_X1 U13546 ( .A1(n17707), .A2(n11964), .ZN(n11991) );
  AND2_X1 U13547 ( .A1(n17703), .A2(n11991), .ZN(n11990) );
  INV_X1 U13548 ( .A(n11967), .ZN(n11970) );
  INV_X1 U13549 ( .A(n11968), .ZN(n11969) );
  NAND2_X1 U13550 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  NAND2_X1 U13551 ( .A1(n11981), .A2(n11971), .ZN(n16450) );
  INV_X1 U13552 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16274) );
  XNOR2_X1 U13553 ( .A(n11979), .B(n16274), .ZN(n15554) );
  OAI21_X1 U13554 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20122), .A(
        n12125), .ZN(n12328) );
  INV_X1 U13555 ( .A(n12328), .ZN(n12326) );
  MUX2_X1 U13556 ( .A(n12326), .B(n12375), .S(n11738), .Z(n12133) );
  MUX2_X1 U13557 ( .A(n12133), .B(P2_EBX_REG_0__SCAN_IN), .S(n20269), .Z(
        n19260) );
  NAND2_X1 U13558 ( .A1(n19260), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14628) );
  NAND3_X1 U13559 ( .A1(n20269), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11972) );
  NAND2_X1 U13560 ( .A1(n11975), .A2(n11972), .ZN(n17358) );
  AND2_X1 U13561 ( .A1(n14628), .A2(n17358), .ZN(n14691) );
  NOR2_X1 U13562 ( .A1(n14628), .A2(n17358), .ZN(n14692) );
  NOR2_X1 U13563 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14692), .ZN(
        n11973) );
  NOR2_X1 U13564 ( .A1(n14691), .A2(n11973), .ZN(n16413) );
  XNOR2_X1 U13565 ( .A(n11975), .B(n11974), .ZN(n15490) );
  XNOR2_X1 U13566 ( .A(n15490), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16412) );
  NAND2_X1 U13567 ( .A1(n16413), .A2(n16412), .ZN(n11978) );
  INV_X1 U13568 ( .A(n15490), .ZN(n11976) );
  NAND2_X1 U13569 ( .A1(n11976), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11977) );
  NAND2_X1 U13570 ( .A1(n11978), .A2(n11977), .ZN(n15553) );
  NAND2_X1 U13571 ( .A1(n11979), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16268) );
  XNOR2_X1 U13572 ( .A(n11981), .B(n11980), .ZN(n11986) );
  INV_X1 U13573 ( .A(n11986), .ZN(n19272) );
  NAND2_X1 U13574 ( .A1(n19272), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11985) );
  AND2_X1 U13575 ( .A1(n16268), .A2(n11985), .ZN(n11982) );
  XNOR2_X1 U13576 ( .A(n11984), .B(n11983), .ZN(n15183) );
  INV_X1 U13577 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16324) );
  XNOR2_X1 U13578 ( .A(n15183), .B(n16324), .ZN(n16316) );
  INV_X1 U13579 ( .A(n11985), .ZN(n11987) );
  XNOR2_X1 U13580 ( .A(n11986), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16271) );
  OR2_X1 U13581 ( .A1(n11987), .A2(n16271), .ZN(n16314) );
  AND2_X1 U13582 ( .A1(n16316), .A2(n16314), .ZN(n11988) );
  NAND2_X1 U13583 ( .A1(n15183), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11989) );
  INV_X1 U13584 ( .A(n11991), .ZN(n11996) );
  AND2_X1 U13585 ( .A1(n15207), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17734) );
  OR2_X1 U13586 ( .A1(n17734), .A2(n11992), .ZN(n17706) );
  NAND2_X1 U13587 ( .A1(n11993), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17704) );
  INV_X1 U13588 ( .A(n17704), .ZN(n11994) );
  NOR2_X1 U13589 ( .A1(n17706), .A2(n11994), .ZN(n11995) );
  NAND2_X1 U13590 ( .A1(n11999), .A2(n11998), .ZN(n12000) );
  NAND2_X1 U13591 ( .A1(n12008), .A2(n12000), .ZN(n17352) );
  NOR2_X1 U13592 ( .A1(n17352), .A2(n11961), .ZN(n12002) );
  INV_X1 U13593 ( .A(n12002), .ZN(n12001) );
  INV_X1 U13594 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17965) );
  NAND2_X1 U13595 ( .A1(n12001), .A2(n17965), .ZN(n17712) );
  NAND2_X1 U13596 ( .A1(n12002), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17713) );
  INV_X1 U13597 ( .A(n19311), .ZN(n12003) );
  INV_X1 U13598 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17979) );
  OR3_X1 U13599 ( .A1(n12003), .A2(n11961), .A3(n17979), .ZN(n17982) );
  AND2_X1 U13600 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U13601 ( .A1(n15261), .A2(n12004), .ZN(n17980) );
  AND2_X1 U13602 ( .A1(n17982), .A2(n17980), .ZN(n17711) );
  NAND2_X1 U13603 ( .A1(n17713), .A2(n17711), .ZN(n12005) );
  INV_X1 U13604 ( .A(n12006), .ZN(n12007) );
  NAND2_X1 U13605 ( .A1(n12008), .A2(n12007), .ZN(n12009) );
  NAND2_X1 U13606 ( .A1(n12024), .A2(n12009), .ZN(n19323) );
  NAND2_X1 U13607 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12010) );
  OR2_X1 U13608 ( .A1(n19323), .A2(n12010), .ZN(n17694) );
  NAND2_X1 U13609 ( .A1(n12038), .A2(n12011), .ZN(n12012) );
  AND2_X1 U13610 ( .A1(n12066), .A2(n12012), .ZN(n19386) );
  NAND2_X1 U13611 ( .A1(n19386), .A2(n12114), .ZN(n17616) );
  INV_X1 U13612 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17845) );
  INV_X1 U13613 ( .A(n12013), .ZN(n12014) );
  XNOR2_X1 U13614 ( .A(n11248), .B(n12014), .ZN(n19356) );
  NAND2_X1 U13615 ( .A1(n19356), .A2(n12114), .ZN(n12015) );
  INV_X1 U13616 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12653) );
  NAND2_X1 U13617 ( .A1(n12015), .A2(n12653), .ZN(n17651) );
  INV_X1 U13618 ( .A(n12016), .ZN(n12018) );
  XNOR2_X1 U13619 ( .A(n12018), .B(n12017), .ZN(n14532) );
  NAND2_X1 U13620 ( .A1(n14532), .A2(n12114), .ZN(n12050) );
  INV_X1 U13621 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17908) );
  NAND2_X1 U13622 ( .A1(n12050), .A2(n17908), .ZN(n17669) );
  INV_X1 U13623 ( .A(n12019), .ZN(n12021) );
  XNOR2_X1 U13624 ( .A(n12021), .B(n12020), .ZN(n19331) );
  NAND2_X1 U13625 ( .A1(n19331), .A2(n12114), .ZN(n12022) );
  INV_X1 U13626 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17928) );
  NAND2_X1 U13627 ( .A1(n12022), .A2(n17928), .ZN(n17917) );
  XNOR2_X1 U13628 ( .A(n12024), .B(n12023), .ZN(n17339) );
  NAND2_X1 U13629 ( .A1(n17339), .A2(n12114), .ZN(n12025) );
  INV_X1 U13630 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17680) );
  NAND2_X1 U13631 ( .A1(n12025), .A2(n17680), .ZN(n17682) );
  AND2_X1 U13632 ( .A1(n17917), .A2(n17682), .ZN(n12026) );
  OR2_X1 U13633 ( .A1(n19323), .A2(n11961), .ZN(n12027) );
  INV_X1 U13634 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17691) );
  NAND2_X1 U13635 ( .A1(n12027), .A2(n17691), .ZN(n17696) );
  NAND3_X1 U13636 ( .A1(n17651), .A2(n12644), .A3(n17696), .ZN(n12028) );
  AOI21_X1 U13637 ( .B1(n17616), .B2(n17845), .A(n12028), .ZN(n12043) );
  INV_X1 U13638 ( .A(n12029), .ZN(n12030) );
  XNOR2_X1 U13639 ( .A(n12031), .B(n12030), .ZN(n19343) );
  NAND2_X1 U13640 ( .A1(n19343), .A2(n12114), .ZN(n12032) );
  XNOR2_X1 U13641 ( .A(n12032), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17662) );
  INV_X1 U13642 ( .A(n12033), .ZN(n12036) );
  INV_X1 U13643 ( .A(n12034), .ZN(n12035) );
  NAND2_X1 U13644 ( .A1(n12036), .A2(n12035), .ZN(n12037) );
  NAND2_X1 U13645 ( .A1(n12038), .A2(n12037), .ZN(n17310) );
  INV_X1 U13646 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17853) );
  NAND2_X1 U13647 ( .A1(n12046), .A2(n17853), .ZN(n17629) );
  INV_X1 U13648 ( .A(n12039), .ZN(n12041) );
  XNOR2_X1 U13649 ( .A(n12041), .B(n12040), .ZN(n19379) );
  NAND2_X1 U13650 ( .A1(n19379), .A2(n12114), .ZN(n12042) );
  INV_X1 U13651 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17866) );
  NAND2_X1 U13652 ( .A1(n12042), .A2(n17866), .ZN(n17641) );
  AND2_X1 U13653 ( .A1(n17629), .A2(n17641), .ZN(n12650) );
  NAND3_X1 U13654 ( .A1(n12043), .A2(n17662), .A3(n12650), .ZN(n12045) );
  XNOR2_X1 U13655 ( .A(n12066), .B(n12044), .ZN(n19395) );
  NAND2_X1 U13656 ( .A1(n19395), .A2(n12114), .ZN(n17620) );
  INV_X1 U13657 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17623) );
  NOR2_X1 U13658 ( .A1(n12045), .A2(n11494), .ZN(n12061) );
  INV_X1 U13659 ( .A(n12046), .ZN(n12047) );
  NAND2_X1 U13660 ( .A1(n12047), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17630) );
  INV_X1 U13661 ( .A(n19379), .ZN(n12048) );
  AND2_X1 U13662 ( .A1(n17630), .A2(n17639), .ZN(n12652) );
  AND2_X1 U13663 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12049) );
  INV_X1 U13664 ( .A(n12050), .ZN(n12051) );
  NAND2_X1 U13665 ( .A1(n12051), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17670) );
  AND2_X1 U13666 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12052) );
  NAND2_X1 U13667 ( .A1(n19331), .A2(n12052), .ZN(n17916) );
  NAND2_X1 U13668 ( .A1(n17670), .A2(n17916), .ZN(n12645) );
  AND2_X1 U13669 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12053) );
  AND2_X1 U13670 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12054) );
  NOR4_X1 U13671 ( .A1(n17652), .A2(n12645), .A3(n12648), .A4(n12643), .ZN(
        n12055) );
  OAI211_X1 U13672 ( .C1(n17616), .C2(n17845), .A(n12652), .B(n12055), .ZN(
        n12056) );
  INV_X1 U13673 ( .A(n12056), .ZN(n12059) );
  INV_X1 U13674 ( .A(n17620), .ZN(n12057) );
  NAND2_X1 U13675 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  XNOR2_X1 U13676 ( .A(n12062), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17611) );
  OAI21_X1 U13677 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n12063), .A(
        n17610), .ZN(n17601) );
  NAND2_X1 U13678 ( .A1(n20269), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12067) );
  INV_X1 U13679 ( .A(n12067), .ZN(n12070) );
  NOR2_X1 U13680 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n12064) );
  NOR2_X1 U13681 ( .A1(n12377), .A2(n12064), .ZN(n12065) );
  NOR2_X2 U13682 ( .A1(n12066), .A2(n12065), .ZN(n12068) );
  INV_X1 U13683 ( .A(n12068), .ZN(n12069) );
  AOI21_X1 U13684 ( .B1(n12070), .B2(n12069), .A(n12075), .ZN(n17304) );
  NAND2_X1 U13685 ( .A1(n17304), .A2(n12114), .ZN(n12071) );
  XNOR2_X1 U13686 ( .A(n12071), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17600) );
  NAND2_X1 U13687 ( .A1(n17601), .A2(n17600), .ZN(n17599) );
  INV_X1 U13688 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12072) );
  NAND2_X1 U13689 ( .A1(n12071), .A2(n12072), .ZN(n12073) );
  INV_X1 U13690 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12276) );
  NOR2_X1 U13691 ( .A1(n12377), .A2(n12276), .ZN(n12077) );
  INV_X1 U13692 ( .A(n12075), .ZN(n12076) );
  INV_X1 U13693 ( .A(n12077), .ZN(n12074) );
  AOI21_X1 U13694 ( .B1(n12077), .B2(n12076), .A(n12081), .ZN(n17282) );
  NAND2_X1 U13695 ( .A1(n17282), .A2(n12114), .ZN(n12078) );
  XNOR2_X1 U13696 ( .A(n12078), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17590) );
  NAND2_X1 U13697 ( .A1(n20269), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U13698 ( .A1(n20269), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12087) );
  NAND2_X1 U13699 ( .A1(n12100), .A2(n12114), .ZN(n12080) );
  XOR2_X1 U13700 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n12080), .Z(
        n17568) );
  INV_X1 U13701 ( .A(n17568), .ZN(n12085) );
  INV_X1 U13702 ( .A(n12081), .ZN(n12083) );
  XNOR2_X1 U13703 ( .A(n12083), .B(n12082), .ZN(n19421) );
  AOI21_X1 U13704 ( .B1(n19421), .B2(n12114), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17581) );
  INV_X1 U13705 ( .A(n17581), .ZN(n12084) );
  NAND2_X1 U13706 ( .A1(n20269), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12095) );
  NAND2_X1 U13707 ( .A1(n20269), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12089) );
  INV_X1 U13708 ( .A(n12089), .ZN(n12090) );
  NAND2_X1 U13709 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NAND2_X1 U13710 ( .A1(n12109), .A2(n12092), .ZN(n19442) );
  INV_X1 U13711 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16407) );
  NOR3_X1 U13712 ( .A1(n19442), .A2(n11961), .A3(n16407), .ZN(n12098) );
  AOI21_X1 U13713 ( .B1(n12099), .B2(n12114), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12093) );
  INV_X1 U13714 ( .A(n12094), .ZN(n12096) );
  XNOR2_X1 U13715 ( .A(n12096), .B(n12095), .ZN(n17264) );
  NAND3_X1 U13716 ( .A1(n12099), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n12113), .ZN(n12104) );
  INV_X1 U13717 ( .A(n12100), .ZN(n12101) );
  INV_X1 U13718 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17768) );
  NOR3_X1 U13719 ( .A1(n12101), .A2(n11961), .A3(n17768), .ZN(n12103) );
  AND2_X1 U13720 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12102) );
  NOR2_X1 U13721 ( .A1(n12103), .A2(n17580), .ZN(n14196) );
  NAND2_X1 U13722 ( .A1(n12107), .A2(n12106), .ZN(n13023) );
  INV_X1 U13723 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12300) );
  NOR2_X1 U13724 ( .A1(n12377), .A2(n12300), .ZN(n12108) );
  XNOR2_X1 U13725 ( .A(n12109), .B(n12108), .ZN(n12112) );
  INV_X1 U13726 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14185) );
  OAI21_X1 U13727 ( .B1(n12112), .B2(n11961), .A(n14185), .ZN(n13022) );
  NAND2_X1 U13728 ( .A1(n13023), .A2(n13022), .ZN(n12626) );
  NAND2_X1 U13729 ( .A1(n20269), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12110) );
  XNOR2_X1 U13730 ( .A(n14464), .B(n12110), .ZN(n19474) );
  AOI21_X1 U13731 ( .B1(n19474), .B2(n12114), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12629) );
  AND2_X1 U13732 ( .A1(n12113), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U13733 ( .A1(n19474), .A2(n12111), .ZN(n12627) );
  INV_X1 U13734 ( .A(n12112), .ZN(n19456) );
  NAND3_X1 U13735 ( .A1(n19456), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12113), .ZN(n13021) );
  NAND2_X1 U13736 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  XNOR2_X1 U13737 ( .A(n12116), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12117) );
  XNOR2_X1 U13738 ( .A(n12118), .B(n12117), .ZN(n12622) );
  NAND2_X1 U13739 ( .A1(n12120), .A2(n12119), .ZN(n12338) );
  NOR2_X1 U13740 ( .A1(n12332), .A2(n12338), .ZN(n12126) );
  INV_X1 U13741 ( .A(n12126), .ZN(n12128) );
  AND2_X1 U13742 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18108), .ZN(
        n12121) );
  INV_X1 U13743 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19492) );
  NAND2_X1 U13744 ( .A1(n19492), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12123) );
  XNOR2_X1 U13745 ( .A(n12327), .B(n12125), .ZN(n12325) );
  AND2_X1 U13746 ( .A1(n12325), .A2(n12126), .ZN(n12127) );
  OAI21_X1 U13747 ( .B1(n12328), .B2(n12128), .A(n14564), .ZN(n12131) );
  INV_X1 U13748 ( .A(n11206), .ZN(n12727) );
  AOI21_X1 U13749 ( .B1(n12130), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19488) );
  AOI21_X1 U13750 ( .B1(n12727), .B2(n19488), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n18206) );
  MUX2_X1 U13751 ( .A(n12131), .B(n18206), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19523) );
  OR2_X1 U13752 ( .A1(n12323), .A2(n12132), .ZN(n12620) );
  NAND2_X1 U13753 ( .A1(n12133), .A2(n12327), .ZN(n12135) );
  NAND2_X1 U13754 ( .A1(n12135), .A2(n12134), .ZN(n12138) );
  NAND3_X1 U13755 ( .A1(n12138), .A2(n12137), .A3(n12136), .ZN(n12140) );
  INV_X1 U13756 ( .A(n12343), .ZN(n12139) );
  AND2_X1 U13757 ( .A1(n19249), .A2(n12819), .ZN(n14470) );
  INV_X1 U13758 ( .A(n14470), .ZN(n19250) );
  NOR2_X1 U13759 ( .A1(n19250), .A2(n12323), .ZN(n15335) );
  NAND2_X1 U13760 ( .A1(n15339), .A2(n15335), .ZN(n12366) );
  OAI21_X1 U13761 ( .B1(n19523), .B2(n12620), .A(n12366), .ZN(n15351) );
  NAND2_X1 U13762 ( .A1(n15351), .A2(n19511), .ZN(n19539) );
  OR2_X1 U13763 ( .A1(n12622), .A2(n18184), .ZN(n12322) );
  NAND2_X1 U13764 ( .A1(n12143), .A2(n12142), .ZN(n12145) );
  INV_X1 U13765 ( .A(n12416), .ZN(n12144) );
  NAND2_X1 U13766 ( .A1(n12145), .A2(n12144), .ZN(n12146) );
  INV_X1 U13767 ( .A(n15565), .ZN(n12155) );
  INV_X1 U13768 ( .A(n12147), .ZN(n12148) );
  XOR2_X1 U13769 ( .A(n12149), .B(n12148), .Z(n16419) );
  XOR2_X1 U13770 ( .A(n12390), .B(n12375), .Z(n12150) );
  NAND2_X1 U13771 ( .A1(n14630), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14629) );
  NOR2_X1 U13772 ( .A1(n12150), .A2(n14629), .ZN(n12151) );
  INV_X1 U13773 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14696) );
  XNOR2_X1 U13774 ( .A(n12150), .B(n14629), .ZN(n14695) );
  NOR2_X1 U13775 ( .A1(n14696), .A2(n14695), .ZN(n14694) );
  NOR2_X1 U13776 ( .A1(n12151), .A2(n14694), .ZN(n12152) );
  XOR2_X1 U13777 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12152), .Z(
        n16418) );
  NOR2_X1 U13778 ( .A1(n16419), .A2(n16418), .ZN(n16417) );
  INV_X1 U13779 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16425) );
  NOR2_X1 U13780 ( .A1(n12152), .A2(n16425), .ZN(n12153) );
  OR2_X1 U13781 ( .A1(n16417), .A2(n12153), .ZN(n12156) );
  XNOR2_X1 U13782 ( .A(n12156), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15564) );
  NAND2_X1 U13783 ( .A1(n12156), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12157) );
  INV_X1 U13784 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16325) );
  INV_X1 U13785 ( .A(n12158), .ZN(n12160) );
  NAND2_X1 U13786 ( .A1(n12160), .A2(n12159), .ZN(n12161) );
  INV_X1 U13787 ( .A(n12167), .ZN(n12165) );
  NAND2_X1 U13788 ( .A1(n12141), .A2(n12419), .ZN(n12163) );
  NAND2_X1 U13789 ( .A1(n12162), .A2(n12163), .ZN(n12171) );
  NAND2_X1 U13790 ( .A1(n12165), .A2(n12164), .ZN(n12178) );
  NAND2_X1 U13791 ( .A1(n12167), .A2(n12171), .ZN(n12166) );
  INV_X1 U13792 ( .A(n12179), .ZN(n12170) );
  OAI21_X1 U13793 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12164), .A(
        n12170), .ZN(n12175) );
  INV_X1 U13794 ( .A(n12181), .ZN(n12172) );
  MUX2_X1 U13795 ( .A(n12172), .B(n16324), .S(n12171), .Z(n12173) );
  OAI21_X1 U13796 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12179), .A(
        n12173), .ZN(n12174) );
  INV_X1 U13797 ( .A(n12176), .ZN(n12177) );
  NAND2_X1 U13798 ( .A1(n16319), .A2(n11190), .ZN(n12180) );
  INV_X1 U13799 ( .A(n12162), .ZN(n12182) );
  XNOR2_X1 U13800 ( .A(n12183), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17738) );
  INV_X1 U13801 ( .A(n12183), .ZN(n12184) );
  NAND2_X1 U13802 ( .A1(n12184), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12185) );
  INV_X1 U13803 ( .A(n12187), .ZN(n12188) );
  NAND2_X1 U13804 ( .A1(n12188), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12189) );
  AND2_X1 U13805 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17931) );
  AND2_X1 U13806 ( .A1(n17931), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17952) );
  AND2_X1 U13807 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12190) );
  AND2_X1 U13808 ( .A1(n17952), .A2(n12190), .ZN(n17925) );
  NAND2_X1 U13809 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12192) );
  AND3_X1 U13810 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17841) );
  AND3_X1 U13811 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U13812 ( .A1(n17841), .A2(n12191), .ZN(n12594) );
  OR2_X1 U13813 ( .A1(n17928), .A2(n12594), .ZN(n12656) );
  NOR2_X1 U13814 ( .A1(n12192), .A2(n12656), .ZN(n17597) );
  AND2_X1 U13815 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17597), .ZN(
        n12193) );
  INV_X1 U13816 ( .A(n17578), .ZN(n12194) );
  NAND2_X1 U13817 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14184) );
  INV_X1 U13818 ( .A(n14184), .ZN(n12195) );
  NAND2_X1 U13819 ( .A1(n13013), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12197) );
  OR2_X1 U13820 ( .A1(n19539), .A2(n12954), .ZN(n18185) );
  NAND2_X1 U13821 ( .A1(n12619), .A2(n18198), .ZN(n12321) );
  INV_X1 U13822 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14472) );
  AOI22_X1 U13823 ( .A1(n12306), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12199) );
  NAND2_X1 U13824 ( .A1(n11777), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12198) );
  OAI211_X1 U13825 ( .C1(n12299), .C2(n14472), .A(n12199), .B(n12198), .ZN(
        n12313) );
  INV_X1 U13826 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12204) );
  NAND2_X1 U13827 ( .A1(n12312), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12203) );
  AOI22_X1 U13828 ( .A1(n12306), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12202) );
  OAI211_X1 U13829 ( .C1(n12309), .C2(n12204), .A(n12203), .B(n12202), .ZN(
        n14909) );
  AOI22_X1 U13830 ( .A1(n12306), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12205) );
  OAI21_X1 U13831 ( .B1(n12309), .B2(n14918), .A(n12205), .ZN(n12206) );
  AOI21_X1 U13832 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12206), .ZN(n14916) );
  NAND2_X1 U13833 ( .A1(n12312), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12208) );
  AOI22_X1 U13834 ( .A1(n12306), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12207) );
  OAI211_X1 U13835 ( .C1(n12309), .C2(n12209), .A(n12208), .B(n12207), .ZN(
        n14924) );
  INV_X1 U13836 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U13837 ( .A1(n12306), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12210) );
  OAI21_X1 U13838 ( .B1(n12309), .B2(n12211), .A(n12210), .ZN(n12212) );
  AOI21_X1 U13839 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12212), .ZN(n14929) );
  OR2_X1 U13840 ( .A1(n12299), .A2(n18037), .ZN(n12217) );
  NAND2_X1 U13841 ( .A1(n12306), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U13842 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12213) );
  OAI211_X1 U13843 ( .C1(n12309), .C2(n19298), .A(n12214), .B(n12213), .ZN(
        n12215) );
  INV_X1 U13844 ( .A(n12215), .ZN(n12216) );
  NAND2_X1 U13845 ( .A1(n12217), .A2(n12216), .ZN(n15087) );
  INV_X1 U13846 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12220) );
  INV_X1 U13847 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17727) );
  OR2_X1 U13848 ( .A1(n12299), .A2(n17727), .ZN(n12219) );
  AOI22_X1 U13849 ( .A1(n12306), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12218) );
  OAI211_X1 U13850 ( .C1(n12309), .C2(n12220), .A(n12219), .B(n12218), .ZN(
        n15194) );
  INV_X1 U13851 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U13852 ( .A1(n12306), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U13853 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12221) );
  OAI211_X1 U13854 ( .C1(n12309), .C2(n12223), .A(n12222), .B(n12221), .ZN(
        n12224) );
  AOI21_X1 U13855 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12224), .ZN(n15590) );
  OR2_X1 U13856 ( .A1(n12299), .A2(n17965), .ZN(n12226) );
  AOI22_X1 U13857 ( .A1(n12306), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12225) );
  OAI211_X1 U13858 ( .C1(n12309), .C2(n12227), .A(n12226), .B(n12225), .ZN(
        n15639) );
  INV_X1 U13859 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U13860 ( .A1(n12306), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12229) );
  NAND2_X1 U13861 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12228) );
  OAI211_X1 U13862 ( .C1(n12309), .C2(n12230), .A(n12229), .B(n12228), .ZN(
        n12231) );
  AOI21_X1 U13863 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12231), .ZN(n15665) );
  NOR2_X2 U13864 ( .A1(n15666), .A2(n15665), .ZN(n15664) );
  INV_X1 U13865 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12234) );
  NAND2_X1 U13866 ( .A1(n12306), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12233) );
  NAND2_X1 U13867 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12232) );
  OAI211_X1 U13868 ( .C1(n12309), .C2(n12234), .A(n12233), .B(n12232), .ZN(
        n12235) );
  AOI21_X1 U13869 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12235), .ZN(n16256) );
  OR2_X1 U13870 ( .A1(n12299), .A2(n17928), .ZN(n12241) );
  INV_X1 U13871 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12237) );
  NOR2_X1 U13872 ( .A1(n12309), .A2(n12237), .ZN(n12239) );
  INV_X1 U13873 ( .A(n12306), .ZN(n12301) );
  INV_X1 U13874 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17924) );
  OAI22_X1 U13875 ( .A1(n12301), .A2(n17924), .B1(n18105), .B2(n11338), .ZN(
        n12238) );
  NOR2_X1 U13876 ( .A1(n12239), .A2(n12238), .ZN(n12240) );
  NAND2_X1 U13877 ( .A1(n12241), .A2(n12240), .ZN(n16364) );
  INV_X1 U13878 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14530) );
  NAND2_X1 U13879 ( .A1(n12306), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U13880 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12242) );
  OAI211_X1 U13881 ( .C1(n12309), .C2(n14530), .A(n12243), .B(n12242), .ZN(
        n12244) );
  AOI21_X1 U13882 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12244), .ZN(n14535) );
  NAND2_X1 U13883 ( .A1(n12306), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U13884 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12245) );
  OAI211_X1 U13885 ( .C1(n12309), .C2(n12247), .A(n12246), .B(n12245), .ZN(
        n12248) );
  AOI21_X1 U13886 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12248), .ZN(n17447) );
  NAND2_X1 U13887 ( .A1(n12306), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U13888 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12249) );
  OAI211_X1 U13889 ( .C1(n12309), .C2(n12251), .A(n12250), .B(n12249), .ZN(
        n12252) );
  AOI21_X1 U13890 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12252), .ZN(n16398) );
  OR2_X1 U13891 ( .A1(n12299), .A2(n17866), .ZN(n12257) );
  INV_X1 U13892 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12253) );
  NOR2_X1 U13893 ( .A1(n12309), .A2(n12253), .ZN(n12255) );
  INV_X1 U13894 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19372) );
  INV_X1 U13895 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n19370) );
  OAI22_X1 U13896 ( .A1(n12301), .A2(n19372), .B1(n18105), .B2(n19370), .ZN(
        n12254) );
  NOR2_X1 U13897 ( .A1(n12255), .A2(n12254), .ZN(n12256) );
  NAND2_X1 U13898 ( .A1(n12257), .A2(n12256), .ZN(n17440) );
  INV_X1 U13899 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12260) );
  OR2_X1 U13900 ( .A1(n12299), .A2(n17853), .ZN(n12259) );
  AOI22_X1 U13901 ( .A1(n12306), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12258) );
  OAI211_X1 U13902 ( .C1(n12309), .C2(n12260), .A(n12259), .B(n12258), .ZN(
        n17312) );
  NAND2_X1 U13903 ( .A1(n12306), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12262) );
  NAND2_X1 U13904 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12261) );
  OAI211_X1 U13905 ( .C1(n12309), .C2(n12263), .A(n12262), .B(n12261), .ZN(
        n12264) );
  AOI21_X1 U13906 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12264), .ZN(n12659) );
  INV_X1 U13907 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U13908 ( .A1(n12306), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12266) );
  NAND2_X1 U13909 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12265) );
  OAI211_X1 U13910 ( .C1(n12309), .C2(n12267), .A(n12266), .B(n12265), .ZN(
        n12268) );
  AOI21_X1 U13911 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12268), .ZN(n17413) );
  INV_X1 U13912 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U13913 ( .A1(n12306), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U13914 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12269) );
  OAI211_X1 U13915 ( .C1(n12309), .C2(n12271), .A(n12270), .B(n12269), .ZN(
        n12272) );
  AOI21_X1 U13916 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12272), .ZN(n17407) );
  INV_X1 U13917 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12275) );
  OR2_X1 U13918 ( .A1(n12299), .A2(n12072), .ZN(n12274) );
  AOI22_X1 U13919 ( .A1(n12306), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12273) );
  OAI211_X1 U13920 ( .C1(n12309), .C2(n12275), .A(n12274), .B(n12273), .ZN(
        n17296) );
  INV_X1 U13921 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17794) );
  OR2_X1 U13922 ( .A1(n12299), .A2(n17794), .ZN(n12280) );
  NOR2_X1 U13923 ( .A1(n12309), .A2(n12276), .ZN(n12278) );
  INV_X1 U13924 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n18302) );
  INV_X1 U13925 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14473) );
  OAI22_X1 U13926 ( .A1(n12301), .A2(n18302), .B1(n18105), .B2(n14473), .ZN(
        n12277) );
  NOR2_X1 U13927 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NAND2_X1 U13928 ( .A1(n12280), .A2(n12279), .ZN(n17280) );
  INV_X1 U13929 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17784) );
  OR2_X1 U13930 ( .A1(n12299), .A2(n17784), .ZN(n12285) );
  INV_X1 U13931 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12281) );
  NOR2_X1 U13932 ( .A1(n12309), .A2(n12281), .ZN(n12283) );
  INV_X1 U13933 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n18303) );
  INV_X1 U13934 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17583) );
  OAI22_X1 U13935 ( .A1(n12301), .A2(n18303), .B1(n18105), .B2(n17583), .ZN(
        n12282) );
  NOR2_X1 U13936 ( .A1(n12283), .A2(n12282), .ZN(n12284) );
  NAND2_X1 U13937 ( .A1(n12285), .A2(n12284), .ZN(n17392) );
  INV_X1 U13938 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U13939 ( .A1(n12306), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12287) );
  NAND2_X1 U13940 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12286) );
  OAI211_X1 U13941 ( .C1(n12309), .C2(n12288), .A(n12287), .B(n12286), .ZN(
        n12289) );
  AOI21_X1 U13942 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12289), .ZN(n17385) );
  INV_X1 U13943 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U13944 ( .A1(n12306), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12291) );
  NAND2_X1 U13945 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12290) );
  OAI211_X1 U13946 ( .C1(n12309), .C2(n12292), .A(n12291), .B(n12290), .ZN(
        n12293) );
  AOI21_X1 U13947 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12293), .ZN(n17271) );
  OR2_X1 U13948 ( .A1(n12299), .A2(n16407), .ZN(n12298) );
  INV_X1 U13949 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12294) );
  NOR2_X1 U13950 ( .A1(n12309), .A2(n12294), .ZN(n12296) );
  INV_X1 U13951 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n18307) );
  INV_X1 U13952 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14204) );
  OAI22_X1 U13953 ( .A1(n12301), .A2(n18307), .B1(n18105), .B2(n14204), .ZN(
        n12295) );
  NOR2_X1 U13954 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  NAND2_X1 U13955 ( .A1(n12298), .A2(n12297), .ZN(n14202) );
  OR2_X1 U13956 ( .A1(n12299), .A2(n14185), .ZN(n12305) );
  NOR2_X1 U13957 ( .A1(n12309), .A2(n12300), .ZN(n12303) );
  INV_X1 U13958 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n18309) );
  INV_X1 U13959 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13017) );
  OAI22_X1 U13960 ( .A1(n12301), .A2(n18309), .B1(n18105), .B2(n13017), .ZN(
        n12302) );
  NOR2_X1 U13961 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  NAND2_X1 U13962 ( .A1(n12305), .A2(n12304), .ZN(n13015) );
  INV_X1 U13963 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U13964 ( .A1(n12306), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U13965 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12307) );
  OAI211_X1 U13966 ( .C1(n12310), .C2(n12309), .A(n12308), .B(n12307), .ZN(
        n12311) );
  AOI21_X1 U13967 ( .B1(n12312), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12311), .ZN(n12637) );
  NOR2_X1 U13968 ( .A1(n18105), .A2(n20103), .ZN(n15499) );
  INV_X1 U13969 ( .A(n15499), .ZN(n18205) );
  NAND2_X1 U13970 ( .A1(n20165), .A2(n18205), .ZN(n19245) );
  OR2_X1 U13971 ( .A1(n19245), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12314) );
  AND2_X1 U13972 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12315) );
  INV_X1 U13973 ( .A(n15498), .ZN(n15358) );
  INV_X1 U13974 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22411) );
  NAND2_X1 U13975 ( .A1(n22411), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U13976 ( .A1(n15358), .A2(n12316), .ZN(n14633) );
  INV_X1 U13977 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17741) );
  INV_X1 U13978 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16332) );
  NAND2_X1 U13979 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n14491), .ZN(
        n14490) );
  INV_X1 U13980 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19358) );
  AND2_X2 U13981 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n14507), .ZN(
        n14508) );
  INV_X1 U13982 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17574) );
  INV_X1 U13983 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14459) );
  AND2_X1 U13984 ( .A1(n20167), .A2(n12317), .ZN(n12603) );
  INV_X1 U13985 ( .A(n14452), .ZN(n19360) );
  NAND2_X1 U13986 ( .A1(n19360), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U13987 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12318) );
  OAI211_X1 U13988 ( .C1(n18181), .C2(n14471), .A(n12597), .B(n12318), .ZN(
        n12319) );
  INV_X1 U13989 ( .A(n12319), .ZN(n12320) );
  NAND4_X1 U13990 ( .A1(n12322), .A2(n12321), .A3(n11504), .A4(n12320), .ZN(
        P2_U2983) );
  OR2_X1 U13991 ( .A1(n12323), .A2(n12819), .ZN(n12369) );
  AOI21_X1 U13992 ( .B1(n12342), .B2(n12954), .A(n12324), .ZN(n12336) );
  OAI211_X1 U13993 ( .C1(n12954), .C2(n12326), .A(n20528), .B(n12325), .ZN(
        n12331) );
  INV_X1 U13994 ( .A(n12327), .ZN(n12329) );
  OAI21_X1 U13995 ( .B1(n12329), .B2(n12328), .A(n11738), .ZN(n12330) );
  OAI211_X1 U13996 ( .C1(n12333), .C2(n12332), .A(n12331), .B(n12330), .ZN(
        n12335) );
  INV_X1 U13997 ( .A(n12338), .ZN(n12334) );
  OAI211_X1 U13998 ( .C1(n12337), .C2(n12336), .A(n12335), .B(n12334), .ZN(
        n12340) );
  AOI21_X1 U13999 ( .B1(n11738), .B2(n12338), .A(n12343), .ZN(n12339) );
  NAND2_X1 U14000 ( .A1(n12340), .A2(n12339), .ZN(n12341) );
  MUX2_X1 U14001 ( .A(n12341), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19251), .Z(n12346) );
  NAND2_X1 U14002 ( .A1(n14682), .A2(n12343), .ZN(n12344) );
  NAND2_X1 U14003 ( .A1(n15472), .A2(n12954), .ZN(n14679) );
  NAND2_X1 U14004 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19531) );
  NAND2_X1 U14005 ( .A1(n18270), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n18316) );
  INV_X2 U14006 ( .A(n18316), .ZN(n18311) );
  INV_X1 U14007 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n18272) );
  NAND2_X1 U14008 ( .A1(n18311), .A2(n18272), .ZN(n18313) );
  NOR2_X1 U14009 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n18099) );
  NAND2_X1 U14010 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n18099), .ZN(n18269) );
  NAND2_X1 U14011 ( .A1(n18308), .A2(n18269), .ZN(n19252) );
  NAND2_X1 U14012 ( .A1(n19531), .A2(n19252), .ZN(n12361) );
  NAND2_X1 U14013 ( .A1(n15332), .A2(n12345), .ZN(n12349) );
  AOI21_X1 U14014 ( .B1(n12346), .B2(n20528), .A(n11725), .ZN(n12347) );
  NAND2_X1 U14015 ( .A1(n14679), .A2(n12347), .ZN(n12348) );
  OAI21_X1 U14016 ( .B1(n14679), .B2(n12349), .A(n12348), .ZN(n12350) );
  INV_X1 U14017 ( .A(n12350), .ZN(n12368) );
  OAI21_X1 U14018 ( .B1(n12352), .B2(n11725), .A(n11727), .ZN(n12360) );
  NAND2_X1 U14019 ( .A1(n12358), .A2(n13007), .ZN(n12353) );
  NAND2_X1 U14020 ( .A1(n12353), .A2(n14470), .ZN(n12583) );
  NAND2_X1 U14021 ( .A1(n12819), .A2(n12357), .ZN(n12569) );
  NAND2_X1 U14022 ( .A1(n12569), .A2(n20528), .ZN(n12354) );
  NAND3_X1 U14023 ( .A1(n12354), .A2(n12584), .A3(n13007), .ZN(n12355) );
  NAND2_X1 U14024 ( .A1(n12355), .A2(n11727), .ZN(n12356) );
  OAI211_X1 U14025 ( .C1(n12358), .C2(n12357), .A(n12583), .B(n12356), .ZN(
        n12359) );
  AOI21_X1 U14026 ( .B1(n12351), .B2(n12360), .A(n12359), .ZN(n12571) );
  INV_X1 U14027 ( .A(n14564), .ZN(n15336) );
  NOR2_X1 U14028 ( .A1(n15336), .A2(n12361), .ZN(n12362) );
  NAND2_X1 U14029 ( .A1(n11169), .A2(n12362), .ZN(n12363) );
  AND2_X1 U14030 ( .A1(n12571), .A2(n12363), .ZN(n15290) );
  MUX2_X1 U14031 ( .A(n11169), .B(n12345), .S(n12819), .Z(n12364) );
  NAND3_X1 U14032 ( .A1(n12364), .A2(n14564), .A3(n19531), .ZN(n12365) );
  AND3_X1 U14033 ( .A1(n15290), .A2(n12366), .A3(n12365), .ZN(n12367) );
  OAI211_X1 U14034 ( .C1(n19523), .C2(n12369), .A(n12368), .B(n12367), .ZN(
        n12370) );
  NAND2_X1 U14035 ( .A1(n11168), .A2(n12819), .ZN(n12372) );
  NAND2_X1 U14036 ( .A1(n12372), .A2(n11773), .ZN(n12373) );
  NOR2_X1 U14037 ( .A1(n13007), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12403) );
  AND2_X1 U14038 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12374) );
  NOR2_X1 U14039 ( .A1(n12403), .A2(n12374), .ZN(n12381) );
  NAND2_X1 U14040 ( .A1(n12402), .A2(n12352), .ZN(n12399) );
  INV_X1 U14041 ( .A(n12382), .ZN(n12378) );
  NAND3_X1 U14042 ( .A1(n12381), .A2(n12399), .A3(n12380), .ZN(n19262) );
  INV_X1 U14043 ( .A(n12998), .ZN(n12383) );
  NOR2_X2 U14044 ( .A1(n12383), .A2(n12382), .ZN(n12401) );
  NAND2_X1 U14045 ( .A1(n12401), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12387) );
  INV_X1 U14046 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19496) );
  NAND2_X1 U14047 ( .A1(n15513), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12384) );
  OAI211_X1 U14048 ( .C1(n12376), .C2(n19496), .A(n12384), .B(n20165), .ZN(
        n12385) );
  INV_X1 U14049 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U14050 ( .A1(n12387), .A2(n12386), .ZN(n19261) );
  NAND2_X1 U14051 ( .A1(n19262), .A2(n19261), .ZN(n12395) );
  AOI22_X1 U14052 ( .A1(n12402), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12403), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12389) );
  NAND2_X1 U14053 ( .A1(n12401), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12388) );
  XNOR2_X1 U14054 ( .A(n12395), .B(n12394), .ZN(n14824) );
  OR2_X1 U14055 ( .A1(n12390), .A2(n12529), .ZN(n12393) );
  NAND2_X1 U14056 ( .A1(n11746), .A2(n13007), .ZN(n12391) );
  MUX2_X1 U14057 ( .A(n12391), .B(n20150), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12392) );
  AND2_X1 U14058 ( .A1(n12393), .A2(n12392), .ZN(n14823) );
  NAND2_X1 U14059 ( .A1(n14824), .A2(n14823), .ZN(n14822) );
  NAND2_X1 U14060 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  NAND2_X1 U14061 ( .A1(n14822), .A2(n12397), .ZN(n12407) );
  OR2_X1 U14062 ( .A1(n12529), .A2(n12398), .ZN(n12400) );
  OAI211_X1 U14063 ( .C1(n20165), .C2(n20146), .A(n12400), .B(n12399), .ZN(
        n12406) );
  XNOR2_X1 U14064 ( .A(n12407), .B(n12406), .ZN(n15485) );
  NAND2_X1 U14065 ( .A1(n11163), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U14066 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12404) );
  AND2_X1 U14067 ( .A1(n12405), .A2(n12404), .ZN(n15484) );
  INV_X1 U14068 ( .A(n12406), .ZN(n12408) );
  NAND2_X1 U14069 ( .A1(n12408), .A2(n12407), .ZN(n12409) );
  NAND2_X1 U14070 ( .A1(n11163), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U14071 ( .A1(n12563), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12413) );
  NAND2_X1 U14072 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12412) );
  OR2_X1 U14073 ( .A1(n12529), .A2(n12410), .ZN(n12411) );
  AOI22_X1 U14074 ( .A1(n11163), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n12563), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U14075 ( .A1(n12379), .A2(n12416), .B1(n12560), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U14076 ( .A1(n12418), .A2(n12417), .ZN(n16277) );
  NAND2_X1 U14077 ( .A1(n16276), .A2(n16277), .ZN(n15181) );
  NAND2_X1 U14078 ( .A1(n11163), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U14079 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12421) );
  OR2_X1 U14080 ( .A1(n12529), .A2(n12419), .ZN(n12420) );
  NOR2_X2 U14081 ( .A1(n15181), .A2(n15182), .ZN(n15180) );
  NOR2_X1 U14082 ( .A1(n15180), .A2(n12424), .ZN(n18058) );
  AOI222_X1 U14083 ( .A1(n11163), .A2(P2_REIP_REG_6__SCAN_IN), .B1(n12560), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(n12563), .C2(
        P2_EAX_REG_6__SCAN_IN), .ZN(n18059) );
  NOR2_X2 U14084 ( .A1(n18058), .A2(n18059), .ZN(n18057) );
  AOI222_X1 U14085 ( .A1(n11163), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n12560), 
        .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12563), .C2(
        P2_EAX_REG_7__SCAN_IN), .ZN(n15198) );
  AOI22_X1 U14086 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U14087 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U14088 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12783), .B1(
        n11871), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U14089 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11211), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12426) );
  NAND4_X1 U14090 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12435) );
  AOI22_X1 U14091 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U14092 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11878), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U14093 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11591), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U14094 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12788), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12430) );
  NAND4_X1 U14095 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12434) );
  INV_X1 U14096 ( .A(n15094), .ZN(n12438) );
  AOI22_X1 U14097 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12437) );
  NAND2_X1 U14098 ( .A1(n11163), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12436) );
  OAI211_X1 U14099 ( .C1(n12529), .C2(n12438), .A(n12437), .B(n12436), .ZN(
        n18033) );
  NAND2_X1 U14100 ( .A1(n11163), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U14101 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U14102 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U14103 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U14104 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U14105 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12439) );
  NAND4_X1 U14106 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12448) );
  AOI22_X1 U14107 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U14108 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U14109 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U14110 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12443) );
  NAND4_X1 U14111 ( .A1(n12446), .A2(n12445), .A3(n12444), .A4(n12443), .ZN(
        n12447) );
  NOR2_X1 U14112 ( .A1(n12448), .A2(n12447), .ZN(n15191) );
  OR2_X1 U14113 ( .A1(n12529), .A2(n15191), .ZN(n12449) );
  AOI22_X1 U14114 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12726), .B1(
        n11870), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U14115 ( .A1(n11871), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U14116 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11206), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U14117 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U14118 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12461) );
  AOI22_X1 U14119 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U14120 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U14121 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U14122 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12456) );
  NAND4_X1 U14123 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n12460) );
  NOR2_X1 U14124 ( .A1(n12461), .A2(n12460), .ZN(n15593) );
  AOI22_X1 U14125 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12463) );
  NAND2_X1 U14126 ( .A1(n11163), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12462) );
  OAI211_X1 U14127 ( .C1(n12529), .C2(n15593), .A(n12463), .B(n12462), .ZN(
        n17990) );
  NAND2_X1 U14128 ( .A1(n11163), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U14129 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U14130 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U14131 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U14132 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U14133 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12464) );
  NAND4_X1 U14134 ( .A1(n12467), .A2(n12466), .A3(n12465), .A4(n12464), .ZN(
        n12473) );
  AOI22_X1 U14135 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U14136 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11878), .B1(
        n11211), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U14137 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U14138 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12468) );
  NAND4_X1 U14139 ( .A1(n12471), .A2(n12470), .A3(n12469), .A4(n12468), .ZN(
        n12472) );
  OR2_X1 U14140 ( .A1(n12473), .A2(n12472), .ZN(n15638) );
  INV_X1 U14141 ( .A(n15638), .ZN(n12474) );
  OR2_X1 U14142 ( .A1(n12529), .A2(n12474), .ZN(n12475) );
  AOI22_X1 U14143 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U14144 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U14145 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11220), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U14146 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11878), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12478) );
  NAND4_X1 U14147 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12487) );
  AOI22_X1 U14148 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U14149 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11211), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U14150 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U14151 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12482) );
  NAND4_X1 U14152 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n12486) );
  INV_X1 U14153 ( .A(n15669), .ZN(n12490) );
  AOI22_X1 U14154 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U14155 ( .A1(n11163), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12488) );
  OAI211_X1 U14156 ( .C1(n12529), .C2(n12490), .A(n12489), .B(n12488), .ZN(
        n17950) );
  AOI22_X1 U14157 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U14158 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U14159 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n11220), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U14160 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U14161 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12500) );
  AOI22_X1 U14162 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U14163 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U14164 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U14165 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U14166 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12499) );
  NOR2_X1 U14167 ( .A1(n12500), .A2(n12499), .ZN(n16252) );
  AOI22_X1 U14168 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U14169 ( .A1(n11163), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12501) );
  OAI211_X1 U14170 ( .C1(n16252), .C2(n12529), .A(n12502), .B(n12501), .ZN(
        n17328) );
  NAND2_X1 U14171 ( .A1(n11163), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U14172 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U14173 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12783), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U14174 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U14175 ( .A1(n11220), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11878), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12503) );
  NAND4_X1 U14177 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12512) );
  AOI22_X1 U14178 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U14179 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11211), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U14180 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11591), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U14181 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12788), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12507) );
  NAND4_X1 U14182 ( .A1(n12510), .A2(n12509), .A3(n12508), .A4(n12507), .ZN(
        n12511) );
  NOR2_X1 U14183 ( .A1(n12512), .A2(n12511), .ZN(n16369) );
  OR2_X1 U14184 ( .A1(n12529), .A2(n16369), .ZN(n12513) );
  AOI22_X1 U14185 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14186 ( .A1(n11163), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12516) );
  NAND2_X1 U14187 ( .A1(n12517), .A2(n12516), .ZN(n16391) );
  INV_X1 U14188 ( .A(n16391), .ZN(n12532) );
  AOI22_X1 U14189 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U14190 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U14191 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U14192 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11873), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12518) );
  NAND4_X1 U14193 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        n12527) );
  AOI22_X1 U14194 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U14195 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11210), .B1(
        n11878), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U14196 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U14197 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U14198 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n12526) );
  OR2_X1 U14199 ( .A1(n12527), .A2(n12526), .ZN(n16374) );
  INV_X1 U14200 ( .A(n16374), .ZN(n12530) );
  AOI22_X1 U14201 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12528) );
  OAI21_X1 U14202 ( .B1(n12530), .B2(n12529), .A(n12528), .ZN(n12531) );
  AOI21_X1 U14203 ( .B1(P2_REIP_REG_15__SCAN_IN), .B2(n11163), .A(n12531), 
        .ZN(n16389) );
  NAND2_X1 U14204 ( .A1(n11163), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U14205 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12533) );
  AND2_X1 U14206 ( .A1(n12534), .A2(n12533), .ZN(n17545) );
  OR2_X2 U14207 ( .A1(n17546), .A2(n17545), .ZN(n17548) );
  NAND2_X1 U14208 ( .A1(n11163), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U14209 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12535) );
  AND2_X1 U14210 ( .A1(n12536), .A2(n12535), .ZN(n17535) );
  NAND2_X1 U14211 ( .A1(n11163), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U14212 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12539) );
  INV_X1 U14213 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U14214 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12541) );
  OAI21_X1 U14215 ( .B1(n12415), .B2(n18298), .A(n12541), .ZN(n17520) );
  NAND2_X1 U14216 ( .A1(n11163), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U14217 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12542) );
  AND2_X1 U14218 ( .A1(n12543), .A2(n12542), .ZN(n17504) );
  NAND2_X1 U14219 ( .A1(n11163), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U14220 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12544) );
  AND2_X1 U14221 ( .A1(n12545), .A2(n12544), .ZN(n17512) );
  OR2_X1 U14222 ( .A1(n17504), .A2(n17512), .ZN(n12546) );
  AOI22_X1 U14223 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12548) );
  NAND2_X1 U14224 ( .A1(n11163), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U14225 ( .A1(n12548), .A2(n12547), .ZN(n17298) );
  AOI22_X1 U14226 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12549) );
  OAI21_X1 U14227 ( .B1(n12415), .B2(n18302), .A(n12549), .ZN(n17284) );
  NAND2_X1 U14228 ( .A1(n11163), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U14229 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12550) );
  AND2_X1 U14230 ( .A1(n12551), .A2(n12550), .ZN(n17481) );
  INV_X1 U14231 ( .A(n17481), .ZN(n12552) );
  NAND2_X1 U14232 ( .A1(n11163), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U14233 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12554) );
  AND2_X1 U14234 ( .A1(n12555), .A2(n12554), .ZN(n17474) );
  NAND2_X1 U14235 ( .A1(n11163), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U14236 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12556) );
  AND2_X1 U14237 ( .A1(n12557), .A2(n12556), .ZN(n17268) );
  AOI22_X1 U14238 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12558) );
  OAI21_X1 U14239 ( .B1(n12415), .B2(n18307), .A(n12558), .ZN(n16403) );
  AOI22_X1 U14240 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12559) );
  OAI21_X1 U14241 ( .B1(n12415), .B2(n18309), .A(n12559), .ZN(n14179) );
  AOI22_X1 U14242 ( .A1(n12560), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n12563), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U14243 ( .A1(n11163), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12561) );
  NAND2_X1 U14244 ( .A1(n12562), .A2(n12561), .ZN(n12983) );
  NAND2_X1 U14245 ( .A1(n12982), .A2(n12983), .ZN(n12987) );
  AOI222_X1 U14246 ( .A1(n11163), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12560), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12563), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n12564) );
  XNOR2_X1 U14247 ( .A(n12987), .B(n12564), .ZN(n14468) );
  NAND2_X1 U14248 ( .A1(n11761), .A2(n12954), .ZN(n12567) );
  AND2_X1 U14249 ( .A1(n12565), .A2(n12566), .ZN(n15282) );
  INV_X1 U14250 ( .A(n15282), .ZN(n15345) );
  NAND2_X1 U14251 ( .A1(n12567), .A2(n15345), .ZN(n12568) );
  NAND2_X1 U14252 ( .A1(n12621), .A2(n12568), .ZN(n18066) );
  NAND2_X1 U14253 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12613) );
  INV_X1 U14254 ( .A(n12569), .ZN(n12570) );
  NAND2_X1 U14255 ( .A1(n12621), .A2(n15341), .ZN(n17877) );
  NOR2_X1 U14256 ( .A1(n18037), .A2(n18046), .ZN(n18024) );
  NAND3_X1 U14257 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18026) );
  NOR2_X1 U14258 ( .A1(n18068), .A2(n18026), .ZN(n12590) );
  NAND2_X1 U14259 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16415) );
  NAND2_X1 U14260 ( .A1(n16425), .A2(n16415), .ZN(n16420) );
  NAND3_X1 U14261 ( .A1(n18024), .A2(n12590), .A3(n16420), .ZN(n12601) );
  NOR2_X1 U14262 ( .A1(n17877), .A2(n12601), .ZN(n12593) );
  OAI21_X1 U14263 ( .B1(n12572), .B2(n12574), .A(n12573), .ZN(n12576) );
  NAND2_X1 U14264 ( .A1(n12576), .A2(n12575), .ZN(n12581) );
  OR2_X1 U14265 ( .A1(n12573), .A2(n11725), .ZN(n12580) );
  INV_X1 U14266 ( .A(n12577), .ZN(n12578) );
  NAND2_X1 U14267 ( .A1(n12578), .A2(n12572), .ZN(n12978) );
  NAND2_X1 U14268 ( .A1(n19249), .A2(n12345), .ZN(n12579) );
  AND4_X1 U14269 ( .A1(n12581), .A2(n12580), .A3(n12978), .A4(n12579), .ZN(
        n12587) );
  NAND2_X1 U14270 ( .A1(n12582), .A2(n12954), .ZN(n15296) );
  NAND2_X1 U14271 ( .A1(n15296), .A2(n12583), .ZN(n12585) );
  NAND2_X1 U14272 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  AND3_X1 U14273 ( .A1(n12588), .A2(n12587), .A3(n12586), .ZN(n15303) );
  NAND2_X1 U14274 ( .A1(n15303), .A2(n15276), .ZN(n12589) );
  NAND2_X1 U14275 ( .A1(n12621), .A2(n12589), .ZN(n18028) );
  OR2_X1 U14276 ( .A1(n16425), .A2(n16415), .ZN(n16421) );
  INV_X1 U14277 ( .A(n12590), .ZN(n12591) );
  NOR2_X1 U14278 ( .A1(n16421), .A2(n12591), .ZN(n18029) );
  NAND2_X1 U14279 ( .A1(n18029), .A2(n18024), .ZN(n12602) );
  NOR2_X1 U14280 ( .A1(n18028), .A2(n12602), .ZN(n12592) );
  NAND2_X1 U14281 ( .A1(n17925), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17837) );
  NOR2_X1 U14282 ( .A1(n17837), .A2(n12594), .ZN(n17827) );
  AND2_X1 U14283 ( .A1(n17827), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12607) );
  AND2_X1 U14284 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12610) );
  NAND2_X1 U14285 ( .A1(n17819), .A2(n12610), .ZN(n12599) );
  NOR2_X1 U14286 ( .A1(n17794), .A2(n12599), .ZN(n17783) );
  INV_X1 U14287 ( .A(n17783), .ZN(n17767) );
  NOR2_X1 U14288 ( .A1(n12613), .A2(n17767), .ZN(n14182) );
  NAND2_X1 U14289 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12595) );
  NOR2_X1 U14290 ( .A1(n14184), .A2(n12595), .ZN(n12615) );
  NAND3_X1 U14291 ( .A1(n14182), .A2(n12615), .A3(n14472), .ZN(n12596) );
  OAI211_X1 U14292 ( .C1(n14468), .C2(n18066), .A(n12597), .B(n12596), .ZN(
        n12598) );
  INV_X1 U14293 ( .A(n12598), .ZN(n12617) );
  NAND2_X1 U14294 ( .A1(n17877), .A2(n18028), .ZN(n17838) );
  INV_X1 U14295 ( .A(n12599), .ZN(n12600) );
  NAND2_X1 U14296 ( .A1(n12600), .A2(n17794), .ZN(n17797) );
  INV_X1 U14297 ( .A(n17877), .ZN(n18030) );
  NAND2_X1 U14298 ( .A1(n18030), .A2(n12601), .ZN(n12606) );
  INV_X1 U14299 ( .A(n18028), .ZN(n17880) );
  NAND2_X1 U14300 ( .A1(n17880), .A2(n12602), .ZN(n12605) );
  INV_X1 U14301 ( .A(n12621), .ZN(n12604) );
  INV_X1 U14302 ( .A(n12603), .ZN(n14452) );
  NAND2_X1 U14303 ( .A1(n12604), .A2(n14452), .ZN(n19497) );
  INV_X1 U14304 ( .A(n12607), .ZN(n12608) );
  NAND2_X1 U14305 ( .A1(n17838), .A2(n12608), .ZN(n12609) );
  NAND2_X1 U14306 ( .A1(n18003), .A2(n12609), .ZN(n17826) );
  INV_X1 U14307 ( .A(n12610), .ZN(n12611) );
  AND2_X1 U14308 ( .A1(n17838), .A2(n12611), .ZN(n12612) );
  NOR2_X1 U14309 ( .A1(n17826), .A2(n12612), .ZN(n17795) );
  AND2_X1 U14310 ( .A1(n17797), .A2(n17795), .ZN(n17782) );
  NAND2_X1 U14311 ( .A1(n17838), .A2(n12613), .ZN(n12614) );
  AND2_X1 U14312 ( .A1(n17782), .A2(n12614), .ZN(n14183) );
  OAI21_X1 U14313 ( .B1(n19502), .B2(n12615), .A(n14183), .ZN(n14440) );
  NAND2_X1 U14314 ( .A1(n14440), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12616) );
  NAND2_X1 U14315 ( .A1(n12621), .A2(n15335), .ZN(n19508) );
  NAND2_X1 U14316 ( .A1(n12619), .A2(n18055), .ZN(n12624) );
  INV_X1 U14317 ( .A(n12620), .ZN(n15342) );
  OR2_X1 U14318 ( .A1(n12622), .A2(n19495), .ZN(n12623) );
  NAND3_X1 U14319 ( .A1(n12625), .A2(n12624), .A3(n12623), .ZN(P2_U3015) );
  NAND2_X1 U14320 ( .A1(n12626), .A2(n13021), .ZN(n12631) );
  INV_X1 U14321 ( .A(n12627), .ZN(n12628) );
  NOR2_X1 U14322 ( .A1(n12629), .A2(n12628), .ZN(n12630) );
  XNOR2_X1 U14323 ( .A(n12631), .B(n12630), .ZN(n14435) );
  INV_X1 U14324 ( .A(n14435), .ZN(n12634) );
  XNOR2_X1 U14325 ( .A(n13016), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n19483) );
  NAND2_X1 U14326 ( .A1(n19360), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14438) );
  NAND2_X1 U14327 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12632) );
  OAI211_X1 U14328 ( .C1(n18181), .C2(n19483), .A(n14438), .B(n12632), .ZN(
        n12633) );
  XNOR2_X1 U14329 ( .A(n13013), .B(n12635), .ZN(n14434) );
  NAND2_X1 U14330 ( .A1(n12636), .A2(n12637), .ZN(n12638) );
  NAND3_X1 U14331 ( .A1(n12641), .A2(n12640), .A3(n11488), .ZN(P2_U2984) );
  INV_X1 U14332 ( .A(n12643), .ZN(n17683) );
  INV_X1 U14333 ( .A(n12645), .ZN(n12646) );
  NAND2_X1 U14334 ( .A1(n12647), .A2(n12646), .ZN(n17663) );
  NAND2_X1 U14335 ( .A1(n17663), .A2(n17662), .ZN(n17661) );
  INV_X1 U14336 ( .A(n12648), .ZN(n12649) );
  INV_X1 U14337 ( .A(n12650), .ZN(n12651) );
  XNOR2_X1 U14338 ( .A(n17619), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17852) );
  NAND2_X2 U14339 ( .A1(n17896), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17878) );
  AOI21_X1 U14340 ( .B1(n17645), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12657) );
  INV_X1 U14341 ( .A(n17598), .ZN(n12655) );
  NOR2_X1 U14342 ( .A1(n12655), .A2(n12656), .ZN(n17624) );
  NAND2_X1 U14343 ( .A1(n12658), .A2(n12659), .ZN(n12660) );
  NAND2_X1 U14344 ( .A1(n17414), .A2(n12660), .ZN(n19384) );
  NOR2_X1 U14345 ( .A1(n19384), .A2(n18190), .ZN(n12663) );
  OAI21_X1 U14346 ( .B1(n14480), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14479), .ZN(n19387) );
  NAND2_X1 U14347 ( .A1(n12603), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n17842) );
  NAND2_X1 U14348 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12661) );
  OAI211_X1 U14349 ( .C1(n18181), .C2(n19387), .A(n17842), .B(n12661), .ZN(
        n12662) );
  AOI211_X1 U14350 ( .C1(n17850), .C2(n18198), .A(n12663), .B(n12662), .ZN(
        n12664) );
  NAND2_X1 U14351 ( .A1(n12665), .A2(n12664), .ZN(P2_U2994) );
  NAND2_X1 U14352 ( .A1(n11729), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U14353 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20147) );
  INV_X1 U14354 ( .A(n20147), .ZN(n12667) );
  NAND2_X1 U14355 ( .A1(n12667), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12675) );
  AOI21_X1 U14356 ( .B1(n12675), .B2(n20145), .A(n20192), .ZN(n12669) );
  INV_X1 U14357 ( .A(n12675), .ZN(n12668) );
  NAND2_X1 U14358 ( .A1(n12668), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20198) );
  AOI22_X1 U14359 ( .A1(n12687), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n12669), .B2(n20198), .ZN(n12670) );
  NOR2_X1 U14360 ( .A1(n12905), .A2(n12866), .ZN(n12671) );
  NAND2_X1 U14361 ( .A1(n12672), .A2(n12671), .ZN(n12696) );
  NAND2_X1 U14362 ( .A1(n20147), .A2(n20146), .ZN(n12674) );
  NAND2_X1 U14363 ( .A1(n12675), .A2(n12674), .ZN(n20058) );
  NOR2_X1 U14364 ( .A1(n20058), .A2(n20192), .ZN(n20050) );
  AOI21_X1 U14365 ( .B1(n12687), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n20050), .ZN(n12680) );
  INV_X1 U14366 ( .A(n12680), .ZN(n12676) );
  INV_X1 U14367 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12842) );
  NOR2_X1 U14368 ( .A1(n12905), .A2(n12842), .ZN(n12678) );
  INV_X1 U14369 ( .A(n12678), .ZN(n12679) );
  AND2_X1 U14370 ( .A1(n12680), .A2(n12679), .ZN(n12681) );
  NAND2_X1 U14371 ( .A1(n12682), .A2(n12681), .ZN(n12683) );
  NAND2_X1 U14372 ( .A1(n12694), .A2(n12683), .ZN(n14893) );
  NOR2_X1 U14373 ( .A1(n20192), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12684) );
  AOI21_X1 U14374 ( .B1(n12687), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12684), .ZN(n12685) );
  NAND2_X1 U14375 ( .A1(n12881), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12690) );
  NAND2_X1 U14376 ( .A1(n12687), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12688) );
  OAI21_X1 U14377 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n20147), .ZN(n20126) );
  OR2_X1 U14378 ( .A1(n20126), .A2(n20192), .ZN(n20162) );
  NAND2_X1 U14379 ( .A1(n12688), .A2(n20162), .ZN(n12689) );
  NAND2_X1 U14380 ( .A1(n14835), .A2(n14834), .ZN(n12693) );
  INV_X1 U14381 ( .A(n14743), .ZN(n12691) );
  NAND2_X1 U14382 ( .A1(n12691), .A2(n12690), .ZN(n12692) );
  NAND2_X1 U14383 ( .A1(n12693), .A2(n12692), .ZN(n14892) );
  NAND2_X1 U14384 ( .A1(n15495), .A2(n15497), .ZN(n15496) );
  NAND2_X1 U14385 ( .A1(n11729), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12695) );
  INV_X1 U14386 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12890) );
  NOR2_X1 U14387 ( .A1(n12905), .A2(n12890), .ZN(n14906) );
  INV_X1 U14388 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U14389 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U14390 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U14391 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11220), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U14392 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U14393 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12709) );
  AOI22_X1 U14394 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U14395 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U14396 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U14397 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12704) );
  NAND4_X1 U14398 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n12704), .ZN(
        n12708) );
  OR2_X1 U14399 ( .A1(n12709), .A2(n12708), .ZN(n17405) );
  AOI22_X1 U14400 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U14401 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U14402 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U14403 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12710) );
  NAND4_X1 U14404 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n12710), .ZN(
        n12719) );
  AOI22_X1 U14405 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U14406 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U14407 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U14408 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12714) );
  NAND4_X1 U14409 ( .A1(n12717), .A2(n12716), .A3(n12715), .A4(n12714), .ZN(
        n12718) );
  OR2_X1 U14410 ( .A1(n12719), .A2(n12718), .ZN(n17424) );
  AOI22_X1 U14411 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U14412 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U14413 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U14414 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12720) );
  NAND4_X1 U14415 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12737) );
  AOI22_X1 U14416 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U14417 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12724) );
  NAND2_X1 U14418 ( .A1(n12725), .A2(n12724), .ZN(n12736) );
  INV_X1 U14419 ( .A(n12726), .ZN(n12728) );
  OAI22_X1 U14420 ( .A1(n12729), .A2(n12728), .B1(n12727), .B2(n12866), .ZN(
        n12735) );
  INV_X1 U14421 ( .A(n12730), .ZN(n12732) );
  OAI22_X1 U14422 ( .A1(n12733), .A2(n12873), .B1(n12732), .B2(n12731), .ZN(
        n12734) );
  NOR4_X1 U14423 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n17429) );
  AOI22_X1 U14424 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U14425 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U14426 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U14427 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U14428 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12747) );
  AOI22_X1 U14429 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U14430 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11878), .B1(
        n11211), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U14431 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U14432 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12742) );
  NAND4_X1 U14433 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12746) );
  NOR2_X1 U14434 ( .A1(n12747), .A2(n12746), .ZN(n17434) );
  OR2_X1 U14435 ( .A1(n17429), .A2(n17434), .ZN(n12758) );
  AOI22_X1 U14436 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U14437 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U14438 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11220), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U14439 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U14440 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12757) );
  AOI22_X1 U14441 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U14442 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11878), .B1(
        n11211), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U14443 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U14444 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12752) );
  NAND4_X1 U14445 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12756) );
  NOR2_X1 U14446 ( .A1(n12757), .A2(n12756), .ZN(n17443) );
  NOR2_X1 U14447 ( .A1(n12758), .A2(n17443), .ZN(n17422) );
  AND2_X1 U14448 ( .A1(n17424), .A2(n17422), .ZN(n12769) );
  AOI22_X1 U14449 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U14450 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U14451 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11220), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U14452 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12759) );
  NAND4_X1 U14453 ( .A1(n12762), .A2(n12761), .A3(n12760), .A4(n12759), .ZN(
        n12768) );
  AOI22_X1 U14454 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U14455 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11878), .B1(
        n11211), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U14456 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11589), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U14457 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12763) );
  NAND4_X1 U14458 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12767) );
  OR2_X1 U14459 ( .A1(n12768), .A2(n12767), .ZN(n16388) );
  AND2_X1 U14460 ( .A1(n12769), .A2(n16388), .ZN(n17415) );
  AOI22_X1 U14461 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U14462 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n11220), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U14463 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U14464 ( .A1(n11870), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12770) );
  NAND4_X1 U14465 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12779) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11878), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U14467 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U14468 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U14469 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12774) );
  NAND4_X1 U14470 ( .A1(n12777), .A2(n12776), .A3(n12775), .A4(n12774), .ZN(
        n12778) );
  NOR2_X1 U14471 ( .A1(n12779), .A2(n12778), .ZN(n17418) );
  INV_X1 U14472 ( .A(n17418), .ZN(n12780) );
  AND2_X1 U14473 ( .A1(n17415), .A2(n12780), .ZN(n17404) );
  AND2_X1 U14474 ( .A1(n17405), .A2(n17404), .ZN(n12781) );
  AND2_X1 U14475 ( .A1(n12781), .A2(n16374), .ZN(n12782) );
  NAND2_X1 U14476 ( .A1(n16367), .A2(n12782), .ZN(n17400) );
  AOI22_X1 U14477 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12726), .B1(
        n11206), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U14478 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12730), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U14479 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11871), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U14480 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11567), .B1(
        n11873), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12784) );
  NAND4_X1 U14481 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12794) );
  AOI22_X1 U14482 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11607), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U14483 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11878), .B1(
        n11211), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U14484 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12788), .B1(
        n11590), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11591), .B1(
        n11592), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12789) );
  NAND4_X1 U14486 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12793) );
  NOR2_X1 U14487 ( .A1(n12794), .A2(n12793), .ZN(n12815) );
  AOI22_X1 U14488 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U14489 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U14490 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12803) );
  INV_X1 U14491 ( .A(n12968), .ZN(n12958) );
  NAND2_X1 U14492 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12800) );
  INV_X1 U14493 ( .A(n12797), .ZN(n12799) );
  NAND2_X1 U14494 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12798) );
  NAND2_X1 U14495 ( .A1(n12799), .A2(n12798), .ZN(n12967) );
  OAI211_X1 U14496 ( .C1(n12958), .C2(n14745), .A(n12800), .B(n12967), .ZN(
        n12801) );
  INV_X1 U14497 ( .A(n12801), .ZN(n12802) );
  NAND4_X1 U14498 ( .A1(n12805), .A2(n12804), .A3(n12803), .A4(n12802), .ZN(
        n12814) );
  AOI22_X1 U14499 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U14500 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U14501 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12810) );
  INV_X1 U14502 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U14503 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12806) );
  INV_X1 U14504 ( .A(n12967), .ZN(n12930) );
  OAI211_X1 U14505 ( .C1(n12958), .C2(n12807), .A(n12806), .B(n12930), .ZN(
        n12808) );
  INV_X1 U14506 ( .A(n12808), .ZN(n12809) );
  NAND4_X1 U14507 ( .A1(n12812), .A2(n12811), .A3(n12810), .A4(n12809), .ZN(
        n12813) );
  NAND2_X1 U14508 ( .A1(n12814), .A2(n12813), .ZN(n12816) );
  XNOR2_X1 U14509 ( .A(n12815), .B(n12816), .ZN(n17401) );
  INV_X1 U14510 ( .A(n12815), .ZN(n12818) );
  INV_X1 U14511 ( .A(n12816), .ZN(n12817) );
  NAND2_X1 U14512 ( .A1(n12818), .A2(n12817), .ZN(n12838) );
  AOI22_X1 U14513 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U14514 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U14515 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U14516 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12822) );
  OAI211_X1 U14517 ( .C1(n12958), .C2(n12823), .A(n12822), .B(n12967), .ZN(
        n12824) );
  INV_X1 U14518 ( .A(n12824), .ZN(n12825) );
  NAND4_X1 U14519 ( .A1(n12828), .A2(n12827), .A3(n12826), .A4(n12825), .ZN(
        n12837) );
  AOI22_X1 U14520 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U14521 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U14522 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U14523 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12829) );
  OAI211_X1 U14524 ( .C1(n12958), .C2(n12830), .A(n12829), .B(n12930), .ZN(
        n12831) );
  INV_X1 U14525 ( .A(n12831), .ZN(n12832) );
  NAND4_X1 U14526 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12836) );
  NAND2_X1 U14527 ( .A1(n12837), .A2(n12836), .ZN(n12858) );
  NOR2_X1 U14528 ( .A1(n12838), .A2(n12858), .ZN(n12840) );
  NAND2_X1 U14529 ( .A1(n12881), .A2(n12820), .ZN(n12839) );
  AOI22_X1 U14530 ( .A1(n12840), .A2(n12954), .B1(n12839), .B2(n12858), .ZN(
        n17396) );
  INV_X1 U14531 ( .A(n12840), .ZN(n12857) );
  AOI22_X1 U14532 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U14533 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U14534 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12845) );
  NAND2_X1 U14535 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12841) );
  OAI211_X1 U14536 ( .C1(n12958), .C2(n12842), .A(n12841), .B(n12967), .ZN(
        n12843) );
  INV_X1 U14537 ( .A(n12843), .ZN(n12844) );
  NAND4_X1 U14538 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12856) );
  AOI22_X1 U14539 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U14540 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U14541 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12852) );
  INV_X1 U14542 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U14543 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12848) );
  OAI211_X1 U14544 ( .C1(n12958), .C2(n12849), .A(n12848), .B(n12930), .ZN(
        n12850) );
  INV_X1 U14545 ( .A(n12850), .ZN(n12851) );
  NAND4_X1 U14546 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12855) );
  NAND2_X1 U14547 ( .A1(n12856), .A2(n12855), .ZN(n12862) );
  NAND2_X1 U14548 ( .A1(n12857), .A2(n12862), .ZN(n12860) );
  NOR2_X1 U14549 ( .A1(n12858), .A2(n12862), .ZN(n12859) );
  NAND2_X1 U14550 ( .A1(n12820), .A2(n12859), .ZN(n12864) );
  NAND3_X1 U14551 ( .A1(n12860), .A2(n12881), .A3(n12864), .ZN(n12863) );
  INV_X1 U14552 ( .A(n12863), .ZN(n12861) );
  NOR2_X1 U14553 ( .A1(n12954), .A2(n12862), .ZN(n17390) );
  INV_X1 U14554 ( .A(n12864), .ZN(n12882) );
  AOI22_X1 U14555 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U14556 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U14557 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12869) );
  NAND2_X1 U14558 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12865) );
  OAI211_X1 U14559 ( .C1(n12958), .C2(n12866), .A(n12865), .B(n12967), .ZN(
        n12867) );
  INV_X1 U14560 ( .A(n12867), .ZN(n12868) );
  NAND4_X1 U14561 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12880) );
  AOI22_X1 U14562 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U14563 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U14564 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12876) );
  NAND2_X1 U14565 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12872) );
  OAI211_X1 U14566 ( .C1(n12958), .C2(n12873), .A(n12872), .B(n12930), .ZN(
        n12874) );
  INV_X1 U14567 ( .A(n12874), .ZN(n12875) );
  NAND4_X1 U14568 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        n12879) );
  AND2_X1 U14569 ( .A1(n12880), .A2(n12879), .ZN(n12883) );
  NAND2_X1 U14570 ( .A1(n12882), .A2(n12883), .ZN(n12906) );
  OAI211_X1 U14571 ( .C1(n12882), .C2(n12883), .A(n12881), .B(n12906), .ZN(
        n12886) );
  INV_X1 U14572 ( .A(n12883), .ZN(n12884) );
  NOR2_X1 U14573 ( .A1(n12954), .A2(n12884), .ZN(n17382) );
  INV_X1 U14574 ( .A(n12886), .ZN(n12887) );
  AOI22_X1 U14575 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U14576 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U14577 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U14578 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12889) );
  OAI211_X1 U14579 ( .C1(n12958), .C2(n12890), .A(n12889), .B(n12967), .ZN(
        n12891) );
  INV_X1 U14580 ( .A(n12891), .ZN(n12892) );
  NAND4_X1 U14581 ( .A1(n12895), .A2(n12894), .A3(n12893), .A4(n12892), .ZN(
        n12904) );
  AOI22_X1 U14582 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U14583 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11213), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U14584 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12900) );
  INV_X1 U14585 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12897) );
  NAND2_X1 U14586 ( .A1(n12937), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12896) );
  OAI211_X1 U14587 ( .C1(n12958), .C2(n12897), .A(n12896), .B(n12930), .ZN(
        n12898) );
  INV_X1 U14588 ( .A(n12898), .ZN(n12899) );
  NAND4_X1 U14589 ( .A1(n12902), .A2(n12901), .A3(n12900), .A4(n12899), .ZN(
        n12903) );
  NAND2_X1 U14590 ( .A1(n12904), .A2(n12903), .ZN(n12907) );
  NOR2_X1 U14591 ( .A1(n12906), .A2(n12907), .ZN(n17369) );
  AOI211_X1 U14592 ( .C1(n12907), .C2(n12906), .A(n12905), .B(n17369), .ZN(
        n12910) );
  INV_X1 U14593 ( .A(n12907), .ZN(n12908) );
  NAND2_X1 U14594 ( .A1(n12819), .A2(n12908), .ZN(n17377) );
  NAND2_X1 U14595 ( .A1(n17368), .A2(n17377), .ZN(n12929) );
  NAND2_X1 U14596 ( .A1(n12912), .A2(n12911), .ZN(n17374) );
  AOI22_X1 U14597 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U14598 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U14599 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U14600 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12913) );
  OAI211_X1 U14601 ( .C1(n12958), .C2(n11621), .A(n12913), .B(n12967), .ZN(
        n12914) );
  INV_X1 U14602 ( .A(n12914), .ZN(n12915) );
  NAND4_X1 U14603 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12927) );
  AOI22_X1 U14604 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11207), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U14605 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U14606 ( .A1(n12969), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12923) );
  INV_X1 U14607 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U14608 ( .A1(n11213), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12919) );
  OAI211_X1 U14609 ( .C1(n12958), .C2(n12920), .A(n12919), .B(n12930), .ZN(
        n12921) );
  INV_X1 U14610 ( .A(n12921), .ZN(n12922) );
  NAND4_X1 U14611 ( .A1(n12925), .A2(n12924), .A3(n12923), .A4(n12922), .ZN(
        n12926) );
  NAND2_X1 U14612 ( .A1(n12927), .A2(n12926), .ZN(n17370) );
  OAI21_X1 U14613 ( .B1(n12958), .B2(n12931), .A(n12930), .ZN(n12936) );
  OAI22_X1 U14614 ( .A1(n12934), .A2(n12933), .B1(n11166), .B2(n12932), .ZN(
        n12935) );
  AOI211_X1 U14615 ( .C1(n12937), .C2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12936), .B(n12935), .ZN(n12941) );
  AOI22_X1 U14616 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U14617 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12939) );
  NAND3_X1 U14618 ( .A1(n12941), .A2(n12940), .A3(n12939), .ZN(n12952) );
  OAI21_X1 U14619 ( .B1(n12958), .B2(n12942), .A(n12967), .ZN(n12947) );
  OAI22_X1 U14620 ( .A1(n15311), .A2(n12945), .B1(n12944), .B2(n12943), .ZN(
        n12946) );
  AOI211_X1 U14621 ( .C1(n11213), .C2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n12947), .B(n12946), .ZN(n12950) );
  AOI22_X1 U14622 ( .A1(n11207), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U14623 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12970), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12948) );
  NAND3_X1 U14624 ( .A1(n12950), .A2(n12949), .A3(n12948), .ZN(n12951) );
  AND2_X1 U14625 ( .A1(n12952), .A2(n12951), .ZN(n12953) );
  NAND3_X1 U14626 ( .A1(n17369), .A2(n12928), .A3(n12954), .ZN(n17364) );
  INV_X1 U14627 ( .A(n12955), .ZN(n12956) );
  OAI21_X1 U14628 ( .B1(n12958), .B2(n12957), .A(n12967), .ZN(n12961) );
  INV_X1 U14629 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16296) );
  INV_X1 U14630 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12959) );
  OAI22_X1 U14631 ( .A1(n11536), .A2(n16296), .B1(n15311), .B2(n12959), .ZN(
        n12960) );
  AOI211_X1 U14632 ( .C1(n11213), .C2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12961), .B(n12960), .ZN(n12964) );
  AOI22_X1 U14633 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U14634 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12962) );
  NAND3_X1 U14635 ( .A1(n12964), .A2(n12963), .A3(n12962), .ZN(n12976) );
  INV_X1 U14636 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12965) );
  NOR2_X1 U14637 ( .A1(n11166), .A2(n12965), .ZN(n12966) );
  AOI211_X1 U14638 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n12968), .A(
        n12967), .B(n12966), .ZN(n12974) );
  AOI22_X1 U14639 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11219), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U14640 ( .A1(n12970), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12969), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U14641 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12937), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12971) );
  NAND4_X1 U14642 ( .A1(n12974), .A2(n12973), .A3(n12972), .A4(n12971), .ZN(
        n12975) );
  XNOR2_X1 U14643 ( .A(n12977), .B(n11486), .ZN(n13008) );
  NAND2_X1 U14644 ( .A1(n15341), .A2(n15472), .ZN(n15291) );
  NAND2_X1 U14645 ( .A1(n15291), .A2(n12978), .ZN(n12979) );
  NAND2_X1 U14646 ( .A1(n12979), .A2(n19511), .ZN(n12981) );
  AND2_X1 U14647 ( .A1(n12573), .A2(n19531), .ZN(n15333) );
  NAND2_X1 U14648 ( .A1(n18168), .A2(n15333), .ZN(n12980) );
  NAND2_X1 U14649 ( .A1(n13008), .A2(n20461), .ZN(n13005) );
  INV_X1 U14650 ( .A(n12982), .ZN(n12985) );
  INV_X1 U14651 ( .A(n12983), .ZN(n12984) );
  NAND2_X1 U14652 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  NAND2_X1 U14653 ( .A1(n20513), .A2(n15513), .ZN(n20515) );
  AND2_X1 U14654 ( .A1(n20513), .A2(n12988), .ZN(n20008) );
  NOR4_X1 U14655 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12992) );
  NOR4_X1 U14656 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12991) );
  NOR4_X1 U14657 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12990) );
  NOR4_X1 U14658 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12989) );
  NAND4_X1 U14659 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        n12997) );
  NOR4_X1 U14660 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12995) );
  NOR4_X1 U14661 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12994) );
  NOR4_X1 U14662 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12993) );
  INV_X1 U14663 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n18274) );
  NAND4_X1 U14664 ( .A1(n12995), .A2(n12994), .A3(n12993), .A4(n18274), .ZN(
        n12996) );
  NAND2_X1 U14665 ( .A1(n20513), .A2(n12998), .ZN(n20009) );
  AOI22_X1 U14666 ( .A1(n15508), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n14661), .ZN(n20014) );
  INV_X1 U14667 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14685) );
  OAI22_X1 U14668 ( .A1(n20009), .A2(n20014), .B1(n14685), .B2(n20513), .ZN(
        n13001) );
  NAND2_X1 U14669 ( .A1(n20008), .A2(n14661), .ZN(n17462) );
  INV_X1 U14670 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n12999) );
  NOR2_X1 U14671 ( .A1(n17462), .A2(n12999), .ZN(n13000) );
  AOI211_X1 U14672 ( .C1(n20005), .C2(BUF1_REG_30__SCAN_IN), .A(n13001), .B(
        n13000), .ZN(n13002) );
  NAND2_X1 U14673 ( .A1(n13005), .A2(n13004), .ZN(P2_U2889) );
  INV_X1 U14674 ( .A(n15472), .ZN(n15346) );
  NAND2_X1 U14675 ( .A1(n15346), .A2(n15282), .ZN(n15289) );
  NAND2_X1 U14676 ( .A1(n15289), .A2(n15276), .ZN(n13006) );
  NAND2_X1 U14677 ( .A1(n13008), .A2(n17419), .ZN(n13012) );
  NAND2_X1 U14678 ( .A1(n17432), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13009) );
  NAND2_X1 U14679 ( .A1(n13012), .A2(n13011), .ZN(P2_U2857) );
  AOI21_X1 U14680 ( .B1(n14207), .B2(n14185), .A(n13013), .ZN(n14178) );
  AOI21_X1 U14681 ( .B1(n11235), .B2(n13017), .A(n13016), .ZN(n14521) );
  NAND2_X1 U14682 ( .A1(n19360), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14186) );
  OAI21_X1 U14683 ( .B1(n18204), .B2(n13017), .A(n14186), .ZN(n13018) );
  AOI21_X1 U14684 ( .B1(n18196), .B2(n14521), .A(n13018), .ZN(n13019) );
  OAI21_X1 U14685 ( .B1(n19457), .B2(n18190), .A(n13019), .ZN(n13020) );
  AOI21_X1 U14686 ( .B1(n14178), .B2(n18198), .A(n13020), .ZN(n13026) );
  XNOR2_X1 U14687 ( .A(n13023), .B(n11499), .ZN(n14176) );
  INV_X1 U14688 ( .A(n14176), .ZN(n13024) );
  NAND2_X1 U14689 ( .A1(n13026), .A2(n13025), .ZN(P2_U2985) );
  NOR2_X4 U14690 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14712) );
  INV_X1 U14691 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13027) );
  NOR2_X4 U14692 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13037) );
  INV_X1 U14693 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U14694 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U14695 ( .A1(n13081), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U14696 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U14697 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13179), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13041) );
  AND2_X2 U14698 ( .A1(n13037), .A2(n14713), .ZN(n13117) );
  AOI22_X1 U14699 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13040) );
  AND2_X4 U14700 ( .A1(n13038), .A2(n14897), .ZN(n13223) );
  AND2_X4 U14701 ( .A1(n14897), .A2(n14713), .ZN(n13105) );
  AOI22_X1 U14702 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U14703 ( .A1(n13081), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U14704 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11224), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U14705 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U14706 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U14707 ( .A1(n13110), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U14708 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11198), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U14709 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U14710 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13179), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U14711 ( .A1(n14249), .A2(n13150), .ZN(n13080) );
  AOI22_X1 U14712 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U14713 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11208), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U14714 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U14715 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U14716 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U14717 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U14718 ( .A1(n13081), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13126), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U14719 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U14720 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U14721 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U14722 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U14723 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11209), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U14724 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U14725 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13081), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U14726 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U14727 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U14728 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11226), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U14729 ( .A1(n13110), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U14730 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11199), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13076) );
  AND2_X2 U14731 ( .A1(n13170), .A2(n14410), .ZN(n14239) );
  NAND2_X1 U14732 ( .A1(n13080), .A2(n13161), .ZN(n13099) );
  AOI22_X1 U14733 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U14734 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U14735 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U14736 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U14737 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U14738 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13087) );
  INV_X1 U14739 ( .A(n13092), .ZN(n13203) );
  NAND2_X1 U14740 ( .A1(n13153), .A2(n13448), .ZN(n13096) );
  NAND2_X1 U14741 ( .A1(n14411), .A2(n14410), .ZN(n13094) );
  NAND2_X1 U14742 ( .A1(n14966), .A2(n13094), .ZN(n13095) );
  NAND2_X1 U14743 ( .A1(n13096), .A2(n13095), .ZN(n13098) );
  INV_X1 U14744 ( .A(n13151), .ZN(n13097) );
  NAND2_X1 U14745 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13103) );
  NAND2_X1 U14746 ( .A1(n13081), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13102) );
  NAND2_X1 U14747 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13101) );
  NAND2_X1 U14748 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13100) );
  NAND2_X1 U14749 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13109) );
  BUF_X4 U14750 ( .A(n13104), .Z(n13945) );
  NAND2_X1 U14751 ( .A1(n13945), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13108) );
  NAND2_X1 U14752 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13107) );
  NAND2_X1 U14753 ( .A1(n13105), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13106) );
  NAND2_X1 U14754 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13113) );
  NAND2_X1 U14755 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13112) );
  NAND2_X1 U14756 ( .A1(n13110), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13111) );
  NAND2_X1 U14757 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13121) );
  NAND2_X1 U14758 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13120) );
  NAND2_X1 U14759 ( .A1(n13116), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13119) );
  NAND2_X1 U14760 ( .A1(n13117), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13118) );
  NAND4_X4 U14761 ( .A1(n13125), .A2(n13124), .A3(n13123), .A4(n13122), .ZN(
        n15025) );
  NAND2_X1 U14762 ( .A1(n13081), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13130) );
  NAND2_X1 U14763 ( .A1(n13126), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13129) );
  NAND2_X1 U14764 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13128) );
  NAND2_X1 U14765 ( .A1(n13945), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13127) );
  NAND2_X1 U14766 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13135) );
  NAND2_X1 U14767 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13134) );
  NAND2_X1 U14768 ( .A1(n13116), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13133) );
  NAND2_X1 U14769 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13132) );
  NAND2_X1 U14770 ( .A1(n13136), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13141) );
  NAND2_X1 U14771 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13140) );
  NAND2_X1 U14772 ( .A1(n13137), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13139) );
  NAND2_X1 U14773 ( .A1(n13105), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13138) );
  NAND2_X1 U14774 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13145) );
  NAND2_X1 U14775 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13144) );
  NAND2_X1 U14776 ( .A1(n13117), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13143) );
  NAND2_X1 U14777 ( .A1(n13110), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13142) );
  NAND2_X1 U14778 ( .A1(n14357), .A2(n15033), .ZN(n13152) );
  XNOR2_X1 U14779 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n14551) );
  NAND3_X1 U14780 ( .A1(n17198), .A2(n13166), .A3(n14999), .ZN(n14707) );
  NAND2_X1 U14781 ( .A1(n14999), .A2(n14411), .ZN(n13154) );
  INV_X1 U14782 ( .A(n13160), .ZN(n13155) );
  NAND2_X1 U14783 ( .A1(n13155), .A2(n13211), .ZN(n13158) );
  INV_X1 U14784 ( .A(n14239), .ZN(n13159) );
  NAND2_X1 U14785 ( .A1(n13160), .A2(n13159), .ZN(n14241) );
  NAND2_X1 U14786 ( .A1(n14241), .A2(n13161), .ZN(n13168) );
  INV_X1 U14787 ( .A(n17198), .ZN(n14361) );
  MUX2_X1 U14788 ( .A(n13165), .B(n14377), .S(n15025), .Z(n13163) );
  NAND2_X1 U14789 ( .A1(n20865), .A2(n22396), .ZN(n14019) );
  MUX2_X1 U14790 ( .A(n14019), .B(n22390), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n13164) );
  INV_X1 U14791 ( .A(n13165), .ZN(n13177) );
  INV_X1 U14792 ( .A(n13166), .ZN(n15017) );
  AND3_X1 U14793 ( .A1(n13159), .A2(n15017), .A3(n13167), .ZN(n13176) );
  OR2_X1 U14794 ( .A1(n13168), .A2(n15026), .ZN(n13175) );
  INV_X1 U14795 ( .A(n13169), .ZN(n13173) );
  NAND2_X1 U14796 ( .A1(n17198), .A2(n14977), .ZN(n14370) );
  NAND2_X1 U14797 ( .A1(n15025), .A2(n13153), .ZN(n13171) );
  NAND4_X1 U14798 ( .A1(n14370), .A2(n20865), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n13171), .ZN(n13172) );
  INV_X1 U14799 ( .A(n13215), .ZN(n13178) );
  AOI22_X1 U14800 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13183) );
  INV_X1 U14801 ( .A(n13223), .ZN(n13196) );
  AOI22_X1 U14803 ( .A1(n13191), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U14804 ( .A1(n13179), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13180) );
  NAND4_X1 U14805 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13189) );
  AOI22_X1 U14806 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13081), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U14807 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U14808 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U14809 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13184) );
  NAND4_X1 U14810 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13188) );
  INV_X1 U14811 ( .A(n13406), .ZN(n13245) );
  AOI22_X1 U14812 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U14813 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13086), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U14814 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13193) );
  INV_X1 U14815 ( .A(n13863), .ZN(n13940) );
  AOI22_X1 U14816 ( .A1(n13940), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13192) );
  NAND4_X1 U14817 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13202) );
  AOI22_X1 U14818 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U14819 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U14820 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U14821 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13197) );
  NAND4_X1 U14822 ( .A1(n13200), .A2(n13199), .A3(n13198), .A4(n13197), .ZN(
        n13201) );
  XNOR2_X1 U14823 ( .A(n13245), .B(n13237), .ZN(n13205) );
  NAND2_X1 U14824 ( .A1(n13205), .A2(n13256), .ZN(n13206) );
  INV_X1 U14825 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13210) );
  AOI21_X1 U14826 ( .B1(n13204), .B2(n13406), .A(n22396), .ZN(n13209) );
  NAND2_X1 U14827 ( .A1(n15130), .A2(n13237), .ZN(n13208) );
  OAI211_X1 U14828 ( .C1(n13489), .C2(n13210), .A(n13209), .B(n13208), .ZN(
        n13254) );
  NAND2_X1 U14829 ( .A1(n14410), .A2(n11221), .ZN(n13403) );
  INV_X1 U14830 ( .A(n13237), .ZN(n13212) );
  NAND2_X1 U14831 ( .A1(n13211), .A2(n13212), .ZN(n13213) );
  NAND2_X1 U14832 ( .A1(n15130), .A2(n13167), .ZN(n13291) );
  AND2_X1 U14833 ( .A1(n13213), .A2(n13291), .ZN(n13214) );
  XNOR2_X1 U14834 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22473) );
  OR2_X1 U14835 ( .A1(n22390), .A2(n22475), .ZN(n13259) );
  OAI21_X1 U14836 ( .B1(n14019), .B2(n22473), .A(n13259), .ZN(n13218) );
  INV_X1 U14837 ( .A(n13218), .ZN(n13219) );
  AOI22_X1 U14838 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U14839 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U14840 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U14841 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13224) );
  NAND4_X1 U14842 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13233) );
  AOI22_X1 U14843 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U14844 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U14845 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13229) );
  AOI22_X1 U14846 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13228) );
  NAND4_X1 U14847 ( .A1(n13231), .A2(n13230), .A3(n13229), .A4(n13228), .ZN(
        n13232) );
  NAND2_X1 U14848 ( .A1(n13256), .A2(n13246), .ZN(n13234) );
  INV_X1 U14849 ( .A(n13252), .ZN(n13236) );
  INV_X1 U14850 ( .A(n13403), .ZN(n13235) );
  NAND2_X1 U14851 ( .A1(n13236), .A2(n13235), .ZN(n13240) );
  NAND2_X1 U14852 ( .A1(n13246), .A2(n13237), .ZN(n13316) );
  OAI211_X1 U14853 ( .C1(n13246), .C2(n13237), .A(n13211), .B(n13316), .ZN(
        n13238) );
  AND3_X1 U14854 ( .A1(n13238), .A2(n14364), .A3(n11183), .ZN(n13239) );
  INV_X1 U14855 ( .A(n13241), .ZN(n13243) );
  NAND2_X1 U14856 ( .A1(n13243), .A2(n13242), .ZN(n13244) );
  INV_X1 U14857 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n22158) );
  INV_X1 U14858 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U14859 ( .A1(n13256), .A2(n13245), .ZN(n13249) );
  INV_X1 U14860 ( .A(n13273), .ZN(n13247) );
  NAND2_X1 U14861 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  OAI211_X1 U14862 ( .C1(n13489), .C2(n13250), .A(n13249), .B(n13248), .ZN(
        n13251) );
  NAND2_X1 U14863 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND2_X1 U14864 ( .A1(n13255), .A2(n13254), .ZN(n13257) );
  NAND2_X1 U14865 ( .A1(n13256), .A2(n13406), .ZN(n13404) );
  INV_X1 U14866 ( .A(n13259), .ZN(n13261) );
  NAND2_X1 U14867 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13265) );
  NAND2_X1 U14868 ( .A1(n18135), .A2(n13265), .ZN(n13267) );
  NAND2_X1 U14869 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22505) );
  INV_X1 U14870 ( .A(n22505), .ZN(n13266) );
  NAND2_X1 U14871 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13266), .ZN(
        n15212) );
  NAND2_X1 U14872 ( .A1(n13267), .A2(n15212), .ZN(n15522) );
  OAI22_X1 U14873 ( .A1(n14019), .A2(n15522), .B1(n22390), .B2(n18135), .ZN(
        n13268) );
  INV_X1 U14874 ( .A(n13268), .ZN(n13269) );
  AOI22_X1 U14875 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U14876 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13276) );
  AOI22_X1 U14877 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13275) );
  NAND4_X1 U14878 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13284) );
  AOI22_X1 U14879 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U14880 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U14881 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U14882 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13279) );
  NAND4_X1 U14883 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  AOI22_X1 U14884 ( .A1(n13481), .A2(n13290), .B1(n13468), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13285) );
  INV_X1 U14885 ( .A(n13286), .ZN(n13288) );
  NAND2_X1 U14886 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  NAND2_X1 U14887 ( .A1(n13323), .A2(n13289), .ZN(n14902) );
  INV_X1 U14888 ( .A(n13290), .ZN(n13315) );
  XNOR2_X1 U14889 ( .A(n13316), .B(n13315), .ZN(n13293) );
  INV_X1 U14890 ( .A(n13291), .ZN(n13292) );
  AOI21_X1 U14891 ( .B1(n13293), .B2(n13211), .A(n13292), .ZN(n13294) );
  OAI21_X1 U14892 ( .B1(n14902), .B2(n13403), .A(n13294), .ZN(n14939) );
  NAND2_X1 U14893 ( .A1(n14940), .A2(n14939), .ZN(n22149) );
  NAND2_X1 U14894 ( .A1(n22149), .A2(n13295), .ZN(n13321) );
  INV_X1 U14895 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n22179) );
  INV_X1 U14896 ( .A(n15212), .ZN(n13297) );
  NAND2_X1 U14897 ( .A1(n13297), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15005) );
  NAND2_X1 U14898 ( .A1(n15212), .A2(n15681), .ZN(n13298) );
  INV_X1 U14899 ( .A(n14019), .ZN(n13300) );
  INV_X1 U14900 ( .A(n22390), .ZN(n13299) );
  AOI22_X1 U14901 ( .A1(n15604), .A2(n13300), .B1(n13299), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U14902 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U14903 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U14904 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U14905 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13303) );
  NAND4_X1 U14906 ( .A1(n13306), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13312) );
  AOI22_X1 U14907 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U14908 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U14909 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U14910 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13307) );
  NAND4_X1 U14911 ( .A1(n13310), .A2(n13309), .A3(n13308), .A4(n13307), .ZN(
        n13311) );
  AOI22_X1 U14912 ( .A1(n13481), .A2(n13338), .B1(n13468), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13313) );
  NAND2_X1 U14913 ( .A1(n13528), .A2(n13235), .ZN(n13320) );
  NAND2_X1 U14914 ( .A1(n13316), .A2(n13315), .ZN(n13339) );
  INV_X1 U14915 ( .A(n13338), .ZN(n13317) );
  XNOR2_X1 U14916 ( .A(n13339), .B(n13317), .ZN(n13318) );
  NAND2_X1 U14917 ( .A1(n13318), .A2(n13211), .ZN(n13319) );
  NAND2_X1 U14918 ( .A1(n13320), .A2(n13319), .ZN(n15170) );
  NAND2_X1 U14919 ( .A1(n13321), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13322) );
  AOI22_X1 U14920 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13816), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U14921 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13945), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U14922 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13327) );
  AOI22_X1 U14923 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13326) );
  NAND4_X1 U14924 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n13335) );
  AOI22_X1 U14925 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U14926 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11227), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13331) );
  AOI22_X1 U14927 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13330) );
  NAND4_X1 U14928 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        n13334) );
  NAND2_X1 U14929 ( .A1(n13481), .A2(n13359), .ZN(n13337) );
  NAND2_X1 U14930 ( .A1(n13468), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13336) );
  NAND2_X1 U14931 ( .A1(n13337), .A2(n13336), .ZN(n13346) );
  XNOR2_X1 U14932 ( .A(n13345), .B(n13346), .ZN(n13548) );
  NAND2_X1 U14933 ( .A1(n13548), .A2(n13235), .ZN(n13342) );
  NAND2_X1 U14934 ( .A1(n13339), .A2(n13338), .ZN(n13361) );
  XNOR2_X1 U14935 ( .A(n13361), .B(n13359), .ZN(n13340) );
  NAND2_X1 U14936 ( .A1(n13340), .A2(n13211), .ZN(n13341) );
  NAND2_X1 U14937 ( .A1(n13342), .A2(n13341), .ZN(n13343) );
  INV_X1 U14938 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n22167) );
  XNOR2_X1 U14939 ( .A(n13343), .B(n22167), .ZN(n20832) );
  NAND2_X1 U14940 ( .A1(n13343), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13344) );
  AOI22_X1 U14941 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U14942 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U14943 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U14944 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13347) );
  NAND4_X1 U14945 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13356) );
  AOI22_X1 U14946 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13354) );
  AOI22_X1 U14947 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U14948 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13352) );
  AOI22_X1 U14949 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13351) );
  NAND4_X1 U14950 ( .A1(n13354), .A2(n13353), .A3(n13352), .A4(n13351), .ZN(
        n13355) );
  NAND2_X1 U14951 ( .A1(n13481), .A2(n13384), .ZN(n13358) );
  NAND2_X1 U14952 ( .A1(n13468), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13357) );
  NAND2_X1 U14953 ( .A1(n13358), .A2(n13357), .ZN(n13368) );
  NAND2_X1 U14954 ( .A1(n13558), .A2(n13235), .ZN(n13364) );
  INV_X1 U14955 ( .A(n13359), .ZN(n13360) );
  OR2_X1 U14956 ( .A1(n13361), .A2(n13360), .ZN(n13383) );
  XNOR2_X1 U14957 ( .A(n13383), .B(n13384), .ZN(n13362) );
  NAND2_X1 U14958 ( .A1(n13362), .A2(n13211), .ZN(n13363) );
  INV_X1 U14959 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n22205) );
  XNOR2_X1 U14960 ( .A(n13365), .B(n22205), .ZN(n20838) );
  NAND2_X1 U14961 ( .A1(n13365), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13366) );
  NAND2_X1 U14962 ( .A1(n20837), .A2(n13366), .ZN(n20845) );
  AOI22_X1 U14963 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U14964 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U14965 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U14966 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13369) );
  NAND4_X1 U14967 ( .A1(n13372), .A2(n13371), .A3(n13370), .A4(n13369), .ZN(
        n13378) );
  AOI22_X1 U14968 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U14969 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13375) );
  AOI22_X1 U14970 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U14971 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13373) );
  NAND4_X1 U14972 ( .A1(n13376), .A2(n13375), .A3(n13374), .A4(n13373), .ZN(
        n13377) );
  AOI22_X1 U14973 ( .A1(n13481), .A2(n13396), .B1(n13468), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U14974 ( .A1(n13382), .A2(n13381), .ZN(n13559) );
  INV_X1 U14975 ( .A(n13383), .ZN(n13385) );
  NAND2_X1 U14976 ( .A1(n13385), .A2(n13384), .ZN(n13395) );
  XNOR2_X1 U14977 ( .A(n13395), .B(n13396), .ZN(n13386) );
  NAND2_X1 U14978 ( .A1(n13386), .A2(n13211), .ZN(n13387) );
  NAND2_X1 U14979 ( .A1(n13388), .A2(n13387), .ZN(n13389) );
  INV_X1 U14980 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n22204) );
  XNOR2_X1 U14981 ( .A(n13389), .B(n22204), .ZN(n20844) );
  NAND2_X1 U14982 ( .A1(n20845), .A2(n20844), .ZN(n20843) );
  NAND2_X1 U14983 ( .A1(n13389), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13390) );
  NAND2_X1 U14984 ( .A1(n13481), .A2(n13406), .ZN(n13392) );
  NAND2_X1 U14985 ( .A1(n13468), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13391) );
  NAND2_X1 U14986 ( .A1(n13392), .A2(n13391), .ZN(n13393) );
  NAND2_X1 U14987 ( .A1(n13572), .A2(n13235), .ZN(n13400) );
  INV_X1 U14988 ( .A(n13395), .ZN(n13397) );
  NAND2_X1 U14989 ( .A1(n13397), .A2(n13396), .ZN(n13408) );
  XNOR2_X1 U14990 ( .A(n13408), .B(n13406), .ZN(n13398) );
  NAND2_X1 U14991 ( .A1(n13398), .A2(n13211), .ZN(n13399) );
  NAND2_X1 U14992 ( .A1(n13400), .A2(n13399), .ZN(n13401) );
  INV_X1 U14993 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n22211) );
  XNOR2_X1 U14994 ( .A(n13401), .B(n22211), .ZN(n20850) );
  NAND2_X1 U14995 ( .A1(n20851), .A2(n20850), .ZN(n20849) );
  NAND2_X1 U14996 ( .A1(n13401), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13402) );
  NOR2_X1 U14997 ( .A1(n13404), .A2(n13403), .ZN(n13405) );
  NAND2_X1 U14998 ( .A1(n13211), .A2(n13406), .ZN(n13407) );
  OR2_X1 U14999 ( .A1(n13408), .A2(n13407), .ZN(n13409) );
  NAND2_X1 U15000 ( .A1(n13412), .A2(n13409), .ZN(n13410) );
  INV_X1 U15001 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n22216) );
  XNOR2_X1 U15002 ( .A(n13410), .B(n22216), .ZN(n16342) );
  NAND2_X1 U15003 ( .A1(n13410), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13411) );
  NAND2_X1 U15004 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16920) );
  INV_X1 U15005 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n22138) );
  NAND2_X1 U15006 ( .A1(n13412), .A2(n22138), .ZN(n13413) );
  NAND2_X1 U15007 ( .A1(n16920), .A2(n13413), .ZN(n16937) );
  INV_X1 U15008 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17182) );
  NAND2_X1 U15009 ( .A1(n13412), .A2(n17182), .ZN(n16936) );
  NAND2_X1 U15010 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U15011 ( .A1(n13412), .A2(n13414), .ZN(n16934) );
  NAND2_X1 U15012 ( .A1(n16936), .A2(n16934), .ZN(n13415) );
  NOR2_X1 U15013 ( .A1(n16937), .A2(n13415), .ZN(n16922) );
  INV_X1 U15014 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U15015 ( .A1(n16955), .A2(n13416), .ZN(n13417) );
  NAND2_X1 U15016 ( .A1(n16922), .A2(n13417), .ZN(n17125) );
  INV_X1 U15017 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17141) );
  NAND2_X1 U15018 ( .A1(n16956), .A2(n17141), .ZN(n17130) );
  NAND2_X1 U15019 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17134) );
  INV_X1 U15020 ( .A(n17134), .ZN(n17140) );
  NAND2_X1 U15021 ( .A1(n17140), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17119) );
  AND2_X1 U15022 ( .A1(n17130), .A2(n17119), .ZN(n13418) );
  NOR2_X1 U15023 ( .A1(n17125), .A2(n13418), .ZN(n13419) );
  NAND2_X1 U15024 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13420) );
  NAND2_X1 U15025 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16900) );
  NAND2_X1 U15026 ( .A1(n16899), .A2(n16900), .ZN(n17126) );
  NAND2_X1 U15027 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16935) );
  INV_X1 U15028 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n22235) );
  INV_X1 U15029 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17177) );
  NAND2_X1 U15030 ( .A1(n22235), .A2(n17177), .ZN(n13421) );
  NAND2_X1 U15031 ( .A1(n16956), .A2(n13421), .ZN(n16932) );
  OAI21_X1 U15032 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n16956), .ZN(n13422) );
  NAND2_X1 U15033 ( .A1(n16918), .A2(n13422), .ZN(n13423) );
  NAND3_X1 U15034 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17058) );
  INV_X1 U15035 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16870) );
  NOR2_X1 U15036 ( .A1(n17058), .A2(n16870), .ZN(n13425) );
  NAND2_X1 U15037 ( .A1(n16869), .A2(n13425), .ZN(n13426) );
  INV_X1 U15038 ( .A(n16869), .ZN(n13429) );
  INV_X1 U15039 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13428) );
  INV_X1 U15040 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13427) );
  INV_X1 U15041 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17095) );
  INV_X1 U15042 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U15043 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16850) );
  AND2_X1 U15044 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17034) );
  NAND2_X1 U15045 ( .A1(n17034), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17012) );
  NAND2_X1 U15046 ( .A1(n13431), .A2(n17012), .ZN(n13433) );
  NAND2_X1 U15047 ( .A1(n16857), .A2(n16955), .ZN(n16831) );
  NOR2_X1 U15048 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16994) );
  NAND2_X1 U15049 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16982) );
  INV_X1 U15050 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16797) );
  INV_X1 U15051 ( .A(n13439), .ZN(n13437) );
  XNOR2_X1 U15052 ( .A(n16955), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13438) );
  INV_X1 U15053 ( .A(n13438), .ZN(n13435) );
  OAI21_X1 U15054 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n16956), .ZN(n13441) );
  AND2_X1 U15055 ( .A1(n13435), .A2(n13441), .ZN(n13436) );
  NAND2_X1 U15056 ( .A1(n13437), .A2(n13436), .ZN(n13446) );
  INV_X1 U15057 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16973) );
  NAND2_X1 U15058 ( .A1(n13412), .A2(n16973), .ZN(n13440) );
  NAND3_X1 U15059 ( .A1(n11175), .A2(n13438), .A3(n13440), .ZN(n13445) );
  INV_X1 U15060 ( .A(n13440), .ZN(n13443) );
  INV_X1 U15061 ( .A(n13441), .ZN(n13442) );
  NAND2_X1 U15062 ( .A1(n11490), .A2(n14716), .ZN(n13444) );
  NAND3_X1 U15063 ( .A1(n13446), .A2(n13445), .A3(n13444), .ZN(n14401) );
  INV_X1 U15064 ( .A(n13447), .ZN(n13450) );
  NAND2_X1 U15065 ( .A1(n13448), .A2(n14977), .ZN(n13449) );
  AND2_X1 U15066 ( .A1(n13448), .A2(n14364), .ZN(n13451) );
  NAND2_X1 U15067 ( .A1(n13161), .A2(n15130), .ZN(n14242) );
  NAND2_X1 U15068 ( .A1(n22390), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22406) );
  NAND2_X1 U15069 ( .A1(n22524), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13474) );
  XNOR2_X1 U15070 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U15071 ( .A1(n13473), .A2(n13471), .ZN(n13453) );
  NAND2_X1 U15072 ( .A1(n22475), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13452) );
  NAND2_X1 U15073 ( .A1(n13453), .A2(n13452), .ZN(n13470) );
  XNOR2_X1 U15074 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U15075 ( .A1(n13470), .A2(n13469), .ZN(n13455) );
  NAND2_X1 U15076 ( .A1(n18135), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13454) );
  NAND2_X1 U15077 ( .A1(n13455), .A2(n13454), .ZN(n13465) );
  XNOR2_X1 U15078 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U15079 ( .A1(n13465), .A2(n13463), .ZN(n13457) );
  NAND2_X1 U15080 ( .A1(n15681), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13456) );
  NAND2_X1 U15081 ( .A1(n13457), .A2(n13456), .ZN(n13462) );
  NAND2_X1 U15082 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18150), .ZN(
        n13461) );
  INV_X1 U15083 ( .A(n14233), .ZN(n13460) );
  NAND2_X1 U15084 ( .A1(n13481), .A2(n13460), .ZN(n13502) );
  OR2_X1 U15085 ( .A1(n13462), .A2(n13461), .ZN(n13467) );
  INV_X1 U15086 ( .A(n13463), .ZN(n13464) );
  XNOR2_X1 U15087 ( .A(n13465), .B(n13464), .ZN(n13466) );
  NOR2_X1 U15088 ( .A1(n13468), .A2(n14232), .ZN(n13496) );
  XOR2_X1 U15089 ( .A(n13470), .B(n13469), .Z(n14229) );
  NAND2_X1 U15090 ( .A1(n14229), .A2(n13481), .ZN(n13487) );
  INV_X1 U15091 ( .A(n13487), .ZN(n13493) );
  AOI21_X1 U15092 ( .B1(n15026), .B2(n14410), .A(n13166), .ZN(n13488) );
  INV_X1 U15093 ( .A(n13488), .ZN(n13492) );
  INV_X1 U15094 ( .A(n13471), .ZN(n13472) );
  XNOR2_X1 U15095 ( .A(n13473), .B(n13472), .ZN(n14230) );
  OAI22_X1 U15096 ( .A1(n22396), .A2(n11183), .B1(n13489), .B2(n14230), .ZN(
        n13480) );
  NOR3_X1 U15097 ( .A1(n11221), .A2(n14230), .A3(n13480), .ZN(n13486) );
  OAI21_X1 U15098 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n22524), .A(
        n13474), .ZN(n13477) );
  INV_X1 U15099 ( .A(n13477), .ZN(n13475) );
  OAI211_X1 U15100 ( .C1(n15130), .C2(n13476), .A(n13488), .B(n13475), .ZN(
        n13479) );
  INV_X1 U15101 ( .A(n13481), .ZN(n13482) );
  OAI21_X1 U15102 ( .B1(n13482), .B2(n13477), .A(n13494), .ZN(n13478) );
  NAND2_X1 U15103 ( .A1(n13479), .A2(n13478), .ZN(n13485) );
  AOI21_X1 U15104 ( .B1(n13481), .B2(n11221), .A(n13480), .ZN(n13484) );
  AOI21_X1 U15105 ( .B1(n13482), .B2(n13235), .A(n14230), .ZN(n13483) );
  OAI22_X1 U15106 ( .A1(n13486), .A2(n13485), .B1(n13484), .B2(n13483), .ZN(
        n13491) );
  OAI211_X1 U15107 ( .C1(n14229), .C2(n13489), .A(n13488), .B(n13487), .ZN(
        n13490) );
  AOI22_X1 U15108 ( .A1(n13493), .A2(n13492), .B1(n13491), .B2(n13490), .ZN(
        n13495) );
  OAI22_X1 U15109 ( .A1(n13496), .A2(n13495), .B1(n14232), .B2(n13494), .ZN(
        n13497) );
  AOI21_X1 U15110 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n22396), .A(
        n13497), .ZN(n13498) );
  INV_X1 U15111 ( .A(n13498), .ZN(n13499) );
  INV_X1 U15112 ( .A(n14428), .ZN(n13503) );
  INV_X1 U15113 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13505) );
  XNOR2_X1 U15114 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15020) );
  AOI21_X1 U15115 ( .B1(n15010), .B2(n15020), .A(n14009), .ZN(n13504) );
  OAI21_X1 U15116 ( .B1(n13519), .B2(n13505), .A(n13504), .ZN(n13506) );
  AOI21_X1 U15117 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13536), .A(
        n13506), .ZN(n13507) );
  NAND2_X1 U15118 ( .A1(n14009), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13527) );
  NAND2_X1 U15119 ( .A1(n13508), .A2(n13527), .ZN(n14936) );
  INV_X1 U15120 ( .A(n14936), .ZN(n13526) );
  NAND2_X1 U15121 ( .A1(n14903), .A2(n13632), .ZN(n13515) );
  INV_X1 U15122 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13512) );
  INV_X1 U15123 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13511) );
  OAI22_X1 U15124 ( .A1(n13519), .A2(n13512), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13511), .ZN(n13513) );
  AOI21_X1 U15125 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13536), .A(
        n13513), .ZN(n13514) );
  NAND2_X1 U15126 ( .A1(n11212), .A2(n14977), .ZN(n13517) );
  NAND2_X1 U15127 ( .A1(n13517), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14844) );
  INV_X1 U15128 ( .A(n13536), .ZN(n13545) );
  NAND2_X1 U15129 ( .A1(n14010), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U15130 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13520) );
  OAI211_X1 U15131 ( .C1(n13545), .C2(n18128), .A(n13521), .B(n13520), .ZN(
        n13522) );
  AOI21_X1 U15132 ( .B1(n11176), .B2(n13632), .A(n13522), .ZN(n13523) );
  OR2_X1 U15133 ( .A1(n14844), .A2(n13523), .ZN(n14845) );
  INV_X1 U15134 ( .A(n13523), .ZN(n14846) );
  OR2_X1 U15135 ( .A1(n14846), .A2(n13982), .ZN(n13524) );
  NAND2_X1 U15136 ( .A1(n14845), .A2(n13524), .ZN(n14884) );
  NAND2_X1 U15137 ( .A1(n14885), .A2(n14884), .ZN(n14935) );
  INV_X1 U15138 ( .A(n14935), .ZN(n13525) );
  NAND2_X1 U15139 ( .A1(n13526), .A2(n13525), .ZN(n14933) );
  NAND2_X1 U15140 ( .A1(n13528), .A2(n13632), .ZN(n13538) );
  INV_X1 U15141 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13534) );
  INV_X1 U15142 ( .A(n13530), .ZN(n13529) );
  INV_X1 U15143 ( .A(n13539), .ZN(n13541) );
  INV_X1 U15144 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13531) );
  NAND2_X1 U15145 ( .A1(n13531), .A2(n13530), .ZN(n13532) );
  NAND2_X1 U15146 ( .A1(n13541), .A2(n13532), .ZN(n15419) );
  AOI22_X1 U15147 ( .A1(n15419), .A2(n15010), .B1(n14009), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13533) );
  OAI21_X1 U15148 ( .B1(n13519), .B2(n13534), .A(n13533), .ZN(n13535) );
  AOI21_X1 U15149 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13536), .A(
        n13535), .ZN(n13537) );
  NAND2_X1 U15150 ( .A1(n15172), .A2(n15173), .ZN(n15252) );
  INV_X1 U15151 ( .A(n15252), .ZN(n13550) );
  INV_X1 U15152 ( .A(n13551), .ZN(n13553) );
  INV_X1 U15153 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13540) );
  NAND2_X1 U15154 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  NAND2_X1 U15155 ( .A1(n13553), .A2(n13542), .ZN(n22260) );
  NAND2_X1 U15156 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13544) );
  NAND2_X1 U15157 ( .A1(n14010), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13543) );
  OAI211_X1 U15158 ( .C1(n13545), .C2(n18150), .A(n13544), .B(n13543), .ZN(
        n13546) );
  MUX2_X1 U15159 ( .A(n22260), .B(n13546), .S(n13982), .Z(n13547) );
  NAND2_X1 U15160 ( .A1(n13550), .A2(n13549), .ZN(n15251) );
  INV_X1 U15161 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n15656) );
  INV_X1 U15162 ( .A(n13560), .ZN(n13555) );
  INV_X1 U15163 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U15164 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  NAND2_X1 U15165 ( .A1(n13555), .A2(n13554), .ZN(n22264) );
  AOI22_X1 U15166 ( .A1(n22264), .A2(n15010), .B1(n14009), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13556) );
  OAI21_X1 U15167 ( .B1(n13519), .B2(n15656), .A(n13556), .ZN(n13557) );
  NAND2_X1 U15168 ( .A1(n13559), .A2(n13632), .ZN(n13565) );
  INV_X1 U15169 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13562) );
  OAI21_X1 U15170 ( .B1(n13560), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13567), .ZN(n22287) );
  AOI22_X1 U15171 ( .A1(n22287), .A2(n13773), .B1(n14009), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13561) );
  OAI21_X1 U15172 ( .B1(n13519), .B2(n13562), .A(n13561), .ZN(n13563) );
  INV_X1 U15173 ( .A(n13563), .ZN(n13564) );
  NAND2_X1 U15174 ( .A1(n15652), .A2(n15659), .ZN(n15658) );
  INV_X1 U15175 ( .A(n15658), .ZN(n13574) );
  INV_X1 U15176 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n15676) );
  NAND2_X1 U15177 ( .A1(n13567), .A2(n13566), .ZN(n13569) );
  INV_X1 U15178 ( .A(n13589), .ZN(n13568) );
  NAND2_X1 U15179 ( .A1(n13569), .A2(n13568), .ZN(n22300) );
  AOI22_X1 U15180 ( .A1(n22300), .A2(n13773), .B1(n14009), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13570) );
  OAI21_X1 U15181 ( .B1(n13519), .B2(n15676), .A(n13570), .ZN(n13571) );
  AOI21_X1 U15182 ( .B1(n13572), .B2(n13632), .A(n13571), .ZN(n15674) );
  INV_X1 U15183 ( .A(n15674), .ZN(n13573) );
  NAND2_X1 U15184 ( .A1(n13574), .A2(n13573), .ZN(n15673) );
  INV_X1 U15185 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n16297) );
  XNOR2_X1 U15186 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13589), .ZN(
        n22306) );
  AOI22_X1 U15187 ( .A1(n13773), .A2(n22306), .B1(n14009), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13575) );
  OAI21_X1 U15188 ( .B1(n13519), .B2(n16297), .A(n13575), .ZN(n13588) );
  AOI22_X1 U15189 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U15190 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U15191 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U15192 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13576) );
  NAND4_X1 U15193 ( .A1(n13579), .A2(n13578), .A3(n13577), .A4(n13576), .ZN(
        n13585) );
  AOI22_X1 U15194 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U15195 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13581) );
  AOI22_X1 U15196 ( .A1(n13940), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13580) );
  NAND4_X1 U15197 ( .A1(n13583), .A2(n13582), .A3(n13581), .A4(n13580), .ZN(
        n13584) );
  NOR2_X1 U15198 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  NOR2_X1 U15199 ( .A1(n13701), .A2(n13586), .ZN(n13587) );
  NOR2_X1 U15200 ( .A1(n13588), .A2(n13587), .ZN(n16262) );
  XOR2_X1 U15201 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13605), .Z(n16382) );
  AOI22_X1 U15202 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U15203 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13592) );
  AOI22_X1 U15204 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13591) );
  AOI22_X1 U15205 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13590) );
  NAND4_X1 U15206 ( .A1(n13593), .A2(n13592), .A3(n13591), .A4(n13590), .ZN(
        n13599) );
  AOI22_X1 U15207 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U15208 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U15209 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U15210 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13594) );
  NAND4_X1 U15211 ( .A1(n13597), .A2(n13596), .A3(n13595), .A4(n13594), .ZN(
        n13598) );
  NOR2_X1 U15212 ( .A1(n13599), .A2(n13598), .ZN(n13601) );
  INV_X1 U15213 ( .A(n14009), .ZN(n13671) );
  INV_X1 U15214 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13600) );
  OAI22_X1 U15215 ( .A1(n13701), .A2(n13601), .B1(n13671), .B2(n13600), .ZN(
        n13603) );
  INV_X1 U15216 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n16339) );
  NOR2_X1 U15217 ( .A1(n13519), .A2(n16339), .ZN(n13602) );
  NOR2_X1 U15218 ( .A1(n13603), .A2(n13602), .ZN(n13604) );
  OAI21_X1 U15219 ( .B1(n16382), .B2(n13982), .A(n13604), .ZN(n16300) );
  XNOR2_X1 U15220 ( .A(n13633), .B(n16965), .ZN(n16964) );
  NAND2_X1 U15221 ( .A1(n16964), .A2(n13773), .ZN(n13620) );
  INV_X1 U15222 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n16361) );
  OAI22_X1 U15223 ( .A1(n13519), .A2(n16361), .B1(n13671), .B2(n16965), .ZN(
        n13618) );
  AOI22_X1 U15224 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U15225 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13607) );
  AOI22_X1 U15226 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13606) );
  NAND4_X1 U15227 ( .A1(n13609), .A2(n13608), .A3(n13607), .A4(n13606), .ZN(
        n13615) );
  AOI22_X1 U15228 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U15229 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U15230 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U15231 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13610) );
  NAND4_X1 U15232 ( .A1(n13613), .A2(n13612), .A3(n13611), .A4(n13610), .ZN(
        n13614) );
  NOR2_X1 U15233 ( .A1(n13615), .A2(n13614), .ZN(n13616) );
  NOR2_X1 U15234 ( .A1(n13701), .A2(n13616), .ZN(n13617) );
  NOR2_X1 U15235 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  NAND2_X1 U15236 ( .A1(n13620), .A2(n13619), .ZN(n16349) );
  AOI22_X1 U15237 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U15238 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U15239 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13622) );
  AOI22_X1 U15240 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13621) );
  NAND4_X1 U15241 ( .A1(n13624), .A2(n13623), .A3(n13622), .A4(n13621), .ZN(
        n13630) );
  AOI22_X1 U15242 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U15243 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13627) );
  AOI22_X1 U15244 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U15245 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13625) );
  NAND4_X1 U15246 ( .A1(n13628), .A2(n13627), .A3(n13626), .A4(n13625), .ZN(
        n13629) );
  OR2_X1 U15247 ( .A1(n13630), .A2(n13629), .ZN(n13631) );
  NAND2_X1 U15248 ( .A1(n13632), .A2(n13631), .ZN(n16704) );
  NOR2_X1 U15249 ( .A1(n13634), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13635) );
  OR2_X1 U15250 ( .A1(n13670), .A2(n13635), .ZN(n22323) );
  INV_X1 U15251 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n16792) );
  INV_X1 U15252 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n22315) );
  OAI22_X1 U15253 ( .A1(n13519), .A2(n16792), .B1(n13671), .B2(n22315), .ZN(
        n13636) );
  AOI21_X1 U15254 ( .B1(n22323), .B2(n13773), .A(n13636), .ZN(n16658) );
  INV_X1 U15255 ( .A(n16658), .ZN(n13637) );
  NAND2_X1 U15256 ( .A1(n13670), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13638) );
  INV_X1 U15257 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16667) );
  XNOR2_X1 U15258 ( .A(n13638), .B(n16667), .ZN(n16941) );
  NAND2_X1 U15259 ( .A1(n16941), .A2(n13773), .ZN(n13653) );
  INV_X1 U15260 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n16784) );
  OAI22_X1 U15261 ( .A1(n13519), .A2(n16784), .B1(n13671), .B2(n16667), .ZN(
        n13651) );
  AOI22_X1 U15262 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U15263 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U15264 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13639) );
  NAND4_X1 U15265 ( .A1(n13642), .A2(n13641), .A3(n13640), .A4(n13639), .ZN(
        n13648) );
  AOI22_X1 U15266 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U15267 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U15268 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U15269 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13643) );
  NAND4_X1 U15270 ( .A1(n13646), .A2(n13645), .A3(n13644), .A4(n13643), .ZN(
        n13647) );
  NOR2_X1 U15271 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  NOR2_X1 U15272 ( .A1(n13701), .A2(n13649), .ZN(n13650) );
  NOR2_X1 U15273 ( .A1(n13651), .A2(n13650), .ZN(n13652) );
  NAND2_X1 U15274 ( .A1(n13653), .A2(n13652), .ZN(n16661) );
  INV_X1 U15275 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16952) );
  XNOR2_X1 U15276 ( .A(n13670), .B(n16952), .ZN(n22329) );
  OR2_X1 U15277 ( .A1(n22329), .A2(n13982), .ZN(n13668) );
  AOI22_X1 U15278 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13816), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13657) );
  AOI22_X1 U15279 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U15280 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U15281 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11227), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13654) );
  NAND4_X1 U15282 ( .A1(n13657), .A2(n13656), .A3(n13655), .A4(n13654), .ZN(
        n13663) );
  AOI22_X1 U15283 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13945), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U15284 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13993), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U15285 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13116), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U15286 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13658) );
  NAND4_X1 U15287 ( .A1(n13661), .A2(n13660), .A3(n13659), .A4(n13658), .ZN(
        n13662) );
  NOR2_X1 U15288 ( .A1(n13663), .A2(n13662), .ZN(n13664) );
  OAI22_X1 U15289 ( .A1(n13701), .A2(n13664), .B1(n13671), .B2(n16952), .ZN(
        n13666) );
  INV_X1 U15290 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n16788) );
  NOR2_X1 U15291 ( .A1(n13519), .A2(n16788), .ZN(n13665) );
  NOR2_X1 U15292 ( .A1(n13666), .A2(n13665), .ZN(n13667) );
  NAND2_X1 U15293 ( .A1(n13668), .A2(n13667), .ZN(n16696) );
  XNOR2_X1 U15294 ( .A(n13697), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16925) );
  NAND2_X1 U15295 ( .A1(n16925), .A2(n13773), .ZN(n13686) );
  INV_X1 U15296 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n16780) );
  INV_X1 U15297 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16926) );
  OAI22_X1 U15298 ( .A1(n13519), .A2(n16780), .B1(n13671), .B2(n16926), .ZN(
        n13684) );
  AOI22_X1 U15299 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13675) );
  AOI22_X1 U15300 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U15301 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13672) );
  NAND4_X1 U15302 ( .A1(n13675), .A2(n13674), .A3(n13673), .A4(n13672), .ZN(
        n13681) );
  AOI22_X1 U15303 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U15304 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13086), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U15305 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U15306 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13676) );
  NAND4_X1 U15307 ( .A1(n13679), .A2(n13678), .A3(n13677), .A4(n13676), .ZN(
        n13680) );
  NOR2_X1 U15308 ( .A1(n13681), .A2(n13680), .ZN(n13682) );
  NOR2_X1 U15309 ( .A1(n13701), .A2(n13682), .ZN(n13683) );
  NOR2_X1 U15310 ( .A1(n13684), .A2(n13683), .ZN(n13685) );
  NAND2_X1 U15311 ( .A1(n13686), .A2(n13685), .ZN(n16646) );
  AOI22_X1 U15312 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13690) );
  AOI22_X1 U15313 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U15314 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U15315 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13687) );
  NAND4_X1 U15316 ( .A1(n13690), .A2(n13689), .A3(n13688), .A4(n13687), .ZN(
        n13696) );
  AOI22_X1 U15317 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13694) );
  AOI22_X1 U15318 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13994), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U15319 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13692) );
  AOI22_X1 U15320 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13691) );
  NAND4_X1 U15321 ( .A1(n13694), .A2(n13693), .A3(n13692), .A4(n13691), .ZN(
        n13695) );
  NOR2_X1 U15322 ( .A1(n13696), .A2(n13695), .ZN(n13702) );
  NAND2_X1 U15323 ( .A1(n14010), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13700) );
  INV_X1 U15324 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n22340) );
  XOR2_X1 U15325 ( .A(n22340), .B(n13717), .Z(n22344) );
  INV_X1 U15326 ( .A(n22344), .ZN(n13698) );
  AOI22_X1 U15327 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n14009), .B1(
        n15010), .B2(n13698), .ZN(n13699) );
  OAI211_X1 U15328 ( .C1(n13702), .C2(n13701), .A(n13700), .B(n13699), .ZN(
        n16777) );
  INV_X1 U15329 ( .A(n13161), .ZN(n14735) );
  AOI22_X1 U15330 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U15331 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U15332 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U15333 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13703) );
  NAND4_X1 U15334 ( .A1(n13706), .A2(n13705), .A3(n13704), .A4(n13703), .ZN(
        n13712) );
  AOI22_X1 U15335 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13710) );
  AOI22_X1 U15336 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U15337 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13708) );
  NAND4_X1 U15338 ( .A1(n13710), .A2(n13709), .A3(n13708), .A4(n13707), .ZN(
        n13711) );
  NOR2_X1 U15339 ( .A1(n13712), .A2(n13711), .ZN(n13716) );
  INV_X1 U15340 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15589) );
  NAND2_X1 U15341 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13713) );
  OAI211_X1 U15342 ( .C1(n13519), .C2(n15589), .A(n13982), .B(n13713), .ZN(
        n13714) );
  INV_X1 U15343 ( .A(n13714), .ZN(n13715) );
  OAI21_X1 U15344 ( .B1(n13979), .B2(n13716), .A(n13715), .ZN(n13722) );
  INV_X1 U15345 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13752) );
  NOR2_X1 U15346 ( .A1(n13719), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13720) );
  OR2_X1 U15347 ( .A1(n13809), .A2(n13720), .ZN(n16888) );
  INV_X1 U15348 ( .A(n16888), .ZN(n22356) );
  NAND2_X1 U15349 ( .A1(n22356), .A2(n15010), .ZN(n13721) );
  AOI22_X1 U15350 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13994), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U15351 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13724) );
  AOI22_X1 U15352 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13723) );
  NAND4_X1 U15353 ( .A1(n13726), .A2(n13725), .A3(n13724), .A4(n13723), .ZN(
        n13734) );
  AOI22_X1 U15354 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U15355 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13728) );
  NAND2_X1 U15356 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13727) );
  AND3_X1 U15357 ( .A1(n13728), .A2(n13727), .A3(n13982), .ZN(n13731) );
  AOI22_X1 U15358 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U15359 ( .A1(n13945), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13729) );
  NAND4_X1 U15360 ( .A1(n13732), .A2(n13731), .A3(n13730), .A4(n13729), .ZN(
        n13733) );
  NAND2_X1 U15361 ( .A1(n13979), .A2(n13982), .ZN(n13828) );
  OAI21_X1 U15362 ( .B1(n13734), .B2(n13733), .A(n13828), .ZN(n13737) );
  NAND2_X1 U15363 ( .A1(n14010), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U15364 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13735) );
  NAND3_X1 U15365 ( .A1(n13737), .A2(n13736), .A3(n13735), .ZN(n13740) );
  INV_X1 U15366 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16616) );
  XNOR2_X1 U15367 ( .A(n13738), .B(n16616), .ZN(n16893) );
  NAND2_X1 U15368 ( .A1(n16893), .A2(n13773), .ZN(n13739) );
  NAND2_X1 U15369 ( .A1(n13740), .A2(n13739), .ZN(n16609) );
  AOI22_X1 U15370 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13744) );
  AOI22_X1 U15371 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U15372 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13741) );
  NAND4_X1 U15373 ( .A1(n13744), .A2(n13743), .A3(n13742), .A4(n13741), .ZN(
        n13750) );
  AOI22_X1 U15374 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13748) );
  AOI22_X1 U15375 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13747) );
  AOI22_X1 U15376 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13746) );
  AOI22_X1 U15377 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13745) );
  NAND4_X1 U15378 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13749) );
  OR2_X1 U15379 ( .A1(n13750), .A2(n13749), .ZN(n13756) );
  INV_X1 U15380 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n16761) );
  XOR2_X1 U15381 ( .A(n13752), .B(n13751), .Z(n20858) );
  INV_X1 U15382 ( .A(n20858), .ZN(n13753) );
  AOI22_X1 U15383 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n14009), .B1(
        n13773), .B2(n13753), .ZN(n13754) );
  OAI21_X1 U15384 ( .B1(n13519), .B2(n16761), .A(n13754), .ZN(n13755) );
  AOI21_X1 U15385 ( .B1(n14003), .B2(n13756), .A(n13755), .ZN(n16625) );
  AOI22_X1 U15386 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U15387 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U15388 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U15389 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13757) );
  NAND4_X1 U15390 ( .A1(n13760), .A2(n13759), .A3(n13758), .A4(n13757), .ZN(
        n13768) );
  NAND2_X1 U15391 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13762) );
  NAND2_X1 U15392 ( .A1(n13987), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13761) );
  AND3_X1 U15393 ( .A1(n13762), .A2(n13982), .A3(n13761), .ZN(n13765) );
  AOI22_X1 U15394 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13764) );
  AOI22_X1 U15395 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13763) );
  NAND4_X1 U15396 ( .A1(n13766), .A2(n13765), .A3(n13764), .A4(n13763), .ZN(
        n13767) );
  OAI21_X1 U15397 ( .B1(n13768), .B2(n13767), .A(n13828), .ZN(n13771) );
  NAND2_X1 U15398 ( .A1(n14010), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n13770) );
  NAND2_X1 U15399 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13769) );
  NAND3_X1 U15400 ( .A1(n13771), .A2(n13770), .A3(n13769), .ZN(n13775) );
  INV_X1 U15401 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16906) );
  XNOR2_X1 U15402 ( .A(n13772), .B(n16906), .ZN(n16908) );
  NAND2_X1 U15403 ( .A1(n16908), .A2(n13773), .ZN(n13774) );
  NAND2_X1 U15404 ( .A1(n13775), .A2(n13774), .ZN(n16634) );
  NOR2_X1 U15405 ( .A1(n16609), .A2(n16607), .ZN(n16608) );
  AOI22_X1 U15406 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13993), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U15407 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13985), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13781) );
  NAND2_X1 U15408 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13778) );
  NAND2_X1 U15409 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13777) );
  AND3_X1 U15410 ( .A1(n13778), .A2(n13777), .A3(n13982), .ZN(n13780) );
  AOI22_X1 U15411 ( .A1(n13940), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11208), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13779) );
  NAND4_X1 U15412 ( .A1(n13782), .A2(n13781), .A3(n13780), .A4(n13779), .ZN(
        n13788) );
  AOI22_X1 U15413 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13816), .B1(
        n13968), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U15414 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13785) );
  AOI22_X1 U15415 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U15416 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13104), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13783) );
  NAND4_X1 U15417 ( .A1(n13786), .A2(n13785), .A3(n13784), .A4(n13783), .ZN(
        n13787) );
  OR2_X1 U15418 ( .A1(n13788), .A2(n13787), .ZN(n13789) );
  NAND2_X1 U15419 ( .A1(n13828), .A2(n13789), .ZN(n13792) );
  INV_X1 U15420 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15581) );
  INV_X1 U15421 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16879) );
  OAI22_X1 U15422 ( .A1(n13519), .A2(n15581), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n16879), .ZN(n13790) );
  INV_X1 U15423 ( .A(n13790), .ZN(n13791) );
  NAND2_X1 U15424 ( .A1(n13792), .A2(n13791), .ZN(n13794) );
  XNOR2_X1 U15425 ( .A(n13809), .B(n16879), .ZN(n16881) );
  NAND2_X1 U15426 ( .A1(n16881), .A2(n15010), .ZN(n13793) );
  NAND2_X1 U15427 ( .A1(n13794), .A2(n13793), .ZN(n16595) );
  AOI22_X1 U15428 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U15429 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13086), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13797) );
  AOI22_X1 U15430 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13796) );
  AOI22_X1 U15431 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13795) );
  NAND4_X1 U15432 ( .A1(n13798), .A2(n13797), .A3(n13796), .A4(n13795), .ZN(
        n13804) );
  AOI22_X1 U15433 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U15434 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13994), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13801) );
  AOI22_X1 U15435 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11209), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U15436 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13799) );
  NAND4_X1 U15437 ( .A1(n13802), .A2(n13801), .A3(n13800), .A4(n13799), .ZN(
        n13803) );
  NOR2_X1 U15438 ( .A1(n13804), .A2(n13803), .ZN(n13808) );
  INV_X1 U15439 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15583) );
  NAND2_X1 U15440 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13805) );
  OAI211_X1 U15441 ( .C1(n13519), .C2(n15583), .A(n13982), .B(n13805), .ZN(
        n13806) );
  INV_X1 U15442 ( .A(n13806), .ZN(n13807) );
  OAI21_X1 U15443 ( .B1(n13979), .B2(n13808), .A(n13807), .ZN(n13814) );
  INV_X1 U15444 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U15445 ( .A1(n13811), .A2(n13810), .ZN(n13812) );
  NAND2_X1 U15446 ( .A1(n13833), .A2(n13812), .ZN(n22385) );
  NAND2_X1 U15447 ( .A1(n13814), .A2(n13813), .ZN(n16740) );
  AOI22_X1 U15448 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13820) );
  AOI22_X1 U15449 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13819) );
  AOI22_X1 U15450 ( .A1(n13986), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U15451 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13817) );
  NAND4_X1 U15452 ( .A1(n13820), .A2(n13819), .A3(n13818), .A4(n13817), .ZN(
        n13830) );
  INV_X1 U15453 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13823) );
  AOI21_X1 U15454 ( .B1(n13963), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n15010), .ZN(n13821) );
  OAI211_X1 U15455 ( .C1(n13190), .C2(n13823), .A(n13822), .B(n13821), .ZN(
        n13824) );
  INV_X1 U15456 ( .A(n13824), .ZN(n13827) );
  AOI22_X1 U15457 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U15458 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13825) );
  NAND3_X1 U15459 ( .A1(n13827), .A2(n13826), .A3(n13825), .ZN(n13829) );
  OAI21_X1 U15460 ( .B1(n13830), .B2(n13829), .A(n13828), .ZN(n13832) );
  AOI22_X1 U15461 ( .A1(n14010), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n22489), .ZN(n13831) );
  XNOR2_X1 U15462 ( .A(n13833), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16583) );
  AOI22_X1 U15463 ( .A1(n13832), .A2(n13831), .B1(n15010), .B2(n16583), .ZN(
        n16579) );
  INV_X1 U15464 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13835) );
  NAND2_X1 U15465 ( .A1(n13836), .A2(n13835), .ZN(n13837) );
  NAND2_X1 U15466 ( .A1(n13896), .A2(n13837), .ZN(n16853) );
  AOI22_X1 U15467 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U15468 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U15469 ( .A1(n13940), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U15470 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13838) );
  NAND4_X1 U15471 ( .A1(n13841), .A2(n13840), .A3(n13839), .A4(n13838), .ZN(
        n13847) );
  AOI22_X1 U15472 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U15473 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U15474 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U15475 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13842) );
  NAND4_X1 U15476 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n13846) );
  NOR2_X1 U15477 ( .A1(n13847), .A2(n13846), .ZN(n13876) );
  AOI22_X1 U15478 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13851) );
  AOI22_X1 U15479 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U15480 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13849) );
  AOI22_X1 U15481 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13848) );
  NAND4_X1 U15482 ( .A1(n13851), .A2(n13850), .A3(n13849), .A4(n13848), .ZN(
        n13857) );
  AOI22_X1 U15483 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U15484 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13086), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U15485 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U15486 ( .A1(n13940), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13852) );
  NAND4_X1 U15487 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  NOR2_X1 U15488 ( .A1(n13857), .A2(n13856), .ZN(n13875) );
  XNOR2_X1 U15489 ( .A(n13876), .B(n13875), .ZN(n13860) );
  AOI21_X1 U15490 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n22489), .A(
        n15010), .ZN(n13859) );
  NAND2_X1 U15491 ( .A1(n14010), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n13858) );
  OAI211_X1 U15492 ( .C1(n13979), .C2(n13860), .A(n13859), .B(n13858), .ZN(
        n13861) );
  INV_X1 U15493 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13862) );
  NOR2_X1 U15494 ( .A1(n13196), .A2(n13862), .ZN(n13866) );
  INV_X1 U15495 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13864) );
  OAI22_X1 U15496 ( .A1(n13190), .A2(n13864), .B1(n13863), .B2(n13250), .ZN(
        n13865) );
  AOI211_X1 U15497 ( .C1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .C2(n11354), .A(
        n13866), .B(n13865), .ZN(n13874) );
  AOI22_X1 U15498 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U15499 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13869) );
  AOI22_X1 U15500 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U15501 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13867) );
  AND4_X1 U15502 ( .A1(n13870), .A2(n13869), .A3(n13868), .A4(n13867), .ZN(
        n13873) );
  AOI22_X1 U15503 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U15504 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13871) );
  NAND4_X1 U15505 ( .A1(n13874), .A2(n13873), .A3(n13872), .A4(n13871), .ZN(
        n13891) );
  NOR2_X1 U15506 ( .A1(n13876), .A2(n13875), .ZN(n13892) );
  XOR2_X1 U15507 ( .A(n13891), .B(n13892), .Z(n13877) );
  NAND2_X1 U15508 ( .A1(n13877), .A2(n14003), .ZN(n13880) );
  INV_X1 U15509 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13895) );
  AOI21_X1 U15510 ( .B1(n13895), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13878) );
  AOI21_X1 U15511 ( .B1(n14010), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13878), .ZN(
        n13879) );
  XNOR2_X1 U15512 ( .A(n13896), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16844) );
  AOI22_X1 U15513 ( .A1(n13880), .A2(n13879), .B1(n15010), .B2(n16844), .ZN(
        n16556) );
  AOI22_X1 U15514 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U15515 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13115), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13883) );
  AOI22_X1 U15516 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U15517 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13881) );
  NAND4_X1 U15518 ( .A1(n13884), .A2(n13883), .A3(n13882), .A4(n13881), .ZN(
        n13890) );
  AOI22_X1 U15519 ( .A1(n13081), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U15520 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U15521 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13885) );
  NAND4_X1 U15522 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13889) );
  NOR2_X1 U15523 ( .A1(n13890), .A2(n13889), .ZN(n13914) );
  NAND2_X1 U15524 ( .A1(n13892), .A2(n13891), .ZN(n13913) );
  XNOR2_X1 U15525 ( .A(n13914), .B(n13913), .ZN(n13893) );
  NOR2_X1 U15526 ( .A1(n13893), .A2(n13979), .ZN(n13902) );
  INV_X1 U15527 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n16721) );
  INV_X1 U15528 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n15972) );
  NOR2_X1 U15529 ( .A1(n15972), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13894) );
  OAI22_X1 U15530 ( .A1(n13519), .A2(n16721), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13894), .ZN(n13901) );
  INV_X1 U15531 ( .A(n13897), .ZN(n13899) );
  INV_X1 U15532 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U15533 ( .A1(n13899), .A2(n13898), .ZN(n13900) );
  NAND2_X1 U15534 ( .A1(n13920), .A2(n13900), .ZN(n16835) );
  OAI22_X1 U15535 ( .A1(n13902), .A2(n13901), .B1(n13982), .B2(n16835), .ZN(
        n16545) );
  AOI22_X1 U15536 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U15537 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13905) );
  AOI22_X1 U15538 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U15539 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13903) );
  NAND4_X1 U15540 ( .A1(n13906), .A2(n13905), .A3(n13904), .A4(n13903), .ZN(
        n13912) );
  AOI22_X1 U15541 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13223), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U15542 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U15543 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U15544 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13907) );
  NAND4_X1 U15545 ( .A1(n13910), .A2(n13909), .A3(n13908), .A4(n13907), .ZN(
        n13911) );
  OR2_X1 U15546 ( .A1(n13912), .A2(n13911), .ZN(n13924) );
  NOR2_X1 U15547 ( .A1(n13914), .A2(n13913), .ZN(n13925) );
  XOR2_X1 U15548 ( .A(n13924), .B(n13925), .Z(n13915) );
  NAND2_X1 U15549 ( .A1(n13915), .A2(n14003), .ZN(n13918) );
  INV_X1 U15550 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13919) );
  AOI21_X1 U15551 ( .B1(n13919), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13916) );
  AOI21_X1 U15552 ( .B1(n14010), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13916), .ZN(
        n13917) );
  XNOR2_X1 U15553 ( .A(n13920), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16824) );
  AOI22_X1 U15554 ( .A1(n13918), .A2(n13917), .B1(n15010), .B2(n16824), .ZN(
        n16530) );
  NAND2_X1 U15555 ( .A1(n16529), .A2(n16530), .ZN(n16517) );
  INV_X1 U15556 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13921) );
  NAND2_X1 U15557 ( .A1(n13922), .A2(n13921), .ZN(n13923) );
  NAND2_X1 U15558 ( .A1(n13958), .A2(n13923), .ZN(n16815) );
  NAND2_X1 U15559 ( .A1(n13925), .A2(n13924), .ZN(n13952) );
  AOI22_X1 U15560 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13816), .B1(
        n13985), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U15561 ( .A1(n11228), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U15562 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U15563 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13926) );
  NAND4_X1 U15564 ( .A1(n13929), .A2(n13928), .A3(n13927), .A4(n13926), .ZN(
        n13935) );
  AOI22_X1 U15565 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13081), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U15566 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13968), .B1(
        n13116), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U15567 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13993), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13930) );
  NAND4_X1 U15568 ( .A1(n13933), .A2(n13932), .A3(n13931), .A4(n13930), .ZN(
        n13934) );
  NOR2_X1 U15569 ( .A1(n13935), .A2(n13934), .ZN(n13953) );
  XNOR2_X1 U15570 ( .A(n13952), .B(n13953), .ZN(n13938) );
  AOI21_X1 U15571 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n22489), .A(
        n15010), .ZN(n13937) );
  NAND2_X1 U15572 ( .A1(n14010), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13936) );
  OAI211_X1 U15573 ( .C1(n13938), .C2(n13979), .A(n13937), .B(n13936), .ZN(
        n13939) );
  XNOR2_X1 U15574 ( .A(n13958), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16514) );
  AOI22_X1 U15575 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11228), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U15576 ( .A1(n13994), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U15577 ( .A1(n11226), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13940), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U15578 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13117), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13941) );
  NAND4_X1 U15579 ( .A1(n13944), .A2(n13943), .A3(n13942), .A4(n13941), .ZN(
        n13951) );
  AOI22_X1 U15580 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13963), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U15581 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13945), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U15582 ( .A1(n13993), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13137), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U15583 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13946) );
  NAND4_X1 U15584 ( .A1(n13949), .A2(n13948), .A3(n13947), .A4(n13946), .ZN(
        n13950) );
  OR2_X1 U15585 ( .A1(n13951), .A2(n13950), .ZN(n13975) );
  NOR2_X1 U15586 ( .A1(n13953), .A2(n13952), .ZN(n13976) );
  XOR2_X1 U15587 ( .A(n13975), .B(n13976), .Z(n13956) );
  INV_X1 U15588 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15585) );
  NOR2_X1 U15589 ( .A1(n15972), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13954) );
  OAI22_X1 U15590 ( .A1(n13519), .A2(n15585), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13954), .ZN(n13955) );
  AOI21_X1 U15591 ( .B1(n13956), .B2(n14003), .A(n13955), .ZN(n13957) );
  INV_X1 U15592 ( .A(n13958), .ZN(n13959) );
  NAND2_X1 U15593 ( .A1(n13959), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13961) );
  INV_X1 U15594 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13960) );
  NAND2_X1 U15595 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  NAND2_X1 U15596 ( .A1(n14014), .A2(n13962), .ZN(n16808) );
  AOI22_X1 U15597 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13988), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U15598 ( .A1(n13086), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13994), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U15599 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U15600 ( .A1(n13131), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11209), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13964) );
  NAND4_X1 U15601 ( .A1(n13967), .A2(n13966), .A3(n13965), .A4(n13964), .ZN(
        n13974) );
  AOI22_X1 U15602 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U15603 ( .A1(n13223), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13971) );
  AOI22_X1 U15604 ( .A1(n13968), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11225), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U15605 ( .A1(n13940), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13969) );
  NAND4_X1 U15606 ( .A1(n13972), .A2(n13971), .A3(n13970), .A4(n13969), .ZN(
        n13973) );
  NOR2_X1 U15607 ( .A1(n13974), .A2(n13973), .ZN(n13984) );
  NAND2_X1 U15608 ( .A1(n13976), .A2(n13975), .ZN(n13983) );
  XNOR2_X1 U15609 ( .A(n13984), .B(n13983), .ZN(n13980) );
  AOI21_X1 U15610 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22489), .A(
        n15010), .ZN(n13978) );
  NAND2_X1 U15611 ( .A1(n14010), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13977) );
  OAI211_X1 U15612 ( .C1(n13980), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        n13981) );
  OAI21_X1 U15613 ( .B1(n13982), .B2(n16808), .A(n13981), .ZN(n16496) );
  INV_X1 U15614 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15579) );
  NOR2_X1 U15615 ( .A1(n13984), .A2(n13983), .ZN(n14002) );
  AOI22_X1 U15616 ( .A1(n13985), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13104), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U15617 ( .A1(n13816), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13986), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U15618 ( .A1(n11225), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13987), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U15619 ( .A1(n13988), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13105), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13989) );
  NAND4_X1 U15620 ( .A1(n13992), .A2(n13991), .A3(n13990), .A4(n13989), .ZN(
        n14000) );
  AOI22_X1 U15621 ( .A1(n13963), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13993), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13998) );
  AOI22_X1 U15622 ( .A1(n11161), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13994), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U15623 ( .A1(n11227), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13110), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13995) );
  NAND4_X1 U15624 ( .A1(n13998), .A2(n13997), .A3(n13996), .A4(n13995), .ZN(
        n13999) );
  NOR2_X1 U15625 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  XNOR2_X1 U15626 ( .A(n14002), .B(n14001), .ZN(n14004) );
  NAND2_X1 U15627 ( .A1(n14004), .A2(n14003), .ZN(n14006) );
  OAI21_X1 U15628 ( .B1(n15972), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n22489), .ZN(n14005) );
  OAI211_X1 U15629 ( .C1(n13519), .C2(n15579), .A(n14006), .B(n14005), .ZN(
        n14008) );
  XNOR2_X1 U15630 ( .A(n14014), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16799) );
  NAND2_X1 U15631 ( .A1(n16799), .A2(n15010), .ZN(n14007) );
  NAND2_X1 U15632 ( .A1(n16495), .A2(n14402), .ZN(n14013) );
  AOI22_X1 U15633 ( .A1(n14010), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14009), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14011) );
  INV_X1 U15634 ( .A(n14011), .ZN(n14012) );
  XNOR2_X2 U15635 ( .A(n14013), .B(n14012), .ZN(n16477) );
  AND2_X1 U15636 ( .A1(n22396), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U15637 ( .A1(n15011), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22393) );
  INV_X2 U15638 ( .A(n16972), .ZN(n20860) );
  INV_X1 U15639 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16801) );
  NAND2_X1 U15640 ( .A1(n22534), .A2(n14019), .ZN(n22128) );
  NAND2_X1 U15641 ( .A1(n22128), .A2(n22396), .ZN(n14016) );
  NAND2_X1 U15642 ( .A1(n22396), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14018) );
  NAND2_X1 U15643 ( .A1(n15972), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14017) );
  AND2_X1 U15644 ( .A1(n14018), .A2(n14017), .ZN(n14877) );
  INV_X1 U15645 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20775) );
  NOR2_X1 U15646 ( .A1(n16939), .A2(n20775), .ZN(n14396) );
  AOI21_X1 U15647 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14396), .ZN(n14020) );
  OAI21_X1 U15648 ( .B1(n15022), .B2(n20856), .A(n14020), .ZN(n14021) );
  OAI21_X1 U15649 ( .B1(n14401), .B2(n22386), .A(n14022), .ZN(P1_U2968) );
  INV_X1 U15650 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21206) );
  INV_X1 U15651 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n21221) );
  NAND3_X1 U15652 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19007) );
  NAND2_X1 U15653 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18795) );
  INV_X1 U15654 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18982) );
  NOR2_X2 U15655 ( .A1(n18983), .A2(n18982), .ZN(n18743) );
  INV_X1 U15656 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21255) );
  NAND2_X1 U15657 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18820) );
  INV_X1 U15658 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18903) );
  INV_X1 U15659 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18961) );
  XOR2_X1 U15660 ( .A(n11351), .B(n14025), .Z(n21407) );
  INV_X1 U15661 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18940) );
  AOI21_X1 U15662 ( .B1(n18937), .B2(n18961), .A(n14025), .ZN(n18970) );
  INV_X1 U15663 ( .A(n18970), .ZN(n21393) );
  INV_X1 U15664 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18885) );
  NOR2_X1 U15665 ( .A1(n14029), .A2(n18885), .ZN(n14027) );
  OAI21_X1 U15666 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n14027), .A(
        n14026), .ZN(n21336) );
  XNOR2_X1 U15667 ( .A(n18885), .B(n14029), .ZN(n21323) );
  OAI21_X1 U15668 ( .B1(n14028), .B2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14029), .ZN(n21314) );
  INV_X1 U15669 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21282) );
  INV_X1 U15670 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21012) );
  NOR2_X1 U15671 ( .A1(n21201), .A2(n21012), .ZN(n18993) );
  NAND3_X1 U15672 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n18993), .ZN(n18779) );
  NOR2_X1 U15673 ( .A1(n18982), .A2(n18779), .ZN(n18744) );
  NAND2_X1 U15674 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18744), .ZN(
        n14033) );
  NOR2_X1 U15675 ( .A1(n21255), .A2(n14033), .ZN(n18818) );
  NAND2_X1 U15676 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18818), .ZN(
        n14031) );
  NOR2_X1 U15677 ( .A1(n21282), .A2(n14031), .ZN(n14030) );
  OAI21_X1 U15678 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14030), .A(
        n18854), .ZN(n21296) );
  XNOR2_X1 U15679 ( .A(n21282), .B(n14031), .ZN(n21288) );
  OAI21_X1 U15680 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18818), .A(
        n14031), .ZN(n21272) );
  AOI21_X1 U15681 ( .B1(n21255), .B2(n14033), .A(n18818), .ZN(n14032) );
  INV_X1 U15682 ( .A(n14032), .ZN(n21259) );
  OAI21_X1 U15683 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18744), .A(
        n14033), .ZN(n21245) );
  AOI21_X1 U15684 ( .B1(n18982), .B2(n18779), .A(n18744), .ZN(n18985) );
  INV_X1 U15685 ( .A(n18985), .ZN(n21235) );
  INV_X1 U15686 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21415) );
  NAND2_X1 U15687 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21415), .ZN(
        n21200) );
  NAND2_X1 U15688 ( .A1(n21259), .A2(n21258), .ZN(n21257) );
  NAND2_X1 U15689 ( .A1(n21199), .A2(n21286), .ZN(n21295) );
  NAND2_X1 U15690 ( .A1(n21296), .A2(n21295), .ZN(n21294) );
  NAND2_X1 U15691 ( .A1(n21199), .A2(n21321), .ZN(n21335) );
  NAND2_X1 U15692 ( .A1(n21336), .A2(n21335), .ZN(n21334) );
  NAND2_X1 U15693 ( .A1(n21199), .A2(n21334), .ZN(n21355) );
  OAI21_X1 U15694 ( .B1(n14034), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14036), .ZN(n21356) );
  NAND2_X1 U15695 ( .A1(n21355), .A2(n21356), .ZN(n21354) );
  NAND2_X1 U15696 ( .A1(n21199), .A2(n21354), .ZN(n21366) );
  AOI21_X1 U15697 ( .B1(n14036), .B2(n18903), .A(n14035), .ZN(n14037) );
  INV_X1 U15698 ( .A(n14037), .ZN(n21367) );
  NAND2_X1 U15699 ( .A1(n21199), .A2(n21365), .ZN(n21381) );
  OAI21_X1 U15700 ( .B1(n14035), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n18937), .ZN(n21382) );
  NAND2_X1 U15701 ( .A1(n21381), .A2(n21382), .ZN(n21380) );
  INV_X1 U15702 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22415) );
  NAND4_X1 U15703 ( .A1(n22113), .A2(n22091), .A3(n22415), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n22096) );
  OAI211_X1 U15704 ( .C1(n21407), .C2(n21406), .A(n21391), .B(n14038), .ZN(
        n14174) );
  OR2_X1 U15705 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n21025) );
  NOR2_X1 U15706 ( .A1(n21025), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n21024) );
  INV_X1 U15707 ( .A(n21024), .ZN(n21032) );
  NOR2_X1 U15708 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n21032), .ZN(n21046) );
  INV_X1 U15709 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n21045) );
  NAND2_X1 U15710 ( .A1(n21046), .A2(n21045), .ZN(n21062) );
  NOR2_X1 U15711 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n21062), .ZN(n21081) );
  INV_X1 U15712 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n21080) );
  NAND2_X1 U15713 ( .A1(n21081), .A2(n21080), .ZN(n21086) );
  NOR2_X1 U15714 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n21086), .ZN(n21111) );
  INV_X1 U15715 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n21110) );
  NAND2_X1 U15716 ( .A1(n21111), .A2(n21110), .ZN(n21117) );
  INV_X1 U15717 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n21140) );
  NAND2_X1 U15718 ( .A1(n21141), .A2(n21140), .ZN(n21146) );
  INV_X1 U15719 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21162) );
  NAND2_X1 U15720 ( .A1(n21163), .A2(n21162), .ZN(n21173) );
  INV_X1 U15721 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n21192) );
  NAND2_X1 U15722 ( .A1(n21193), .A2(n21192), .ZN(n21205) );
  INV_X1 U15723 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n21218) );
  NAND2_X1 U15724 ( .A1(n21219), .A2(n21218), .ZN(n21232) );
  INV_X1 U15725 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21246) );
  NAND2_X1 U15726 ( .A1(n21247), .A2(n21246), .ZN(n21254) );
  NOR2_X1 U15727 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n21254), .ZN(n21274) );
  INV_X1 U15728 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n21273) );
  NAND2_X1 U15729 ( .A1(n21274), .A2(n21273), .ZN(n21281) );
  NOR2_X1 U15730 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n21281), .ZN(n21298) );
  INV_X1 U15731 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n21297) );
  NAND2_X1 U15732 ( .A1(n21298), .A2(n21297), .ZN(n21307) );
  NOR2_X1 U15733 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n21307), .ZN(n21319) );
  INV_X1 U15734 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21326) );
  NAND2_X1 U15735 ( .A1(n21319), .A2(n21326), .ZN(n21330) );
  NOR2_X1 U15736 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n21330), .ZN(n21345) );
  INV_X1 U15737 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21346) );
  NAND2_X1 U15738 ( .A1(n21345), .A2(n21346), .ZN(n21360) );
  NOR2_X1 U15739 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n21360), .ZN(n21371) );
  INV_X1 U15740 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n21376) );
  NAND2_X1 U15741 ( .A1(n21371), .A2(n21376), .ZN(n21387) );
  NOR2_X1 U15742 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n21387), .ZN(n14165) );
  NAND2_X2 U15743 ( .A1(n21622), .A2(n21609), .ZN(n21005) );
  NOR2_X2 U15744 ( .A1(n21651), .A2(n14042), .ZN(n16134) );
  NAND2_X2 U15745 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21640) );
  INV_X2 U15746 ( .A(n14126), .ZN(n18547) );
  NOR2_X2 U15747 ( .A1(n21651), .A2(n14041), .ZN(n16155) );
  NOR2_X2 U15748 ( .A1(n21005), .A2(n14040), .ZN(n14107) );
  NOR2_X2 U15749 ( .A1(n21640), .A2(n14041), .ZN(n18475) );
  AOI22_X1 U15750 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14039) );
  OAI21_X1 U15751 ( .B1(n14125), .B2(n18690), .A(n14039), .ZN(n14049) );
  NOR2_X2 U15752 ( .A1(n21640), .A2(n14042), .ZN(n14067) );
  BUF_X2 U15753 ( .A(n14067), .Z(n18672) );
  AOI22_X1 U15754 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14047) );
  BUF_X2 U15755 ( .A(n14068), .Z(n18622) );
  NOR2_X2 U15756 ( .A1(n21651), .A2(n21638), .ZN(n14079) );
  AOI22_X1 U15757 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n21034), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14046) );
  NOR2_X2 U15758 ( .A1(n21638), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n21628) );
  NOR2_X2 U15759 ( .A1(n21656), .A2(n21015), .ZN(n18424) );
  NOR2_X2 U15760 ( .A1(n14043), .A2(n14042), .ZN(n16190) );
  BUF_X4 U15761 ( .A(n16190), .Z(n18716) );
  AOI22_X1 U15762 ( .A1(n21637), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14045) );
  INV_X4 U15763 ( .A(n11234), .ZN(n18674) );
  BUF_X2 U15764 ( .A(n14102), .Z(n18558) );
  AOI22_X1 U15765 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14044) );
  NAND4_X1 U15766 ( .A1(n14047), .A2(n14046), .A3(n14045), .A4(n14044), .ZN(
        n14048) );
  AOI22_X1 U15767 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U15768 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14062) );
  INV_X1 U15769 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U15770 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14053) );
  OAI21_X1 U15771 ( .B1(n14125), .B2(n14054), .A(n14053), .ZN(n14060) );
  AOI22_X1 U15772 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14058) );
  AOI22_X1 U15773 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U15774 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14056) );
  BUF_X2 U15775 ( .A(n14102), .Z(n18673) );
  AOI22_X1 U15776 ( .A1(n18673), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14055) );
  NAND4_X1 U15777 ( .A1(n14058), .A2(n14057), .A3(n14056), .A4(n14055), .ZN(
        n14059) );
  AOI211_X1 U15778 ( .C1(n18717), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n14060), .B(n14059), .ZN(n14061) );
  NAND3_X1 U15779 ( .A1(n14063), .A2(n14062), .A3(n14061), .ZN(n19196) );
  NAND2_X1 U15780 ( .A1(n19855), .A2(n19905), .ZN(n21424) );
  AOI22_X1 U15781 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U15782 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14077) );
  INV_X1 U15783 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14074) );
  INV_X1 U15784 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18710) );
  AOI22_X1 U15785 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n21637), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14065) );
  OAI21_X1 U15786 ( .B1(n14125), .B2(n18710), .A(n14065), .ZN(n14066) );
  INV_X1 U15787 ( .A(n14066), .ZN(n14073) );
  AOI22_X1 U15788 ( .A1(n16155), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U15789 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14071) );
  AOI22_X1 U15790 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14090), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U15791 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14069) );
  INV_X1 U15792 ( .A(n14075), .ZN(n14076) );
  NAND3_X2 U15793 ( .A1(n14078), .A2(n14077), .A3(n14076), .ZN(n21521) );
  NOR2_X1 U15794 ( .A1(n21424), .A2(n18687), .ZN(n14140) );
  AOI22_X1 U15795 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16190), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U15796 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14088) );
  INV_X1 U15797 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18546) );
  AOI22_X1 U15798 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14080) );
  OAI21_X1 U15799 ( .B1(n14125), .B2(n18546), .A(n14080), .ZN(n14086) );
  AOI22_X1 U15800 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U15801 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U15802 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U15803 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14081) );
  NAND4_X1 U15804 ( .A1(n14084), .A2(n14083), .A3(n14082), .A4(n14081), .ZN(
        n14085) );
  AOI211_X1 U15805 ( .C1(n18711), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n14086), .B(n14085), .ZN(n14087) );
  NAND3_X1 U15806 ( .A1(n14089), .A2(n14088), .A3(n14087), .ZN(n21486) );
  INV_X2 U15807 ( .A(n21486), .ZN(n19692) );
  AOI22_X1 U15808 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14101) );
  AOI22_X1 U15809 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14100) );
  INV_X1 U15810 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U15811 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14091) );
  OAI21_X1 U15812 ( .B1(n14125), .B2(n18350), .A(n14091), .ZN(n14098) );
  AOI22_X1 U15813 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U15814 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U15815 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U15816 ( .A1(n18673), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14093) );
  NAND4_X1 U15817 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14097) );
  NAND2_X1 U15818 ( .A1(n19692), .A2(n19652), .ZN(n16112) );
  AOI22_X1 U15819 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U15820 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U15821 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U15822 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14103) );
  NAND4_X1 U15823 ( .A1(n14106), .A2(n14105), .A3(n14104), .A4(n14103), .ZN(
        n14113) );
  AOI22_X1 U15824 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U15825 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14110) );
  AOI22_X1 U15826 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14107), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U15827 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14108) );
  NAND4_X1 U15828 ( .A1(n14111), .A2(n14110), .A3(n14109), .A4(n14108), .ZN(
        n14112) );
  AOI22_X1 U15829 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18711), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U15830 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14116) );
  AOI22_X1 U15831 ( .A1(n14107), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U15832 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18708), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14114) );
  NAND4_X1 U15833 ( .A1(n14117), .A2(n14116), .A3(n14115), .A4(n14114), .ZN(
        n14123) );
  AOI22_X1 U15834 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18707), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U15835 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14120) );
  AOI22_X1 U15836 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U15837 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14118) );
  NAND4_X1 U15838 ( .A1(n14121), .A2(n14120), .A3(n14119), .A4(n14118), .ZN(
        n14122) );
  NAND2_X1 U15839 ( .A1(n19813), .A2(n19773), .ZN(n21619) );
  NAND2_X1 U15840 ( .A1(n20937), .A2(n19905), .ZN(n16103) );
  AOI22_X1 U15841 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U15842 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18711), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14135) );
  INV_X1 U15843 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18323) );
  AOI22_X1 U15844 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14124) );
  OAI21_X1 U15845 ( .B1(n14125), .B2(n18323), .A(n14124), .ZN(n14133) );
  AOI22_X1 U15846 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U15847 ( .A1(n14126), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U15848 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14129) );
  AOI22_X1 U15849 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14128) );
  NAND4_X1 U15850 ( .A1(n14131), .A2(n14130), .A3(n14129), .A4(n14128), .ZN(
        n14132) );
  AOI211_X1 U15851 ( .C1(n18621), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n14133), .B(n14132), .ZN(n14134) );
  NAND3_X1 U15852 ( .A1(n14136), .A2(n14135), .A3(n14134), .ZN(n18318) );
  INV_X2 U15853 ( .A(n19652), .ZN(n21487) );
  NAND3_X2 U15854 ( .A1(n19733), .A2(n14148), .A3(n16123), .ZN(n16240) );
  OR2_X2 U15855 ( .A1(n16240), .A2(n19813), .ZN(n16119) );
  NOR2_X2 U15856 ( .A1(n14137), .A2(n19773), .ZN(n16113) );
  NAND2_X1 U15857 ( .A1(n21487), .A2(n16115), .ZN(n14141) );
  NAND2_X1 U15858 ( .A1(n16119), .A2(n14139), .ZN(n22059) );
  NOR2_X1 U15859 ( .A1(n20937), .A2(n14139), .ZN(n22089) );
  OAI21_X1 U15860 ( .B1(n16103), .B2(n18697), .A(n20947), .ZN(n18087) );
  OR2_X2 U15861 ( .A1(n18087), .A2(n20948), .ZN(n14149) );
  AOI21_X1 U15862 ( .B1(n14140), .B2(n18321), .A(n14149), .ZN(n16102) );
  INV_X1 U15863 ( .A(n16102), .ZN(n21621) );
  NAND2_X1 U15864 ( .A1(n19813), .A2(n21486), .ZN(n16127) );
  AOI21_X1 U15865 ( .B1(n16127), .B2(n14141), .A(n19773), .ZN(n14147) );
  NOR2_X1 U15866 ( .A1(n18687), .A2(n21607), .ZN(n21429) );
  NAND2_X1 U15867 ( .A1(n19855), .A2(n19196), .ZN(n16104) );
  NOR2_X1 U15868 ( .A1(n21429), .A2(n16104), .ZN(n16114) );
  NOR2_X1 U15869 ( .A1(n18687), .A2(n16123), .ZN(n14143) );
  NAND2_X1 U15870 ( .A1(n16103), .A2(n19813), .ZN(n16120) );
  INV_X1 U15871 ( .A(n16120), .ZN(n14142) );
  OAI22_X1 U15872 ( .A1(n19733), .A2(n14143), .B1(n16123), .B2(n14142), .ZN(
        n14144) );
  AOI211_X1 U15873 ( .C1(n21607), .C2(n19733), .A(n16114), .B(n14144), .ZN(
        n14146) );
  NAND2_X1 U15874 ( .A1(n21487), .A2(n18318), .ZN(n21620) );
  NAND4_X1 U15875 ( .A1(n19813), .A2(n19905), .A3(n16112), .A4(n21620), .ZN(
        n14145) );
  OR2_X2 U15876 ( .A1(n21621), .A2(n21642), .ZN(n21617) );
  NOR2_X4 U15877 ( .A1(n21617), .A2(n16240), .ZN(n21616) );
  NOR2_X1 U15878 ( .A1(n22113), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n22093) );
  NAND2_X1 U15879 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n22093), .ZN(n22088) );
  AOI22_X1 U15880 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n22069), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21622), .ZN(n16109) );
  INV_X1 U15881 ( .A(n16109), .ZN(n14157) );
  NAND2_X1 U15882 ( .A1(n19617), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16107) );
  OAI22_X1 U15883 ( .A1(n21033), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n22076), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14155) );
  OAI22_X1 U15884 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n22080), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14152), .ZN(n14158) );
  NOR2_X1 U15885 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n22080), .ZN(
        n14153) );
  NAND2_X1 U15886 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14152), .ZN(
        n14159) );
  AOI22_X1 U15887 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14158), .B1(
        n14153), .B2(n14159), .ZN(n16108) );
  NAND2_X1 U15888 ( .A1(n14156), .A2(n14155), .ZN(n14154) );
  OAI211_X1 U15889 ( .C1(n14156), .C2(n14155), .A(n16108), .B(n14154), .ZN(
        n16122) );
  XNOR2_X1 U15890 ( .A(n16107), .B(n14157), .ZN(n14161) );
  AOI21_X1 U15891 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14159), .A(
        n14158), .ZN(n14160) );
  OAI21_X1 U15892 ( .B1(n16122), .B2(n14161), .A(n16110), .ZN(n16129) );
  NAND2_X1 U15893 ( .A1(n20942), .A2(n19196), .ZN(n14164) );
  NAND2_X1 U15894 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n20941) );
  NAND2_X1 U15895 ( .A1(n20941), .A2(n22415), .ZN(n14162) );
  NOR2_X1 U15896 ( .A1(n14165), .A2(n21385), .ZN(n21389) );
  INV_X1 U15897 ( .A(n21389), .ZN(n14167) );
  INV_X1 U15898 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22419) );
  INV_X1 U15899 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22440) );
  NOR2_X1 U15900 ( .A1(n22440), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n22437) );
  INV_X1 U15901 ( .A(n22437), .ZN(n22444) );
  AOI21_X1 U15902 ( .B1(n19239), .B2(n22444), .A(n19229), .ZN(n20936) );
  OAI211_X1 U15903 ( .C1(n20936), .C2(n20937), .A(n20941), .B(n22415), .ZN(
        n14163) );
  INV_X1 U15904 ( .A(n14163), .ZN(n22090) );
  AOI211_X4 U15905 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20937), .A(n22090), .B(
        n14164), .ZN(n21420) );
  AND2_X1 U15906 ( .A1(n21419), .A2(n14165), .ZN(n21404) );
  NOR2_X1 U15907 ( .A1(n21420), .A2(n21404), .ZN(n14166) );
  MUX2_X1 U15908 ( .A(n14167), .B(n14166), .S(P3_EBX_REG_30__SCAN_IN), .Z(
        n14173) );
  INV_X1 U15909 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21612) );
  NAND2_X1 U15910 ( .A1(n21612), .A2(n22091), .ZN(n22102) );
  NOR2_X1 U15911 ( .A1(n22102), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18696) );
  NOR2_X1 U15912 ( .A1(n22100), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19628) );
  AND2_X1 U15913 ( .A1(n22093), .A2(n19628), .ZN(n22108) );
  NOR4_X2 U15914 ( .A1(n22043), .A2(n20942), .A3(n21391), .A4(n22108), .ZN(
        n21416) );
  INV_X1 U15915 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21940) );
  INV_X1 U15916 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21898) );
  NOR2_X1 U15917 ( .A1(n21940), .A2(n21898), .ZN(n14169) );
  INV_X1 U15918 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21862) );
  INV_X1 U15919 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21359) );
  INV_X1 U15920 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21965) );
  INV_X1 U15921 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21242) );
  INV_X1 U15922 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n21126) );
  INV_X1 U15923 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19225) );
  INV_X1 U15924 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n21060) );
  NAND3_X1 U15925 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n21052) );
  NOR2_X1 U15926 ( .A1(n21060), .A2(n21052), .ZN(n21065) );
  NAND2_X1 U15927 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n21065), .ZN(n21064) );
  NOR2_X1 U15928 ( .A1(n19225), .A2(n21064), .ZN(n21089) );
  NAND2_X1 U15929 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21089), .ZN(n21125) );
  NOR2_X1 U15930 ( .A1(n21126), .A2(n21125), .ZN(n21101) );
  NAND4_X1 U15931 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_11__SCAN_IN), .A4(n21101), .ZN(n21185) );
  NAND3_X1 U15932 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_14__SCAN_IN), 
        .A3(P3_REIP_REG_12__SCAN_IN), .ZN(n21198) );
  NAND2_X1 U15933 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n21231) );
  NOR4_X1 U15934 ( .A1(n21242), .A2(n21185), .A3(n21198), .A4(n21231), .ZN(
        n21267) );
  INV_X1 U15935 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19232) );
  NAND2_X1 U15936 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n21268) );
  NOR2_X1 U15937 ( .A1(n19232), .A2(n21268), .ZN(n21280) );
  INV_X1 U15938 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21291) );
  INV_X1 U15939 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21680) );
  NOR2_X1 U15940 ( .A1(n21291), .A2(n21680), .ZN(n21304) );
  NAND4_X1 U15941 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n21267), .A3(n21280), 
        .A4(n21304), .ZN(n21305) );
  NOR2_X1 U15942 ( .A1(n21965), .A2(n21305), .ZN(n21338) );
  NAND2_X1 U15943 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21338), .ZN(n21348) );
  NOR2_X1 U15944 ( .A1(n21359), .A2(n21348), .ZN(n14170) );
  NAND2_X1 U15945 ( .A1(n14170), .A2(n21306), .ZN(n21344) );
  NOR2_X1 U15946 ( .A1(n21862), .A2(n21344), .ZN(n21372) );
  NAND2_X1 U15947 ( .A1(n21349), .A2(n21306), .ZN(n21418) );
  INV_X1 U15948 ( .A(n21418), .ZN(n21373) );
  AOI21_X1 U15949 ( .B1(n14169), .B2(n21372), .A(n21373), .ZN(n21400) );
  AOI22_X1 U15950 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21399), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n21400), .ZN(n14171) );
  NAND2_X1 U15951 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21364), .ZN(n21374) );
  NOR3_X1 U15952 ( .A1(n21940), .A2(n21898), .A3(n21374), .ZN(n21410) );
  INV_X1 U15953 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19235) );
  NAND2_X1 U15954 ( .A1(n21410), .A2(n19235), .ZN(n21402) );
  NAND3_X1 U15955 ( .A1(n14174), .A2(n14173), .A3(n14172), .ZN(P3_U2641) );
  NOR2_X1 U15956 ( .A1(n14176), .A2(n19495), .ZN(n14177) );
  AOI21_X1 U15957 ( .B1(n14178), .B2(n18055), .A(n14177), .ZN(n14195) );
  NOR2_X1 U15958 ( .A1(n14180), .A2(n14179), .ZN(n14181) );
  INV_X1 U15959 ( .A(n14182), .ZN(n16404) );
  INV_X1 U15960 ( .A(n14183), .ZN(n17759) );
  NOR2_X1 U15961 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17757) );
  NOR2_X1 U15962 ( .A1(n17759), .A2(n17757), .ZN(n16408) );
  OAI21_X1 U15963 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16404), .A(
        n16408), .ZN(n14189) );
  NOR2_X1 U15964 ( .A1(n16404), .A2(n14184), .ZN(n14436) );
  NAND2_X1 U15965 ( .A1(n14436), .A2(n14185), .ZN(n14187) );
  NAND2_X1 U15966 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  INV_X1 U15967 ( .A(n14191), .ZN(n14192) );
  OAI21_X1 U15968 ( .B1(n19457), .B2(n18061), .A(n14192), .ZN(n14193) );
  NAND2_X1 U15969 ( .A1(n14195), .A2(n14194), .ZN(P2_U3017) );
  INV_X1 U15970 ( .A(n17570), .ZN(n14197) );
  NAND2_X1 U15971 ( .A1(n14197), .A2(n14196), .ZN(n14198) );
  INV_X1 U15972 ( .A(n11244), .ZN(n14200) );
  INV_X1 U15973 ( .A(n18190), .ZN(n18199) );
  INV_X1 U15974 ( .A(n14202), .ZN(n14203) );
  XNOR2_X1 U15975 ( .A(n14201), .B(n14203), .ZN(n19445) );
  NAND2_X1 U15976 ( .A1(n14520), .A2(n14204), .ZN(n14205) );
  NAND2_X1 U15977 ( .A1(n11235), .A2(n14205), .ZN(n19452) );
  NOR2_X1 U15978 ( .A1(n14452), .A2(n18307), .ZN(n16406) );
  AOI21_X1 U15979 ( .B1(n18174), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16406), .ZN(n14206) );
  OAI21_X1 U15980 ( .B1(n18181), .B2(n19452), .A(n14206), .ZN(n14208) );
  INV_X1 U15981 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17557) );
  NOR2_X1 U15982 ( .A1(n17565), .A2(n17557), .ZN(n17556) );
  NAND2_X1 U15983 ( .A1(n16955), .A2(n17012), .ZN(n16820) );
  NAND2_X1 U15984 ( .A1(n13431), .A2(n16820), .ZN(n14214) );
  INV_X1 U15985 ( .A(n14214), .ZN(n14212) );
  NOR2_X1 U15986 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17033) );
  NOR3_X1 U15987 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14213) );
  NAND3_X1 U15988 ( .A1(n14214), .A2(n17033), .A3(n14213), .ZN(n14215) );
  INV_X1 U15989 ( .A(n17000), .ZN(n14218) );
  NAND2_X1 U15990 ( .A1(n14218), .A2(n20853), .ZN(n14221) );
  INV_X1 U15991 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16508) );
  INV_X1 U15992 ( .A(n16939), .ZN(n22241) );
  NAND2_X1 U15993 ( .A1(n22241), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16992) );
  OAI21_X1 U15994 ( .B1(n16966), .B2(n16508), .A(n16992), .ZN(n14219) );
  AOI21_X1 U15995 ( .B1(n20859), .B2(n16514), .A(n14219), .ZN(n14220) );
  NAND3_X1 U15996 ( .A1(n11507), .A2(n14221), .A3(n14220), .ZN(P1_U2971) );
  INV_X1 U15997 ( .A(n14222), .ZN(n14226) );
  NOR2_X1 U15998 ( .A1(n13161), .A2(n15017), .ZN(n17199) );
  NAND2_X1 U15999 ( .A1(n17199), .A2(n14364), .ZN(n14404) );
  INV_X1 U16000 ( .A(n14404), .ZN(n14223) );
  OR2_X1 U16001 ( .A1(n18145), .A2(n14223), .ZN(n16467) );
  NOR2_X1 U16002 ( .A1(n14359), .A2(n13204), .ZN(n14224) );
  NOR2_X1 U16003 ( .A1(n16467), .A2(n14224), .ZN(n14225) );
  NAND2_X1 U16004 ( .A1(n14226), .A2(n14225), .ZN(n14247) );
  NAND2_X1 U16005 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22129) );
  INV_X1 U16006 ( .A(n22129), .ZN(n22389) );
  OR2_X1 U16007 ( .A1(n18156), .A2(n22389), .ZN(n14405) );
  NOR2_X1 U16008 ( .A1(n14551), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n14944) );
  INV_X1 U16009 ( .A(n14944), .ZN(n18155) );
  NAND2_X1 U16010 ( .A1(n15026), .A2(n18155), .ZN(n15024) );
  INV_X1 U16011 ( .A(n15024), .ZN(n14227) );
  OAI211_X1 U16012 ( .C1(n14405), .C2(n14227), .A(n15025), .B(n14428), .ZN(
        n14228) );
  NAND2_X1 U16013 ( .A1(n14228), .A2(n16472), .ZN(n14237) );
  AND2_X1 U16014 ( .A1(n14230), .A2(n14229), .ZN(n14231) );
  NAND2_X1 U16015 ( .A1(n14232), .A2(n14231), .ZN(n14234) );
  AND2_X1 U16016 ( .A1(n14234), .A2(n14233), .ZN(n16471) );
  AOI21_X1 U16017 ( .B1(n11221), .B2(n18155), .A(n22389), .ZN(n14235) );
  NAND2_X1 U16018 ( .A1(n16471), .A2(n14235), .ZN(n14236) );
  MUX2_X1 U16019 ( .A(n14237), .B(n14236), .S(n13153), .Z(n14245) );
  AOI21_X1 U16020 ( .B1(n14239), .B2(n11221), .A(n15130), .ZN(n14240) );
  NAND2_X1 U16021 ( .A1(n14241), .A2(n14240), .ZN(n14368) );
  NAND4_X1 U16022 ( .A1(n14368), .A2(n14364), .A3(n14362), .A4(n14242), .ZN(
        n14243) );
  NAND2_X1 U16023 ( .A1(n14238), .A2(n14243), .ZN(n14724) );
  NAND3_X1 U16024 ( .A1(n16466), .A2(n14735), .A3(n11221), .ZN(n14244) );
  NAND3_X1 U16025 ( .A1(n14245), .A2(n14724), .A3(n14244), .ZN(n14246) );
  INV_X1 U16026 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U16027 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14250) );
  NAND2_X1 U16028 ( .A1(n14345), .A2(n14250), .ZN(n14252) );
  NAND2_X1 U16029 ( .A1(n15033), .A2(n14248), .ZN(n14251) );
  NAND2_X1 U16030 ( .A1(n14252), .A2(n14251), .ZN(n14253) );
  NAND2_X1 U16031 ( .A1(n14254), .A2(n14253), .ZN(n14255) );
  MUX2_X1 U16032 ( .A(n14351), .B(n14345), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14816) );
  OR2_X1 U16033 ( .A1(n14347), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U16034 ( .A1(n14345), .A2(n22158), .ZN(n14258) );
  INV_X1 U16035 ( .A(n14256), .ZN(n14625) );
  INV_X1 U16036 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n15031) );
  NAND2_X1 U16037 ( .A1(n15033), .A2(n15031), .ZN(n14257) );
  NAND3_X1 U16038 ( .A1(n14258), .A2(n14351), .A3(n14257), .ZN(n14259) );
  NAND2_X1 U16039 ( .A1(n14260), .A2(n14259), .ZN(n14949) );
  MUX2_X1 U16040 ( .A(n14344), .B(n14256), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n14261) );
  OAI21_X1 U16041 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14814), .A(
        n14261), .ZN(n15374) );
  OR2_X1 U16042 ( .A1(n14347), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n14265) );
  NAND2_X1 U16043 ( .A1(n14345), .A2(n22167), .ZN(n14263) );
  INV_X1 U16044 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n16074) );
  NAND2_X1 U16045 ( .A1(n15033), .A2(n16074), .ZN(n14262) );
  NAND3_X1 U16046 ( .A1(n14263), .A2(n14351), .A3(n14262), .ZN(n14264) );
  NAND2_X1 U16047 ( .A1(n14265), .A2(n14264), .ZN(n15257) );
  NAND2_X1 U16048 ( .A1(n15258), .A2(n15257), .ZN(n15256) );
  INV_X1 U16049 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20829) );
  NAND2_X1 U16050 ( .A1(n15033), .A2(n20829), .ZN(n14267) );
  NAND2_X1 U16051 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14266) );
  NAND3_X1 U16052 ( .A1(n14267), .A2(n14345), .A3(n14266), .ZN(n14268) );
  OAI21_X1 U16053 ( .B1(n14344), .B2(P1_EBX_REG_5__SCAN_IN), .A(n14268), .ZN(
        n20823) );
  NAND2_X1 U16054 ( .A1(n14270), .A2(n14269), .ZN(n20825) );
  OR2_X1 U16055 ( .A1(n14347), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n14274) );
  NAND2_X1 U16056 ( .A1(n14345), .A2(n22204), .ZN(n14272) );
  INV_X1 U16057 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n22275) );
  NAND2_X1 U16058 ( .A1(n15033), .A2(n22275), .ZN(n14271) );
  NAND3_X1 U16059 ( .A1(n14272), .A2(n14351), .A3(n14271), .ZN(n14273) );
  INV_X1 U16060 ( .A(n14814), .ZN(n14321) );
  NAND2_X1 U16061 ( .A1(n22211), .A2(n14321), .ZN(n14276) );
  MUX2_X1 U16062 ( .A(n14344), .B(n14351), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n14275) );
  NAND2_X1 U16063 ( .A1(n14276), .A2(n14275), .ZN(n20816) );
  OR2_X1 U16064 ( .A1(n14347), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U16065 ( .A1(n14345), .A2(n22216), .ZN(n14278) );
  INV_X1 U16066 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n22303) );
  NAND2_X1 U16067 ( .A1(n15033), .A2(n22303), .ZN(n14277) );
  NAND3_X1 U16068 ( .A1(n14278), .A2(n14256), .A3(n14277), .ZN(n14279) );
  NAND2_X1 U16069 ( .A1(n14280), .A2(n14279), .ZN(n16265) );
  MUX2_X1 U16070 ( .A(n14344), .B(n14351), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n14281) );
  OAI21_X1 U16071 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n14814), .A(
        n14281), .ZN(n16304) );
  OR2_X1 U16072 ( .A1(n14347), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14286) );
  NAND2_X1 U16073 ( .A1(n14345), .A2(n22235), .ZN(n14284) );
  INV_X1 U16074 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n16363) );
  NAND2_X1 U16075 ( .A1(n15033), .A2(n16363), .ZN(n14283) );
  NAND3_X1 U16076 ( .A1(n14284), .A2(n14351), .A3(n14283), .ZN(n14285) );
  INV_X1 U16077 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16063) );
  NAND2_X1 U16078 ( .A1(n15033), .A2(n16063), .ZN(n14288) );
  NAND2_X1 U16079 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14287) );
  NAND3_X1 U16080 ( .A1(n14288), .A2(n14345), .A3(n14287), .ZN(n14289) );
  OAI21_X1 U16081 ( .B1(n14344), .B2(P1_EBX_REG_11__SCAN_IN), .A(n14289), .ZN(
        n16706) );
  OR2_X1 U16082 ( .A1(n14347), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n14294) );
  NAND2_X1 U16083 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14290) );
  NAND2_X1 U16084 ( .A1(n14345), .A2(n14290), .ZN(n14292) );
  INV_X1 U16085 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n22325) );
  NAND2_X1 U16086 ( .A1(n15033), .A2(n22325), .ZN(n14291) );
  NAND2_X1 U16087 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  NAND2_X1 U16088 ( .A1(n14294), .A2(n14293), .ZN(n16698) );
  MUX2_X1 U16089 ( .A(n14344), .B(n14351), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14296) );
  OR2_X1 U16090 ( .A1(n14814), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14295) );
  OR2_X1 U16091 ( .A1(n14347), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U16092 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14297) );
  NAND2_X1 U16093 ( .A1(n14345), .A2(n14297), .ZN(n14299) );
  INV_X1 U16094 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16693) );
  NAND2_X1 U16095 ( .A1(n15033), .A2(n16693), .ZN(n14298) );
  NAND2_X1 U16096 ( .A1(n14299), .A2(n14298), .ZN(n14300) );
  NOR2_X2 U16097 ( .A1(n16665), .A2(n16649), .ZN(n16648) );
  MUX2_X1 U16098 ( .A(n14344), .B(n14256), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14302) );
  OAI21_X1 U16099 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14814), .A(
        n14302), .ZN(n17149) );
  OR2_X1 U16100 ( .A1(n14347), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U16101 ( .A1(n14345), .A2(n17141), .ZN(n14305) );
  INV_X1 U16102 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16692) );
  NAND2_X1 U16103 ( .A1(n15033), .A2(n16692), .ZN(n14304) );
  NAND3_X1 U16104 ( .A1(n14305), .A2(n14351), .A3(n14304), .ZN(n14306) );
  NAND2_X1 U16105 ( .A1(n14307), .A2(n14306), .ZN(n16637) );
  MUX2_X1 U16106 ( .A(n14344), .B(n14351), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14309) );
  OR2_X1 U16107 ( .A1(n14814), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14308) );
  NAND2_X1 U16108 ( .A1(n14309), .A2(n14308), .ZN(n16631) );
  INV_X1 U16109 ( .A(n16631), .ZN(n14310) );
  OR2_X1 U16110 ( .A1(n14347), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U16111 ( .A1(n14345), .A2(n16870), .ZN(n14312) );
  INV_X1 U16112 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16052) );
  NAND2_X1 U16113 ( .A1(n15033), .A2(n16052), .ZN(n14311) );
  NAND3_X1 U16114 ( .A1(n14312), .A2(n14351), .A3(n14311), .ZN(n14313) );
  MUX2_X1 U16115 ( .A(n14344), .B(n14256), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14315) );
  OAI21_X1 U16116 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14814), .A(
        n14315), .ZN(n17097) );
  OR2_X1 U16117 ( .A1(n14347), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U16118 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14316) );
  NAND2_X1 U16119 ( .A1(n14345), .A2(n14316), .ZN(n14318) );
  INV_X1 U16120 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n16690) );
  NAND2_X1 U16121 ( .A1(n15033), .A2(n16690), .ZN(n14317) );
  NAND2_X1 U16122 ( .A1(n14318), .A2(n14317), .ZN(n14319) );
  NAND2_X1 U16123 ( .A1(n14320), .A2(n14319), .ZN(n16600) );
  NAND2_X1 U16124 ( .A1(n17100), .A2(n16600), .ZN(n16599) );
  MUX2_X1 U16125 ( .A(n14344), .B(n14351), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14323) );
  NAND2_X1 U16126 ( .A1(n14321), .A2(n13427), .ZN(n14322) );
  NAND2_X1 U16127 ( .A1(n14323), .A2(n14322), .ZN(n17069) );
  OR2_X1 U16128 ( .A1(n14347), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14328) );
  NAND2_X1 U16129 ( .A1(n14351), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14324) );
  NAND2_X1 U16130 ( .A1(n14345), .A2(n14324), .ZN(n14326) );
  INV_X1 U16131 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16045) );
  NAND2_X1 U16132 ( .A1(n15033), .A2(n16045), .ZN(n14325) );
  NAND2_X1 U16133 ( .A1(n14326), .A2(n14325), .ZN(n14327) );
  AND2_X1 U16134 ( .A1(n14328), .A2(n14327), .ZN(n16582) );
  MUX2_X1 U16135 ( .A(n14344), .B(n14351), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14329) );
  OAI21_X1 U16136 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14814), .A(
        n14329), .ZN(n16570) );
  OR2_X1 U16137 ( .A1(n14347), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U16138 ( .A1(n14345), .A2(n14330), .ZN(n14332) );
  INV_X1 U16139 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n16687) );
  NAND2_X1 U16140 ( .A1(n15033), .A2(n16687), .ZN(n14331) );
  NAND3_X1 U16141 ( .A1(n14332), .A2(n14351), .A3(n14331), .ZN(n14333) );
  NAND2_X1 U16142 ( .A1(n14334), .A2(n14333), .ZN(n16562) );
  MUX2_X1 U16143 ( .A(n14344), .B(n14256), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14336) );
  OR2_X1 U16144 ( .A1(n14814), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14335) );
  AND2_X1 U16145 ( .A1(n14336), .A2(n14335), .ZN(n16542) );
  NAND2_X1 U16146 ( .A1(n16560), .A2(n16542), .ZN(n16541) );
  OR2_X1 U16147 ( .A1(n14347), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14340) );
  INV_X1 U16148 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17014) );
  NAND2_X1 U16149 ( .A1(n14345), .A2(n17014), .ZN(n14338) );
  INV_X1 U16150 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16036) );
  NAND2_X1 U16151 ( .A1(n15033), .A2(n16036), .ZN(n14337) );
  NAND3_X1 U16152 ( .A1(n14338), .A2(n14351), .A3(n14337), .ZN(n14339) );
  AND2_X1 U16153 ( .A1(n14340), .A2(n14339), .ZN(n16533) );
  OR2_X2 U16154 ( .A1(n16541), .A2(n16533), .ZN(n16531) );
  INV_X1 U16155 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15848) );
  NAND2_X1 U16156 ( .A1(n15033), .A2(n15848), .ZN(n14342) );
  NAND2_X1 U16157 ( .A1(n14256), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14341) );
  NAND3_X1 U16158 ( .A1(n14342), .A2(n14345), .A3(n14341), .ZN(n14343) );
  OAI21_X1 U16159 ( .B1(n14344), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14343), .ZN(
        n16520) );
  OAI21_X1 U16160 ( .B1(n14866), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14351), .ZN(
        n14349) );
  INV_X1 U16161 ( .A(n14345), .ZN(n14346) );
  NOR2_X1 U16162 ( .A1(n14346), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14348) );
  OAI22_X1 U16163 ( .A1(n14349), .A2(n14348), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14347), .ZN(n16505) );
  INV_X1 U16164 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16032) );
  NAND2_X1 U16165 ( .A1(n15033), .A2(n16032), .ZN(n14350) );
  OAI21_X1 U16166 ( .B1(n14814), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14350), .ZN(n16487) );
  MUX2_X1 U16167 ( .A(n14350), .B(n16487), .S(n14351), .Z(n16498) );
  AOI22_X1 U16168 ( .A1(n14814), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14866), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16488) );
  NAND2_X1 U16169 ( .A1(n16497), .A2(n16488), .ZN(n14352) );
  AOI22_X1 U16170 ( .A1(n14814), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14866), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14354) );
  INV_X1 U16171 ( .A(n14354), .ZN(n14355) );
  NAND2_X1 U16172 ( .A1(n14357), .A2(n13211), .ZN(n14358) );
  OAI21_X1 U16173 ( .B1(n14359), .B2(n14409), .A(n14358), .ZN(n14360) );
  NAND2_X1 U16174 ( .A1(n14362), .A2(n14361), .ZN(n14366) );
  OAI22_X1 U16175 ( .A1(n13448), .A2(n14363), .B1(n14364), .B2(n15130), .ZN(
        n14365) );
  AOI21_X1 U16176 ( .B1(n14366), .B2(n11221), .A(n14365), .ZN(n14369) );
  NAND2_X1 U16177 ( .A1(n13165), .A2(n13166), .ZN(n14367) );
  AND3_X1 U16178 ( .A1(n14369), .A2(n14368), .A3(n14367), .ZN(n14709) );
  OAI211_X1 U16179 ( .C1(n14706), .C2(n15025), .A(n14709), .B(n14370), .ZN(
        n14371) );
  INV_X1 U16180 ( .A(n14363), .ZN(n16475) );
  NAND2_X1 U16181 ( .A1(n14372), .A2(n16475), .ZN(n18127) );
  INV_X1 U16182 ( .A(n18127), .ZN(n17202) );
  NAND2_X1 U16183 ( .A1(n14378), .A2(n17202), .ZN(n17157) );
  NAND2_X1 U16184 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n22203) );
  INV_X1 U16185 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n22148) );
  NOR2_X1 U16186 ( .A1(n22158), .A2(n22148), .ZN(n22161) );
  INV_X1 U16187 ( .A(n22161), .ZN(n22165) );
  NOR2_X1 U16188 ( .A1(n22203), .A2(n22165), .ZN(n22183) );
  NOR2_X1 U16189 ( .A1(n22216), .A2(n22211), .ZN(n22219) );
  AND3_X1 U16190 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n22219), .ZN(n22220) );
  NAND4_X1 U16191 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n22183), .A4(n22220), .ZN(
        n17173) );
  NAND2_X1 U16192 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n22137) );
  NOR2_X1 U16193 ( .A1(n17173), .A2(n22137), .ZN(n17164) );
  NAND2_X1 U16194 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17109) );
  NOR3_X1 U16195 ( .A1(n16870), .A2(n17119), .A3(n17109), .ZN(n17051) );
  NAND2_X1 U16196 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17051), .ZN(
        n14373) );
  NOR2_X1 U16197 ( .A1(n17058), .A2(n14373), .ZN(n14374) );
  AND2_X1 U16198 ( .A1(n17164), .A2(n14374), .ZN(n14390) );
  INV_X1 U16199 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14389) );
  NAND2_X1 U16200 ( .A1(n17081), .A2(n14389), .ZN(n14376) );
  INV_X1 U16201 ( .A(n14378), .ZN(n14375) );
  NAND2_X1 U16202 ( .A1(n14375), .A2(n16939), .ZN(n14864) );
  NOR2_X1 U16203 ( .A1(n14377), .A2(n13161), .ZN(n17201) );
  AND2_X1 U16204 ( .A1(n17201), .A2(n15033), .ZN(n16468) );
  NAND2_X1 U16205 ( .A1(n14378), .A2(n16468), .ZN(n22151) );
  NOR2_X1 U16206 ( .A1(n22205), .A2(n22203), .ZN(n22181) );
  OAI21_X1 U16207 ( .B1(n14389), .B2(n22148), .A(n22158), .ZN(n22162) );
  NAND2_X1 U16208 ( .A1(n22181), .A2(n22162), .ZN(n22186) );
  NOR2_X1 U16209 ( .A1(n22204), .A2(n22186), .ZN(n22200) );
  NAND2_X1 U16210 ( .A1(n22219), .A2(n22200), .ZN(n22224) );
  INV_X1 U16211 ( .A(n22224), .ZN(n14380) );
  AND2_X1 U16212 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14379) );
  NAND2_X1 U16213 ( .A1(n14380), .A2(n14379), .ZN(n17050) );
  OR2_X1 U16214 ( .A1(n17050), .A2(n17177), .ZN(n17174) );
  NOR2_X1 U16215 ( .A1(n17182), .A2(n17174), .ZN(n17108) );
  NAND2_X1 U16216 ( .A1(n17051), .A2(n17108), .ZN(n17078) );
  INV_X1 U16217 ( .A(n17078), .ZN(n17057) );
  NAND2_X1 U16218 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17057), .ZN(
        n14381) );
  NOR2_X1 U16219 ( .A1(n17058), .A2(n14381), .ZN(n14391) );
  NAND2_X1 U16220 ( .A1(n14391), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14382) );
  NAND2_X1 U16221 ( .A1(n22225), .A2(n14382), .ZN(n14383) );
  OAI211_X1 U16222 ( .C1(n22221), .C2(n14390), .A(n22182), .B(n14383), .ZN(
        n17043) );
  INV_X1 U16223 ( .A(n17157), .ZN(n17165) );
  NAND2_X1 U16224 ( .A1(n17165), .A2(n17012), .ZN(n14386) );
  INV_X1 U16225 ( .A(n17034), .ZN(n14384) );
  NAND2_X1 U16226 ( .A1(n17081), .A2(n14384), .ZN(n14385) );
  OAI211_X1 U16227 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n22151), .A(
        n14386), .B(n14385), .ZN(n14387) );
  OR2_X1 U16228 ( .A1(n17043), .A2(n14387), .ZN(n17026) );
  NAND2_X1 U16229 ( .A1(n22221), .A2(n22151), .ZN(n17054) );
  NOR2_X1 U16230 ( .A1(n17026), .A2(n17054), .ZN(n17003) );
  INV_X1 U16231 ( .A(n16982), .ZN(n16993) );
  NAND2_X1 U16232 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14388) );
  NOR2_X1 U16233 ( .A1(n17026), .A2(n14388), .ZN(n17002) );
  AOI21_X1 U16234 ( .B1(n16993), .B2(n17002), .A(n17003), .ZN(n16985) );
  AOI21_X1 U16235 ( .B1(n16797), .B2(n17054), .A(n16985), .ZN(n16974) );
  OAI21_X1 U16236 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17003), .A(
        n16974), .ZN(n14397) );
  NAND2_X1 U16237 ( .A1(n22160), .A2(n14390), .ZN(n14393) );
  NAND2_X1 U16238 ( .A1(n22225), .A2(n14391), .ZN(n14392) );
  NAND2_X1 U16239 ( .A1(n14393), .A2(n14392), .ZN(n17032) );
  NOR2_X1 U16240 ( .A1(n17012), .A2(n17014), .ZN(n14394) );
  NAND2_X1 U16241 ( .A1(n17032), .A2(n14394), .ZN(n17001) );
  OR3_X1 U16242 ( .A1(n17001), .A2(n16797), .A3(n16982), .ZN(n16976) );
  NOR3_X1 U16243 ( .A1(n16976), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16973), .ZN(n14395) );
  AOI211_X1 U16244 ( .C1(n14397), .C2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14396), .B(n14395), .ZN(n14398) );
  OAI21_X1 U16245 ( .B1(n14401), .B2(n22226), .A(n14400), .ZN(P1_U3000) );
  INV_X1 U16246 ( .A(n16803), .ZN(n16681) );
  NAND2_X1 U16247 ( .A1(n16474), .A2(n15026), .ZN(n14620) );
  OAI21_X1 U16248 ( .B1(n14405), .B2(n14866), .A(n14404), .ZN(n14406) );
  NAND2_X1 U16249 ( .A1(n14406), .A2(n16472), .ZN(n14407) );
  NOR2_X1 U16250 ( .A1(n14409), .A2(n22406), .ZN(n14413) );
  NOR2_X1 U16251 ( .A1(n11182), .A2(n11183), .ZN(n14412) );
  NAND4_X1 U16252 ( .A1(n17198), .A2(n14413), .A3(n14412), .A4(n14411), .ZN(
        n14841) );
  OR2_X1 U16253 ( .A1(n14841), .A2(n15017), .ZN(n14414) );
  NAND2_X1 U16254 ( .A1(n13159), .A2(n11182), .ZN(n14882) );
  NOR4_X1 U16255 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14419) );
  NOR4_X1 U16256 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14418) );
  NOR4_X1 U16257 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14417) );
  NOR4_X1 U16258 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14416) );
  AND4_X1 U16259 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        n14424) );
  NOR4_X1 U16260 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n14422) );
  NOR4_X1 U16261 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14421) );
  NOR4_X1 U16262 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14420) );
  INV_X1 U16263 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20721) );
  AND4_X1 U16264 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n20721), .ZN(
        n14423) );
  NAND2_X1 U16265 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  AND2_X2 U16266 ( .A1(n14425), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14954)
         );
  INV_X1 U16267 ( .A(n14954), .ZN(n14784) );
  NOR3_X4 U16268 ( .A1(n16770), .A2(n14428), .A3(n14784), .ZN(n16774) );
  MUX2_X1 U16269 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14954), .Z(
        n16779) );
  AOI22_X1 U16270 ( .A1(n16774), .A2(BUF1_REG_30__SCAN_IN), .B1(n16773), .B2(
        n16779), .ZN(n14427) );
  INV_X1 U16271 ( .A(n14427), .ZN(n14432) );
  NOR2_X1 U16272 ( .A1(n14428), .A2(n14954), .ZN(n14429) );
  NAND2_X1 U16273 ( .A1(n16791), .A2(n14429), .ZN(n16763) );
  AOI22_X1 U16274 ( .A1(n16771), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16770), .ZN(n14430) );
  INV_X1 U16275 ( .A(n14430), .ZN(n14431) );
  NOR2_X1 U16276 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  OAI21_X1 U16277 ( .B1(n16681), .B2(n16782), .A(n14433), .ZN(P1_U2874) );
  NAND2_X1 U16278 ( .A1(n14434), .A2(n18055), .ZN(n14445) );
  OR2_X1 U16279 ( .A1(n14435), .A2(n19495), .ZN(n14444) );
  NAND3_X1 U16280 ( .A1(n14436), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12635), .ZN(n14437) );
  OAI211_X1 U16281 ( .C1(n19476), .C2(n18066), .A(n14438), .B(n14437), .ZN(
        n14439) );
  OAI21_X1 U16282 ( .B1(n19478), .B2(n18061), .A(n14441), .ZN(n14442) );
  INV_X1 U16283 ( .A(n14442), .ZN(n14443) );
  NAND3_X1 U16284 ( .A1(n14445), .A2(n14444), .A3(n14443), .ZN(P2_U3016) );
  INV_X1 U16285 ( .A(n13150), .ZN(n15140) );
  AND2_X1 U16286 ( .A1(n16791), .A2(n15140), .ZN(n14446) );
  NAND2_X1 U16287 ( .A1(n16477), .A2(n14446), .ZN(n14451) );
  AOI22_X1 U16288 ( .A1(n16774), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16770), .ZN(n14447) );
  INV_X1 U16289 ( .A(DATAI_31_), .ZN(n15907) );
  NOR2_X1 U16290 ( .A1(n16763), .A2(n15907), .ZN(n14448) );
  NOR2_X1 U16291 ( .A1(n14449), .A2(n14448), .ZN(n14450) );
  NAND2_X1 U16292 ( .A1(n14451), .A2(n14450), .ZN(P1_U2873) );
  NAND2_X1 U16293 ( .A1(n18168), .A2(n11738), .ZN(n14463) );
  NAND2_X1 U16294 ( .A1(n22411), .A2(n19531), .ZN(n14460) );
  NAND4_X1 U16295 ( .A1(n19251), .A2(n20103), .A3(n22411), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19518) );
  NAND2_X1 U16296 ( .A1(n19518), .A2(n14452), .ZN(n14453) );
  NAND2_X1 U16297 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20103), .ZN(n19521) );
  NOR3_X1 U16298 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n20165), .A3(n19521), 
        .ZN(n19524) );
  OR2_X1 U16299 ( .A1(n14453), .A2(n19524), .ZN(n14454) );
  INV_X2 U16300 ( .A(n19371), .ZN(n19471) );
  NAND2_X1 U16301 ( .A1(n15332), .A2(n22411), .ZN(n14455) );
  NAND2_X1 U16302 ( .A1(n14470), .A2(n14455), .ZN(n14457) );
  INV_X1 U16303 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14462) );
  NAND3_X1 U16304 ( .A1(n19249), .A2(n14460), .A3(n14462), .ZN(n14456) );
  NAND2_X1 U16305 ( .A1(n14457), .A2(n14456), .ZN(n14458) );
  INV_X1 U16306 ( .A(n19470), .ZN(n19409) );
  OAI22_X1 U16307 ( .A1(n19409), .A2(n14462), .B1(n19443), .B2(n14459), .ZN(
        n14466) );
  INV_X1 U16308 ( .A(n14460), .ZN(n14461) );
  NOR3_X1 U16309 ( .A1(n14464), .A2(P2_EBX_REG_30__SCAN_IN), .A3(n19441), .ZN(
        n14465) );
  AOI211_X1 U16310 ( .C1(n19471), .C2(P2_REIP_REG_31__SCAN_IN), .A(n14466), 
        .B(n14465), .ZN(n14467) );
  OAI21_X1 U16311 ( .B1(n16442), .B2(n19477), .A(n14467), .ZN(n14522) );
  AND3_X1 U16312 ( .A1(n15332), .A2(n14470), .A3(n22411), .ZN(n15360) );
  AOI21_X1 U16313 ( .B1(n17583), .B2(n14475), .A(n11345), .ZN(n17586) );
  INV_X1 U16314 ( .A(n17586), .ZN(n19427) );
  NAND2_X1 U16315 ( .A1(n14514), .A2(n14473), .ZN(n14474) );
  NAND2_X1 U16316 ( .A1(n14475), .A2(n14474), .ZN(n17593) );
  INV_X1 U16317 ( .A(n14479), .ZN(n14476) );
  AOI21_X1 U16318 ( .B1(n14476), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14477) );
  OR2_X1 U16319 ( .A1(n14477), .A2(n14512), .ZN(n19417) );
  INV_X1 U16320 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14478) );
  XNOR2_X1 U16321 ( .A(n14479), .B(n14478), .ZN(n19403) );
  INV_X1 U16322 ( .A(n19403), .ZN(n14511) );
  INV_X1 U16323 ( .A(n14480), .ZN(n14484) );
  INV_X1 U16324 ( .A(n14508), .ZN(n14482) );
  INV_X1 U16325 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U16326 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U16327 ( .A1(n14484), .A2(n14483), .ZN(n17634) );
  INV_X1 U16328 ( .A(n17634), .ZN(n14510) );
  AOI21_X1 U16329 ( .B1(n14505), .B2(n19358), .A(n14507), .ZN(n19355) );
  INV_X1 U16330 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17673) );
  INV_X1 U16331 ( .A(n14503), .ZN(n14485) );
  AOI21_X1 U16332 ( .B1(n17673), .B2(n14485), .A(n14506), .ZN(n17675) );
  OAI21_X1 U16333 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n14500), .A(
        n14504), .ZN(n17686) );
  INV_X1 U16334 ( .A(n17686), .ZN(n17336) );
  OAI21_X1 U16335 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n14496), .A(
        n14499), .ZN(n17716) );
  OAI21_X1 U16336 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n14492), .A(
        n14497), .ZN(n17729) );
  AOI21_X1 U16337 ( .B1(n17741), .B2(n14490), .A(n14494), .ZN(n17744) );
  AOI21_X1 U16338 ( .B1(n16332), .B2(n14488), .A(n14491), .ZN(n16335) );
  INV_X1 U16339 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17748) );
  NAND2_X1 U16340 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14487) );
  AOI21_X1 U16341 ( .B1(n17748), .B2(n14487), .A(n14489), .ZN(n17750) );
  OAI22_X1 U16342 ( .A1(n19251), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14486) );
  INV_X1 U16343 ( .A(n14486), .ZN(n19259) );
  AOI22_X1 U16344 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14696), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19251), .ZN(n15646) );
  NOR2_X1 U16345 ( .A1(n19259), .A2(n15646), .ZN(n15645) );
  OAI21_X1 U16346 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n14487), .ZN(n15481) );
  NAND2_X1 U16347 ( .A1(n15645), .A2(n15481), .ZN(n16445) );
  NOR2_X1 U16348 ( .A1(n17750), .A2(n16445), .ZN(n19279) );
  OAI21_X1 U16349 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14489), .A(
        n14488), .ZN(n19278) );
  NAND2_X1 U16350 ( .A1(n19279), .A2(n19278), .ZN(n15178) );
  NOR2_X1 U16351 ( .A1(n16335), .A2(n15178), .ZN(n19289) );
  OAI21_X1 U16352 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n14491), .A(
        n14490), .ZN(n19291) );
  NAND2_X1 U16353 ( .A1(n19289), .A2(n19291), .ZN(n15200) );
  NOR2_X1 U16354 ( .A1(n17744), .A2(n15200), .ZN(n19302) );
  INV_X1 U16355 ( .A(n14492), .ZN(n14493) );
  OAI21_X1 U16356 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n14494), .A(
        n14493), .ZN(n19304) );
  NAND2_X1 U16357 ( .A1(n19302), .A2(n19304), .ZN(n15262) );
  INV_X1 U16358 ( .A(n15262), .ZN(n14495) );
  NAND2_X1 U16359 ( .A1(n17729), .A2(n14495), .ZN(n19315) );
  AOI21_X1 U16360 ( .B1(n19313), .B2(n14497), .A(n14496), .ZN(n19316) );
  NOR2_X1 U16361 ( .A1(n19315), .A2(n19316), .ZN(n17342) );
  AND2_X1 U16362 ( .A1(n17716), .A2(n17342), .ZN(n17341) );
  NAND2_X1 U16363 ( .A1(n14499), .A2(n14498), .ZN(n14502) );
  INV_X1 U16364 ( .A(n14500), .ZN(n14501) );
  NAND2_X1 U16365 ( .A1(n14502), .A2(n14501), .ZN(n19325) );
  NAND2_X1 U16366 ( .A1(n17341), .A2(n19325), .ZN(n17335) );
  NOR2_X1 U16367 ( .A1(n17336), .A2(n17335), .ZN(n17334) );
  AOI21_X1 U16368 ( .B1(n11338), .B2(n14504), .A(n14503), .ZN(n18195) );
  INV_X1 U16369 ( .A(n18195), .ZN(n19334) );
  NAND2_X1 U16370 ( .A1(n17334), .A2(n19334), .ZN(n14529) );
  NOR2_X1 U16371 ( .A1(n17675), .A2(n14529), .ZN(n19340) );
  OAI21_X1 U16372 ( .B1(n14506), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14505), .ZN(n19342) );
  NAND2_X1 U16373 ( .A1(n19340), .A2(n19342), .ZN(n19353) );
  NOR2_X1 U16374 ( .A1(n19355), .A2(n19353), .ZN(n19367) );
  INV_X1 U16375 ( .A(n14507), .ZN(n14509) );
  AOI21_X1 U16376 ( .B1(n19370), .B2(n14509), .A(n14508), .ZN(n17647) );
  INV_X1 U16377 ( .A(n17647), .ZN(n19368) );
  NAND2_X1 U16378 ( .A1(n19367), .A2(n19368), .ZN(n17307) );
  NOR2_X1 U16379 ( .A1(n14510), .A2(n17307), .ZN(n19388) );
  NAND2_X1 U16380 ( .A1(n19388), .A2(n19387), .ZN(n19400) );
  OAI21_X1 U16381 ( .B1(n14511), .B2(n19400), .A(n14531), .ZN(n19416) );
  NAND2_X1 U16382 ( .A1(n19417), .A2(n19416), .ZN(n19415) );
  NAND2_X1 U16383 ( .A1(n14531), .A2(n19415), .ZN(n17294) );
  OR2_X1 U16384 ( .A1(n14512), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14513) );
  NAND2_X1 U16385 ( .A1(n14514), .A2(n14513), .ZN(n17603) );
  NAND2_X1 U16386 ( .A1(n11185), .A2(n19425), .ZN(n19435) );
  INV_X1 U16387 ( .A(n14518), .ZN(n14517) );
  NAND2_X1 U16388 ( .A1(n14515), .A2(n17574), .ZN(n14516) );
  NAND2_X1 U16389 ( .A1(n14517), .A2(n14516), .ZN(n19436) );
  NAND2_X1 U16390 ( .A1(n11185), .A2(n19434), .ZN(n17266) );
  OR2_X1 U16391 ( .A1(n14518), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14519) );
  NAND2_X1 U16392 ( .A1(n14520), .A2(n14519), .ZN(n17558) );
  INV_X1 U16393 ( .A(n14521), .ZN(n19465) );
  NAND2_X1 U16394 ( .A1(n11185), .A2(n19463), .ZN(n19482) );
  INV_X1 U16395 ( .A(n19518), .ZN(n19481) );
  NAND2_X1 U16396 ( .A1(n19481), .A2(n11185), .ZN(n14528) );
  NOR2_X1 U16397 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14524) );
  NOR4_X1 U16398 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14523) );
  NAND4_X1 U16399 ( .A1(n14524), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14523), .ZN(n14527) );
  NOR2_X1 U16400 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14527), .ZN(n19565)
         );
  INV_X1 U16401 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20935) );
  INV_X1 U16402 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22785) );
  NOR4_X1 U16403 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20935), .A4(n22785), .ZN(n14526) );
  NOR4_X1 U16404 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14525) );
  NAND3_X1 U16405 ( .A1(n14954), .A2(n14526), .A3(n14525), .ZN(U214) );
  OR2_X1 U16406 ( .A1(n15507), .A2(n14527), .ZN(n20869) );
  INV_X2 U16407 ( .A(U214), .ZN(n20920) );
  AOI211_X1 U16408 ( .C1(n17675), .C2(n14529), .A(n19340), .B(n14528), .ZN(
        n14541) );
  OAI22_X1 U16409 ( .A1(n19409), .A2(n14530), .B1(n19443), .B2(n17673), .ZN(
        n14540) );
  INV_X1 U16410 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n18295) );
  NAND2_X1 U16411 ( .A1(n19481), .A2(n11184), .ZN(n17330) );
  AOI22_X1 U16412 ( .A1(n14532), .A2(n19473), .B1(n17675), .B2(n17354), .ZN(
        n14533) );
  OAI211_X1 U16413 ( .C1(n18295), .C2(n19371), .A(n14533), .B(n14452), .ZN(
        n14539) );
  NAND2_X1 U16414 ( .A1(n14534), .A2(n14535), .ZN(n14536) );
  NAND2_X1 U16415 ( .A1(n11382), .A2(n14536), .ZN(n17911) );
  XNOR2_X1 U16416 ( .A(n14537), .B(n16389), .ZN(n20013) );
  OAI22_X1 U16417 ( .A1(n17911), .A2(n19477), .B1(n20013), .B2(n19475), .ZN(
        n14538) );
  OR4_X1 U16418 ( .A1(n14541), .A2(n14540), .A3(n14539), .A4(n14538), .ZN(
        P2_U2840) );
  INV_X1 U16419 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n14542) );
  OAI21_X1 U16420 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n14542), .A(HOLD), .ZN(
        n14546) );
  INV_X1 U16421 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n14552) );
  OAI21_X1 U16422 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n14552), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n14553) );
  OAI21_X1 U16423 ( .B1(n14552), .B2(n14542), .A(n14546), .ZN(n14543) );
  INV_X1 U16424 ( .A(NA), .ZN(n22452) );
  NAND4_X1 U16425 ( .A1(n22389), .A2(P1_STATE_REG_0__SCAN_IN), .A3(n14543), 
        .A4(n22452), .ZN(n14545) );
  OAI21_X1 U16426 ( .B1(n14552), .B2(n22129), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n22422) );
  OAI211_X1 U16427 ( .C1(n22452), .C2(P1_STATE_REG_1__SCAN_IN), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n22422), .ZN(n14544) );
  OAI211_X1 U16428 ( .C1(n14546), .C2(n14553), .A(n14545), .B(n14544), .ZN(
        P1_U3196) );
  NAND2_X1 U16429 ( .A1(HOLD), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22423) );
  NAND2_X1 U16430 ( .A1(HOLD), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U16431 ( .A1(n14547), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n22425) );
  INV_X1 U16432 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22426) );
  NAND2_X1 U16433 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22389), .ZN(n14548) );
  OAI21_X1 U16434 ( .B1(n22425), .B2(n22426), .A(n14548), .ZN(n14549) );
  INV_X1 U16435 ( .A(n14549), .ZN(n14550) );
  OAI211_X1 U16436 ( .C1(n14551), .C2(n22423), .A(n18155), .B(n14550), .ZN(
        P1_U3195) );
  AND2_X1 U16437 ( .A1(n14553), .A2(n22784), .ZN(n22410) );
  INV_X1 U16438 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20720) );
  OAI221_X1 U16439 ( .B1(n20720), .B2(BS16), .C1(n22426), .C2(BS16), .A(n22410), .ZN(n22408) );
  OAI21_X1 U16440 ( .B1(n22410), .B2(n15972), .A(n22408), .ZN(P1_U2805) );
  INV_X1 U16441 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n14555) );
  INV_X1 U16442 ( .A(n14553), .ZN(n14554) );
  INV_X2 U16443 ( .A(n22784), .ZN(n22787) );
  AOI21_X1 U16444 ( .B1(n14555), .B2(n14554), .A(n22787), .ZN(P1_U2802) );
  INV_X1 U16445 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n14557) );
  OAI21_X1 U16446 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20720), .A(n22426), 
        .ZN(n14556) );
  AOI22_X1 U16447 ( .A1(n14557), .A2(n14556), .B1(n22787), .B2(
        P1_CODEFETCH_REG_SCAN_IN), .ZN(P1_U2804) );
  INV_X1 U16448 ( .A(n19531), .ZN(n19514) );
  NAND2_X1 U16449 ( .A1(n19514), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n14570) );
  OAI22_X1 U16450 ( .A1(NA), .A2(n14570), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n14560) );
  INV_X1 U16451 ( .A(n14560), .ZN(n14558) );
  INV_X1 U16452 ( .A(HOLD), .ZN(n22442) );
  AOI21_X1 U16453 ( .B1(n14558), .B2(n18272), .A(n22442), .ZN(n14559) );
  AOI21_X1 U16454 ( .B1(n14560), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n14559), .ZN(n14563) );
  NAND2_X1 U16455 ( .A1(n14570), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n22433) );
  INV_X1 U16456 ( .A(n22433), .ZN(n14562) );
  INV_X1 U16457 ( .A(n18099), .ZN(n14561) );
  OAI21_X1 U16458 ( .B1(n14561), .B2(n22452), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n22432) );
  OAI22_X1 U16459 ( .A1(n14563), .A2(n18270), .B1(n14562), .B2(n22432), .ZN(
        P2_U3211) );
  NAND2_X1 U16460 ( .A1(n14564), .A2(n19511), .ZN(n14566) );
  OR2_X1 U16461 ( .A1(n12351), .A2(n14566), .ZN(n19276) );
  INV_X1 U16462 ( .A(n19276), .ZN(n19268) );
  INV_X1 U16463 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14568) );
  NOR2_X1 U16464 ( .A1(n20192), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14575) );
  INV_X1 U16465 ( .A(n14575), .ZN(n14567) );
  OAI211_X1 U16466 ( .C1(n19268), .C2(n14568), .A(n14567), .B(n14578), .ZN(
        P2_U2814) );
  NAND2_X1 U16467 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n14574) );
  NOR2_X1 U16468 ( .A1(n22442), .A2(n18272), .ZN(n14573) );
  INV_X1 U16469 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n14569) );
  NOR2_X1 U16470 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n14569), .ZN(n18100) );
  INV_X1 U16471 ( .A(n14570), .ZN(n14571) );
  AOI211_X1 U16472 ( .C1(n18100), .C2(HOLD), .A(n14571), .B(n19252), .ZN(
        n14572) );
  OAI21_X1 U16473 ( .B1(n14574), .B2(n14573), .A(n14572), .ZN(P2_U3210) );
  INV_X1 U16474 ( .A(n12573), .ZN(n14577) );
  INV_X1 U16475 ( .A(n18168), .ZN(n19244) );
  OAI21_X1 U16476 ( .B1(n14575), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19244), 
        .ZN(n14576) );
  OAI21_X1 U16477 ( .B1(n14577), .B2(n19244), .A(n14576), .ZN(P2_U3612) );
  INV_X1 U16478 ( .A(n14578), .ZN(n14580) );
  OAI21_X1 U16479 ( .B1(n19514), .B2(n14578), .A(n14701), .ZN(n14602) );
  INV_X1 U16480 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14582) );
  NOR2_X1 U16481 ( .A1(n12819), .A2(n19514), .ZN(n14579) );
  NAND2_X1 U16482 ( .A1(n14580), .A2(n14579), .ZN(n14702) );
  AOI22_X1 U16483 ( .A1(n15508), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14661), .ZN(n20365) );
  NOR2_X1 U16484 ( .A1(n14702), .A2(n20365), .ZN(n14653) );
  AOI21_X1 U16485 ( .B1(n14687), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14653), .ZN(
        n14581) );
  OAI21_X1 U16486 ( .B1(n14602), .B2(n14582), .A(n14581), .ZN(P2_U2955) );
  INV_X1 U16487 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U16488 ( .A1(n15508), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15507), .ZN(n20414) );
  NOR2_X1 U16489 ( .A1(n14702), .A2(n20414), .ZN(n14676) );
  AOI21_X1 U16490 ( .B1(n14687), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14676), .ZN(
        n14583) );
  OAI21_X1 U16491 ( .B1(n14602), .B2(n14584), .A(n14583), .ZN(P2_U2954) );
  INV_X1 U16492 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14587) );
  INV_X1 U16493 ( .A(n14702), .ZN(n14618) );
  AOI22_X1 U16494 ( .A1(n15508), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15507), .ZN(n20032) );
  INV_X1 U16495 ( .A(n20032), .ZN(n14585) );
  NAND2_X1 U16496 ( .A1(n14618), .A2(n14585), .ZN(n14612) );
  NAND2_X1 U16497 ( .A1(n14687), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n14586) );
  OAI211_X1 U16498 ( .C1(n14602), .C2(n14587), .A(n14612), .B(n14586), .ZN(
        P2_U2975) );
  INV_X1 U16499 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n14592) );
  INV_X1 U16500 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20894) );
  OR2_X1 U16501 ( .A1(n15507), .A2(n20894), .ZN(n14589) );
  NAND2_X1 U16502 ( .A1(n15507), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14588) );
  AND2_X1 U16503 ( .A1(n14589), .A2(n14588), .ZN(n20020) );
  INV_X1 U16504 ( .A(n20020), .ZN(n14590) );
  NAND2_X1 U16505 ( .A1(n14618), .A2(n14590), .ZN(n14604) );
  NAND2_X1 U16506 ( .A1(n14687), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n14591) );
  OAI211_X1 U16507 ( .C1(n14602), .C2(n14592), .A(n14604), .B(n14591), .ZN(
        P2_U2979) );
  INV_X1 U16508 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n14595) );
  INV_X1 U16509 ( .A(n20014), .ZN(n14593) );
  NAND2_X1 U16510 ( .A1(n14618), .A2(n14593), .ZN(n14606) );
  NAND2_X1 U16511 ( .A1(n14687), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n14594) );
  OAI211_X1 U16512 ( .C1(n14602), .C2(n14595), .A(n14606), .B(n14594), .ZN(
        P2_U2981) );
  INV_X1 U16513 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n14601) );
  INV_X1 U16514 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14596) );
  OR2_X1 U16515 ( .A1(n15507), .A2(n14596), .ZN(n14598) );
  NAND2_X1 U16516 ( .A1(n15507), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14597) );
  AND2_X1 U16517 ( .A1(n14598), .A2(n14597), .ZN(n20026) );
  INV_X1 U16518 ( .A(n20026), .ZN(n14599) );
  NAND2_X1 U16519 ( .A1(n14618), .A2(n14599), .ZN(n14610) );
  NAND2_X1 U16520 ( .A1(n14687), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n14600) );
  OAI211_X1 U16521 ( .C1(n14602), .C2(n14601), .A(n14610), .B(n14600), .ZN(
        P2_U2977) );
  INV_X1 U16522 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18260) );
  NAND2_X1 U16523 ( .A1(n14636), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14603) );
  MUX2_X1 U16524 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n15507), .Z(n20023) );
  NAND2_X1 U16525 ( .A1(n14618), .A2(n20023), .ZN(n14608) );
  OAI211_X1 U16526 ( .C1(n18260), .C2(n14701), .A(n14603), .B(n14608), .ZN(
        P2_U2978) );
  INV_X1 U16527 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n17460) );
  NAND2_X1 U16528 ( .A1(n14636), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14605) );
  OAI211_X1 U16529 ( .C1(n14701), .C2(n17460), .A(n14605), .B(n14604), .ZN(
        P2_U2964) );
  NAND2_X1 U16530 ( .A1(n14636), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14607) );
  OAI211_X1 U16531 ( .C1(n14701), .C2(n14685), .A(n14607), .B(n14606), .ZN(
        P2_U2966) );
  INV_X1 U16532 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14856) );
  NAND2_X1 U16533 ( .A1(n14636), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14609) );
  OAI211_X1 U16534 ( .C1(n14856), .C2(n14701), .A(n14609), .B(n14608), .ZN(
        P2_U2963) );
  INV_X1 U16535 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n17476) );
  NAND2_X1 U16536 ( .A1(n14636), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14611) );
  OAI211_X1 U16537 ( .C1(n14701), .C2(n17476), .A(n14611), .B(n14610), .ZN(
        P2_U2962) );
  INV_X1 U16538 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n17491) );
  NAND2_X1 U16539 ( .A1(n14636), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14613) );
  OAI211_X1 U16540 ( .C1(n14701), .C2(n17491), .A(n14613), .B(n14612), .ZN(
        P2_U2960) );
  INV_X1 U16541 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n17454) );
  NAND2_X1 U16542 ( .A1(n14636), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14619) );
  INV_X1 U16543 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14614) );
  OR2_X1 U16544 ( .A1(n15507), .A2(n14614), .ZN(n14616) );
  NAND2_X1 U16545 ( .A1(n14661), .A2(BUF2_REG_13__SCAN_IN), .ZN(n14615) );
  AND2_X1 U16546 ( .A1(n14616), .A2(n14615), .ZN(n20019) );
  INV_X1 U16547 ( .A(n20019), .ZN(n14617) );
  NAND2_X1 U16548 ( .A1(n14618), .A2(n14617), .ZN(n14689) );
  OAI211_X1 U16549 ( .C1(n14701), .C2(n17454), .A(n14619), .B(n14689), .ZN(
        P2_U2965) );
  INV_X1 U16550 ( .A(n22534), .ZN(n22494) );
  AND2_X1 U16551 ( .A1(n22494), .A2(n18164), .ZN(n16461) );
  NOR2_X1 U16552 ( .A1(n16461), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14627)
         );
  NAND2_X1 U16553 ( .A1(n16472), .A2(n14840), .ZN(n14621) );
  NOR2_X1 U16554 ( .A1(n16465), .A2(n22406), .ZN(n14622) );
  OAI21_X1 U16555 ( .B1(n13166), .B2(n14625), .A(n22127), .ZN(n14626) );
  OAI21_X1 U16556 ( .B1(n14627), .B2(n22127), .A(n14626), .ZN(P1_U3487) );
  OAI21_X1 U16557 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19260), .A(
        n14628), .ZN(n19494) );
  INV_X1 U16558 ( .A(n19494), .ZN(n14632) );
  OAI21_X1 U16559 ( .B1(n14630), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14629), .ZN(n19509) );
  NAND2_X1 U16560 ( .A1(n12603), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19506) );
  OAI21_X1 U16561 ( .B1(n18185), .B2(n19509), .A(n19506), .ZN(n14631) );
  AOI21_X1 U16562 ( .B1(n18200), .B2(n14632), .A(n14631), .ZN(n14635) );
  OAI21_X1 U16563 ( .B1(n18174), .B2(n14633), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14634) );
  OAI211_X1 U16564 ( .C1(n18190), .C2(n15304), .A(n14635), .B(n14634), .ZN(
        P2_U3014) );
  INV_X1 U16565 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14638) );
  AOI22_X1 U16566 ( .A1(n15508), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14661), .ZN(n20213) );
  NOR2_X1 U16567 ( .A1(n14702), .A2(n20213), .ZN(n14673) );
  AOI21_X1 U16568 ( .B1(n14687), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14673), .ZN(
        n14637) );
  OAI21_X1 U16569 ( .B1(n14704), .B2(n14638), .A(n14637), .ZN(P2_U2973) );
  INV_X1 U16570 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16571 ( .A1(n15508), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15507), .ZN(n20466) );
  NOR2_X1 U16572 ( .A1(n14702), .A2(n20466), .ZN(n14641) );
  AOI21_X1 U16573 ( .B1(n14687), .B2(P2_EAX_REG_1__SCAN_IN), .A(n14641), .ZN(
        n14639) );
  OAI21_X1 U16574 ( .B1(n14704), .B2(n14640), .A(n14639), .ZN(P2_U2968) );
  INV_X1 U16575 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14643) );
  AOI21_X1 U16576 ( .B1(n14687), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14641), .ZN(
        n14642) );
  OAI21_X1 U16577 ( .B1(n14704), .B2(n14643), .A(n14642), .ZN(P2_U2953) );
  INV_X1 U16578 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n14645) );
  AOI22_X1 U16579 ( .A1(n15508), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n15507), .ZN(n20031) );
  NOR2_X1 U16580 ( .A1(n14702), .A2(n20031), .ZN(n14670) );
  AOI21_X1 U16581 ( .B1(n14687), .B2(P2_EAX_REG_25__SCAN_IN), .A(n14670), .ZN(
        n14644) );
  OAI21_X1 U16582 ( .B1(n14704), .B2(n14645), .A(n14644), .ZN(P2_U2961) );
  INV_X1 U16583 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14647) );
  AOI22_X1 U16584 ( .A1(n15508), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14661), .ZN(n20268) );
  NOR2_X1 U16585 ( .A1(n14702), .A2(n20268), .ZN(n14648) );
  AOI21_X1 U16586 ( .B1(n14687), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14648), .ZN(
        n14646) );
  OAI21_X1 U16587 ( .B1(n14704), .B2(n14647), .A(n14646), .ZN(P2_U2972) );
  INV_X1 U16588 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14650) );
  AOI21_X1 U16589 ( .B1(n14687), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14648), .ZN(
        n14649) );
  OAI21_X1 U16590 ( .B1(n14704), .B2(n14650), .A(n14649), .ZN(P2_U2957) );
  INV_X1 U16591 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14652) );
  AOI22_X1 U16592 ( .A1(n15508), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14661), .ZN(n20317) );
  NOR2_X1 U16593 ( .A1(n14702), .A2(n20317), .ZN(n14656) );
  AOI21_X1 U16594 ( .B1(n14687), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14656), .ZN(
        n14651) );
  OAI21_X1 U16595 ( .B1(n14704), .B2(n14652), .A(n14651), .ZN(P2_U2956) );
  INV_X1 U16596 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14655) );
  AOI21_X1 U16597 ( .B1(n14687), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14653), .ZN(
        n14654) );
  OAI21_X1 U16598 ( .B1(n14704), .B2(n14655), .A(n14654), .ZN(P2_U2970) );
  INV_X1 U16599 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14658) );
  AOI21_X1 U16600 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n14687), .A(n14656), .ZN(
        n14657) );
  OAI21_X1 U16601 ( .B1(n14704), .B2(n14658), .A(n14657), .ZN(P2_U2971) );
  INV_X1 U16602 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14660) );
  AOI22_X1 U16603 ( .A1(n15508), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14661), .ZN(n20037) );
  NOR2_X1 U16604 ( .A1(n14702), .A2(n20037), .ZN(n14664) );
  AOI21_X1 U16605 ( .B1(n14687), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14664), .ZN(
        n14659) );
  OAI21_X1 U16606 ( .B1(n14704), .B2(n14660), .A(n14659), .ZN(P2_U2974) );
  INV_X1 U16607 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14663) );
  AOI22_X1 U16608 ( .A1(n15508), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14661), .ZN(n20526) );
  NOR2_X1 U16609 ( .A1(n14702), .A2(n20526), .ZN(n14667) );
  AOI21_X1 U16610 ( .B1(n14687), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14667), .ZN(
        n14662) );
  OAI21_X1 U16611 ( .B1(n14704), .B2(n14663), .A(n14662), .ZN(P2_U2952) );
  INV_X1 U16612 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14666) );
  AOI21_X1 U16613 ( .B1(n14687), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14664), .ZN(
        n14665) );
  OAI21_X1 U16614 ( .B1(n14704), .B2(n14666), .A(n14665), .ZN(P2_U2959) );
  INV_X1 U16615 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14669) );
  AOI21_X1 U16616 ( .B1(n14687), .B2(P2_EAX_REG_0__SCAN_IN), .A(n14667), .ZN(
        n14668) );
  OAI21_X1 U16617 ( .B1(n14704), .B2(n14669), .A(n14668), .ZN(P2_U2967) );
  INV_X1 U16618 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n14672) );
  AOI21_X1 U16619 ( .B1(n14687), .B2(P2_EAX_REG_9__SCAN_IN), .A(n14670), .ZN(
        n14671) );
  OAI21_X1 U16620 ( .B1(n14704), .B2(n14672), .A(n14671), .ZN(P2_U2976) );
  INV_X1 U16621 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14675) );
  AOI21_X1 U16622 ( .B1(n14687), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14673), .ZN(
        n14674) );
  OAI21_X1 U16623 ( .B1(n14704), .B2(n14675), .A(n14674), .ZN(P2_U2958) );
  INV_X1 U16624 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14678) );
  AOI21_X1 U16625 ( .B1(n14687), .B2(P2_EAX_REG_2__SCAN_IN), .A(n14676), .ZN(
        n14677) );
  OAI21_X1 U16626 ( .B1(n14704), .B2(n14678), .A(n14677), .ZN(P2_U2969) );
  INV_X1 U16627 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n17549) );
  NOR2_X1 U16628 ( .A1(n14679), .A2(n12351), .ZN(n15292) );
  NAND2_X1 U16629 ( .A1(n15292), .A2(n19511), .ZN(n14680) );
  NAND2_X1 U16630 ( .A1(n14680), .A2(n14701), .ZN(n14681) );
  NAND2_X1 U16631 ( .A1(n18238), .A2(n14682), .ZN(n14862) );
  NOR2_X1 U16632 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18205), .ZN(n18257) );
  AOI22_X1 U16633 ( .A1(n18257), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14683) );
  OAI21_X1 U16634 ( .B1(n17549), .B2(n14862), .A(n14683), .ZN(P2_U2934) );
  AOI22_X1 U16635 ( .A1(n18257), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14684) );
  OAI21_X1 U16636 ( .B1(n14685), .B2(n14862), .A(n14684), .ZN(P2_U2921) );
  INV_X1 U16637 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U16638 ( .A1(n18257), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14686) );
  OAI21_X1 U16639 ( .B1(n17538), .B2(n14862), .A(n14686), .ZN(P2_U2933) );
  INV_X1 U16640 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U16641 ( .A1(n14687), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14688) );
  OAI211_X1 U16642 ( .C1(n14704), .C2(n14690), .A(n14689), .B(n14688), .ZN(
        P2_U2980) );
  INV_X1 U16643 ( .A(n17360), .ZN(n14833) );
  NOR2_X1 U16644 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  XOR2_X1 U16645 ( .A(n14693), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n14831) );
  AOI21_X1 U16646 ( .B1(n14696), .B2(n14695), .A(n14694), .ZN(n14825) );
  INV_X1 U16647 ( .A(n14825), .ZN(n14697) );
  NAND2_X1 U16648 ( .A1(n12603), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14826) );
  OAI21_X1 U16649 ( .B1(n18185), .B2(n14697), .A(n14826), .ZN(n14699) );
  MUX2_X1 U16650 ( .A(n18196), .B(n18174), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14698) );
  AOI211_X1 U16651 ( .C1(n18200), .C2(n14831), .A(n14699), .B(n14698), .ZN(
        n14700) );
  OAI21_X1 U16652 ( .B1(n14833), .B2(n18190), .A(n14700), .ZN(P2_U3013) );
  INV_X1 U16653 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14703) );
  AOI22_X1 U16654 ( .A1(n15508), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15507), .ZN(n20011) );
  INV_X1 U16655 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n20012) );
  OAI222_X1 U16656 ( .A1(n14704), .A2(n14703), .B1(n14702), .B2(n20011), .C1(
        n14701), .C2(n20012), .ZN(P2_U2982) );
  AND3_X1 U16657 ( .A1(n18156), .A2(n14707), .A3(n14706), .ZN(n14708) );
  AND2_X1 U16658 ( .A1(n14709), .A2(n14708), .ZN(n14711) );
  NAND2_X1 U16659 ( .A1(n14711), .A2(n14710), .ZN(n17228) );
  INV_X1 U16660 ( .A(n17228), .ZN(n17207) );
  NOR2_X1 U16661 ( .A1(n18127), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17219) );
  INV_X1 U16662 ( .A(n17219), .ZN(n17203) );
  INV_X1 U16663 ( .A(n14712), .ZN(n14714) );
  INV_X1 U16664 ( .A(n14713), .ZN(n14717) );
  NAND3_X1 U16665 ( .A1(n14735), .A2(n14714), .A3(n14717), .ZN(n14715) );
  OAI211_X1 U16666 ( .C1(n11222), .C2(n17207), .A(n17203), .B(n14715), .ZN(
        n18129) );
  INV_X1 U16667 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U16668 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n14716), .B2(n22148), .ZN(
        n17211) );
  NAND2_X1 U16669 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17209) );
  NOR2_X1 U16670 ( .A1(n17211), .A2(n17209), .ZN(n14719) );
  NOR3_X1 U16671 ( .A1(n14712), .A2(n14713), .A3(n17230), .ZN(n14718) );
  AOI211_X1 U16672 ( .C1(n18129), .C2(n20865), .A(n14719), .B(n14718), .ZN(
        n14734) );
  INV_X1 U16673 ( .A(n14720), .ZN(n14728) );
  NAND2_X1 U16674 ( .A1(n18127), .A2(n18156), .ZN(n14722) );
  AND2_X1 U16675 ( .A1(n16472), .A2(n14944), .ZN(n14721) );
  NAND3_X1 U16676 ( .A1(n14722), .A2(n22129), .A3(n14721), .ZN(n14726) );
  NOR2_X1 U16677 ( .A1(n14363), .A2(n13153), .ZN(n14723) );
  AOI21_X1 U16678 ( .B1(n16468), .B2(n16466), .A(n14723), .ZN(n14725) );
  AND3_X1 U16679 ( .A1(n14726), .A2(n14725), .A3(n14724), .ZN(n14727) );
  NAND2_X1 U16680 ( .A1(n14728), .A2(n14727), .ZN(n18151) );
  NAND2_X1 U16681 ( .A1(n18151), .A2(n14840), .ZN(n14732) );
  INV_X1 U16682 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22387) );
  NAND2_X1 U16683 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22395) );
  NOR3_X1 U16684 ( .A1(n22387), .A2(n22396), .A3(n22395), .ZN(n14730) );
  NOR2_X1 U16685 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15600), .ZN(n14729) );
  NOR2_X1 U16686 ( .A1(n14730), .A2(n14729), .ZN(n14731) );
  NAND2_X1 U16687 ( .A1(n14732), .A2(n14731), .ZN(n17233) );
  INV_X1 U16688 ( .A(n17233), .ZN(n14738) );
  NAND2_X1 U16689 ( .A1(n14738), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14733) );
  OAI21_X1 U16690 ( .B1(n14734), .B2(n14738), .A(n14733), .ZN(P1_U3473) );
  AOI22_X1 U16691 ( .A1(n11176), .A2(n17228), .B1(n14735), .B2(n18128), .ZN(
        n18126) );
  OAI21_X1 U16692 ( .B1(n18126), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n18164), 
        .ZN(n14736) );
  AOI22_X1 U16693 ( .A1(n14736), .A2(n17209), .B1(n18128), .B2(n22400), .ZN(
        n14739) );
  AOI21_X1 U16694 ( .B1(n17202), .B2(n20865), .A(n14738), .ZN(n14737) );
  OAI22_X1 U16695 ( .A1(n14739), .A2(n14738), .B1(n14737), .B2(n18128), .ZN(
        P1_U3474) );
  INV_X1 U16696 ( .A(n15211), .ZN(n14960) );
  OR2_X1 U16697 ( .A1(n14740), .A2(n14960), .ZN(n14741) );
  XNOR2_X1 U16698 ( .A(n14741), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n22251) );
  INV_X1 U16699 ( .A(n14710), .ZN(n18138) );
  NAND4_X1 U16700 ( .A1(n22251), .A2(n20865), .A3(n18138), .A4(n17233), .ZN(
        n14742) );
  OAI21_X1 U16701 ( .B1(n18150), .B2(n17233), .A(n14742), .ZN(P1_U3468) );
  AND2_X1 U16702 ( .A1(n20165), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14744) );
  OAI211_X1 U16703 ( .C1(n12819), .C2(n14745), .A(n11732), .B(n14744), .ZN(
        n14746) );
  INV_X1 U16704 ( .A(n14746), .ZN(n14747) );
  MUX2_X1 U16705 ( .A(n15304), .B(n11578), .S(n17432), .Z(n14748) );
  OAI21_X1 U16706 ( .B1(n20519), .B2(n17452), .A(n14748), .ZN(P2_U2887) );
  INV_X1 U16707 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20719) );
  NOR2_X1 U16708 ( .A1(n13211), .A2(n22129), .ZN(n14749) );
  NOR2_X2 U16709 ( .A1(n14809), .A2(n15026), .ZN(n14798) );
  INV_X1 U16710 ( .A(n14798), .ZN(n14753) );
  INV_X1 U16711 ( .A(DATAI_15_), .ZN(n15930) );
  NOR2_X1 U16712 ( .A1(n14954), .A2(n15930), .ZN(n14750) );
  AOI21_X1 U16713 ( .B1(n14954), .B2(BUF1_REG_15__SCAN_IN), .A(n14750), .ZN(
        n16778) );
  INV_X1 U16714 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14751) );
  OAI222_X1 U16715 ( .A1(n14808), .A2(n20719), .B1(n14753), .B2(n16778), .C1(
        n14752), .C2(n14751), .ZN(P1_U2967) );
  NAND2_X1 U16716 ( .A1(n14798), .A2(n16779), .ZN(n14792) );
  NAND2_X1 U16717 ( .A1(n14809), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n14754) );
  OAI211_X1 U16718 ( .C1(n16780), .C2(n14808), .A(n14792), .B(n14754), .ZN(
        P1_U2966) );
  MUX2_X1 U16719 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14954), .Z(
        n16790) );
  NAND2_X1 U16720 ( .A1(n14798), .A2(n16790), .ZN(n14773) );
  NAND2_X1 U16721 ( .A1(n14809), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14755) );
  OAI211_X1 U16722 ( .C1(n16792), .C2(n14808), .A(n14773), .B(n14755), .ZN(
        P1_U2963) );
  MUX2_X1 U16723 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14954), .Z(
        n16787) );
  NAND2_X1 U16724 ( .A1(n14798), .A2(n16787), .ZN(n14794) );
  NAND2_X1 U16725 ( .A1(n14809), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14756) );
  OAI211_X1 U16726 ( .C1(n16788), .C2(n14808), .A(n14794), .B(n14756), .ZN(
        P1_U2964) );
  MUX2_X1 U16727 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14954), .Z(
        n16783) );
  NAND2_X1 U16728 ( .A1(n14798), .A2(n16783), .ZN(n14771) );
  NAND2_X1 U16729 ( .A1(n14809), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n14757) );
  OAI211_X1 U16730 ( .C1(n16784), .C2(n14808), .A(n14771), .B(n14757), .ZN(
        P1_U2965) );
  INV_X1 U16731 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20883) );
  NAND2_X1 U16732 ( .A1(n14954), .A2(n20883), .ZN(n14758) );
  OAI21_X1 U16733 ( .B1(n14954), .B2(DATAI_6_), .A(n14758), .ZN(n16736) );
  INV_X1 U16734 ( .A(n16736), .ZN(n14976) );
  NAND2_X1 U16735 ( .A1(n14798), .A2(n14976), .ZN(n14779) );
  NAND2_X1 U16736 ( .A1(n14809), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n14759) );
  OAI211_X1 U16737 ( .C1(n13562), .C2(n14808), .A(n14779), .B(n14759), .ZN(
        P1_U2958) );
  INV_X1 U16738 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20704) );
  MUX2_X1 U16739 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n14954), .Z(
        n16746) );
  NAND2_X1 U16740 ( .A1(n14798), .A2(n16746), .ZN(n14775) );
  NAND2_X1 U16741 ( .A1(n14809), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14760) );
  OAI211_X1 U16742 ( .C1(n20704), .C2(n14808), .A(n14775), .B(n14760), .ZN(
        P1_U2956) );
  MUX2_X1 U16743 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n14954), .Z(
        n16743) );
  NAND2_X1 U16744 ( .A1(n14798), .A2(n16743), .ZN(n14777) );
  NAND2_X1 U16745 ( .A1(n14809), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14761) );
  OAI211_X1 U16746 ( .C1(n15656), .C2(n14808), .A(n14777), .B(n14761), .ZN(
        P1_U2957) );
  MUX2_X1 U16747 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14954), .Z(
        n16724) );
  NAND2_X1 U16748 ( .A1(n14798), .A2(n16724), .ZN(n14803) );
  NAND2_X1 U16749 ( .A1(n14809), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14762) );
  OAI211_X1 U16750 ( .C1(n14808), .C2(n16721), .A(n14803), .B(n14762), .ZN(
        P1_U2946) );
  INV_X1 U16751 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14948) );
  NAND2_X1 U16752 ( .A1(n14784), .A2(DATAI_2_), .ZN(n14764) );
  NAND2_X1 U16753 ( .A1(n14954), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14763) );
  AND2_X1 U16754 ( .A1(n14764), .A2(n14763), .ZN(n14964) );
  INV_X1 U16755 ( .A(n14964), .ZN(n16757) );
  NAND2_X1 U16756 ( .A1(n14798), .A2(n16757), .ZN(n14797) );
  NAND2_X1 U16757 ( .A1(n14809), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14765) );
  OAI211_X1 U16758 ( .C1(n14948), .C2(n14808), .A(n14797), .B(n14765), .ZN(
        P1_U2939) );
  NAND2_X1 U16759 ( .A1(n14784), .A2(DATAI_3_), .ZN(n14767) );
  NAND2_X1 U16760 ( .A1(n14954), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14766) );
  AND2_X1 U16761 ( .A1(n14767), .A2(n14766), .ZN(n15177) );
  INV_X1 U16762 ( .A(n15177), .ZN(n16753) );
  NAND2_X1 U16763 ( .A1(n14798), .A2(n16753), .ZN(n14805) );
  NAND2_X1 U16764 ( .A1(n14809), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14768) );
  OAI211_X1 U16765 ( .C1(n14808), .C2(n15589), .A(n14805), .B(n14768), .ZN(
        P1_U2940) );
  INV_X1 U16766 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20699) );
  MUX2_X1 U16767 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n14954), .Z(
        n16772) );
  NAND2_X1 U16768 ( .A1(n14798), .A2(n16772), .ZN(n14783) );
  NAND2_X1 U16769 ( .A1(n14809), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14769) );
  OAI211_X1 U16770 ( .C1(n20699), .C2(n14808), .A(n14783), .B(n14769), .ZN(
        P1_U2952) );
  INV_X1 U16771 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15577) );
  NAND2_X1 U16772 ( .A1(n14809), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14770) );
  OAI211_X1 U16773 ( .C1(n14808), .C2(n15577), .A(n14771), .B(n14770), .ZN(
        P1_U2950) );
  INV_X1 U16774 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15897) );
  NAND2_X1 U16775 ( .A1(n14809), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14772) );
  OAI211_X1 U16776 ( .C1(n15897), .C2(n14808), .A(n14773), .B(n14772), .ZN(
        P1_U2948) );
  NAND2_X1 U16777 ( .A1(n14809), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14774) );
  OAI211_X1 U16778 ( .C1(n14808), .C2(n15581), .A(n14775), .B(n14774), .ZN(
        P1_U2941) );
  NAND2_X1 U16779 ( .A1(n14809), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14776) );
  OAI211_X1 U16780 ( .C1(n14808), .C2(n15583), .A(n14777), .B(n14776), .ZN(
        P1_U2942) );
  INV_X1 U16781 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n16735) );
  NAND2_X1 U16782 ( .A1(n14809), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14778) );
  OAI211_X1 U16783 ( .C1(n14808), .C2(n16735), .A(n14779), .B(n14778), .ZN(
        P1_U2943) );
  INV_X1 U16784 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15571) );
  INV_X1 U16785 ( .A(DATAI_7_), .ZN(n15942) );
  NAND2_X1 U16786 ( .A1(n14954), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14780) );
  OAI21_X1 U16787 ( .B1(n14954), .B2(n15942), .A(n14780), .ZN(n16731) );
  NAND2_X1 U16788 ( .A1(n14798), .A2(n16731), .ZN(n14807) );
  NAND2_X1 U16789 ( .A1(n14809), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14781) );
  OAI211_X1 U16790 ( .C1(n15571), .C2(n14808), .A(n14807), .B(n14781), .ZN(
        P1_U2944) );
  INV_X1 U16791 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15569) );
  NAND2_X1 U16792 ( .A1(n14809), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14782) );
  OAI211_X1 U16793 ( .C1(n15569), .C2(n14808), .A(n14783), .B(n14782), .ZN(
        P1_U2937) );
  NAND2_X1 U16794 ( .A1(n14784), .A2(DATAI_1_), .ZN(n14786) );
  NAND2_X1 U16795 ( .A1(n14954), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14785) );
  AND2_X1 U16796 ( .A1(n14786), .A2(n14785), .ZN(n16764) );
  INV_X1 U16797 ( .A(n16764), .ZN(n14787) );
  NAND2_X1 U16798 ( .A1(n14798), .A2(n14787), .ZN(n14790) );
  NAND2_X1 U16799 ( .A1(n14809), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14788) );
  OAI211_X1 U16800 ( .C1(n16761), .C2(n14808), .A(n14790), .B(n14788), .ZN(
        P1_U2938) );
  NAND2_X1 U16801 ( .A1(n14809), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14789) );
  OAI211_X1 U16802 ( .C1(n13512), .C2(n14808), .A(n14790), .B(n14789), .ZN(
        P1_U2953) );
  NAND2_X1 U16803 ( .A1(n14809), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14791) );
  OAI211_X1 U16804 ( .C1(n14808), .C2(n15579), .A(n14792), .B(n14791), .ZN(
        P1_U2951) );
  NAND2_X1 U16805 ( .A1(n14809), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14793) );
  OAI211_X1 U16806 ( .C1(n14808), .C2(n15585), .A(n14794), .B(n14793), .ZN(
        P1_U2949) );
  INV_X1 U16807 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n16089) );
  MUX2_X1 U16808 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n14954), .Z(
        n16728) );
  NAND2_X1 U16809 ( .A1(n14798), .A2(n16728), .ZN(n14801) );
  NAND2_X1 U16810 ( .A1(n14809), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14795) );
  OAI211_X1 U16811 ( .C1(n16089), .C2(n14808), .A(n14801), .B(n14795), .ZN(
        P1_U2945) );
  NAND2_X1 U16812 ( .A1(n14809), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14796) );
  OAI211_X1 U16813 ( .C1(n13505), .C2(n14808), .A(n14797), .B(n14796), .ZN(
        P1_U2954) );
  INV_X1 U16814 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15899) );
  MUX2_X1 U16815 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14954), .Z(
        n16718) );
  NAND2_X1 U16816 ( .A1(n14798), .A2(n16718), .ZN(n14811) );
  NAND2_X1 U16817 ( .A1(n14809), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14799) );
  OAI211_X1 U16818 ( .C1(n15899), .C2(n14808), .A(n14811), .B(n14799), .ZN(
        P1_U2947) );
  NAND2_X1 U16819 ( .A1(n14809), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14800) );
  OAI211_X1 U16820 ( .C1(n16297), .C2(n14808), .A(n14801), .B(n14800), .ZN(
        P1_U2960) );
  NAND2_X1 U16821 ( .A1(n14809), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14802) );
  OAI211_X1 U16822 ( .C1(n16339), .C2(n14808), .A(n14803), .B(n14802), .ZN(
        P1_U2961) );
  NAND2_X1 U16823 ( .A1(n14809), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n14804) );
  OAI211_X1 U16824 ( .C1(n13534), .C2(n14808), .A(n14805), .B(n14804), .ZN(
        P1_U2955) );
  NAND2_X1 U16825 ( .A1(n14809), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n14806) );
  OAI211_X1 U16826 ( .C1(n15676), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        P1_U2959) );
  NAND2_X1 U16827 ( .A1(n14809), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14810) );
  OAI211_X1 U16828 ( .C1(n16361), .C2(n14808), .A(n14811), .B(n14810), .ZN(
        P1_U2962) );
  OR2_X1 U16829 ( .A1(n14812), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14813) );
  NAND2_X1 U16830 ( .A1(n13241), .A2(n14813), .ZN(n14874) );
  OR2_X1 U16831 ( .A1(n14814), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14815) );
  NAND2_X1 U16832 ( .A1(n14816), .A2(n14815), .ZN(n15364) );
  OAI21_X1 U16833 ( .B1(n22225), .B2(n17081), .A(n14389), .ZN(n14863) );
  INV_X1 U16834 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14817) );
  OR2_X1 U16835 ( .A1(n16939), .A2(n14817), .ZN(n14875) );
  OAI211_X1 U16836 ( .C1(n22245), .C2(n15364), .A(n14863), .B(n14875), .ZN(
        n14818) );
  INV_X1 U16837 ( .A(n14818), .ZN(n14821) );
  INV_X1 U16838 ( .A(n14864), .ZN(n14819) );
  OAI21_X1 U16839 ( .B1(n14819), .B2(n17165), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14820) );
  OAI211_X1 U16840 ( .C1(n14874), .C2(n22226), .A(n14821), .B(n14820), .ZN(
        P1_U3031) );
  OAI21_X1 U16841 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n20458) );
  AOI22_X1 U16842 ( .A1(n18055), .A2(n14825), .B1(n19500), .B2(n20458), .ZN(
        n14827) );
  OAI211_X1 U16843 ( .C1(n19497), .C2(n14696), .A(n14827), .B(n14826), .ZN(
        n14830) );
  INV_X1 U16844 ( .A(n16415), .ZN(n14828) );
  AOI211_X1 U16845 ( .C1(n14696), .C2(n19496), .A(n14828), .B(n19502), .ZN(
        n14829) );
  AOI211_X1 U16846 ( .C1(n14831), .C2(n14175), .A(n14830), .B(n14829), .ZN(
        n14832) );
  OAI21_X1 U16847 ( .B1(n14833), .B2(n18061), .A(n14832), .ZN(P2_U3045) );
  INV_X1 U16848 ( .A(n20255), .ZN(n18214) );
  NOR2_X1 U16849 ( .A1(n17411), .A2(n14836), .ZN(n14837) );
  AOI21_X1 U16850 ( .B1(n17360), .B2(n17411), .A(n14837), .ZN(n14838) );
  OAI21_X1 U16851 ( .B1(n18214), .B2(n17452), .A(n14838), .ZN(P2_U2886) );
  INV_X1 U16852 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n16393) );
  AOI22_X1 U16853 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n18266), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n18265), .ZN(n14839) );
  OAI21_X1 U16854 ( .B1(n16393), .B2(n14862), .A(n14839), .ZN(P2_U2935) );
  NAND3_X1 U16855 ( .A1(n16468), .A2(n14840), .A3(n16466), .ZN(n14843) );
  OR2_X1 U16856 ( .A1(n14841), .A2(n14866), .ZN(n14842) );
  INV_X1 U16857 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14848) );
  NAND2_X2 U16858 ( .A1(n20830), .A2(n11182), .ZN(n20805) );
  INV_X1 U16859 ( .A(n14844), .ZN(n14847) );
  OAI21_X1 U16860 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(n15369) );
  OAI222_X1 U16861 ( .A1(n15364), .A2(n20820), .B1(n14848), .B2(n20830), .C1(
        n20805), .C2(n15369), .ZN(P1_U2872) );
  INV_X1 U16862 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n17523) );
  AOI22_X1 U16863 ( .A1(n18266), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14849) );
  OAI21_X1 U16864 ( .B1(n17523), .B2(n14862), .A(n14849), .ZN(P2_U2931) );
  AOI22_X1 U16865 ( .A1(n18266), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14850) );
  OAI21_X1 U16866 ( .B1(n17491), .B2(n14862), .A(n14850), .ZN(P2_U2927) );
  INV_X1 U16867 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U16868 ( .A1(n18266), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14851) );
  OAI21_X1 U16869 ( .B1(n17497), .B2(n14862), .A(n14851), .ZN(P2_U2928) );
  INV_X1 U16870 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n17506) );
  AOI22_X1 U16871 ( .A1(n18266), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14852) );
  OAI21_X1 U16872 ( .B1(n17506), .B2(n14862), .A(n14852), .ZN(P2_U2929) );
  AOI22_X1 U16873 ( .A1(n18266), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14853) );
  OAI21_X1 U16874 ( .B1(n17454), .B2(n14862), .A(n14853), .ZN(P2_U2922) );
  AOI22_X1 U16875 ( .A1(n18266), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14854) );
  OAI21_X1 U16876 ( .B1(n17460), .B2(n14862), .A(n14854), .ZN(P2_U2923) );
  AOI22_X1 U16877 ( .A1(n18266), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14855) );
  OAI21_X1 U16878 ( .B1(n14856), .B2(n14862), .A(n14855), .ZN(P2_U2924) );
  AOI22_X1 U16879 ( .A1(n18266), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14857) );
  OAI21_X1 U16880 ( .B1(n17476), .B2(n14862), .A(n14857), .ZN(P2_U2925) );
  INV_X1 U16881 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U16882 ( .A1(n18266), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14858) );
  OAI21_X1 U16883 ( .B1(n17485), .B2(n14862), .A(n14858), .ZN(P2_U2926) );
  INV_X1 U16884 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14860) );
  AOI22_X1 U16885 ( .A1(n18266), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14859) );
  OAI21_X1 U16886 ( .B1(n14860), .B2(n14862), .A(n14859), .ZN(P2_U2930) );
  INV_X1 U16887 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n17529) );
  AOI22_X1 U16888 ( .A1(n18257), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14861) );
  OAI21_X1 U16889 ( .B1(n17529), .B2(n14862), .A(n14861), .ZN(P2_U2932) );
  AOI21_X1 U16890 ( .B1(n14864), .B2(n14863), .A(n22148), .ZN(n14869) );
  INV_X1 U16891 ( .A(n17054), .ZN(n17114) );
  NOR3_X1 U16892 ( .A1(n17114), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14865), .ZN(n14868) );
  INV_X1 U16893 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20722) );
  NOR2_X1 U16894 ( .A1(n16939), .A2(n20722), .ZN(n14886) );
  XNOR2_X1 U16895 ( .A(n15463), .B(n14866), .ZN(n14896) );
  NOR2_X1 U16896 ( .A1(n22245), .A2(n14896), .ZN(n14867) );
  NOR4_X1 U16897 ( .A1(n14869), .A2(n14868), .A3(n14886), .A4(n14867), .ZN(
        n14873) );
  OR2_X1 U16898 ( .A1(n14870), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14889) );
  NAND3_X1 U16899 ( .A1(n14889), .A2(n14871), .A3(n22239), .ZN(n14872) );
  NAND2_X1 U16900 ( .A1(n14873), .A2(n14872), .ZN(P1_U3030) );
  INV_X1 U16901 ( .A(n14874), .ZN(n14880) );
  INV_X1 U16902 ( .A(n14875), .ZN(n14879) );
  INV_X1 U16903 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14876) );
  AOI21_X1 U16904 ( .B1(n16966), .B2(n14877), .A(n14876), .ZN(n14878) );
  AOI211_X1 U16905 ( .C1(n14880), .C2(n20853), .A(n14879), .B(n14878), .ZN(
        n14881) );
  OAI21_X1 U16906 ( .B1(n16972), .B2(n15369), .A(n14881), .ZN(P1_U2999) );
  INV_X1 U16907 ( .A(n16772), .ZN(n14883) );
  OAI222_X1 U16908 ( .A1(n16794), .A2(n14883), .B1(n16791), .B2(n20699), .C1(
        n16782), .C2(n15369), .ZN(P1_U2904) );
  OAI21_X1 U16909 ( .B1(n14885), .B2(n14884), .A(n14935), .ZN(n15471) );
  AOI21_X1 U16910 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14886), .ZN(n14887) );
  OAI21_X1 U16911 ( .B1(n20856), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14887), .ZN(n14888) );
  INV_X1 U16912 ( .A(n14888), .ZN(n14891) );
  NAND3_X1 U16913 ( .A1(n14889), .A2(n14871), .A3(n20853), .ZN(n14890) );
  OAI211_X1 U16914 ( .C1(n15471), .C2(n16972), .A(n14891), .B(n14890), .ZN(
        P1_U2998) );
  MUX2_X1 U16915 ( .A(n16440), .B(n14894), .S(n17432), .Z(n14895) );
  OAI21_X1 U16916 ( .B1(n20409), .B2(n17452), .A(n14895), .ZN(P2_U2885) );
  OAI222_X1 U16917 ( .A1(n15471), .A2(n16782), .B1(n16794), .B2(n16764), .C1(
        n16791), .C2(n13512), .ZN(P1_U2903) );
  OAI222_X1 U16918 ( .A1(n14896), .A2(n20820), .B1(n14248), .B2(n20830), .C1(
        n15471), .C2(n20805), .ZN(P1_U2871) );
  NOR2_X1 U16919 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22401) );
  INV_X1 U16920 ( .A(n22401), .ZN(n18159) );
  INV_X1 U16921 ( .A(n14897), .ZN(n14898) );
  OAI21_X1 U16922 ( .B1(n14898), .B2(n14712), .A(n18150), .ZN(n14899) );
  NAND2_X1 U16923 ( .A1(n14899), .A2(n22387), .ZN(n17193) );
  OR2_X1 U16924 ( .A1(n22396), .A2(n22395), .ZN(n14900) );
  AOI21_X1 U16925 ( .B1(n17193), .B2(n22387), .A(n14900), .ZN(n14901) );
  OR2_X1 U16926 ( .A1(n15139), .A2(n14901), .ZN(n18165) );
  NAND2_X1 U16927 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15600), .ZN(n17195) );
  NAND2_X1 U16928 ( .A1(n18165), .A2(n17195), .ZN(n16459) );
  NAND2_X1 U16929 ( .A1(n18165), .A2(n22494), .ZN(n16454) );
  NAND2_X1 U16930 ( .A1(n11223), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22482) );
  XNOR2_X1 U16931 ( .A(n14902), .B(n22482), .ZN(n14904) );
  OAI222_X1 U16932 ( .A1(n16459), .A2(n17208), .B1(n18165), .B2(n18135), .C1(
        n16454), .C2(n14904), .ZN(P1_U3476) );
  OR2_X1 U16933 ( .A1(n14907), .A2(n14906), .ZN(n14908) );
  NAND2_X1 U16934 ( .A1(n14905), .A2(n14908), .ZN(n20313) );
  OR2_X1 U16935 ( .A1(n14910), .A2(n14909), .ZN(n14911) );
  AND2_X1 U16936 ( .A1(n14911), .A2(n14915), .ZN(n18170) );
  INV_X1 U16937 ( .A(n18170), .ZN(n19275) );
  NOR2_X1 U16938 ( .A1(n19275), .A2(n17432), .ZN(n14912) );
  AOI21_X1 U16939 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n17432), .A(n14912), .ZN(
        n14913) );
  OAI21_X1 U16940 ( .B1(n20313), .B2(n17452), .A(n14913), .ZN(P2_U2883) );
  XOR2_X1 U16941 ( .A(n14905), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14920)
         );
  AOI21_X1 U16942 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14917) );
  INV_X1 U16943 ( .A(n14917), .ZN(n16331) );
  MUX2_X1 U16944 ( .A(n14918), .B(n16331), .S(n17411), .Z(n14919) );
  OAI21_X1 U16945 ( .B1(n14920), .B2(n17452), .A(n14919), .ZN(P2_U2882) );
  NOR2_X1 U16946 ( .A1(n14905), .A2(n11621), .ZN(n14922) );
  OAI211_X1 U16947 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14922), .A(
        n14921), .B(n17419), .ZN(n14927) );
  OAI21_X1 U16948 ( .B1(n14924), .B2(n14914), .A(n14923), .ZN(n19292) );
  INV_X1 U16949 ( .A(n19292), .ZN(n14925) );
  NAND2_X1 U16950 ( .A1(n14925), .A2(n17411), .ZN(n14926) );
  OAI211_X1 U16951 ( .C1(n17411), .C2(n12209), .A(n14927), .B(n14926), .ZN(
        P2_U2881) );
  XOR2_X1 U16952 ( .A(n14921), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14932)
         );
  AOI21_X1 U16953 ( .B1(n14929), .B2(n14923), .A(n14928), .ZN(n14930) );
  INV_X1 U16954 ( .A(n14930), .ZN(n18043) );
  MUX2_X1 U16955 ( .A(n12211), .B(n18043), .S(n17411), .Z(n14931) );
  OAI21_X1 U16956 ( .B1(n14932), .B2(n17452), .A(n14931), .ZN(P2_U2880) );
  INV_X1 U16957 ( .A(n14933), .ZN(n14934) );
  AOI21_X1 U16958 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n15019) );
  INV_X1 U16959 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20724) );
  NOR2_X1 U16960 ( .A1(n16939), .A2(n20724), .ZN(n22154) );
  AOI21_X1 U16961 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n22154), .ZN(n14937) );
  OAI21_X1 U16962 ( .B1(n20856), .B2(n15020), .A(n14937), .ZN(n14938) );
  AOI21_X1 U16963 ( .B1(n15019), .B2(n20860), .A(n14938), .ZN(n14942) );
  OR2_X1 U16964 ( .A1(n14940), .A2(n14939), .ZN(n22150) );
  NAND3_X1 U16965 ( .A1(n22150), .A2(n22149), .A3(n20853), .ZN(n14941) );
  NAND2_X1 U16966 ( .A1(n14942), .A2(n14941), .ZN(P1_U2997) );
  NAND2_X1 U16967 ( .A1(n14943), .A2(n14808), .ZN(n14945) );
  NAND2_X1 U16968 ( .A1(n20697), .A2(n15025), .ZN(n15588) );
  NOR2_X1 U16969 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22395), .ZN(n20708) );
  NOR2_X4 U16970 ( .A1(n20697), .A2(n22130), .ZN(n20711) );
  AOI22_X1 U16971 ( .A1(n20708), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14946) );
  OAI21_X1 U16972 ( .B1(n16761), .B2(n15588), .A(n14946), .ZN(P1_U2919) );
  AOI22_X1 U16973 ( .A1(n22130), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14947) );
  OAI21_X1 U16974 ( .B1(n14948), .B2(n15588), .A(n14947), .ZN(P1_U2918) );
  INV_X1 U16975 ( .A(n15019), .ZN(n14953) );
  OAI21_X1 U16976 ( .B1(n14950), .B2(n14949), .A(n15373), .ZN(n22152) );
  INV_X1 U16977 ( .A(n22152), .ZN(n14951) );
  AOI22_X1 U16978 ( .A1(n14951), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14952) );
  OAI21_X1 U16979 ( .B1(n14953), .B2(n20805), .A(n14952), .ZN(P1_U2870) );
  OAI222_X1 U16980 ( .A1(n14953), .A2(n16782), .B1(n16794), .B2(n14964), .C1(
        n16791), .C2(n13505), .ZN(P1_U2902) );
  INV_X1 U16981 ( .A(DATAI_26_), .ZN(n14956) );
  NAND2_X1 U16982 ( .A1(n14954), .A2(n20860), .ZN(n15137) );
  INV_X1 U16983 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20922) );
  OR2_X1 U16984 ( .A1(n15137), .A2(n20922), .ZN(n14955) );
  INV_X1 U16985 ( .A(n22602), .ZN(n15444) );
  INV_X1 U16986 ( .A(n15079), .ZN(n14957) );
  INV_X1 U16987 ( .A(DATAI_18_), .ZN(n14959) );
  INV_X1 U16988 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20905) );
  OR2_X1 U16989 ( .A1(n15137), .A2(n20905), .ZN(n14958) );
  OAI21_X1 U16990 ( .B1(n15138), .B2(n14959), .A(n14958), .ZN(n22596) );
  NOR2_X1 U16991 ( .A1(n17208), .A2(n14960), .ZN(n22538) );
  INV_X1 U16992 ( .A(n14961), .ZN(n14962) );
  NAND2_X1 U16993 ( .A1(n14962), .A2(n11176), .ZN(n22484) );
  INV_X1 U16994 ( .A(n22484), .ZN(n15213) );
  INV_X1 U16995 ( .A(n15005), .ZN(n22774) );
  AOI21_X1 U16996 ( .B1(n22538), .B2(n15213), .A(n22774), .ZN(n14968) );
  NOR2_X1 U16997 ( .A1(n15681), .A2(n22505), .ZN(n14970) );
  INV_X1 U16998 ( .A(n14970), .ZN(n14963) );
  OAI22_X1 U16999 ( .A1(n14968), .A2(n22534), .B1(n14963), .B2(n22489), .ZN(
        n22776) );
  INV_X1 U17000 ( .A(n22776), .ZN(n15006) );
  NOR2_X1 U17001 ( .A1(n15602), .A2(n14964), .ZN(n17236) );
  NOR2_X1 U17002 ( .A1(n15141), .A2(n14966), .ZN(n22595) );
  INV_X1 U17003 ( .A(n22595), .ZN(n22599) );
  OAI22_X1 U17004 ( .A1(n15006), .A2(n22605), .B1(n15005), .B2(n22599), .ZN(
        n14967) );
  AOI21_X1 U17005 ( .B1(n22778), .B2(n22596), .A(n14967), .ZN(n14972) );
  OAI211_X1 U17006 ( .C1(n15081), .C2(n22482), .A(n22494), .B(n14968), .ZN(
        n14969) );
  OAI211_X1 U17007 ( .C1(n22494), .C2(n14970), .A(n14969), .B(n22492), .ZN(
        n22779) );
  NAND2_X1 U17008 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14971) );
  OAI211_X1 U17009 ( .C1(n15444), .C2(n22782), .A(n14972), .B(n14971), .ZN(
        P1_U3155) );
  INV_X1 U17010 ( .A(DATAI_30_), .ZN(n14974) );
  INV_X1 U17011 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20930) );
  OR2_X1 U17012 ( .A1(n15137), .A2(n20930), .ZN(n14973) );
  OAI21_X2 U17013 ( .B1(n15138), .B2(n14974), .A(n14973), .ZN(n22709) );
  INV_X1 U17014 ( .A(n22709), .ZN(n22680) );
  INV_X1 U17015 ( .A(DATAI_22_), .ZN(n14975) );
  INV_X1 U17016 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20913) );
  OAI22_X1 U17017 ( .A1(n14975), .A2(n15138), .B1(n20913), .B2(n15137), .ZN(
        n22698) );
  NAND2_X1 U17018 ( .A1(n15139), .A2(n14976), .ZN(n22706) );
  OAI22_X1 U17019 ( .A1(n15006), .A2(n22706), .B1(n15005), .B2(n22705), .ZN(
        n14978) );
  AOI21_X1 U17020 ( .B1(n22778), .B2(n22698), .A(n14978), .ZN(n14980) );
  NAND2_X1 U17021 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14979) );
  OAI211_X1 U17022 ( .C1(n22680), .C2(n22782), .A(n14980), .B(n14979), .ZN(
        P1_U3159) );
  INV_X1 U17023 ( .A(DATAI_27_), .ZN(n14982) );
  INV_X1 U17024 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20924) );
  OR2_X1 U17025 ( .A1(n15137), .A2(n20924), .ZN(n14981) );
  INV_X1 U17026 ( .A(n22624), .ZN(n15440) );
  INV_X1 U17027 ( .A(DATAI_19_), .ZN(n14984) );
  INV_X1 U17028 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20907) );
  OR2_X1 U17029 ( .A1(n15137), .A2(n20907), .ZN(n14983) );
  OAI21_X1 U17030 ( .B1(n15138), .B2(n14984), .A(n14983), .ZN(n22618) );
  NOR2_X1 U17031 ( .A1(n15602), .A2(n15177), .ZN(n17244) );
  NOR2_X1 U17032 ( .A1(n15141), .A2(n14249), .ZN(n22617) );
  INV_X1 U17033 ( .A(n22617), .ZN(n22621) );
  OAI22_X1 U17034 ( .A1(n15006), .A2(n22627), .B1(n15005), .B2(n22621), .ZN(
        n14985) );
  AOI21_X1 U17035 ( .B1(n22778), .B2(n22618), .A(n14985), .ZN(n14987) );
  NAND2_X1 U17036 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14986) );
  OAI211_X1 U17037 ( .C1(n15440), .C2(n22782), .A(n14987), .B(n14986), .ZN(
        P1_U3156) );
  INV_X1 U17038 ( .A(DATAI_28_), .ZN(n14989) );
  INV_X1 U17039 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20926) );
  OR2_X1 U17040 ( .A1(n15137), .A2(n20926), .ZN(n14988) );
  OAI21_X1 U17041 ( .B1(n15138), .B2(n14989), .A(n14988), .ZN(n22646) );
  INV_X1 U17042 ( .A(n22646), .ZN(n22630) );
  INV_X1 U17043 ( .A(DATAI_20_), .ZN(n14991) );
  INV_X1 U17044 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20909) );
  OR2_X1 U17045 ( .A1(n15137), .A2(n20909), .ZN(n14990) );
  OAI21_X1 U17046 ( .B1(n15138), .B2(n14991), .A(n14990), .ZN(n22640) );
  NAND2_X1 U17047 ( .A1(n15139), .A2(n16746), .ZN(n22649) );
  NOR2_X1 U17048 ( .A1(n15141), .A2(n13204), .ZN(n22639) );
  OAI22_X1 U17049 ( .A1(n15006), .A2(n22649), .B1(n15005), .B2(n22643), .ZN(
        n14992) );
  AOI21_X1 U17050 ( .B1(n22778), .B2(n22640), .A(n14992), .ZN(n14994) );
  NAND2_X1 U17051 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14993) );
  OAI211_X1 U17052 ( .C1(n22630), .C2(n22782), .A(n14994), .B(n14993), .ZN(
        P1_U3157) );
  INV_X1 U17053 ( .A(DATAI_29_), .ZN(n14996) );
  INV_X1 U17054 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20928) );
  OR2_X1 U17055 ( .A1(n15137), .A2(n20928), .ZN(n14995) );
  OAI21_X1 U17056 ( .B1(n15138), .B2(n14996), .A(n14995), .ZN(n22668) );
  INV_X1 U17057 ( .A(n22668), .ZN(n22652) );
  INV_X1 U17058 ( .A(DATAI_21_), .ZN(n14998) );
  INV_X1 U17059 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20911) );
  OR2_X1 U17060 ( .A1(n15137), .A2(n20911), .ZN(n14997) );
  OAI21_X1 U17061 ( .B1(n15138), .B2(n14998), .A(n14997), .ZN(n22662) );
  NAND2_X1 U17062 ( .A1(n15139), .A2(n16743), .ZN(n22671) );
  NOR2_X1 U17063 ( .A1(n15141), .A2(n14999), .ZN(n22661) );
  INV_X1 U17064 ( .A(n22661), .ZN(n22665) );
  OAI22_X1 U17065 ( .A1(n15006), .A2(n22671), .B1(n15005), .B2(n22665), .ZN(
        n15000) );
  AOI21_X1 U17066 ( .B1(n22778), .B2(n22662), .A(n15000), .ZN(n15002) );
  NAND2_X1 U17067 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n15001) );
  OAI211_X1 U17068 ( .C1(n22652), .C2(n22782), .A(n15002), .B(n15001), .ZN(
        P1_U3158) );
  INV_X1 U17069 ( .A(DATAI_25_), .ZN(n16722) );
  INV_X1 U17070 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20919) );
  OR2_X1 U17071 ( .A1(n15137), .A2(n20919), .ZN(n15003) );
  INV_X1 U17072 ( .A(n22582), .ZN(n15451) );
  INV_X1 U17073 ( .A(DATAI_17_), .ZN(n16762) );
  INV_X1 U17074 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20903) );
  OR2_X1 U17075 ( .A1(n15137), .A2(n20903), .ZN(n15004) );
  OAI21_X1 U17076 ( .B1(n15138), .B2(n16762), .A(n15004), .ZN(n22576) );
  NOR2_X1 U17077 ( .A1(n15602), .A2(n16764), .ZN(n15622) );
  NOR2_X1 U17078 ( .A1(n15141), .A2(n15026), .ZN(n22575) );
  INV_X1 U17079 ( .A(n22575), .ZN(n22579) );
  OAI22_X1 U17080 ( .A1(n15006), .A2(n22585), .B1(n15005), .B2(n22579), .ZN(
        n15007) );
  AOI21_X1 U17081 ( .B1(n22778), .B2(n22576), .A(n15007), .ZN(n15009) );
  NAND2_X1 U17082 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n15008) );
  OAI211_X1 U17083 ( .C1(n15451), .C2(n22782), .A(n15009), .B(n15008), .ZN(
        P1_U3154) );
  NOR3_X1 U17084 ( .A1(n22396), .A2(n15600), .A3(n18159), .ZN(n15014) );
  AND2_X1 U17085 ( .A1(n15011), .A2(n15010), .ZN(n18160) );
  INV_X1 U17086 ( .A(n18160), .ZN(n15012) );
  NAND2_X1 U17087 ( .A1(n15012), .A2(n16939), .ZN(n15013) );
  OR2_X1 U17088 ( .A1(n15014), .A2(n15013), .ZN(n15015) );
  INV_X1 U17089 ( .A(n15035), .ZN(n15016) );
  NAND2_X1 U17090 ( .A1(n15016), .A2(n16475), .ZN(n22254) );
  NAND2_X1 U17091 ( .A1(n16584), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15021) );
  NOR2_X1 U17092 ( .A1(n15035), .A2(n15017), .ZN(n15018) );
  OR2_X1 U17093 ( .A1(n22360), .A2(n15018), .ZN(n22270) );
  NAND2_X1 U17094 ( .A1(n15019), .A2(n22270), .ZN(n15041) );
  INV_X1 U17095 ( .A(n15020), .ZN(n15039) );
  INV_X1 U17096 ( .A(n15021), .ZN(n15023) );
  INV_X1 U17097 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16678) );
  AND2_X1 U17098 ( .A1(n22129), .A2(n15972), .ZN(n15032) );
  NAND2_X1 U17099 ( .A1(n15024), .A2(n15032), .ZN(n15028) );
  OAI211_X1 U17100 ( .C1(n15026), .C2(n16678), .A(n15028), .B(n15025), .ZN(
        n15027) );
  NOR2_X2 U17101 ( .A1(n15035), .A2(n15027), .ZN(n22376) );
  OR2_X1 U17102 ( .A1(n15028), .A2(n15130), .ZN(n15029) );
  NAND2_X1 U17103 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n16302) );
  OAI211_X1 U17104 ( .C1(P1_REIP_REG_1__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n22333), .B(n16302), .ZN(n15030) );
  OAI21_X1 U17105 ( .B1(n22342), .B2(n15031), .A(n15030), .ZN(n15038) );
  INV_X1 U17106 ( .A(n15032), .ZN(n18154) );
  NAND3_X1 U17107 ( .A1(n15033), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n18154), 
        .ZN(n15034) );
  NAND2_X1 U17108 ( .A1(n16584), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22370) );
  INV_X1 U17109 ( .A(n16584), .ZN(n22279) );
  AOI22_X1 U17110 ( .A1(n22355), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n22279), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n15036) );
  OAI21_X1 U17111 ( .B1(n22377), .B2(n22152), .A(n15036), .ZN(n15037) );
  AOI211_X1 U17112 ( .C1(n15039), .C2(n22357), .A(n15038), .B(n15037), .ZN(
        n15040) );
  OAI211_X1 U17113 ( .C1(n22254), .C2(n17208), .A(n15041), .B(n15040), .ZN(
        P1_U2838) );
  INV_X1 U17114 ( .A(n22482), .ZN(n15042) );
  NAND3_X1 U17115 ( .A1(n15083), .A2(n22494), .A3(n15042), .ZN(n15044) );
  NOR3_X1 U17116 ( .A1(n15681), .A2(n22475), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22523) );
  INV_X1 U17117 ( .A(n22523), .ZN(n15045) );
  INV_X1 U17118 ( .A(n22492), .ZN(n15043) );
  AOI21_X1 U17119 ( .B1(n15044), .B2(n15045), .A(n15043), .ZN(n15126) );
  INV_X1 U17120 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15054) );
  INV_X1 U17121 ( .A(n22698), .ZN(n22713) );
  AND2_X1 U17122 ( .A1(n17229), .A2(n17208), .ZN(n22519) );
  NAND2_X1 U17123 ( .A1(n22519), .A2(n15213), .ZN(n15047) );
  NOR2_X1 U17124 ( .A1(n22524), .A2(n15045), .ZN(n15162) );
  INV_X1 U17125 ( .A(n15162), .ZN(n15046) );
  NAND2_X1 U17126 ( .A1(n15047), .A2(n15046), .ZN(n15048) );
  NAND2_X1 U17127 ( .A1(n15048), .A2(n22494), .ZN(n15050) );
  NAND2_X1 U17128 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22523), .ZN(n15049) );
  NAND2_X1 U17129 ( .A1(n15050), .A2(n15049), .ZN(n15163) );
  INV_X1 U17130 ( .A(n22706), .ZN(n22691) );
  AOI22_X1 U17131 ( .A1(n15163), .A2(n22691), .B1(n22697), .B2(n15162), .ZN(
        n15051) );
  OAI21_X1 U17132 ( .B1(n22551), .B2(n22713), .A(n15051), .ZN(n15052) );
  AOI21_X1 U17133 ( .B1(n22749), .B2(n22709), .A(n15052), .ZN(n15053) );
  OAI21_X1 U17134 ( .B1(n15126), .B2(n15054), .A(n15053), .ZN(P1_U3127) );
  INV_X1 U17135 ( .A(n15434), .ZN(n15099) );
  NOR3_X1 U17136 ( .A1(n15681), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15060) );
  INV_X1 U17137 ( .A(n15060), .ZN(n15517) );
  NOR2_X1 U17138 ( .A1(n22524), .A2(n15517), .ZN(n22742) );
  AOI21_X1 U17139 ( .B1(n22519), .B2(n15099), .A(n22742), .ZN(n15057) );
  INV_X1 U17140 ( .A(n15057), .ZN(n15055) );
  AOI22_X1 U17141 ( .A1(n15055), .A2(n22494), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15060), .ZN(n22514) );
  INV_X1 U17142 ( .A(n22742), .ZN(n15075) );
  OAI22_X1 U17143 ( .A1(n22514), .A2(n22706), .B1(n22705), .B2(n15075), .ZN(
        n15056) );
  AOI21_X1 U17144 ( .B1(n22750), .B2(n22698), .A(n15056), .ZN(n15062) );
  NAND2_X1 U17145 ( .A1(n15427), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15080) );
  OAI211_X1 U17146 ( .C1(n15058), .C2(n15080), .A(n22494), .B(n15057), .ZN(
        n15059) );
  OAI211_X1 U17147 ( .C1(n22494), .C2(n15060), .A(n15059), .B(n22492), .ZN(
        n22744) );
  NAND2_X1 U17148 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n15061) );
  OAI211_X1 U17149 ( .C1(n22680), .C2(n22747), .A(n15062), .B(n15061), .ZN(
        P1_U3111) );
  OAI22_X1 U17150 ( .A1(n22514), .A2(n22649), .B1(n22643), .B2(n15075), .ZN(
        n15063) );
  AOI21_X1 U17151 ( .B1(n22750), .B2(n22640), .A(n15063), .ZN(n15065) );
  NAND2_X1 U17152 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n15064) );
  OAI211_X1 U17153 ( .C1(n22630), .C2(n22747), .A(n15065), .B(n15064), .ZN(
        P1_U3109) );
  OAI22_X1 U17154 ( .A1(n22514), .A2(n22671), .B1(n22665), .B2(n15075), .ZN(
        n15066) );
  AOI21_X1 U17155 ( .B1(n22750), .B2(n22662), .A(n15066), .ZN(n15068) );
  NAND2_X1 U17156 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n15067) );
  OAI211_X1 U17157 ( .C1(n22652), .C2(n22747), .A(n15068), .B(n15067), .ZN(
        P1_U3110) );
  OAI22_X1 U17158 ( .A1(n22514), .A2(n22585), .B1(n22579), .B2(n15075), .ZN(
        n15069) );
  AOI21_X1 U17159 ( .B1(n22750), .B2(n22576), .A(n15069), .ZN(n15071) );
  NAND2_X1 U17160 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15070) );
  OAI211_X1 U17161 ( .C1(n15451), .C2(n22747), .A(n15071), .B(n15070), .ZN(
        P1_U3106) );
  OAI22_X1 U17162 ( .A1(n22514), .A2(n22627), .B1(n22621), .B2(n15075), .ZN(
        n15072) );
  AOI21_X1 U17163 ( .B1(n22750), .B2(n22618), .A(n15072), .ZN(n15074) );
  NAND2_X1 U17164 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15073) );
  OAI211_X1 U17165 ( .C1(n15440), .C2(n22747), .A(n15074), .B(n15073), .ZN(
        P1_U3108) );
  OAI22_X1 U17166 ( .A1(n22514), .A2(n22605), .B1(n22599), .B2(n15075), .ZN(
        n15076) );
  AOI21_X1 U17167 ( .B1(n22750), .B2(n22596), .A(n15076), .ZN(n15078) );
  NAND2_X1 U17168 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n15077) );
  OAI211_X1 U17169 ( .C1(n15444), .C2(n22747), .A(n15078), .B(n15077), .ZN(
        P1_U3107) );
  INV_X1 U17170 ( .A(n17229), .ZN(n15425) );
  OR2_X1 U17171 ( .A1(n14902), .A2(n15079), .ZN(n15377) );
  MUX2_X1 U17172 ( .A(n15217), .B(n13528), .S(n15972), .Z(n15084) );
  OR2_X1 U17173 ( .A1(n15081), .A2(n15080), .ZN(n15100) );
  INV_X1 U17174 ( .A(n15100), .ZN(n15082) );
  NOR3_X1 U17175 ( .A1(n15084), .A2(n15083), .A3(n15082), .ZN(n15085) );
  OAI222_X1 U17176 ( .A1(n18165), .A2(n15681), .B1(n16459), .B2(n15425), .C1(
        n16454), .C2(n15085), .ZN(P1_U3475) );
  INV_X1 U17177 ( .A(n15086), .ZN(n15091) );
  INV_X1 U17178 ( .A(n15087), .ZN(n15089) );
  INV_X1 U17179 ( .A(n14928), .ZN(n15088) );
  NAND2_X1 U17180 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  NAND2_X1 U17181 ( .A1(n15091), .A2(n15090), .ZN(n19305) );
  INV_X1 U17182 ( .A(n15092), .ZN(n15093) );
  OAI211_X1 U17183 ( .C1(n15095), .C2(n15094), .A(n15093), .B(n17419), .ZN(
        n15097) );
  NAND2_X1 U17184 ( .A1(n17432), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15096) );
  OAI211_X1 U17185 ( .C1(n19305), .C2(n17432), .A(n15097), .B(n15096), .ZN(
        P2_U2879) );
  INV_X1 U17186 ( .A(n22640), .ZN(n22644) );
  NOR3_X1 U17187 ( .A1(n18135), .A2(n15681), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15105) );
  INV_X1 U17188 ( .A(n15105), .ZN(n22542) );
  NOR2_X1 U17189 ( .A1(n22524), .A2(n22542), .ZN(n22766) );
  AOI21_X1 U17190 ( .B1(n22538), .B2(n15099), .A(n22766), .ZN(n15104) );
  NAND3_X1 U17191 ( .A1(n15100), .A2(n22494), .A3(n15104), .ZN(n15101) );
  OAI211_X1 U17192 ( .C1(n22494), .C2(n15105), .A(n22492), .B(n15101), .ZN(
        n22769) );
  NAND2_X1 U17193 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15109) );
  INV_X1 U17194 ( .A(n15104), .ZN(n15106) );
  AOI22_X1 U17195 ( .A1(n15106), .A2(n22494), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15105), .ZN(n22556) );
  INV_X1 U17196 ( .A(n22766), .ZN(n15122) );
  OAI22_X1 U17197 ( .A1(n22556), .A2(n22649), .B1(n22643), .B2(n15122), .ZN(
        n15107) );
  AOI21_X1 U17198 ( .B1(n22535), .B2(n22646), .A(n15107), .ZN(n15108) );
  OAI211_X1 U17199 ( .C1(n22644), .C2(n15684), .A(n15109), .B(n15108), .ZN(
        P1_U3141) );
  INV_X1 U17200 ( .A(n22596), .ZN(n22600) );
  NAND2_X1 U17201 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n15112) );
  OAI22_X1 U17202 ( .A1(n22556), .A2(n22605), .B1(n22599), .B2(n15122), .ZN(
        n15110) );
  AOI21_X1 U17203 ( .B1(n22535), .B2(n22602), .A(n15110), .ZN(n15111) );
  OAI211_X1 U17204 ( .C1(n22600), .C2(n15684), .A(n15112), .B(n15111), .ZN(
        P1_U3139) );
  INV_X1 U17205 ( .A(n22662), .ZN(n22666) );
  NAND2_X1 U17206 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n15115) );
  OAI22_X1 U17207 ( .A1(n22556), .A2(n22671), .B1(n22665), .B2(n15122), .ZN(
        n15113) );
  AOI21_X1 U17208 ( .B1(n22535), .B2(n22668), .A(n15113), .ZN(n15114) );
  OAI211_X1 U17209 ( .C1(n22666), .C2(n15684), .A(n15115), .B(n15114), .ZN(
        P1_U3142) );
  INV_X1 U17210 ( .A(n22576), .ZN(n22580) );
  NAND2_X1 U17211 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n15118) );
  OAI22_X1 U17212 ( .A1(n22556), .A2(n22585), .B1(n22579), .B2(n15122), .ZN(
        n15116) );
  AOI21_X1 U17213 ( .B1(n22535), .B2(n22582), .A(n15116), .ZN(n15117) );
  OAI211_X1 U17214 ( .C1(n22580), .C2(n15684), .A(n15118), .B(n15117), .ZN(
        P1_U3138) );
  NAND2_X1 U17215 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n15121) );
  OAI22_X1 U17216 ( .A1(n22556), .A2(n22706), .B1(n22705), .B2(n15122), .ZN(
        n15119) );
  AOI21_X1 U17217 ( .B1(n22535), .B2(n22709), .A(n15119), .ZN(n15120) );
  OAI211_X1 U17218 ( .C1(n15684), .C2(n22713), .A(n15121), .B(n15120), .ZN(
        P1_U3143) );
  INV_X1 U17219 ( .A(n22618), .ZN(n22622) );
  NAND2_X1 U17220 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n15125) );
  OAI22_X1 U17221 ( .A1(n22556), .A2(n22627), .B1(n22621), .B2(n15122), .ZN(
        n15123) );
  AOI21_X1 U17222 ( .B1(n22535), .B2(n22624), .A(n15123), .ZN(n15124) );
  OAI211_X1 U17223 ( .C1(n22622), .C2(n15684), .A(n15125), .B(n15124), .ZN(
        P1_U3140) );
  INV_X1 U17224 ( .A(DATAI_16_), .ZN(n15128) );
  INV_X1 U17225 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20901) );
  OR2_X1 U17226 ( .A1(n15137), .A2(n20901), .ZN(n15127) );
  OAI21_X1 U17227 ( .B1(n15138), .B2(n15128), .A(n15127), .ZN(n22561) );
  INV_X1 U17228 ( .A(n22561), .ZN(n22544) );
  INV_X1 U17229 ( .A(DATAI_24_), .ZN(n15129) );
  INV_X1 U17230 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20917) );
  OAI22_X1 U17231 ( .A1(n15129), .A2(n15138), .B1(n20917), .B2(n15137), .ZN(
        n22552) );
  NAND2_X1 U17232 ( .A1(n22749), .A2(n22552), .ZN(n15132) );
  NAND2_X1 U17233 ( .A1(n15139), .A2(n16772), .ZN(n22555) );
  INV_X1 U17234 ( .A(n22555), .ZN(n22560) );
  NOR2_X1 U17235 ( .A1(n15141), .A2(n15130), .ZN(n22559) );
  AOI22_X1 U17236 ( .A1(n15163), .A2(n22560), .B1(n22559), .B2(n15162), .ZN(
        n15131) );
  OAI211_X1 U17237 ( .C1(n22544), .C2(n22551), .A(n15132), .B(n15131), .ZN(
        n15133) );
  AOI21_X1 U17238 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n15133), .ZN(n15134) );
  INV_X1 U17239 ( .A(n15134), .ZN(P1_U3121) );
  INV_X1 U17240 ( .A(DATAI_23_), .ZN(n15136) );
  INV_X1 U17241 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20915) );
  OR2_X1 U17242 ( .A1(n15137), .A2(n20915), .ZN(n15135) );
  OAI21_X1 U17243 ( .B1(n15138), .B2(n15136), .A(n15135), .ZN(n22777) );
  INV_X1 U17244 ( .A(n22777), .ZN(n22757) );
  INV_X1 U17245 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20932) );
  OAI22_X1 U17246 ( .A1(n15907), .A2(n15138), .B1(n20932), .B2(n15137), .ZN(
        n22760) );
  NAND2_X1 U17247 ( .A1(n22749), .A2(n22760), .ZN(n15143) );
  NAND2_X1 U17248 ( .A1(n15139), .A2(n16731), .ZN(n22764) );
  INV_X1 U17249 ( .A(n22764), .ZN(n22775) );
  AOI22_X1 U17250 ( .A1(n15163), .A2(n22775), .B1(n22773), .B2(n15162), .ZN(
        n15142) );
  OAI211_X1 U17251 ( .C1(n22757), .C2(n22551), .A(n15143), .B(n15142), .ZN(
        n15144) );
  AOI21_X1 U17252 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n15144), .ZN(n15145) );
  INV_X1 U17253 ( .A(n15145), .ZN(P1_U3128) );
  NAND2_X1 U17254 ( .A1(n22749), .A2(n22646), .ZN(n15147) );
  INV_X1 U17255 ( .A(n22649), .ZN(n15608) );
  AOI22_X1 U17256 ( .A1(n15163), .A2(n15608), .B1(n22639), .B2(n15162), .ZN(
        n15146) );
  OAI211_X1 U17257 ( .C1(n22644), .C2(n22551), .A(n15147), .B(n15146), .ZN(
        n15148) );
  AOI21_X1 U17258 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15148), .ZN(n15149) );
  INV_X1 U17259 ( .A(n15149), .ZN(P1_U3125) );
  NAND2_X1 U17260 ( .A1(n22749), .A2(n22624), .ZN(n15151) );
  AOI22_X1 U17261 ( .A1(n15163), .A2(n17244), .B1(n22617), .B2(n15162), .ZN(
        n15150) );
  OAI211_X1 U17262 ( .C1(n22622), .C2(n22551), .A(n15151), .B(n15150), .ZN(
        n15152) );
  AOI21_X1 U17263 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n15152), .ZN(n15153) );
  INV_X1 U17264 ( .A(n15153), .ZN(P1_U3124) );
  NAND2_X1 U17265 ( .A1(n22749), .A2(n22668), .ZN(n15155) );
  INV_X1 U17266 ( .A(n22671), .ZN(n15613) );
  AOI22_X1 U17267 ( .A1(n15163), .A2(n15613), .B1(n22661), .B2(n15162), .ZN(
        n15154) );
  OAI211_X1 U17268 ( .C1(n22666), .C2(n22551), .A(n15155), .B(n15154), .ZN(
        n15156) );
  AOI21_X1 U17269 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15156), .ZN(n15157) );
  INV_X1 U17270 ( .A(n15157), .ZN(P1_U3126) );
  NAND2_X1 U17271 ( .A1(n22749), .A2(n22602), .ZN(n15159) );
  AOI22_X1 U17272 ( .A1(n15163), .A2(n17236), .B1(n22595), .B2(n15162), .ZN(
        n15158) );
  OAI211_X1 U17273 ( .C1(n22600), .C2(n22551), .A(n15159), .B(n15158), .ZN(
        n15160) );
  AOI21_X1 U17274 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15160), .ZN(n15161) );
  INV_X1 U17275 ( .A(n15161), .ZN(P1_U3123) );
  NAND2_X1 U17276 ( .A1(n22749), .A2(n22582), .ZN(n15165) );
  AOI22_X1 U17277 ( .A1(n15163), .A2(n15622), .B1(n22575), .B2(n15162), .ZN(
        n15164) );
  OAI211_X1 U17278 ( .C1(n22580), .C2(n22551), .A(n15165), .B(n15164), .ZN(
        n15166) );
  AOI21_X1 U17279 ( .B1(n15167), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n15166), .ZN(n15168) );
  INV_X1 U17280 ( .A(n15168), .ZN(P1_U3122) );
  OAI21_X1 U17281 ( .B1(n15171), .B2(n15170), .A(n11174), .ZN(n22173) );
  XOR2_X1 U17282 ( .A(n15173), .B(n15172), .Z(n15415) );
  INV_X1 U17283 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20726) );
  NOR2_X1 U17284 ( .A1(n16939), .A2(n20726), .ZN(n22175) );
  AOI21_X1 U17285 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n22175), .ZN(n15174) );
  OAI21_X1 U17286 ( .B1(n20856), .B2(n15419), .A(n15174), .ZN(n15175) );
  AOI21_X1 U17287 ( .B1(n15415), .B2(n20860), .A(n15175), .ZN(n15176) );
  OAI21_X1 U17288 ( .B1(n22173), .B2(n22386), .A(n15176), .ZN(P1_U2996) );
  INV_X1 U17289 ( .A(n15415), .ZN(n15375) );
  OAI222_X1 U17290 ( .A1(n15375), .A2(n16782), .B1(n16794), .B2(n15177), .C1(
        n16791), .C2(n13534), .ZN(P1_U2901) );
  NAND2_X1 U17291 ( .A1(n11185), .A2(n15178), .ZN(n15179) );
  XNOR2_X1 U17292 ( .A(n16335), .B(n15179), .ZN(n15189) );
  AOI21_X1 U17293 ( .B1(n15182), .B2(n15181), .A(n15180), .ZN(n20254) );
  NAND2_X1 U17294 ( .A1(n20254), .A2(n19459), .ZN(n15187) );
  INV_X1 U17295 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U17296 ( .A1(n15183), .A2(n19473), .B1(P2_EBX_REG_5__SCAN_IN), .B2(
        n19470), .ZN(n15184) );
  OAI211_X1 U17297 ( .C1(n18281), .C2(n19371), .A(n15184), .B(n14452), .ZN(
        n15185) );
  AOI21_X1 U17298 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19472), .A(
        n15185), .ZN(n15186) );
  OAI211_X1 U17299 ( .C1(n19477), .C2(n16331), .A(n15187), .B(n15186), .ZN(
        n15188) );
  AOI21_X1 U17300 ( .B1(n15189), .B2(n19481), .A(n15188), .ZN(n15190) );
  INV_X1 U17301 ( .A(n15190), .ZN(P2_U2850) );
  OAI211_X1 U17302 ( .C1(n15092), .C2(n12698), .A(n17419), .B(n15192), .ZN(
        n15196) );
  OAI21_X1 U17303 ( .B1(n15086), .B2(n15194), .A(n15193), .ZN(n18006) );
  INV_X1 U17304 ( .A(n18006), .ZN(n15270) );
  NAND2_X1 U17305 ( .A1(n15270), .A2(n17411), .ZN(n15195) );
  OAI211_X1 U17306 ( .C1(n17411), .C2(n12220), .A(n15196), .B(n15195), .ZN(
        P2_U2878) );
  AOI21_X1 U17307 ( .B1(n15199), .B2(n15198), .A(n15197), .ZN(n20035) );
  INV_X1 U17308 ( .A(n20035), .ZN(n15210) );
  NAND2_X1 U17309 ( .A1(n11185), .A2(n15200), .ZN(n15201) );
  XNOR2_X1 U17310 ( .A(n17744), .B(n15201), .ZN(n15202) );
  NAND2_X1 U17311 ( .A1(n15202), .A2(n19481), .ZN(n15209) );
  AOI21_X1 U17312 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19472), .A(
        n12603), .ZN(n15203) );
  OAI21_X1 U17313 ( .B1(n19409), .B2(n12211), .A(n15203), .ZN(n15204) );
  AOI21_X1 U17314 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n19471), .A(n15204), .ZN(
        n15205) );
  OAI21_X1 U17315 ( .B1(n18043), .B2(n19477), .A(n15205), .ZN(n15206) );
  AOI21_X1 U17316 ( .B1(n19473), .B2(n15207), .A(n15206), .ZN(n15208) );
  OAI211_X1 U17317 ( .C1(n19475), .C2(n15210), .A(n15209), .B(n15208), .ZN(
        P2_U2848) );
  NOR2_X1 U17318 ( .A1(n22505), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15220) );
  INV_X1 U17319 ( .A(n15217), .ZN(n15215) );
  OR2_X1 U17320 ( .A1(n17208), .A2(n15211), .ZN(n22502) );
  INV_X1 U17321 ( .A(n22502), .ZN(n15214) );
  NOR2_X1 U17322 ( .A1(n15212), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17258) );
  AOI21_X1 U17323 ( .B1(n15214), .B2(n15213), .A(n17258), .ZN(n15218) );
  OAI211_X1 U17324 ( .C1(n15215), .C2(n15972), .A(n22494), .B(n15218), .ZN(
        n15216) );
  OAI211_X1 U17325 ( .C1(n22494), .C2(n15220), .A(n15216), .B(n22492), .ZN(
        n17257) );
  NAND2_X1 U17326 ( .A1(n22618), .A2(n22693), .ZN(n15224) );
  INV_X1 U17327 ( .A(n15218), .ZN(n15219) );
  NAND2_X1 U17328 ( .A1(n15219), .A2(n22494), .ZN(n15222) );
  NAND2_X1 U17329 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15220), .ZN(n15221) );
  NAND2_X1 U17330 ( .A1(n15222), .A2(n15221), .ZN(n17259) );
  AOI22_X1 U17331 ( .A1(n17244), .A2(n17259), .B1(n22617), .B2(n17258), .ZN(
        n15223) );
  OAI211_X1 U17332 ( .C1(n15440), .C2(n22735), .A(n15224), .B(n15223), .ZN(
        n15225) );
  AOI21_X1 U17333 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15225), .ZN(n15226) );
  INV_X1 U17334 ( .A(n15226), .ZN(P1_U3092) );
  NAND2_X1 U17335 ( .A1(n22693), .A2(n22662), .ZN(n15228) );
  AOI22_X1 U17336 ( .A1(n17259), .A2(n15613), .B1(n22661), .B2(n17258), .ZN(
        n15227) );
  OAI211_X1 U17337 ( .C1(n22652), .C2(n22735), .A(n15228), .B(n15227), .ZN(
        n15229) );
  AOI21_X1 U17338 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15229), .ZN(n15230) );
  INV_X1 U17339 ( .A(n15230), .ZN(P1_U3094) );
  INV_X1 U17340 ( .A(n22552), .ZN(n22564) );
  NAND2_X1 U17341 ( .A1(n22693), .A2(n22561), .ZN(n15232) );
  AOI22_X1 U17342 ( .A1(n17259), .A2(n22560), .B1(n22559), .B2(n17258), .ZN(
        n15231) );
  OAI211_X1 U17343 ( .C1(n22735), .C2(n22564), .A(n15232), .B(n15231), .ZN(
        n15233) );
  AOI21_X1 U17344 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n15233), .ZN(n15234) );
  INV_X1 U17345 ( .A(n15234), .ZN(P1_U3089) );
  NAND2_X1 U17346 ( .A1(n22596), .A2(n22693), .ZN(n15236) );
  AOI22_X1 U17347 ( .A1(n17236), .A2(n17259), .B1(n22595), .B2(n17258), .ZN(
        n15235) );
  OAI211_X1 U17348 ( .C1(n15444), .C2(n22735), .A(n15236), .B(n15235), .ZN(
        n15237) );
  AOI21_X1 U17349 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n15237), .ZN(n15238) );
  INV_X1 U17350 ( .A(n15238), .ZN(P1_U3091) );
  NAND2_X1 U17351 ( .A1(n22693), .A2(n22576), .ZN(n15240) );
  AOI22_X1 U17352 ( .A1(n15622), .A2(n17259), .B1(n22575), .B2(n17258), .ZN(
        n15239) );
  OAI211_X1 U17353 ( .C1(n15451), .C2(n22735), .A(n15240), .B(n15239), .ZN(
        n15241) );
  AOI21_X1 U17354 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n15241), .ZN(n15242) );
  INV_X1 U17355 ( .A(n15242), .ZN(P1_U3090) );
  INV_X1 U17356 ( .A(n22760), .ZN(n22783) );
  NAND2_X1 U17357 ( .A1(n22693), .A2(n22777), .ZN(n15244) );
  AOI22_X1 U17358 ( .A1(n17259), .A2(n22775), .B1(n22773), .B2(n17258), .ZN(
        n15243) );
  OAI211_X1 U17359 ( .C1(n22735), .C2(n22783), .A(n15244), .B(n15243), .ZN(
        n15245) );
  AOI21_X1 U17360 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n15245), .ZN(n15246) );
  INV_X1 U17361 ( .A(n15246), .ZN(P1_U3096) );
  NAND2_X1 U17362 ( .A1(n22693), .A2(n22640), .ZN(n15248) );
  AOI22_X1 U17363 ( .A1(n17259), .A2(n15608), .B1(n22639), .B2(n17258), .ZN(
        n15247) );
  OAI211_X1 U17364 ( .C1(n22630), .C2(n22735), .A(n15248), .B(n15247), .ZN(
        n15249) );
  AOI21_X1 U17365 ( .B1(n17257), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n15249), .ZN(n15250) );
  INV_X1 U17366 ( .A(n15250), .ZN(P1_U3093) );
  INV_X1 U17367 ( .A(n16746), .ZN(n15255) );
  NAND2_X1 U17368 ( .A1(n15252), .A2(n15253), .ZN(n15254) );
  AND2_X1 U17369 ( .A1(n15251), .A2(n15254), .ZN(n22257) );
  INV_X1 U17370 ( .A(n22257), .ZN(n15260) );
  OAI222_X1 U17371 ( .A1(n16794), .A2(n15255), .B1(n16791), .B2(n20704), .C1(
        n16782), .C2(n15260), .ZN(P1_U2900) );
  OR2_X1 U17372 ( .A1(n15258), .A2(n15257), .ZN(n15259) );
  NAND2_X1 U17373 ( .A1(n15256), .A2(n15259), .ZN(n22246) );
  OAI222_X1 U17374 ( .A1(n22246), .A2(n20820), .B1(n16074), .B2(n20830), .C1(
        n20805), .C2(n15260), .ZN(P1_U2868) );
  INV_X1 U17375 ( .A(n15261), .ZN(n15273) );
  NAND2_X1 U17376 ( .A1(n11185), .A2(n15262), .ZN(n15263) );
  XOR2_X1 U17377 ( .A(n17729), .B(n15263), .Z(n15264) );
  NAND2_X1 U17378 ( .A1(n15264), .A2(n19481), .ZN(n15272) );
  AOI21_X1 U17379 ( .B1(n15266), .B2(n18032), .A(n17989), .ZN(n20029) );
  AOI22_X1 U17380 ( .A1(n19471), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n19459), 
        .B2(n20029), .ZN(n15268) );
  AOI21_X1 U17381 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19472), .A(
        n12603), .ZN(n15267) );
  OAI211_X1 U17382 ( .C1(n12220), .C2(n19409), .A(n15268), .B(n15267), .ZN(
        n15269) );
  AOI21_X1 U17383 ( .B1(n15270), .B2(n19461), .A(n15269), .ZN(n15271) );
  OAI211_X1 U17384 ( .C1(n15273), .C2(n19441), .A(n15272), .B(n15271), .ZN(
        P2_U2846) );
  INV_X1 U17385 ( .A(n15303), .ZN(n15309) );
  INV_X1 U17386 ( .A(n12130), .ZN(n15275) );
  NAND2_X1 U17387 ( .A1(n11168), .A2(n15275), .ZN(n15281) );
  NAND2_X1 U17388 ( .A1(n11773), .A2(n15276), .ZN(n15315) );
  INV_X1 U17389 ( .A(n11542), .ZN(n15278) );
  NAND2_X1 U17390 ( .A1(n15278), .A2(n15277), .ZN(n15310) );
  INV_X1 U17391 ( .A(n15310), .ZN(n15279) );
  AOI21_X1 U17392 ( .B1(n15315), .B2(n15311), .A(n15279), .ZN(n15280) );
  AND2_X1 U17393 ( .A1(n15281), .A2(n15280), .ZN(n15284) );
  OR2_X1 U17394 ( .A1(n15341), .A2(n15282), .ZN(n15320) );
  AOI22_X1 U17395 ( .A1(n15320), .A2(n15310), .B1(n12130), .B2(n11168), .ZN(
        n15283) );
  MUX2_X1 U17396 ( .A(n15284), .B(n15283), .S(n11713), .Z(n15286) );
  NAND2_X1 U17397 ( .A1(n15286), .A2(n15285), .ZN(n15287) );
  AOI21_X1 U17398 ( .B1(n11196), .B2(n15309), .A(n15287), .ZN(n18079) );
  NAND2_X1 U17399 ( .A1(n15331), .A2(n15333), .ZN(n15288) );
  AND4_X1 U17400 ( .A1(n15291), .A2(n15290), .A3(n15289), .A4(n15288), .ZN(
        n15294) );
  NAND2_X1 U17401 ( .A1(n15292), .A2(n15332), .ZN(n15293) );
  NAND2_X1 U17402 ( .A1(n15294), .A2(n15293), .ZN(n15474) );
  MUX2_X1 U17403 ( .A(n11713), .B(n18079), .S(n15474), .Z(n15330) );
  INV_X1 U17404 ( .A(n12371), .ZN(n15300) );
  NAND2_X1 U17405 ( .A1(n17360), .A2(n15309), .ZN(n15299) );
  INV_X1 U17406 ( .A(n12565), .ZN(n15295) );
  AND2_X1 U17407 ( .A1(n15296), .A2(n15295), .ZN(n15301) );
  INV_X1 U17408 ( .A(n15301), .ZN(n15297) );
  OAI21_X1 U17409 ( .B1(n11543), .B2(n11541), .A(n15297), .ZN(n15298) );
  OAI211_X1 U17410 ( .C1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15300), .A(
        n15299), .B(n15298), .ZN(n18074) );
  MUX2_X1 U17411 ( .A(n15301), .B(n15300), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15302) );
  OAI21_X1 U17412 ( .B1(n15304), .B2(n15303), .A(n15302), .ZN(n15473) );
  OR2_X1 U17413 ( .A1(n20122), .A2(n15473), .ZN(n15305) );
  OAI21_X1 U17414 ( .B1(n18074), .B2(n15305), .A(n20150), .ZN(n15308) );
  NAND2_X1 U17415 ( .A1(n18074), .A2(n15305), .ZN(n15307) );
  INV_X1 U17416 ( .A(n15474), .ZN(n15306) );
  AOI21_X1 U17417 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15323) );
  NAND2_X1 U17418 ( .A1(n12677), .A2(n15309), .ZN(n15322) );
  AND2_X1 U17419 ( .A1(n15311), .A2(n15310), .ZN(n15314) );
  INV_X1 U17420 ( .A(n15314), .ZN(n15319) );
  NOR2_X1 U17421 ( .A1(n15312), .A2(n12130), .ZN(n15313) );
  NAND2_X1 U17422 ( .A1(n12371), .A2(n15313), .ZN(n15317) );
  NAND2_X1 U17423 ( .A1(n15315), .A2(n15314), .ZN(n15316) );
  NAND2_X1 U17424 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  AOI21_X1 U17425 ( .B1(n15320), .B2(n15319), .A(n15318), .ZN(n15321) );
  NAND2_X1 U17426 ( .A1(n15322), .A2(n15321), .ZN(n15649) );
  MUX2_X1 U17427 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15649), .S(
        n15474), .Z(n15328) );
  AOI222_X1 U17428 ( .A1(n15323), .A2(n20146), .B1(n15323), .B2(n15649), .C1(
        n20146), .C2(n15328), .ZN(n15327) );
  OR2_X1 U17429 ( .A1(n15327), .A2(n15330), .ZN(n15324) );
  NAND2_X1 U17430 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15324), .ZN(
        n15325) );
  NAND2_X1 U17431 ( .A1(n18108), .A2(n15325), .ZN(n15326) );
  AOI21_X1 U17432 ( .B1(n15330), .B2(n15327), .A(n15326), .ZN(n15357) );
  INV_X1 U17433 ( .A(n15328), .ZN(n15329) );
  NOR2_X1 U17434 ( .A1(n15330), .A2(n15329), .ZN(n15356) );
  INV_X1 U17435 ( .A(n15331), .ZN(n15334) );
  NOR3_X1 U17436 ( .A1(n15334), .A2(n15333), .A3(n15332), .ZN(n19537) );
  OAI21_X1 U17437 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19537), .ZN(n15354) );
  INV_X1 U17438 ( .A(n15335), .ZN(n15338) );
  NAND2_X1 U17439 ( .A1(n11761), .A2(n15336), .ZN(n15337) );
  OAI21_X1 U17440 ( .B1(n15339), .B2(n15338), .A(n15337), .ZN(n15340) );
  AOI21_X1 U17441 ( .B1(n15346), .B2(n15341), .A(n15340), .ZN(n15344) );
  NAND2_X1 U17442 ( .A1(n19523), .A2(n15342), .ZN(n15343) );
  OAI211_X1 U17443 ( .C1(n15346), .C2(n15345), .A(n15344), .B(n15343), .ZN(
        n19538) );
  INV_X1 U17444 ( .A(n19488), .ZN(n15347) );
  NAND2_X1 U17445 ( .A1(n19490), .A2(n15347), .ZN(n15348) );
  NOR2_X1 U17446 ( .A1(n11181), .A2(n15348), .ZN(n15350) );
  NOR3_X1 U17447 ( .A1(n19538), .A2(n15351), .A3(n15350), .ZN(n15353) );
  OR2_X1 U17448 ( .A1(n15474), .A2(n19492), .ZN(n15352) );
  NAND3_X1 U17449 ( .A1(n15354), .A2(n15353), .A3(n15352), .ZN(n15355) );
  NAND2_X1 U17450 ( .A1(n18105), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15359) );
  OAI21_X1 U17451 ( .B1(n19520), .B2(n15359), .A(n15358), .ZN(n15362) );
  NAND2_X1 U17452 ( .A1(n15360), .A2(n11169), .ZN(n15361) );
  OAI21_X1 U17453 ( .B1(n19527), .B2(n19251), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15363) );
  NOR2_X1 U17454 ( .A1(n19251), .A2(n18205), .ZN(n18104) );
  INV_X1 U17455 ( .A(n18104), .ZN(n19522) );
  NAND2_X1 U17456 ( .A1(n15363), .A2(n19522), .ZN(P2_U3593) );
  INV_X1 U17457 ( .A(n22254), .ZN(n15468) );
  INV_X1 U17458 ( .A(n15364), .ZN(n15365) );
  AOI22_X1 U17459 ( .A1(n22359), .A2(n15365), .B1(n22376), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n15368) );
  NAND2_X1 U17460 ( .A1(n22339), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15367) );
  OAI21_X1 U17461 ( .B1(n22357), .B2(n22355), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15366) );
  NAND3_X1 U17462 ( .A1(n15368), .A2(n15367), .A3(n15366), .ZN(n15371) );
  INV_X1 U17463 ( .A(n22270), .ZN(n15470) );
  NOR2_X1 U17464 ( .A1(n15369), .A2(n15470), .ZN(n15370) );
  AOI211_X1 U17465 ( .C1(n15468), .C2(n11176), .A(n15371), .B(n15370), .ZN(
        n15372) );
  INV_X1 U17466 ( .A(n15372), .ZN(P1_U2840) );
  XOR2_X1 U17467 ( .A(n15374), .B(n15373), .Z(n22176) );
  INV_X1 U17468 ( .A(n22176), .ZN(n15376) );
  INV_X1 U17469 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n15418) );
  OAI222_X1 U17470 ( .A1(n15376), .A2(n20820), .B1(n20830), .B2(n15418), .C1(
        n20805), .C2(n15375), .ZN(P1_U2869) );
  NOR3_X1 U17471 ( .A1(n18135), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15383) );
  INV_X1 U17472 ( .A(n15386), .ZN(n15380) );
  INV_X1 U17473 ( .A(n15383), .ZN(n15599) );
  NOR2_X1 U17474 ( .A1(n22524), .A2(n15599), .ZN(n17250) );
  INV_X1 U17475 ( .A(n17250), .ZN(n15378) );
  OAI21_X1 U17476 ( .B1(n22502), .B2(n15434), .A(n15378), .ZN(n15382) );
  INV_X1 U17477 ( .A(n15382), .ZN(n15379) );
  OAI211_X1 U17478 ( .C1(n15380), .C2(n15972), .A(n22494), .B(n15379), .ZN(
        n15381) );
  OAI211_X1 U17479 ( .C1(n22494), .C2(n15383), .A(n15381), .B(n22492), .ZN(
        n17249) );
  NAND2_X1 U17480 ( .A1(n15382), .A2(n22494), .ZN(n15385) );
  NAND2_X1 U17481 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15383), .ZN(n15384) );
  NAND2_X1 U17482 ( .A1(n15385), .A2(n15384), .ZN(n17251) );
  AOI22_X1 U17483 ( .A1(n17236), .A2(n17251), .B1(n22595), .B2(n17250), .ZN(
        n15388) );
  NAND2_X1 U17484 ( .A1(n22737), .A2(n22596), .ZN(n15387) );
  OAI211_X1 U17485 ( .C1(n15632), .C2(n15444), .A(n15388), .B(n15387), .ZN(
        n15389) );
  AOI21_X1 U17486 ( .B1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n17249), .A(
        n15389), .ZN(n15390) );
  INV_X1 U17487 ( .A(n15390), .ZN(P1_U3075) );
  AOI22_X1 U17488 ( .A1(n15622), .A2(n17251), .B1(n22575), .B2(n17250), .ZN(
        n15392) );
  NAND2_X1 U17489 ( .A1(n22737), .A2(n22576), .ZN(n15391) );
  OAI211_X1 U17490 ( .C1(n15632), .C2(n15451), .A(n15392), .B(n15391), .ZN(
        n15393) );
  AOI21_X1 U17491 ( .B1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17249), .A(
        n15393), .ZN(n15394) );
  INV_X1 U17492 ( .A(n15394), .ZN(P1_U3074) );
  AOI22_X1 U17493 ( .A1(n17251), .A2(n22560), .B1(n22559), .B2(n17250), .ZN(
        n15396) );
  NAND2_X1 U17494 ( .A1(n22737), .A2(n22561), .ZN(n15395) );
  OAI211_X1 U17495 ( .C1(n15632), .C2(n22564), .A(n15396), .B(n15395), .ZN(
        n15397) );
  AOI21_X1 U17496 ( .B1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B2(n17249), .A(
        n15397), .ZN(n15398) );
  INV_X1 U17497 ( .A(n15398), .ZN(P1_U3073) );
  AOI22_X1 U17498 ( .A1(n17251), .A2(n15608), .B1(n22639), .B2(n17250), .ZN(
        n15400) );
  NAND2_X1 U17499 ( .A1(n22737), .A2(n22640), .ZN(n15399) );
  OAI211_X1 U17500 ( .C1(n15632), .C2(n22630), .A(n15400), .B(n15399), .ZN(
        n15401) );
  AOI21_X1 U17501 ( .B1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n17249), .A(
        n15401), .ZN(n15402) );
  INV_X1 U17502 ( .A(n15402), .ZN(P1_U3077) );
  AOI22_X1 U17503 ( .A1(n17244), .A2(n17251), .B1(n22617), .B2(n17250), .ZN(
        n15404) );
  NAND2_X1 U17504 ( .A1(n22737), .A2(n22618), .ZN(n15403) );
  OAI211_X1 U17505 ( .C1(n15632), .C2(n15440), .A(n15404), .B(n15403), .ZN(
        n15405) );
  AOI21_X1 U17506 ( .B1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n17249), .A(
        n15405), .ZN(n15406) );
  INV_X1 U17507 ( .A(n15406), .ZN(P1_U3076) );
  AOI22_X1 U17508 ( .A1(n17251), .A2(n22775), .B1(n22773), .B2(n17250), .ZN(
        n15408) );
  NAND2_X1 U17509 ( .A1(n22737), .A2(n22777), .ZN(n15407) );
  OAI211_X1 U17510 ( .C1(n15632), .C2(n22783), .A(n15408), .B(n15407), .ZN(
        n15409) );
  AOI21_X1 U17511 ( .B1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17249), .A(
        n15409), .ZN(n15410) );
  INV_X1 U17512 ( .A(n15410), .ZN(P1_U3080) );
  AOI22_X1 U17513 ( .A1(n17251), .A2(n15613), .B1(n22661), .B2(n17250), .ZN(
        n15412) );
  NAND2_X1 U17514 ( .A1(n22737), .A2(n22662), .ZN(n15411) );
  OAI211_X1 U17515 ( .C1(n15632), .C2(n22652), .A(n15412), .B(n15411), .ZN(
        n15413) );
  AOI21_X1 U17516 ( .B1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B2(n17249), .A(
        n15413), .ZN(n15414) );
  INV_X1 U17517 ( .A(n15414), .ZN(P1_U3078) );
  NAND2_X1 U17518 ( .A1(n15415), .A2(n22270), .ZN(n15424) );
  XOR2_X1 U17519 ( .A(n20726), .B(n16302), .Z(n15422) );
  AOI22_X1 U17520 ( .A1(n22355), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n22279), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n15417) );
  NAND2_X1 U17521 ( .A1(n22359), .A2(n22176), .ZN(n15416) );
  OAI211_X1 U17522 ( .C1(n22342), .C2(n15418), .A(n15417), .B(n15416), .ZN(
        n15421) );
  NOR2_X1 U17523 ( .A1(n22384), .A2(n15419), .ZN(n15420) );
  AOI211_X1 U17524 ( .C1(n15422), .C2(n22333), .A(n15421), .B(n15420), .ZN(
        n15423) );
  OAI211_X1 U17525 ( .C1(n15425), .C2(n22254), .A(n15424), .B(n15423), .ZN(
        P1_U2837) );
  INV_X1 U17526 ( .A(n14902), .ZN(n15426) );
  NOR3_X1 U17527 ( .A1(n15429), .A2(n22534), .A3(n15972), .ZN(n15430) );
  NOR3_X1 U17528 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15435) );
  NAND2_X1 U17529 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15439) );
  INV_X1 U17530 ( .A(n17208), .ZN(n15433) );
  OR2_X1 U17531 ( .A1(n17229), .A2(n15433), .ZN(n22485) );
  INV_X1 U17532 ( .A(n15435), .ZN(n22462) );
  NOR2_X1 U17533 ( .A1(n22524), .A2(n22462), .ZN(n22675) );
  INV_X1 U17534 ( .A(n22675), .ZN(n15458) );
  OAI21_X1 U17535 ( .B1(n22485), .B2(n15434), .A(n15458), .ZN(n15436) );
  AOI22_X1 U17536 ( .A1(n15436), .A2(n22494), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15435), .ZN(n22674) );
  OAI22_X1 U17537 ( .A1(n22674), .A2(n22627), .B1(n22621), .B2(n15458), .ZN(
        n15437) );
  AOI21_X1 U17538 ( .B1(n22722), .B2(n22618), .A(n15437), .ZN(n15438) );
  OAI211_X1 U17539 ( .C1(n15440), .C2(n15462), .A(n15439), .B(n15438), .ZN(
        P1_U3044) );
  NAND2_X1 U17540 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15443) );
  OAI22_X1 U17541 ( .A1(n22674), .A2(n22605), .B1(n22599), .B2(n15458), .ZN(
        n15441) );
  AOI21_X1 U17542 ( .B1(n22722), .B2(n22596), .A(n15441), .ZN(n15442) );
  OAI211_X1 U17543 ( .C1(n15444), .C2(n15462), .A(n15443), .B(n15442), .ZN(
        P1_U3043) );
  NAND2_X1 U17544 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15447) );
  OAI22_X1 U17545 ( .A1(n22674), .A2(n22671), .B1(n22665), .B2(n15458), .ZN(
        n15445) );
  AOI21_X1 U17546 ( .B1(n22722), .B2(n22662), .A(n15445), .ZN(n15446) );
  OAI211_X1 U17547 ( .C1(n22652), .C2(n15462), .A(n15447), .B(n15446), .ZN(
        P1_U3046) );
  NAND2_X1 U17548 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15450) );
  OAI22_X1 U17549 ( .A1(n22674), .A2(n22585), .B1(n22579), .B2(n15458), .ZN(
        n15448) );
  AOI21_X1 U17550 ( .B1(n22722), .B2(n22576), .A(n15448), .ZN(n15449) );
  OAI211_X1 U17551 ( .C1(n15451), .C2(n15462), .A(n15450), .B(n15449), .ZN(
        P1_U3042) );
  NAND2_X1 U17552 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15454) );
  OAI22_X1 U17553 ( .A1(n22674), .A2(n22649), .B1(n22643), .B2(n15458), .ZN(
        n15452) );
  AOI21_X1 U17554 ( .B1(n22722), .B2(n22640), .A(n15452), .ZN(n15453) );
  OAI211_X1 U17555 ( .C1(n22630), .C2(n15462), .A(n15454), .B(n15453), .ZN(
        P1_U3045) );
  NAND2_X1 U17556 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n15457) );
  INV_X1 U17557 ( .A(n22773), .ZN(n22755) );
  OAI22_X1 U17558 ( .A1(n22674), .A2(n22764), .B1(n22755), .B2(n15458), .ZN(
        n15455) );
  AOI21_X1 U17559 ( .B1(n22722), .B2(n22777), .A(n15455), .ZN(n15456) );
  OAI211_X1 U17560 ( .C1(n22783), .C2(n15462), .A(n15457), .B(n15456), .ZN(
        P1_U3048) );
  NAND2_X1 U17561 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15461) );
  INV_X1 U17562 ( .A(n22559), .ZN(n22543) );
  OAI22_X1 U17563 ( .A1(n22674), .A2(n22555), .B1(n22543), .B2(n15458), .ZN(
        n15459) );
  AOI21_X1 U17564 ( .B1(n22722), .B2(n22561), .A(n15459), .ZN(n15460) );
  OAI211_X1 U17565 ( .C1(n22564), .C2(n15462), .A(n15461), .B(n15460), .ZN(
        P1_U3041) );
  INV_X1 U17566 ( .A(n11222), .ZN(n22518) );
  AOI22_X1 U17567 ( .A1(n22355), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n22279), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n15465) );
  NAND2_X1 U17568 ( .A1(n22359), .A2(n15463), .ZN(n15464) );
  OAI211_X1 U17569 ( .C1(n22384), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15465), .B(n15464), .ZN(n15467) );
  OAI22_X1 U17570 ( .A1(n22373), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n22342), 
        .B2(n14248), .ZN(n15466) );
  AOI211_X1 U17571 ( .C1(n22518), .C2(n15468), .A(n15467), .B(n15466), .ZN(
        n15469) );
  OAI21_X1 U17572 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(P1_U2839) );
  NOR2_X1 U17573 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U17574 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19259), .B2(n11185), .ZN(n15647) );
  AOI222_X1 U17575 ( .A1(n15473), .A2(n18078), .B1(n19529), .B2(n19269), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15647), .ZN(n15479) );
  NAND2_X1 U17576 ( .A1(n15474), .A2(n19511), .ZN(n15477) );
  INV_X1 U17577 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19540) );
  NOR2_X1 U17578 ( .A1(n19522), .A2(n19540), .ZN(n15475) );
  AOI21_X1 U17579 ( .B1(n19251), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n15475), 
        .ZN(n15476) );
  NAND2_X1 U17580 ( .A1(n15477), .A2(n15476), .ZN(n19493) );
  INV_X1 U17581 ( .A(n19493), .ZN(n18076) );
  NAND2_X1 U17582 ( .A1(n18076), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15478) );
  OAI21_X1 U17583 ( .B1(n15479), .B2(n18076), .A(n15478), .ZN(P2_U3601) );
  INV_X1 U17584 ( .A(n15481), .ZN(n16438) );
  NOR2_X1 U17585 ( .A1(n11184), .A2(n15645), .ZN(n15482) );
  INV_X1 U17586 ( .A(n15482), .ZN(n15480) );
  AOI221_X1 U17587 ( .B1(n16438), .B2(n15482), .C1(n15481), .C2(n15480), .A(
        n19518), .ZN(n15483) );
  INV_X1 U17588 ( .A(n15483), .ZN(n15494) );
  OR2_X1 U17589 ( .A1(n15485), .A2(n15484), .ZN(n15487) );
  NAND2_X1 U17590 ( .A1(n15487), .A2(n15486), .ZN(n20408) );
  AOI22_X1 U17591 ( .A1(n19470), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19472), .ZN(n15489) );
  NAND2_X1 U17592 ( .A1(n19471), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n15488) );
  OAI211_X1 U17593 ( .C1(n19441), .C2(n15490), .A(n15489), .B(n15488), .ZN(
        n15492) );
  NOR2_X1 U17594 ( .A1(n16440), .A2(n19477), .ZN(n15491) );
  AOI211_X1 U17595 ( .C1(n19459), .C2(n20408), .A(n15492), .B(n15491), .ZN(
        n15493) );
  OAI211_X1 U17596 ( .C1(n19276), .C2(n20409), .A(n15494), .B(n15493), .ZN(
        P2_U2853) );
  OR2_X1 U17597 ( .A1(n20255), .A2(n22411), .ZN(n20178) );
  NAND3_X1 U17598 ( .A1(n20150), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20051) );
  OAI21_X1 U17599 ( .B1(n15710), .B2(n20178), .A(n20051), .ZN(n15505) );
  NOR2_X1 U17600 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18105), .ZN(n19247) );
  NOR2_X1 U17601 ( .A1(n15498), .A2(n19247), .ZN(n19528) );
  NOR2_X1 U17602 ( .A1(n15499), .A2(n19528), .ZN(n15500) );
  NAND2_X1 U17603 ( .A1(n20165), .A2(n15500), .ZN(n20180) );
  INV_X1 U17604 ( .A(n15500), .ZN(n15501) );
  NOR2_X1 U17605 ( .A1(n20122), .A2(n20051), .ZN(n20544) );
  INV_X1 U17606 ( .A(n20544), .ZN(n20042) );
  AND2_X1 U17607 ( .A1(n20192), .A2(n20042), .ZN(n15503) );
  OAI22_X1 U17608 ( .A1(n15509), .A2(n20180), .B1(n20525), .B2(n15503), .ZN(
        n15504) );
  NAND2_X1 U17609 ( .A1(n15505), .A2(n15504), .ZN(n20546) );
  INV_X1 U17610 ( .A(n20546), .ZN(n20422) );
  INV_X1 U17611 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15516) );
  INV_X1 U17612 ( .A(n20163), .ZN(n15506) );
  AOI22_X1 U17613 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20531), .ZN(n20188) );
  INV_X1 U17614 ( .A(n20532), .ZN(n20212) );
  INV_X1 U17615 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19569) );
  INV_X1 U17616 ( .A(n20531), .ZN(n20211) );
  AOI22_X1 U17617 ( .A1(n20538), .A2(n20191), .B1(n20552), .B2(n20185), .ZN(
        n15515) );
  INV_X1 U17618 ( .A(n15509), .ZN(n15510) );
  OAI21_X1 U17619 ( .B1(n15510), .B2(n20544), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15511) );
  OAI21_X1 U17620 ( .B1(n20051), .B2(n20192), .A(n15511), .ZN(n20545) );
  NOR2_X2 U17621 ( .A1(n15513), .A2(n20527), .ZN(n20190) );
  AOI22_X1 U17622 ( .A1(n20545), .A2(n15512), .B1(n20190), .B2(n20544), .ZN(
        n15514) );
  OAI211_X1 U17623 ( .C1(n20422), .C2(n15516), .A(n15515), .B(n15514), .ZN(
        P2_U3159) );
  NOR2_X1 U17624 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15517), .ZN(
        n22690) );
  INV_X1 U17625 ( .A(n22747), .ZN(n15518) );
  OAI21_X1 U17626 ( .B1(n15518), .B2(n22693), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15519) );
  AOI21_X1 U17627 ( .B1(n22519), .B2(n11222), .A(n22690), .ZN(n15521) );
  NAND2_X1 U17628 ( .A1(n15519), .A2(n15521), .ZN(n15520) );
  NOR2_X1 U17629 ( .A1(n15522), .A2(n22489), .ZN(n22540) );
  NAND2_X1 U17630 ( .A1(n22693), .A2(n22602), .ZN(n15526) );
  OR2_X1 U17631 ( .A1(n15521), .A2(n22534), .ZN(n15524) );
  NAND2_X1 U17632 ( .A1(n15604), .A2(n22473), .ZN(n22546) );
  INV_X1 U17633 ( .A(n22546), .ZN(n22539) );
  AND2_X1 U17634 ( .A1(n15522), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22521) );
  NAND2_X1 U17635 ( .A1(n22539), .A2(n22521), .ZN(n15523) );
  NAND2_X1 U17636 ( .A1(n15524), .A2(n15523), .ZN(n22692) );
  AOI22_X1 U17637 ( .A1(n22692), .A2(n17236), .B1(n22595), .B2(n22690), .ZN(
        n15525) );
  OAI211_X1 U17638 ( .C1(n22747), .C2(n22600), .A(n15526), .B(n15525), .ZN(
        n15527) );
  AOI21_X1 U17639 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n15527), .ZN(n15528) );
  INV_X1 U17640 ( .A(n15528), .ZN(P1_U3099) );
  NAND2_X1 U17641 ( .A1(n22693), .A2(n22760), .ZN(n15530) );
  AOI22_X1 U17642 ( .A1(n22692), .A2(n22775), .B1(n22773), .B2(n22690), .ZN(
        n15529) );
  OAI211_X1 U17643 ( .C1(n22747), .C2(n22757), .A(n15530), .B(n15529), .ZN(
        n15531) );
  AOI21_X1 U17644 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15531), .ZN(n15532) );
  INV_X1 U17645 ( .A(n15532), .ZN(P1_U3104) );
  NAND2_X1 U17646 ( .A1(n22693), .A2(n22552), .ZN(n15534) );
  AOI22_X1 U17647 ( .A1(n22692), .A2(n22560), .B1(n22559), .B2(n22690), .ZN(
        n15533) );
  OAI211_X1 U17648 ( .C1(n22747), .C2(n22544), .A(n15534), .B(n15533), .ZN(
        n15535) );
  AOI21_X1 U17649 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n15535), .ZN(n15536) );
  INV_X1 U17650 ( .A(n15536), .ZN(P1_U3097) );
  NAND2_X1 U17651 ( .A1(n22693), .A2(n22624), .ZN(n15538) );
  AOI22_X1 U17652 ( .A1(n22692), .A2(n17244), .B1(n22617), .B2(n22690), .ZN(
        n15537) );
  OAI211_X1 U17653 ( .C1(n22747), .C2(n22622), .A(n15538), .B(n15537), .ZN(
        n15539) );
  AOI21_X1 U17654 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n15539), .ZN(n15540) );
  INV_X1 U17655 ( .A(n15540), .ZN(P1_U3100) );
  NAND2_X1 U17656 ( .A1(n22693), .A2(n22668), .ZN(n15542) );
  AOI22_X1 U17657 ( .A1(n22692), .A2(n15613), .B1(n22661), .B2(n22690), .ZN(
        n15541) );
  OAI211_X1 U17658 ( .C1(n22747), .C2(n22666), .A(n15542), .B(n15541), .ZN(
        n15543) );
  AOI21_X1 U17659 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15543), .ZN(n15544) );
  INV_X1 U17660 ( .A(n15544), .ZN(P1_U3102) );
  NAND2_X1 U17661 ( .A1(n22693), .A2(n22646), .ZN(n15546) );
  AOI22_X1 U17662 ( .A1(n22692), .A2(n15608), .B1(n22639), .B2(n22690), .ZN(
        n15545) );
  OAI211_X1 U17663 ( .C1(n22747), .C2(n22644), .A(n15546), .B(n15545), .ZN(
        n15547) );
  AOI21_X1 U17664 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n15547), .ZN(n15548) );
  INV_X1 U17665 ( .A(n15548), .ZN(P1_U3101) );
  NAND2_X1 U17666 ( .A1(n22693), .A2(n22582), .ZN(n15550) );
  AOI22_X1 U17667 ( .A1(n22692), .A2(n15622), .B1(n22575), .B2(n22690), .ZN(
        n15549) );
  OAI211_X1 U17668 ( .C1(n22747), .C2(n22580), .A(n15550), .B(n15549), .ZN(
        n15551) );
  AOI21_X1 U17669 ( .B1(n22694), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n15551), .ZN(n15552) );
  INV_X1 U17670 ( .A(n15552), .ZN(P1_U3098) );
  XNOR2_X1 U17671 ( .A(n15554), .B(n15553), .ZN(n17747) );
  INV_X1 U17672 ( .A(n19497), .ZN(n15555) );
  AOI21_X1 U17673 ( .B1(n17880), .B2(n16415), .A(n15555), .ZN(n16426) );
  NAND2_X1 U17674 ( .A1(n17880), .A2(n16425), .ZN(n16416) );
  OAI211_X1 U17675 ( .C1(n16420), .C2(n17877), .A(n16426), .B(n16416), .ZN(
        n16273) );
  INV_X1 U17676 ( .A(n16273), .ZN(n15557) );
  INV_X1 U17677 ( .A(n16420), .ZN(n18025) );
  OAI21_X1 U17678 ( .B1(n17877), .B2(n18025), .A(n16421), .ZN(n15556) );
  NAND2_X1 U17679 ( .A1(n15556), .A2(n17838), .ZN(n18023) );
  MUX2_X1 U17680 ( .A(n15557), .B(n18023), .S(n16274), .Z(n15561) );
  INV_X1 U17681 ( .A(n20263), .ZN(n20358) );
  INV_X1 U17682 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n18277) );
  NOR2_X1 U17683 ( .A1(n18277), .A2(n14452), .ZN(n15559) );
  AOI21_X1 U17684 ( .B1(n19500), .B2(n20358), .A(n15559), .ZN(n15560) );
  NAND2_X1 U17685 ( .A1(n15561), .A2(n15560), .ZN(n15562) );
  AOI21_X1 U17686 ( .B1(n11196), .B2(n19504), .A(n15562), .ZN(n15567) );
  NAND2_X1 U17687 ( .A1(n15565), .A2(n15564), .ZN(n17751) );
  NAND3_X1 U17688 ( .A1(n15563), .A2(n17751), .A3(n18055), .ZN(n15566) );
  OAI211_X1 U17689 ( .C1(n17747), .C2(n19495), .A(n15567), .B(n15566), .ZN(
        P2_U3043) );
  AOI22_X1 U17690 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20711), .B1(n20708), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15568) );
  OAI21_X1 U17691 ( .B1(n15569), .B2(n15588), .A(n15568), .ZN(P1_U2920) );
  AOI22_X1 U17692 ( .A1(n20708), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15570) );
  OAI21_X1 U17693 ( .B1(n15571), .B2(n15588), .A(n15570), .ZN(P1_U2913) );
  AOI22_X1 U17694 ( .A1(n22130), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15572) );
  OAI21_X1 U17695 ( .B1(n16735), .B2(n15588), .A(n15572), .ZN(P1_U2914) );
  AOI22_X1 U17696 ( .A1(n22130), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15573) );
  OAI21_X1 U17697 ( .B1(n16721), .B2(n15588), .A(n15573), .ZN(P1_U2911) );
  AOI22_X1 U17698 ( .A1(n22130), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15574) );
  OAI21_X1 U17699 ( .B1(n15897), .B2(n15588), .A(n15574), .ZN(P1_U2909) );
  AOI22_X1 U17700 ( .A1(n22130), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15575) );
  OAI21_X1 U17701 ( .B1(n15899), .B2(n15588), .A(n15575), .ZN(P1_U2910) );
  AOI22_X1 U17702 ( .A1(n22130), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15576) );
  OAI21_X1 U17703 ( .B1(n15577), .B2(n15588), .A(n15576), .ZN(P1_U2907) );
  AOI22_X1 U17704 ( .A1(n22130), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15578) );
  OAI21_X1 U17705 ( .B1(n15579), .B2(n15588), .A(n15578), .ZN(P1_U2906) );
  AOI22_X1 U17706 ( .A1(n22130), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15580) );
  OAI21_X1 U17707 ( .B1(n15581), .B2(n15588), .A(n15580), .ZN(P1_U2916) );
  AOI22_X1 U17708 ( .A1(n22130), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15582) );
  OAI21_X1 U17709 ( .B1(n15583), .B2(n15588), .A(n15582), .ZN(P1_U2915) );
  AOI22_X1 U17710 ( .A1(n22130), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15584) );
  OAI21_X1 U17711 ( .B1(n15585), .B2(n15588), .A(n15584), .ZN(P1_U2908) );
  AOI22_X1 U17712 ( .A1(n22130), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15586) );
  OAI21_X1 U17713 ( .B1(n16089), .B2(n15588), .A(n15586), .ZN(P1_U2912) );
  AOI22_X1 U17714 ( .A1(n22130), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15587) );
  OAI21_X1 U17715 ( .B1(n15589), .B2(n15588), .A(n15587), .ZN(P1_U2917) );
  AND2_X1 U17716 ( .A1(n15193), .A2(n15590), .ZN(n15591) );
  OR2_X1 U17717 ( .A1(n15591), .A2(n15640), .ZN(n17987) );
  NOR2_X1 U17718 ( .A1(n17987), .A2(n17432), .ZN(n15595) );
  AOI211_X1 U17719 ( .C1(n15593), .C2(n15192), .A(n17452), .B(n15592), .ZN(
        n15594) );
  AOI211_X1 U17720 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n17432), .A(n15595), .B(
        n15594), .ZN(n15596) );
  INV_X1 U17721 ( .A(n15596), .ZN(P2_U2877) );
  OAI21_X1 U17722 ( .B1(n22728), .B2(n17252), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15598) );
  OAI21_X1 U17723 ( .B1(n22518), .B2(n22502), .A(n15598), .ZN(n15601) );
  INV_X1 U17724 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n15600) );
  NOR2_X1 U17725 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15599), .ZN(
        n17242) );
  AOI21_X1 U17726 ( .B1(n15601), .B2(n15600), .A(n17242), .ZN(n15603) );
  INV_X1 U17727 ( .A(n22548), .ZN(n22507) );
  INV_X1 U17728 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15612) );
  NAND2_X1 U17729 ( .A1(n11222), .A2(n22494), .ZN(n15607) );
  INV_X1 U17730 ( .A(n15604), .ZN(n15605) );
  NAND2_X1 U17731 ( .A1(n15605), .A2(n22473), .ZN(n22464) );
  INV_X1 U17732 ( .A(n22540), .ZN(n15606) );
  OAI22_X1 U17733 ( .A1(n22502), .A2(n15607), .B1(n22464), .B2(n15606), .ZN(
        n17243) );
  AOI22_X1 U17734 ( .A1(n15608), .A2(n17243), .B1(n17242), .B2(n22639), .ZN(
        n15609) );
  OAI21_X1 U17735 ( .B1(n15632), .B2(n22644), .A(n15609), .ZN(n15610) );
  AOI21_X1 U17736 ( .B1(n22728), .B2(n22646), .A(n15610), .ZN(n15611) );
  OAI21_X1 U17737 ( .B1(n17235), .B2(n15612), .A(n15611), .ZN(P1_U3069) );
  INV_X1 U17738 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U17739 ( .A1(n15613), .A2(n17243), .B1(n17242), .B2(n22661), .ZN(
        n15614) );
  OAI21_X1 U17740 ( .B1(n15632), .B2(n22666), .A(n15614), .ZN(n15615) );
  AOI21_X1 U17741 ( .B1(n22728), .B2(n22668), .A(n15615), .ZN(n15616) );
  OAI21_X1 U17742 ( .B1(n17235), .B2(n15617), .A(n15616), .ZN(P1_U3070) );
  INV_X1 U17743 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15621) );
  AOI22_X1 U17744 ( .A1(n22560), .A2(n17243), .B1(n17242), .B2(n22559), .ZN(
        n15618) );
  OAI21_X1 U17745 ( .B1(n15632), .B2(n22544), .A(n15618), .ZN(n15619) );
  AOI21_X1 U17746 ( .B1(n22728), .B2(n22552), .A(n15619), .ZN(n15620) );
  OAI21_X1 U17747 ( .B1(n17235), .B2(n15621), .A(n15620), .ZN(P1_U3065) );
  INV_X1 U17748 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U17749 ( .A1(n15622), .A2(n17243), .B1(n17242), .B2(n22575), .ZN(
        n15623) );
  OAI21_X1 U17750 ( .B1(n15632), .B2(n22580), .A(n15623), .ZN(n15624) );
  AOI21_X1 U17751 ( .B1(n22728), .B2(n22582), .A(n15624), .ZN(n15625) );
  OAI21_X1 U17752 ( .B1(n17235), .B2(n15626), .A(n15625), .ZN(P1_U3066) );
  INV_X1 U17753 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U17754 ( .A1(n22691), .A2(n17243), .B1(n17242), .B2(n22697), .ZN(
        n15627) );
  OAI21_X1 U17755 ( .B1(n15632), .B2(n22713), .A(n15627), .ZN(n15628) );
  AOI21_X1 U17756 ( .B1(n22728), .B2(n22709), .A(n15628), .ZN(n15629) );
  OAI21_X1 U17757 ( .B1(n17235), .B2(n15630), .A(n15629), .ZN(P1_U3071) );
  INV_X1 U17758 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U17759 ( .A1(n22775), .A2(n17243), .B1(n17242), .B2(n22773), .ZN(
        n15631) );
  OAI21_X1 U17760 ( .B1(n15632), .B2(n22757), .A(n15631), .ZN(n15633) );
  AOI21_X1 U17761 ( .B1(n22728), .B2(n22760), .A(n15633), .ZN(n15634) );
  OAI21_X1 U17762 ( .B1(n17235), .B2(n15635), .A(n15634), .ZN(P1_U3072) );
  INV_X1 U17763 ( .A(n15636), .ZN(n15637) );
  OAI211_X1 U17764 ( .C1(n15592), .C2(n15638), .A(n15637), .B(n17419), .ZN(
        n15644) );
  OR2_X1 U17765 ( .A1(n15640), .A2(n15639), .ZN(n15641) );
  NAND2_X1 U17766 ( .A1(n15666), .A2(n15641), .ZN(n17971) );
  INV_X1 U17767 ( .A(n17971), .ZN(n15642) );
  NAND2_X1 U17768 ( .A1(n15642), .A2(n17411), .ZN(n15643) );
  OAI211_X1 U17769 ( .C1(n17411), .C2(n12227), .A(n15644), .B(n15643), .ZN(
        P2_U2876) );
  AOI211_X1 U17770 ( .C1(n19259), .C2(n15646), .A(n11184), .B(n15645), .ZN(
        n17353) );
  AOI21_X1 U17771 ( .B1(n11184), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17353), .ZN(n18072) );
  INV_X1 U17772 ( .A(n18072), .ZN(n15648) );
  NOR2_X1 U17773 ( .A1(n15647), .A2(n18105), .ZN(n18073) );
  AOI222_X1 U17774 ( .A1(n15649), .A2(n18078), .B1(n19529), .B2(n18220), .C1(
        n15648), .C2(n18073), .ZN(n15651) );
  NAND2_X1 U17775 ( .A1(n18076), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15650) );
  OAI21_X1 U17776 ( .B1(n15651), .B2(n18076), .A(n15650), .ZN(P2_U3599) );
  AND2_X1 U17777 ( .A1(n15251), .A2(n15653), .ZN(n15654) );
  NOR2_X1 U17778 ( .A1(n15652), .A2(n15654), .ZN(n22271) );
  INV_X1 U17779 ( .A(n22271), .ZN(n15657) );
  INV_X1 U17780 ( .A(n16743), .ZN(n15655) );
  OAI222_X1 U17781 ( .A1(n15657), .A2(n16782), .B1(n16791), .B2(n15656), .C1(
        n15655), .C2(n16794), .ZN(P1_U2899) );
  OR2_X1 U17782 ( .A1(n15652), .A2(n15659), .ZN(n15660) );
  AND2_X1 U17783 ( .A1(n15658), .A2(n15660), .ZN(n22284) );
  INV_X1 U17784 ( .A(n22284), .ZN(n15663) );
  OAI222_X1 U17785 ( .A1(n16794), .A2(n16736), .B1(n16791), .B2(n13562), .C1(
        n16782), .C2(n15663), .ZN(P1_U2898) );
  NAND2_X1 U17786 ( .A1(n20825), .A2(n15661), .ZN(n15662) );
  NAND2_X1 U17787 ( .A1(n20817), .A2(n15662), .ZN(n22276) );
  OAI222_X1 U17788 ( .A1(n22276), .A2(n20820), .B1(n22275), .B2(n20830), .C1(
        n20805), .C2(n15663), .ZN(P1_U2866) );
  INV_X1 U17789 ( .A(n15664), .ZN(n16257) );
  NAND2_X1 U17790 ( .A1(n15666), .A2(n15665), .ZN(n15667) );
  AND2_X1 U17791 ( .A1(n16257), .A2(n15667), .ZN(n19327) );
  INV_X1 U17792 ( .A(n19327), .ZN(n15672) );
  OAI211_X1 U17793 ( .C1(n15636), .C2(n15669), .A(n15668), .B(n17419), .ZN(
        n15671) );
  NAND2_X1 U17794 ( .A1(n17432), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15670) );
  OAI211_X1 U17795 ( .C1(n15672), .C2(n17432), .A(n15671), .B(n15670), .ZN(
        P2_U2875) );
  NAND2_X1 U17796 ( .A1(n15658), .A2(n15674), .ZN(n15675) );
  AND2_X1 U17797 ( .A1(n15673), .A2(n15675), .ZN(n22298) );
  INV_X1 U17798 ( .A(n22298), .ZN(n15678) );
  INV_X1 U17799 ( .A(n16731), .ZN(n15677) );
  OAI222_X1 U17800 ( .A1(n15678), .A2(n16782), .B1(n16794), .B2(n15677), .C1(
        n15676), .C2(n16791), .ZN(P1_U2897) );
  AOI21_X1 U17801 ( .B1(n22782), .B2(n15684), .A(n15972), .ZN(n15679) );
  AOI21_X1 U17802 ( .B1(n22538), .B2(n22518), .A(n15679), .ZN(n15680) );
  NOR2_X1 U17803 ( .A1(n15680), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15683) );
  NOR3_X1 U17804 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15681), .A3(
        n22505), .ZN(n15688) );
  INV_X1 U17805 ( .A(n22473), .ZN(n15682) );
  NAND2_X1 U17806 ( .A1(n15682), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15685) );
  NAND2_X1 U17807 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15685), .ZN(n22525) );
  NAND2_X1 U17808 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n15691) );
  NAND3_X1 U17809 ( .A1(n22538), .A2(n22518), .A3(n22494), .ZN(n15687) );
  INV_X1 U17810 ( .A(n15685), .ZN(n22520) );
  NAND2_X1 U17811 ( .A1(n22520), .A2(n22540), .ZN(n15686) );
  AND2_X1 U17812 ( .A1(n15687), .A2(n15686), .ZN(n22707) );
  INV_X1 U17813 ( .A(n15688), .ZN(n22704) );
  OAI22_X1 U17814 ( .A1(n22585), .A2(n22707), .B1(n22579), .B2(n22704), .ZN(
        n15689) );
  AOI21_X1 U17815 ( .B1(n22768), .B2(n22582), .A(n15689), .ZN(n15690) );
  OAI211_X1 U17816 ( .C1(n22580), .C2(n22782), .A(n15691), .B(n15690), .ZN(
        P1_U3146) );
  NAND2_X1 U17817 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n15694) );
  OAI22_X1 U17818 ( .A1(n22627), .A2(n22707), .B1(n22621), .B2(n22704), .ZN(
        n15692) );
  AOI21_X1 U17819 ( .B1(n22768), .B2(n22624), .A(n15692), .ZN(n15693) );
  OAI211_X1 U17820 ( .C1(n22622), .C2(n22782), .A(n15694), .B(n15693), .ZN(
        P1_U3148) );
  NAND2_X1 U17821 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n15697) );
  OAI22_X1 U17822 ( .A1(n22707), .A2(n22671), .B1(n22665), .B2(n22704), .ZN(
        n15695) );
  AOI21_X1 U17823 ( .B1(n22768), .B2(n22668), .A(n15695), .ZN(n15696) );
  OAI211_X1 U17824 ( .C1(n22666), .C2(n22782), .A(n15697), .B(n15696), .ZN(
        P1_U3150) );
  NAND2_X1 U17825 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n15700) );
  OAI22_X1 U17826 ( .A1(n22707), .A2(n22764), .B1(n22755), .B2(n22704), .ZN(
        n15698) );
  AOI21_X1 U17827 ( .B1(n22768), .B2(n22760), .A(n15698), .ZN(n15699) );
  OAI211_X1 U17828 ( .C1(n22757), .C2(n22782), .A(n15700), .B(n15699), .ZN(
        P1_U3152) );
  NAND2_X1 U17829 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n15703) );
  OAI22_X1 U17830 ( .A1(n22605), .A2(n22707), .B1(n22599), .B2(n22704), .ZN(
        n15701) );
  AOI21_X1 U17831 ( .B1(n22768), .B2(n22602), .A(n15701), .ZN(n15702) );
  OAI211_X1 U17832 ( .C1(n22600), .C2(n22782), .A(n15703), .B(n15702), .ZN(
        P1_U3147) );
  NAND2_X1 U17833 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n15706) );
  OAI22_X1 U17834 ( .A1(n22707), .A2(n22649), .B1(n22643), .B2(n22704), .ZN(
        n15704) );
  AOI21_X1 U17835 ( .B1(n22768), .B2(n22646), .A(n15704), .ZN(n15705) );
  OAI211_X1 U17836 ( .C1(n22644), .C2(n22782), .A(n15706), .B(n15705), .ZN(
        P1_U3149) );
  NAND2_X1 U17837 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n15709) );
  OAI22_X1 U17838 ( .A1(n22707), .A2(n22555), .B1(n22543), .B2(n22704), .ZN(
        n15707) );
  AOI21_X1 U17839 ( .B1(n22768), .B2(n22552), .A(n15707), .ZN(n15708) );
  OAI211_X1 U17840 ( .C1(n22544), .C2(n22782), .A(n15709), .B(n15708), .ZN(
        P1_U3145) );
  NAND2_X1 U17841 ( .A1(n20255), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n18209) );
  NAND3_X1 U17842 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20038) );
  OAI21_X1 U17843 ( .B1(n15710), .B2(n18209), .A(n20038), .ZN(n15715) );
  INV_X1 U17844 ( .A(n20195), .ZN(n15712) );
  INV_X1 U17845 ( .A(n20198), .ZN(n20529) );
  NAND2_X1 U17846 ( .A1(n20199), .A2(n20529), .ZN(n15711) );
  OAI211_X1 U17847 ( .C1(n15713), .C2(n20180), .A(n15712), .B(n15711), .ZN(
        n15714) );
  NAND2_X1 U17848 ( .A1(n15715), .A2(n15714), .ZN(n20534) );
  INV_X1 U17849 ( .A(n20534), .ZN(n20470) );
  INV_X1 U17850 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15724) );
  OAI21_X1 U17851 ( .B1(n15716), .B2(n20529), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15717) );
  OAI21_X1 U17852 ( .B1(n20038), .B2(n20192), .A(n15717), .ZN(n20530) );
  INV_X1 U17853 ( .A(n20190), .ZN(n16288) );
  NAND2_X1 U17854 ( .A1(n20255), .A2(n19269), .ZN(n20100) );
  INV_X1 U17855 ( .A(n20100), .ZN(n15718) );
  INV_X1 U17856 ( .A(n20144), .ZN(n15719) );
  AOI22_X1 U17857 ( .A1(n20533), .A2(n20191), .B1(n20471), .B2(n20185), .ZN(
        n15721) );
  OAI21_X1 U17858 ( .B1(n16288), .B2(n20198), .A(n15721), .ZN(n15722) );
  AOI21_X1 U17859 ( .B1(n20530), .B2(n15512), .A(n15722), .ZN(n15723) );
  OAI21_X1 U17860 ( .B1(n20470), .B2(n15724), .A(n15723), .ZN(P2_U3175) );
  XOR2_X1 U17861 ( .A(DATAI_30_), .B(keyinput_2), .Z(n15728) );
  XNOR2_X1 U17862 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .ZN(n15727) );
  XNOR2_X1 U17863 ( .A(DATAI_29_), .B(keyinput_3), .ZN(n15726) );
  XNOR2_X1 U17864 ( .A(DATAI_31_), .B(keyinput_1), .ZN(n15725) );
  NOR4_X1 U17865 ( .A1(n15728), .A2(n15727), .A3(n15726), .A4(n15725), .ZN(
        n15731) );
  XOR2_X1 U17866 ( .A(DATAI_25_), .B(keyinput_7), .Z(n15730) );
  XNOR2_X1 U17867 ( .A(DATAI_28_), .B(keyinput_4), .ZN(n15729) );
  NOR3_X1 U17868 ( .A1(n15731), .A2(n15730), .A3(n15729), .ZN(n15736) );
  INV_X1 U17869 ( .A(keyinput_8), .ZN(n15732) );
  XNOR2_X1 U17870 ( .A(n15732), .B(DATAI_24_), .ZN(n15735) );
  XNOR2_X1 U17871 ( .A(DATAI_27_), .B(keyinput_5), .ZN(n15734) );
  XNOR2_X1 U17872 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n15733) );
  NAND4_X1 U17873 ( .A1(n15736), .A2(n15735), .A3(n15734), .A4(n15733), .ZN(
        n15739) );
  XOR2_X1 U17874 ( .A(DATAI_23_), .B(keyinput_9), .Z(n15738) );
  XNOR2_X1 U17875 ( .A(n14975), .B(keyinput_10), .ZN(n15737) );
  NAND3_X1 U17876 ( .A1(n15739), .A2(n15738), .A3(n15737), .ZN(n15743) );
  XOR2_X1 U17877 ( .A(DATAI_19_), .B(keyinput_13), .Z(n15742) );
  XNOR2_X1 U17878 ( .A(DATAI_20_), .B(keyinput_12), .ZN(n15741) );
  XNOR2_X1 U17879 ( .A(DATAI_21_), .B(keyinput_11), .ZN(n15740) );
  NAND4_X1 U17880 ( .A1(n15743), .A2(n15742), .A3(n15741), .A4(n15740), .ZN(
        n15746) );
  XNOR2_X1 U17881 ( .A(DATAI_17_), .B(keyinput_15), .ZN(n15745) );
  XNOR2_X1 U17882 ( .A(DATAI_18_), .B(keyinput_14), .ZN(n15744) );
  NAND3_X1 U17883 ( .A1(n15746), .A2(n15745), .A3(n15744), .ZN(n15750) );
  XNOR2_X1 U17884 ( .A(DATAI_16_), .B(keyinput_16), .ZN(n15749) );
  XNOR2_X1 U17885 ( .A(n15930), .B(keyinput_17), .ZN(n15748) );
  XOR2_X1 U17886 ( .A(DATAI_14_), .B(keyinput_18), .Z(n15747) );
  AOI211_X1 U17887 ( .C1(n15750), .C2(n15749), .A(n15748), .B(n15747), .ZN(
        n15754) );
  XNOR2_X1 U17888 ( .A(DATAI_13_), .B(keyinput_19), .ZN(n15753) );
  XOR2_X1 U17889 ( .A(DATAI_11_), .B(keyinput_21), .Z(n15752) );
  XNOR2_X1 U17890 ( .A(DATAI_12_), .B(keyinput_20), .ZN(n15751) );
  OAI211_X1 U17891 ( .C1(n15754), .C2(n15753), .A(n15752), .B(n15751), .ZN(
        n15757) );
  XOR2_X1 U17892 ( .A(DATAI_10_), .B(keyinput_22), .Z(n15756) );
  XNOR2_X1 U17893 ( .A(DATAI_9_), .B(keyinput_23), .ZN(n15755) );
  AOI21_X1 U17894 ( .B1(n15757), .B2(n15756), .A(n15755), .ZN(n15760) );
  XNOR2_X1 U17895 ( .A(n15942), .B(keyinput_25), .ZN(n15759) );
  XOR2_X1 U17896 ( .A(DATAI_8_), .B(keyinput_24), .Z(n15758) );
  NOR3_X1 U17897 ( .A1(n15760), .A2(n15759), .A3(n15758), .ZN(n15764) );
  XOR2_X1 U17898 ( .A(DATAI_6_), .B(keyinput_26), .Z(n15763) );
  XOR2_X1 U17899 ( .A(DATAI_4_), .B(keyinput_28), .Z(n15762) );
  XNOR2_X1 U17900 ( .A(DATAI_5_), .B(keyinput_27), .ZN(n15761) );
  OAI211_X1 U17901 ( .C1(n15764), .C2(n15763), .A(n15762), .B(n15761), .ZN(
        n15767) );
  XNOR2_X1 U17902 ( .A(DATAI_3_), .B(keyinput_29), .ZN(n15766) );
  XNOR2_X1 U17903 ( .A(DATAI_2_), .B(keyinput_30), .ZN(n15765) );
  NAND3_X1 U17904 ( .A1(n15767), .A2(n15766), .A3(n15765), .ZN(n15776) );
  XOR2_X1 U17905 ( .A(DATAI_1_), .B(keyinput_31), .Z(n15775) );
  XOR2_X1 U17906 ( .A(HOLD), .B(keyinput_33), .Z(n15770) );
  XNOR2_X1 U17907 ( .A(READY1), .B(keyinput_36), .ZN(n15769) );
  XNOR2_X1 U17908 ( .A(DATAI_0_), .B(keyinput_32), .ZN(n15768) );
  NOR3_X1 U17909 ( .A1(n15770), .A2(n15769), .A3(n15768), .ZN(n15773) );
  XOR2_X1 U17910 ( .A(BS16), .B(keyinput_35), .Z(n15772) );
  XOR2_X1 U17911 ( .A(NA), .B(keyinput_34), .Z(n15771) );
  NAND3_X1 U17912 ( .A1(n15773), .A2(n15772), .A3(n15771), .ZN(n15774) );
  AOI21_X1 U17913 ( .B1(n15776), .B2(n15775), .A(n15774), .ZN(n15779) );
  XOR2_X1 U17914 ( .A(READY2), .B(keyinput_37), .Z(n15778) );
  XNOR2_X1 U17915 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_38), .ZN(
        n15777) );
  NOR3_X1 U17916 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n15783) );
  XOR2_X1 U17917 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_39), .Z(n15782) );
  XOR2_X1 U17918 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_40), .Z(n15781)
         );
  XOR2_X1 U17919 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_41), .Z(n15780) );
  OAI211_X1 U17920 ( .C1(n15783), .C2(n15782), .A(n15781), .B(n15780), .ZN(
        n15786) );
  XNOR2_X1 U17921 ( .A(P1_D_C_N_REG_SCAN_IN), .B(keyinput_42), .ZN(n15785) );
  XNOR2_X1 U17922 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .ZN(
        n15784) );
  AOI21_X1 U17923 ( .B1(n15786), .B2(n15785), .A(n15784), .ZN(n15790) );
  XNOR2_X1 U17924 ( .A(n15972), .B(keyinput_44), .ZN(n15789) );
  XNOR2_X1 U17925 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_46), .ZN(n15788) );
  XNOR2_X1 U17926 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_45), .ZN(n15787) );
  NOR4_X1 U17927 ( .A1(n15790), .A2(n15789), .A3(n15788), .A4(n15787), .ZN(
        n15796) );
  XOR2_X1 U17928 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .Z(n15795) );
  INV_X1 U17929 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20799) );
  XNOR2_X1 U17930 ( .A(n20799), .B(keyinput_49), .ZN(n15793) );
  INV_X1 U17931 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20802) );
  XNOR2_X1 U17932 ( .A(n20802), .B(keyinput_48), .ZN(n15792) );
  INV_X1 U17933 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20794) );
  XNOR2_X1 U17934 ( .A(n20794), .B(keyinput_50), .ZN(n15791) );
  NOR3_X1 U17935 ( .A1(n15793), .A2(n15792), .A3(n15791), .ZN(n15794) );
  OAI21_X1 U17936 ( .B1(n15796), .B2(n15795), .A(n15794), .ZN(n15804) );
  INV_X1 U17937 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20789) );
  XNOR2_X1 U17938 ( .A(n20789), .B(keyinput_51), .ZN(n15803) );
  XOR2_X1 U17939 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_55), .Z(n15802) );
  XOR2_X1 U17940 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .Z(n15800) );
  XOR2_X1 U17941 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_54), .Z(n15799) );
  XOR2_X1 U17942 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .Z(n15798) );
  XOR2_X1 U17943 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .Z(n15797) );
  NOR4_X1 U17944 ( .A1(n15800), .A2(n15799), .A3(n15798), .A4(n15797), .ZN(
        n15801) );
  NAND4_X1 U17945 ( .A1(n15804), .A2(n15803), .A3(n15802), .A4(n15801), .ZN(
        n15807) );
  XOR2_X1 U17946 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_58), .Z(n15806) );
  XNOR2_X1 U17947 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_57), .ZN(n15805)
         );
  NAND3_X1 U17948 ( .A1(n15807), .A2(n15806), .A3(n15805), .ZN(n15816) );
  XOR2_X1 U17949 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_59), .Z(n15815) );
  XOR2_X1 U17950 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_61), .Z(n15810) );
  XOR2_X1 U17951 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_63), .Z(n15809) );
  XNOR2_X1 U17952 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_60), .ZN(n15808)
         );
  NOR3_X1 U17953 ( .A1(n15810), .A2(n15809), .A3(n15808), .ZN(n15813) );
  XOR2_X1 U17954 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_64), .Z(n15812) );
  XOR2_X1 U17955 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_62), .Z(n15811) );
  NAND3_X1 U17956 ( .A1(n15813), .A2(n15812), .A3(n15811), .ZN(n15814) );
  AOI21_X1 U17957 ( .B1(n15816), .B2(n15815), .A(n15814), .ZN(n15819) );
  XOR2_X1 U17958 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_65), .Z(n15818) );
  XNOR2_X1 U17959 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_66), .ZN(n15817)
         );
  NOR3_X1 U17960 ( .A1(n15819), .A2(n15818), .A3(n15817), .ZN(n15823) );
  XNOR2_X1 U17961 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_67), .ZN(n15822)
         );
  XOR2_X1 U17962 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_69), .Z(n15821) );
  XNOR2_X1 U17963 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_68), .ZN(n15820)
         );
  OAI211_X1 U17964 ( .C1(n15823), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        n15831) );
  XOR2_X1 U17965 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_70), .Z(n15830) );
  INV_X1 U17966 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n22317) );
  OAI22_X1 U17967 ( .A1(n22317), .A2(keyinput_72), .B1(n16950), .B2(
        keyinput_71), .ZN(n15824) );
  AOI221_X1 U17968 ( .B1(n22317), .B2(keyinput_72), .C1(keyinput_71), .C2(
        n16950), .A(n15824), .ZN(n15828) );
  INV_X1 U17969 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20731) );
  OAI22_X1 U17970 ( .A1(n20731), .A2(keyinput_75), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(keyinput_74), .ZN(n15825) );
  AOI221_X1 U17971 ( .B1(n20731), .B2(keyinput_75), .C1(keyinput_74), .C2(
        P1_REIP_REG_9__SCAN_IN), .A(n15825), .ZN(n15827) );
  XOR2_X1 U17972 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .Z(n15826) );
  NAND3_X1 U17973 ( .A1(n15828), .A2(n15827), .A3(n15826), .ZN(n15829) );
  AOI21_X1 U17974 ( .B1(n15831), .B2(n15830), .A(n15829), .ZN(n15835) );
  XOR2_X1 U17975 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_78), .Z(n15834) );
  XOR2_X1 U17976 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_76), .Z(n15833) );
  XOR2_X1 U17977 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_77), .Z(n15832) );
  NOR4_X1 U17978 ( .A1(n15835), .A2(n15834), .A3(n15833), .A4(n15832), .ZN(
        n15838) );
  XOR2_X1 U17979 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_79), .Z(n15837) );
  XOR2_X1 U17980 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_80), .Z(n15836) );
  OAI21_X1 U17981 ( .B1(n15838), .B2(n15837), .A(n15836), .ZN(n15841) );
  XNOR2_X1 U17982 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_81), .ZN(n15840)
         );
  XNOR2_X1 U17983 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_82), .ZN(n15839)
         );
  AOI21_X1 U17984 ( .B1(n15841), .B2(n15840), .A(n15839), .ZN(n15844) );
  XOR2_X1 U17985 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_83), .Z(n15843) );
  XOR2_X1 U17986 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .Z(n15842) );
  NOR3_X1 U17987 ( .A1(n15844), .A2(n15843), .A3(n15842), .ZN(n15847) );
  XOR2_X1 U17988 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_85), .Z(n15846) );
  XNOR2_X1 U17989 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_86), .ZN(n15845)
         );
  NOR3_X1 U17990 ( .A1(n15847), .A2(n15846), .A3(n15845), .ZN(n15852) );
  XNOR2_X1 U17991 ( .A(n15848), .B(keyinput_88), .ZN(n15851) );
  XNOR2_X1 U17992 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_87), .ZN(n15850)
         );
  XNOR2_X1 U17993 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_89), .ZN(n15849)
         );
  NOR4_X1 U17994 ( .A1(n15852), .A2(n15851), .A3(n15850), .A4(n15849), .ZN(
        n15856) );
  XNOR2_X1 U17995 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .ZN(n15855)
         );
  XNOR2_X1 U17996 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_91), .ZN(n15854)
         );
  XNOR2_X1 U17997 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_92), .ZN(n15853)
         );
  OAI211_X1 U17998 ( .C1(n15856), .C2(n15855), .A(n15854), .B(n15853), .ZN(
        n15859) );
  XNOR2_X1 U17999 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_93), .ZN(n15858)
         );
  XOR2_X1 U18000 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_94), .Z(n15857) );
  AOI21_X1 U18001 ( .B1(n15859), .B2(n15858), .A(n15857), .ZN(n15862) );
  XNOR2_X1 U18002 ( .A(n16690), .B(keyinput_95), .ZN(n15861) );
  XNOR2_X1 U18003 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_96), .ZN(n15860)
         );
  NOR3_X1 U18004 ( .A1(n15862), .A2(n15861), .A3(n15860), .ZN(n15866) );
  XNOR2_X1 U18005 ( .A(n16052), .B(keyinput_97), .ZN(n15865) );
  XOR2_X1 U18006 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .Z(n15864) );
  XNOR2_X1 U18007 ( .A(n16692), .B(keyinput_99), .ZN(n15863) );
  OAI211_X1 U18008 ( .C1(n15866), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        n15872) );
  XNOR2_X1 U18009 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_100), .ZN(n15871)
         );
  XOR2_X1 U18010 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_102), .Z(n15869) );
  XNOR2_X1 U18011 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n15868)
         );
  XNOR2_X1 U18012 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n15867)
         );
  NAND3_X1 U18013 ( .A1(n15869), .A2(n15868), .A3(n15867), .ZN(n15870) );
  AOI21_X1 U18014 ( .B1(n15872), .B2(n15871), .A(n15870), .ZN(n15875) );
  XNOR2_X1 U18015 ( .A(n16063), .B(keyinput_104), .ZN(n15874) );
  XNOR2_X1 U18016 ( .A(n16363), .B(keyinput_105), .ZN(n15873) );
  OAI21_X1 U18017 ( .B1(n15875), .B2(n15874), .A(n15873), .ZN(n15878) );
  XOR2_X1 U18018 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_106), .Z(n15877) );
  XNOR2_X1 U18019 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n15876)
         );
  AOI21_X1 U18020 ( .B1(n15878), .B2(n15877), .A(n15876), .ZN(n15882) );
  XNOR2_X1 U18021 ( .A(n22275), .B(keyinput_109), .ZN(n15881) );
  XNOR2_X1 U18022 ( .A(n20829), .B(keyinput_110), .ZN(n15880) );
  XOR2_X1 U18023 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .Z(n15879) );
  NOR4_X1 U18024 ( .A1(n15882), .A2(n15881), .A3(n15880), .A4(n15879), .ZN(
        n15886) );
  XNOR2_X1 U18025 ( .A(n16074), .B(keyinput_111), .ZN(n15885) );
  XOR2_X1 U18026 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .Z(n15884) );
  XOR2_X1 U18027 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_113), .Z(n15883) );
  OAI211_X1 U18028 ( .C1(n15886), .C2(n15885), .A(n15884), .B(n15883), .ZN(
        n15889) );
  XNOR2_X1 U18029 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_114), .ZN(n15888)
         );
  XNOR2_X1 U18030 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_115), .ZN(n15887)
         );
  AOI21_X1 U18031 ( .B1(n15889), .B2(n15888), .A(n15887), .ZN(n15892) );
  XNOR2_X1 U18032 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_116), .ZN(n15891)
         );
  XNOR2_X1 U18033 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n15890)
         );
  OAI21_X1 U18034 ( .B1(n15892), .B2(n15891), .A(n15890), .ZN(n15895) );
  XOR2_X1 U18035 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_118), .Z(n15894) );
  XNOR2_X1 U18036 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_119), .ZN(n15893)
         );
  AOI21_X1 U18037 ( .B1(n15895), .B2(n15894), .A(n15893), .ZN(n15903) );
  AOI22_X1 U18038 ( .A1(n16721), .A2(keyinput_122), .B1(keyinput_120), .B2(
        n15897), .ZN(n15896) );
  OAI221_X1 U18039 ( .B1(n16721), .B2(keyinput_122), .C1(n15897), .C2(
        keyinput_120), .A(n15896), .ZN(n15902) );
  AOI22_X1 U18040 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_123), .B1(n15899), .B2(keyinput_121), .ZN(n15898) );
  OAI221_X1 U18041 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_123), .C1(
        n15899), .C2(keyinput_121), .A(n15898), .ZN(n15901) );
  XNOR2_X1 U18042 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .ZN(n15900)
         );
  NOR4_X1 U18043 ( .A1(n15903), .A2(n15902), .A3(n15901), .A4(n15900), .ZN(
        n15906) );
  XNOR2_X1 U18044 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .ZN(n15905)
         );
  XNOR2_X1 U18045 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .ZN(n15904)
         );
  OAI21_X1 U18046 ( .B1(n15906), .B2(n15905), .A(n15904), .ZN(n16101) );
  XNOR2_X1 U18047 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_127), .ZN(n16100)
         );
  XOR2_X1 U18048 ( .A(DATAI_30_), .B(keyinput_130), .Z(n15911) );
  XOR2_X1 U18049 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_128), .Z(n15910) );
  XNOR2_X1 U18050 ( .A(n15907), .B(keyinput_129), .ZN(n15909) );
  XNOR2_X1 U18051 ( .A(DATAI_29_), .B(keyinput_131), .ZN(n15908) );
  NAND4_X1 U18052 ( .A1(n15911), .A2(n15910), .A3(n15909), .A4(n15908), .ZN(
        n15914) );
  XOR2_X1 U18053 ( .A(DATAI_26_), .B(keyinput_134), .Z(n15913) );
  XNOR2_X1 U18054 ( .A(DATAI_27_), .B(keyinput_133), .ZN(n15912) );
  NAND3_X1 U18055 ( .A1(n15914), .A2(n15913), .A3(n15912), .ZN(n15919) );
  XNOR2_X1 U18056 ( .A(DATAI_24_), .B(keyinput_136), .ZN(n15918) );
  XNOR2_X1 U18057 ( .A(DATAI_28_), .B(keyinput_132), .ZN(n15916) );
  XNOR2_X1 U18058 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n15915) );
  NAND2_X1 U18059 ( .A1(n15916), .A2(n15915), .ZN(n15917) );
  NOR3_X1 U18060 ( .A1(n15919), .A2(n15918), .A3(n15917), .ZN(n15922) );
  XOR2_X1 U18061 ( .A(DATAI_23_), .B(keyinput_137), .Z(n15921) );
  XNOR2_X1 U18062 ( .A(DATAI_22_), .B(keyinput_138), .ZN(n15920) );
  NOR3_X1 U18063 ( .A1(n15922), .A2(n15921), .A3(n15920), .ZN(n15926) );
  XOR2_X1 U18064 ( .A(DATAI_19_), .B(keyinput_141), .Z(n15925) );
  XOR2_X1 U18065 ( .A(DATAI_20_), .B(keyinput_140), .Z(n15924) );
  XOR2_X1 U18066 ( .A(DATAI_21_), .B(keyinput_139), .Z(n15923) );
  NOR4_X1 U18067 ( .A1(n15926), .A2(n15925), .A3(n15924), .A4(n15923), .ZN(
        n15929) );
  XOR2_X1 U18068 ( .A(DATAI_18_), .B(keyinput_142), .Z(n15928) );
  XNOR2_X1 U18069 ( .A(DATAI_17_), .B(keyinput_143), .ZN(n15927) );
  NOR3_X1 U18070 ( .A1(n15929), .A2(n15928), .A3(n15927), .ZN(n15934) );
  XNOR2_X1 U18071 ( .A(DATAI_16_), .B(keyinput_144), .ZN(n15933) );
  XNOR2_X1 U18072 ( .A(n15930), .B(keyinput_145), .ZN(n15932) );
  XOR2_X1 U18073 ( .A(DATAI_14_), .B(keyinput_146), .Z(n15931) );
  OAI211_X1 U18074 ( .C1(n15934), .C2(n15933), .A(n15932), .B(n15931), .ZN(
        n15938) );
  XOR2_X1 U18075 ( .A(DATAI_13_), .B(keyinput_147), .Z(n15937) );
  XNOR2_X1 U18076 ( .A(DATAI_12_), .B(keyinput_148), .ZN(n15936) );
  XNOR2_X1 U18077 ( .A(DATAI_11_), .B(keyinput_149), .ZN(n15935) );
  AOI211_X1 U18078 ( .C1(n15938), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        n15941) );
  XNOR2_X1 U18079 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n15940) );
  XNOR2_X1 U18080 ( .A(DATAI_9_), .B(keyinput_151), .ZN(n15939) );
  OAI21_X1 U18081 ( .B1(n15941), .B2(n15940), .A(n15939), .ZN(n15945) );
  XNOR2_X1 U18082 ( .A(n15942), .B(keyinput_153), .ZN(n15944) );
  XNOR2_X1 U18083 ( .A(DATAI_8_), .B(keyinput_152), .ZN(n15943) );
  NAND3_X1 U18084 ( .A1(n15945), .A2(n15944), .A3(n15943), .ZN(n15949) );
  XOR2_X1 U18085 ( .A(DATAI_6_), .B(keyinput_154), .Z(n15948) );
  XOR2_X1 U18086 ( .A(DATAI_4_), .B(keyinput_156), .Z(n15947) );
  XNOR2_X1 U18087 ( .A(DATAI_5_), .B(keyinput_155), .ZN(n15946) );
  AOI211_X1 U18088 ( .C1(n15949), .C2(n15948), .A(n15947), .B(n15946), .ZN(
        n15952) );
  XOR2_X1 U18089 ( .A(DATAI_3_), .B(keyinput_157), .Z(n15951) );
  XOR2_X1 U18090 ( .A(DATAI_2_), .B(keyinput_158), .Z(n15950) );
  NOR3_X1 U18091 ( .A1(n15952), .A2(n15951), .A3(n15950), .ZN(n15961) );
  XOR2_X1 U18092 ( .A(DATAI_1_), .B(keyinput_159), .Z(n15960) );
  XOR2_X1 U18093 ( .A(BS16), .B(keyinput_163), .Z(n15955) );
  XNOR2_X1 U18094 ( .A(DATAI_0_), .B(keyinput_160), .ZN(n15954) );
  XNOR2_X1 U18095 ( .A(READY1), .B(keyinput_164), .ZN(n15953) );
  NAND3_X1 U18096 ( .A1(n15955), .A2(n15954), .A3(n15953), .ZN(n15958) );
  XOR2_X1 U18097 ( .A(HOLD), .B(keyinput_161), .Z(n15957) );
  XNOR2_X1 U18098 ( .A(NA), .B(keyinput_162), .ZN(n15956) );
  NOR3_X1 U18099 ( .A1(n15958), .A2(n15957), .A3(n15956), .ZN(n15959) );
  OAI21_X1 U18100 ( .B1(n15961), .B2(n15960), .A(n15959), .ZN(n15964) );
  XOR2_X1 U18101 ( .A(READY2), .B(keyinput_165), .Z(n15963) );
  XNOR2_X1 U18102 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_166), .ZN(
        n15962) );
  NAND3_X1 U18103 ( .A1(n15964), .A2(n15963), .A3(n15962), .ZN(n15968) );
  XNOR2_X1 U18104 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_167), .ZN(n15967) );
  XOR2_X1 U18105 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_169), .Z(n15966) );
  XNOR2_X1 U18106 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_168), .ZN(n15965) );
  AOI211_X1 U18107 ( .C1(n15968), .C2(n15967), .A(n15966), .B(n15965), .ZN(
        n15971) );
  XOR2_X1 U18108 ( .A(P1_D_C_N_REG_SCAN_IN), .B(keyinput_170), .Z(n15970) );
  XOR2_X1 U18109 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_171), .Z(
        n15969) );
  OAI21_X1 U18110 ( .B1(n15971), .B2(n15970), .A(n15969), .ZN(n15976) );
  XOR2_X1 U18111 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_173), .Z(n15975) );
  XNOR2_X1 U18112 ( .A(n15972), .B(keyinput_172), .ZN(n15974) );
  XNOR2_X1 U18113 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_174), .ZN(n15973) );
  NAND4_X1 U18114 ( .A1(n15976), .A2(n15975), .A3(n15974), .A4(n15973), .ZN(
        n15982) );
  XOR2_X1 U18115 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_175), .Z(n15981) );
  XNOR2_X1 U18116 ( .A(n20802), .B(keyinput_176), .ZN(n15979) );
  XNOR2_X1 U18117 ( .A(n20794), .B(keyinput_178), .ZN(n15978) );
  XNOR2_X1 U18118 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_177), .ZN(
        n15977) );
  NAND3_X1 U18119 ( .A1(n15979), .A2(n15978), .A3(n15977), .ZN(n15980) );
  AOI21_X1 U18120 ( .B1(n15982), .B2(n15981), .A(n15980), .ZN(n15990) );
  XNOR2_X1 U18121 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .ZN(n15989)
         );
  XNOR2_X1 U18122 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .ZN(n15988)
         );
  XOR2_X1 U18123 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_180), .Z(n15986)
         );
  XNOR2_X1 U18124 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .ZN(n15985)
         );
  XNOR2_X1 U18125 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_179), .ZN(
        n15984) );
  XNOR2_X1 U18126 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_182), .ZN(n15983)
         );
  NAND4_X1 U18127 ( .A1(n15986), .A2(n15985), .A3(n15984), .A4(n15983), .ZN(
        n15987) );
  NOR4_X1 U18128 ( .A1(n15990), .A2(n15989), .A3(n15988), .A4(n15987), .ZN(
        n15993) );
  XNOR2_X1 U18129 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .ZN(n15992)
         );
  XNOR2_X1 U18130 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .ZN(n15991)
         );
  NOR3_X1 U18131 ( .A1(n15993), .A2(n15992), .A3(n15991), .ZN(n16002) );
  XNOR2_X1 U18132 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .ZN(n16001)
         );
  XOR2_X1 U18133 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_192), .Z(n15996)
         );
  XNOR2_X1 U18134 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_190), .ZN(n15995)
         );
  XNOR2_X1 U18135 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_188), .ZN(n15994)
         );
  NAND3_X1 U18136 ( .A1(n15996), .A2(n15995), .A3(n15994), .ZN(n15999) );
  XOR2_X1 U18137 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_189), .Z(n15998)
         );
  XNOR2_X1 U18138 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .ZN(n15997)
         );
  NOR3_X1 U18139 ( .A1(n15999), .A2(n15998), .A3(n15997), .ZN(n16000) );
  OAI21_X1 U18140 ( .B1(n16002), .B2(n16001), .A(n16000), .ZN(n16005) );
  XNOR2_X1 U18141 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_193), .ZN(n16004)
         );
  XNOR2_X1 U18142 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_194), .ZN(n16003)
         );
  NAND3_X1 U18143 ( .A1(n16005), .A2(n16004), .A3(n16003), .ZN(n16009) );
  XOR2_X1 U18144 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_195), .Z(n16008)
         );
  XOR2_X1 U18145 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_197), .Z(n16007)
         );
  XNOR2_X1 U18146 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_196), .ZN(n16006)
         );
  AOI211_X1 U18147 ( .C1(n16009), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        n16018) );
  XNOR2_X1 U18148 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_198), .ZN(n16017)
         );
  OAI22_X1 U18149 ( .A1(n20731), .A2(keyinput_203), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_199), .ZN(n16010) );
  AOI221_X1 U18150 ( .B1(n20731), .B2(keyinput_203), .C1(keyinput_199), .C2(
        P1_REIP_REG_12__SCAN_IN), .A(n16010), .ZN(n16016) );
  INV_X1 U18151 ( .A(keyinput_201), .ZN(n16014) );
  XNOR2_X1 U18152 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_200), .ZN(n16013)
         );
  INV_X1 U18153 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20734) );
  INV_X1 U18154 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20735) );
  AOI22_X1 U18155 ( .A1(n20734), .A2(keyinput_202), .B1(n20735), .B2(
        keyinput_201), .ZN(n16011) );
  OAI21_X1 U18156 ( .B1(n20734), .B2(keyinput_202), .A(n16011), .ZN(n16012) );
  AOI211_X1 U18157 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n16014), .A(n16013), 
        .B(n16012), .ZN(n16015) );
  OAI211_X1 U18158 ( .C1(n16018), .C2(n16017), .A(n16016), .B(n16015), .ZN(
        n16022) );
  XNOR2_X1 U18159 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_205), .ZN(n16021)
         );
  XNOR2_X1 U18160 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_204), .ZN(n16020)
         );
  XNOR2_X1 U18161 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_206), .ZN(n16019)
         );
  NAND4_X1 U18162 ( .A1(n16022), .A2(n16021), .A3(n16020), .A4(n16019), .ZN(
        n16025) );
  XOR2_X1 U18163 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_207), .Z(n16024) );
  XOR2_X1 U18164 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_208), .Z(n16023) );
  AOI21_X1 U18165 ( .B1(n16025), .B2(n16024), .A(n16023), .ZN(n16028) );
  XNOR2_X1 U18166 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .ZN(n16027)
         );
  XNOR2_X1 U18167 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_210), .ZN(n16026)
         );
  OAI21_X1 U18168 ( .B1(n16028), .B2(n16027), .A(n16026), .ZN(n16031) );
  XOR2_X1 U18169 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_211), .Z(n16030) );
  XNOR2_X1 U18170 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .ZN(n16029)
         );
  NAND3_X1 U18171 ( .A1(n16031), .A2(n16030), .A3(n16029), .ZN(n16035) );
  XNOR2_X1 U18172 ( .A(n16032), .B(keyinput_214), .ZN(n16034) );
  XNOR2_X1 U18173 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n16033)
         );
  NAND3_X1 U18174 ( .A1(n16035), .A2(n16034), .A3(n16033), .ZN(n16040) );
  XNOR2_X1 U18175 ( .A(n16036), .B(keyinput_217), .ZN(n16039) );
  XNOR2_X1 U18176 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_215), .ZN(n16038)
         );
  XNOR2_X1 U18177 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_216), .ZN(n16037)
         );
  NAND4_X1 U18178 ( .A1(n16040), .A2(n16039), .A3(n16038), .A4(n16037), .ZN(
        n16044) );
  XNOR2_X1 U18179 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .ZN(n16043)
         );
  XNOR2_X1 U18180 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .ZN(n16042)
         );
  XNOR2_X1 U18181 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_220), .ZN(n16041)
         );
  AOI211_X1 U18182 ( .C1(n16044), .C2(n16043), .A(n16042), .B(n16041), .ZN(
        n16048) );
  XNOR2_X1 U18183 ( .A(n16045), .B(keyinput_221), .ZN(n16047) );
  XOR2_X1 U18184 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_222), .Z(n16046) );
  OAI21_X1 U18185 ( .B1(n16048), .B2(n16047), .A(n16046), .ZN(n16051) );
  XOR2_X1 U18186 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_224), .Z(n16050) );
  XNOR2_X1 U18187 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_223), .ZN(n16049)
         );
  NAND3_X1 U18188 ( .A1(n16051), .A2(n16050), .A3(n16049), .ZN(n16056) );
  XNOR2_X1 U18189 ( .A(n16052), .B(keyinput_225), .ZN(n16055) );
  XOR2_X1 U18190 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_226), .Z(n16054) );
  XNOR2_X1 U18191 ( .A(n16692), .B(keyinput_227), .ZN(n16053) );
  AOI211_X1 U18192 ( .C1(n16056), .C2(n16055), .A(n16054), .B(n16053), .ZN(
        n16062) );
  XOR2_X1 U18193 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_228), .Z(n16061) );
  XOR2_X1 U18194 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_230), .Z(n16059) );
  XNOR2_X1 U18195 ( .A(n22325), .B(keyinput_231), .ZN(n16058) );
  XNOR2_X1 U18196 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n16057)
         );
  NOR3_X1 U18197 ( .A1(n16059), .A2(n16058), .A3(n16057), .ZN(n16060) );
  OAI21_X1 U18198 ( .B1(n16062), .B2(n16061), .A(n16060), .ZN(n16066) );
  XNOR2_X1 U18199 ( .A(n16063), .B(keyinput_232), .ZN(n16065) );
  XNOR2_X1 U18200 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_233), .ZN(n16064)
         );
  AOI21_X1 U18201 ( .B1(n16066), .B2(n16065), .A(n16064), .ZN(n16069) );
  XNOR2_X1 U18202 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n16068)
         );
  XNOR2_X1 U18203 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .ZN(n16067)
         );
  OAI21_X1 U18204 ( .B1(n16069), .B2(n16068), .A(n16067), .ZN(n16073) );
  XNOR2_X1 U18205 ( .A(n22275), .B(keyinput_237), .ZN(n16072) );
  XOR2_X1 U18206 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .Z(n16071) );
  XNOR2_X1 U18207 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .ZN(n16070)
         );
  NAND4_X1 U18208 ( .A1(n16073), .A2(n16072), .A3(n16071), .A4(n16070), .ZN(
        n16078) );
  XNOR2_X1 U18209 ( .A(n16074), .B(keyinput_239), .ZN(n16077) );
  XNOR2_X1 U18210 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_241), .ZN(n16076)
         );
  XNOR2_X1 U18211 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .ZN(n16075)
         );
  AOI211_X1 U18212 ( .C1(n16078), .C2(n16077), .A(n16076), .B(n16075), .ZN(
        n16081) );
  XNOR2_X1 U18213 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .ZN(n16080)
         );
  XNOR2_X1 U18214 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .ZN(n16079)
         );
  OAI21_X1 U18215 ( .B1(n16081), .B2(n16080), .A(n16079), .ZN(n16084) );
  XOR2_X1 U18216 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .Z(n16083) );
  XOR2_X1 U18217 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .Z(n16082) );
  AOI21_X1 U18218 ( .B1(n16084), .B2(n16083), .A(n16082), .ZN(n16087) );
  XNOR2_X1 U18219 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .ZN(n16086)
         );
  XNOR2_X1 U18220 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n16085)
         );
  OAI21_X1 U18221 ( .B1(n16087), .B2(n16086), .A(n16085), .ZN(n16094) );
  OAI22_X1 U18222 ( .A1(n16089), .A2(keyinput_251), .B1(P1_EAX_REG_26__SCAN_IN), .B2(keyinput_249), .ZN(n16088) );
  AOI221_X1 U18223 ( .B1(n16089), .B2(keyinput_251), .C1(keyinput_249), .C2(
        P1_EAX_REG_26__SCAN_IN), .A(n16088), .ZN(n16093) );
  XOR2_X1 U18224 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_252), .Z(n16092) );
  OAI22_X1 U18225 ( .A1(n16721), .A2(keyinput_250), .B1(keyinput_248), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n16090) );
  AOI221_X1 U18226 ( .B1(n16721), .B2(keyinput_250), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput_248), .A(n16090), .ZN(n16091) );
  NAND4_X1 U18227 ( .A1(n16094), .A2(n16093), .A3(n16092), .A4(n16091), .ZN(
        n16097) );
  XNOR2_X1 U18228 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .ZN(n16096)
         );
  XOR2_X1 U18229 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .Z(n16095) );
  AOI21_X1 U18230 ( .B1(n16097), .B2(n16096), .A(n16095), .ZN(n16099) );
  XOR2_X1 U18231 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .Z(n16098) );
  AOI211_X1 U18232 ( .C1(n16101), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        n16251) );
  NAND2_X1 U18233 ( .A1(n20937), .A2(n16105), .ZN(n21618) );
  NAND2_X1 U18234 ( .A1(n21619), .A2(n21618), .ZN(n16242) );
  AOI21_X2 U18235 ( .B1(n16102), .B2(n16242), .A(n21642), .ZN(n21888) );
  NAND2_X1 U18236 ( .A1(n16104), .A2(n16103), .ZN(n20939) );
  NOR2_X4 U18237 ( .A1(n21911), .A2(n20937), .ZN(n22117) );
  OAI21_X1 U18238 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19617), .A(
        n16107), .ZN(n16121) );
  NAND2_X1 U18239 ( .A1(n16109), .A2(n16108), .ZN(n16111) );
  OAI211_X1 U18240 ( .C1(n21607), .C2(n19733), .A(n16113), .B(n16112), .ZN(
        n16118) );
  AOI221_X1 U18241 ( .B1(n16115), .B2(n19905), .C1(n16115), .C2(n21607), .A(
        n16114), .ZN(n16116) );
  INV_X1 U18242 ( .A(n16116), .ZN(n16117) );
  AOI221_X1 U18243 ( .B1(n16120), .B2(n16119), .C1(n16118), .C2(n16119), .A(
        n16117), .ZN(n18088) );
  OAI21_X1 U18244 ( .B1(n16122), .B2(n16121), .A(n22063), .ZN(n22118) );
  NOR2_X1 U18245 ( .A1(n19855), .A2(n22118), .ZN(n16124) );
  INV_X1 U18246 ( .A(n22116), .ZN(n22061) );
  OAI211_X1 U18247 ( .C1(n16124), .C2(n22061), .A(n16123), .B(n19813), .ZN(
        n16125) );
  OAI211_X1 U18248 ( .C1(n19733), .C2(n22116), .A(n18088), .B(n16125), .ZN(
        n16126) );
  INV_X1 U18249 ( .A(n16126), .ZN(n16132) );
  INV_X1 U18250 ( .A(n16127), .ZN(n16130) );
  XNOR2_X1 U18251 ( .A(n20937), .B(n19813), .ZN(n16128) );
  OAI21_X1 U18252 ( .B1(n16128), .B2(n20936), .A(n20941), .ZN(n22060) );
  OR3_X1 U18253 ( .A1(n16130), .A2(n16129), .A3(n22060), .ZN(n16131) );
  NAND2_X1 U18254 ( .A1(n16132), .A2(n16131), .ZN(n16133) );
  INV_X1 U18255 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16207) );
  AOI22_X1 U18256 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16138) );
  AOI22_X1 U18257 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16137) );
  AOI22_X1 U18258 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16136) );
  AOI22_X1 U18259 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16135) );
  NAND4_X1 U18260 ( .A1(n16138), .A2(n16137), .A3(n16136), .A4(n16135), .ZN(
        n16144) );
  AOI22_X1 U18261 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16142) );
  AOI22_X1 U18262 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16141) );
  AOI22_X1 U18263 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16140) );
  AOI22_X1 U18264 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16139) );
  NAND4_X1 U18265 ( .A1(n16142), .A2(n16141), .A3(n16140), .A4(n16139), .ZN(
        n16143) );
  AOI22_X1 U18266 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16148) );
  AOI22_X1 U18267 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U18268 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U18269 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16145) );
  NAND4_X1 U18270 ( .A1(n16148), .A2(n16147), .A3(n16146), .A4(n16145), .ZN(
        n16154) );
  AOI22_X1 U18271 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16152) );
  AOI22_X1 U18272 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18524), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16151) );
  AOI22_X1 U18273 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16150) );
  AOI22_X1 U18274 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18408), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16149) );
  NAND4_X1 U18275 ( .A1(n16152), .A2(n16151), .A3(n16150), .A4(n16149), .ZN(
        n16153) );
  AOI22_X1 U18276 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16165) );
  AOI22_X1 U18277 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16164) );
  INV_X1 U18278 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18535) );
  AOI22_X1 U18279 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16156) );
  OAI21_X1 U18280 ( .B1(n11234), .B2(n18535), .A(n16156), .ZN(n16162) );
  AOI22_X1 U18281 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16160) );
  AOI22_X1 U18282 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16159) );
  AOI22_X1 U18283 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U18284 ( .A1(n14107), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16157) );
  NAND4_X1 U18285 ( .A1(n16160), .A2(n16159), .A3(n16158), .A4(n16157), .ZN(
        n16161) );
  AOI211_X1 U18286 ( .C1(n18717), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n16162), .B(n16161), .ZN(n16163) );
  NAND3_X1 U18287 ( .A1(n16165), .A2(n16164), .A3(n16163), .ZN(n16228) );
  AOI22_X1 U18288 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14107), .ZN(n16169) );
  AOI22_X1 U18289 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U18290 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18673), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n18674), .ZN(n16167) );
  AOI22_X1 U18291 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21637), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16166) );
  NAND4_X1 U18292 ( .A1(n16169), .A2(n16168), .A3(n16167), .A4(n16166), .ZN(
        n16175) );
  AOI22_X1 U18293 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11165), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18548), .ZN(n16173) );
  AOI22_X1 U18294 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21034), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16172) );
  AOI22_X1 U18295 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16171) );
  AOI22_X1 U18296 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n16190), .ZN(n16170) );
  NAND4_X1 U18297 ( .A1(n16173), .A2(n16172), .A3(n16171), .A4(n16170), .ZN(
        n16174) );
  NOR2_X2 U18298 ( .A1(n16175), .A2(n16174), .ZN(n21598) );
  AOI22_X1 U18299 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16179) );
  AOI22_X1 U18300 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16178) );
  AOI22_X1 U18301 ( .A1(n21637), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16177) );
  AOI22_X1 U18302 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16176) );
  NAND4_X1 U18303 ( .A1(n16179), .A2(n16178), .A3(n16177), .A4(n16176), .ZN(
        n16185) );
  AOI22_X1 U18304 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U18305 ( .A1(n14107), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16182) );
  AOI22_X1 U18306 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U18307 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16180) );
  NAND4_X1 U18308 ( .A1(n16183), .A2(n16182), .A3(n16181), .A4(n16180), .ZN(
        n16184) );
  AOI22_X1 U18309 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16189) );
  AOI22_X1 U18310 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16188) );
  AOI22_X1 U18311 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16187) );
  AOI22_X1 U18312 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16186) );
  NAND4_X1 U18313 ( .A1(n16189), .A2(n16188), .A3(n16187), .A4(n16186), .ZN(
        n16196) );
  AOI22_X1 U18314 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14107), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16194) );
  AOI22_X1 U18315 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16190), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U18316 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16192) );
  AOI22_X1 U18317 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16191) );
  NAND4_X1 U18318 ( .A1(n16194), .A2(n16193), .A3(n16192), .A4(n16191), .ZN(
        n16195) );
  OAI21_X1 U18319 ( .B1(n21598), .B2(n21599), .A(n21482), .ZN(n16211) );
  AND2_X1 U18320 ( .A1(n16228), .A2(n16211), .ZN(n16219) );
  AOI22_X1 U18321 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16200) );
  AOI22_X1 U18322 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16199) );
  AOI22_X1 U18323 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16198) );
  AOI22_X1 U18324 ( .A1(n18673), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16197) );
  NAND4_X1 U18325 ( .A1(n16200), .A2(n16199), .A3(n16198), .A4(n16197), .ZN(
        n16206) );
  AOI22_X1 U18326 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16204) );
  AOI22_X1 U18327 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16203) );
  AOI22_X1 U18328 ( .A1(n14107), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16202) );
  AOI22_X1 U18329 ( .A1(n18397), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16201) );
  NAND4_X1 U18330 ( .A1(n16204), .A2(n16203), .A3(n16202), .A4(n16201), .ZN(
        n16205) );
  NAND2_X1 U18331 ( .A1(n16219), .A2(n16234), .ZN(n16208) );
  NOR2_X1 U18332 ( .A1(n21467), .A2(n16208), .ZN(n18736) );
  XOR2_X1 U18333 ( .A(n21932), .B(n18736), .Z(n18735) );
  XOR2_X1 U18334 ( .A(n16207), .B(n18735), .Z(n16222) );
  XOR2_X1 U18335 ( .A(n21467), .B(n16208), .Z(n16209) );
  NAND2_X1 U18336 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16209), .ZN(
        n16221) );
  XOR2_X1 U18337 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n16209), .Z(
        n19090) );
  XOR2_X1 U18338 ( .A(n16228), .B(n16211), .Z(n16210) );
  NAND2_X1 U18339 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16210), .ZN(
        n16217) );
  XOR2_X1 U18340 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n16210), .Z(
        n19116) );
  OAI21_X1 U18341 ( .B1(n21599), .B2(n16227), .A(n16211), .ZN(n16212) );
  NAND2_X1 U18342 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n16212), .ZN(
        n16216) );
  INV_X1 U18343 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21698) );
  XNOR2_X1 U18344 ( .A(n21698), .B(n16212), .ZN(n19127) );
  INV_X1 U18345 ( .A(n21599), .ZN(n19131) );
  INV_X1 U18346 ( .A(n21598), .ZN(n16215) );
  AOI21_X1 U18347 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16215), .A(
        n19131), .ZN(n16214) );
  INV_X1 U18348 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21767) );
  NOR2_X1 U18349 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16215), .ZN(
        n16213) );
  AOI221_X1 U18350 ( .B1(n19131), .B2(n16215), .C1(n16214), .C2(n21767), .A(
        n16213), .ZN(n19126) );
  NAND2_X1 U18351 ( .A1(n19127), .A2(n19126), .ZN(n19125) );
  NAND2_X1 U18352 ( .A1(n16216), .A2(n19125), .ZN(n19115) );
  NAND2_X1 U18353 ( .A1(n19116), .A2(n19115), .ZN(n19114) );
  NAND2_X1 U18354 ( .A1(n16217), .A2(n19114), .ZN(n16218) );
  NAND2_X1 U18355 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n16218), .ZN(
        n16220) );
  INV_X1 U18356 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21725) );
  XNOR2_X1 U18357 ( .A(n21725), .B(n16218), .ZN(n19105) );
  XOR2_X1 U18358 ( .A(n16234), .B(n16219), .Z(n19104) );
  NAND2_X1 U18359 ( .A1(n19105), .A2(n19104), .ZN(n19103) );
  NAND2_X1 U18360 ( .A1(n16220), .A2(n19103), .ZN(n19089) );
  NAND2_X1 U18361 ( .A1(n19090), .A2(n19089), .ZN(n19088) );
  NAND2_X1 U18362 ( .A1(n16221), .A2(n19088), .ZN(n18734) );
  XNOR2_X1 U18363 ( .A(n16222), .B(n18734), .ZN(n19075) );
  NAND2_X1 U18364 ( .A1(n22043), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19079) );
  OAI21_X1 U18365 ( .B1(n21950), .B2(n16207), .A(n19079), .ZN(n16249) );
  XOR2_X1 U18366 ( .A(n16234), .B(n16233), .Z(n16231) );
  NAND2_X1 U18367 ( .A1(n21598), .A2(n21482), .ZN(n16223) );
  OR2_X1 U18368 ( .A1(n21698), .A2(n16224), .ZN(n16226) );
  NAND2_X1 U18369 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21598), .ZN(
        n16225) );
  INV_X1 U18370 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21694) );
  XNOR2_X1 U18371 ( .A(n21694), .B(n21598), .ZN(n19134) );
  NAND2_X1 U18372 ( .A1(n16225), .A2(n19133), .ZN(n19122) );
  NAND2_X1 U18373 ( .A1(n19123), .A2(n19122), .ZN(n19121) );
  NAND2_X1 U18374 ( .A1(n16226), .A2(n19121), .ZN(n19111) );
  XNOR2_X1 U18375 ( .A(n16228), .B(n16227), .ZN(n16229) );
  XOR2_X1 U18376 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n16229), .Z(
        n19112) );
  NAND2_X1 U18377 ( .A1(n19111), .A2(n19112), .ZN(n19110) );
  NAND2_X1 U18378 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16229), .ZN(
        n16230) );
  NAND2_X1 U18379 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n16231), .ZN(
        n16232) );
  NAND2_X1 U18380 ( .A1(n16234), .A2(n16233), .ZN(n16239) );
  XOR2_X1 U18381 ( .A(n16239), .B(n21467), .Z(n16237) );
  INV_X1 U18382 ( .A(n16237), .ZN(n16235) );
  NAND2_X1 U18383 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19084), .ZN(
        n19083) );
  NAND2_X1 U18384 ( .A1(n16237), .A2(n16236), .ZN(n16238) );
  NAND2_X1 U18385 ( .A1(n19083), .A2(n16238), .ZN(n18730) );
  XOR2_X1 U18386 ( .A(n21934), .B(n21932), .Z(n18727) );
  XOR2_X1 U18387 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n18727), .Z(
        n18729) );
  XOR2_X1 U18388 ( .A(n18730), .B(n18729), .Z(n19071) );
  NOR2_X4 U18389 ( .A1(n19855), .A2(n21911), .ZN(n22119) );
  NAND2_X1 U18390 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21707) );
  NAND2_X1 U18391 ( .A1(n16241), .A2(n16240), .ZN(n21646) );
  NOR2_X1 U18392 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n22022), .ZN(
        n21685) );
  NOR2_X1 U18393 ( .A1(n21998), .A2(n21685), .ZN(n21699) );
  INV_X1 U18394 ( .A(n21699), .ZN(n21740) );
  AOI21_X1 U18395 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21708) );
  OAI22_X1 U18396 ( .A1(n21707), .A2(n21740), .B1(n16106), .B2(n21708), .ZN(
        n21710) );
  INV_X1 U18397 ( .A(n21710), .ZN(n21727) );
  NAND3_X1 U18398 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16243) );
  NOR2_X1 U18399 ( .A1(n21727), .A2(n16243), .ZN(n16245) );
  INV_X1 U18400 ( .A(n21888), .ZN(n21791) );
  NAND2_X1 U18401 ( .A1(n21791), .A2(n21767), .ZN(n21986) );
  INV_X1 U18402 ( .A(n21986), .ZN(n21871) );
  NOR2_X1 U18403 ( .A1(n16243), .A2(n21707), .ZN(n21739) );
  NOR2_X1 U18404 ( .A1(n21708), .A2(n16243), .ZN(n21738) );
  OAI22_X1 U18405 ( .A1(n21739), .A2(n21998), .B1(n21738), .B2(n16106), .ZN(
        n16244) );
  OR2_X1 U18406 ( .A1(n21871), .A2(n16244), .ZN(n21728) );
  MUX2_X1 U18407 ( .A(n16245), .B(n21728), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n16246) );
  AOI21_X1 U18408 ( .B1(n19071), .B2(n22119), .A(n16246), .ZN(n16247) );
  NOR2_X1 U18409 ( .A1(n16247), .A2(n22044), .ZN(n16248) );
  AOI211_X1 U18410 ( .C1(n21853), .C2(n19075), .A(n16249), .B(n16248), .ZN(
        n16250) );
  XNOR2_X1 U18411 ( .A(n16251), .B(n16250), .ZN(P3_U2856) );
  INV_X1 U18412 ( .A(n15668), .ZN(n16254) );
  INV_X1 U18413 ( .A(n16253), .ZN(n16368) );
  OAI211_X1 U18414 ( .C1(n16254), .C2(n11464), .A(n17419), .B(n16368), .ZN(
        n16261) );
  AND2_X1 U18415 ( .A1(n16257), .A2(n16256), .ZN(n16258) );
  OR2_X1 U18416 ( .A1(n16255), .A2(n16258), .ZN(n17937) );
  INV_X1 U18417 ( .A(n17937), .ZN(n16259) );
  NAND2_X1 U18418 ( .A1(n16259), .A2(n17411), .ZN(n16260) );
  OAI211_X1 U18419 ( .C1(n17411), .C2(n12234), .A(n16261), .B(n16260), .ZN(
        P2_U2874) );
  AND2_X1 U18420 ( .A1(n15673), .A2(n16262), .ZN(n16264) );
  OR2_X1 U18421 ( .A1(n16264), .A2(n16263), .ZN(n22307) );
  OR2_X1 U18422 ( .A1(n20819), .A2(n16265), .ZN(n16266) );
  AND2_X1 U18423 ( .A1(n16305), .A2(n16266), .ZN(n22302) );
  AOI22_X1 U18424 ( .A1(n22302), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n16267) );
  OAI21_X1 U18425 ( .B1(n22307), .B2(n20805), .A(n16267), .ZN(P1_U2864) );
  NAND2_X1 U18426 ( .A1(n16269), .A2(n16268), .ZN(n16270) );
  XOR2_X1 U18427 ( .A(n16271), .B(n16270), .Z(n18171) );
  INV_X1 U18428 ( .A(n18171), .ZN(n16281) );
  XNOR2_X1 U18429 ( .A(n16272), .B(n16325), .ZN(n18169) );
  OR2_X1 U18430 ( .A1(n16274), .A2(n18023), .ZN(n16323) );
  AOI21_X1 U18431 ( .B1(n16274), .B2(n17838), .A(n16273), .ZN(n16320) );
  NAND2_X1 U18432 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19360), .ZN(n16275) );
  OAI221_X1 U18433 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16323), .C1(
        n16325), .C2(n16320), .A(n16275), .ZN(n16279) );
  XNOR2_X1 U18434 ( .A(n16276), .B(n16277), .ZN(n20310) );
  OAI22_X1 U18435 ( .A1(n20310), .A2(n18066), .B1(n18061), .B2(n19275), .ZN(
        n16278) );
  AOI211_X1 U18436 ( .C1(n18169), .C2(n18055), .A(n16279), .B(n16278), .ZN(
        n16280) );
  OAI21_X1 U18437 ( .B1(n16281), .B2(n19495), .A(n16280), .ZN(P2_U3042) );
  OAI21_X1 U18438 ( .B1(n20603), .B2(n20602), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16282) );
  NAND2_X1 U18439 ( .A1(n16282), .A2(n20167), .ZN(n16293) );
  INV_X1 U18440 ( .A(n16293), .ZN(n16286) );
  INV_X1 U18441 ( .A(n20058), .ZN(n16283) );
  NAND3_X1 U18442 ( .A1(n16283), .A2(n20145), .A3(n20126), .ZN(n16292) );
  INV_X1 U18443 ( .A(n11926), .ZN(n16290) );
  INV_X1 U18444 ( .A(n20180), .ZN(n20196) );
  NAND2_X1 U18445 ( .A1(n20145), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20132) );
  INV_X1 U18446 ( .A(n20601), .ZN(n16287) );
  AOI21_X1 U18447 ( .B1(n16287), .B2(n20192), .A(n20525), .ZN(n16284) );
  AOI21_X1 U18448 ( .B1(n16290), .B2(n20196), .A(n16284), .ZN(n16285) );
  OAI22_X1 U18449 ( .A1(n20207), .A2(n20615), .B1(n16288), .B2(n16287), .ZN(
        n16289) );
  AOI21_X1 U18450 ( .B1(n20602), .B2(n20191), .A(n16289), .ZN(n16295) );
  OAI21_X1 U18451 ( .B1(n16290), .B2(n20601), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16291) );
  NAND2_X1 U18452 ( .A1(n20604), .A2(n15512), .ZN(n16294) );
  OAI211_X1 U18453 ( .C1(n20608), .C2(n16296), .A(n16295), .B(n16294), .ZN(
        P2_U3087) );
  INV_X1 U18454 ( .A(n16728), .ZN(n16298) );
  OAI222_X1 U18455 ( .A1(n22307), .A2(n16782), .B1(n16794), .B2(n16298), .C1(
        n16297), .C2(n16791), .ZN(P1_U2896) );
  NOR2_X1 U18456 ( .A1(n16263), .A2(n16300), .ZN(n16301) );
  OR2_X1 U18457 ( .A1(n16299), .A2(n16301), .ZN(n16381) );
  INV_X1 U18458 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22295) );
  INV_X1 U18459 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n22273) );
  NOR2_X1 U18460 ( .A1(n20726), .A2(n16302), .ZN(n22250) );
  NAND2_X1 U18461 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22250), .ZN(n22262) );
  NOR2_X1 U18462 ( .A1(n22273), .A2(n22262), .ZN(n22278) );
  NAND3_X1 U18463 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22333), .A3(n22278), 
        .ZN(n22290) );
  NOR2_X1 U18464 ( .A1(n22295), .A2(n22290), .ZN(n22301) );
  NAND2_X1 U18465 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22301), .ZN(n16356) );
  NAND2_X1 U18466 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22278), .ZN(n22280) );
  OR3_X1 U18467 ( .A1(n22295), .A2(n20731), .A3(n22280), .ZN(n16352) );
  AOI21_X1 U18468 ( .B1(n22333), .B2(n16352), .A(n22279), .ZN(n22311) );
  NAND2_X1 U18469 ( .A1(n16584), .A2(n16461), .ZN(n16666) );
  NAND2_X1 U18470 ( .A1(n16305), .A2(n16304), .ZN(n16306) );
  AND2_X1 U18471 ( .A1(n16303), .A2(n16306), .ZN(n22230) );
  INV_X1 U18472 ( .A(n22230), .ZN(n16308) );
  INV_X1 U18473 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n16307) );
  OAI22_X1 U18474 ( .A1(n16308), .A2(n22377), .B1(n22342), .B2(n16307), .ZN(
        n16309) );
  AOI211_X1 U18475 ( .C1(n22355), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n22353), .B(n16309), .ZN(n16310) );
  OAI221_X1 U18476 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n16356), .C1(n20734), 
        .C2(n22311), .A(n16310), .ZN(n16311) );
  AOI21_X1 U18477 ( .B1(n16382), .B2(n22357), .A(n16311), .ZN(n16312) );
  OAI21_X1 U18478 ( .B1(n16381), .B2(n22379), .A(n16312), .ZN(P1_U2831) );
  AOI22_X1 U18479 ( .A1(n22230), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n16313) );
  OAI21_X1 U18480 ( .B1(n16381), .B2(n20805), .A(n16313), .ZN(P1_U2863) );
  AND2_X1 U18481 ( .A1(n16315), .A2(n16314), .ZN(n16317) );
  XNOR2_X1 U18482 ( .A(n16317), .B(n16316), .ZN(n16338) );
  OR2_X1 U18483 ( .A1(n16318), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16330) );
  NAND3_X1 U18484 ( .A1(n16330), .A2(n18055), .A3(n16319), .ZN(n16329) );
  INV_X1 U18485 ( .A(n16320), .ZN(n16321) );
  AOI22_X1 U18486 ( .A1(n12603), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16321), .ZN(n16322) );
  OAI21_X1 U18487 ( .B1(n16331), .B2(n18061), .A(n16322), .ZN(n16327) );
  AOI221_X1 U18488 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16325), .C2(n16324), .A(
        n16323), .ZN(n16326) );
  AOI211_X1 U18489 ( .C1(n19500), .C2(n20254), .A(n16327), .B(n16326), .ZN(
        n16328) );
  OAI211_X1 U18490 ( .C1(n16338), .C2(n19495), .A(n16329), .B(n16328), .ZN(
        P2_U3041) );
  NAND3_X1 U18491 ( .A1(n16330), .A2(n18198), .A3(n16319), .ZN(n16337) );
  NOR2_X1 U18492 ( .A1(n18190), .A2(n16331), .ZN(n16334) );
  OAI22_X1 U18493 ( .A1(n16332), .A2(n18204), .B1(n18281), .B2(n14452), .ZN(
        n16333) );
  AOI211_X1 U18494 ( .C1(n18196), .C2(n16335), .A(n16334), .B(n16333), .ZN(
        n16336) );
  OAI211_X1 U18495 ( .C1(n16338), .C2(n18184), .A(n16337), .B(n16336), .ZN(
        P2_U3009) );
  INV_X1 U18496 ( .A(n16724), .ZN(n16340) );
  OAI222_X1 U18497 ( .A1(n16381), .A2(n16782), .B1(n16794), .B2(n16340), .C1(
        n16339), .C2(n16791), .ZN(P1_U2895) );
  OAI21_X1 U18498 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n22212) );
  INV_X1 U18499 ( .A(n22307), .ZN(n16346) );
  AOI22_X1 U18500 ( .A1(n20857), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n22241), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n16344) );
  OAI21_X1 U18501 ( .B1(n20856), .B2(n22306), .A(n16344), .ZN(n16345) );
  AOI21_X1 U18502 ( .B1(n16346), .B2(n20860), .A(n16345), .ZN(n16347) );
  OAI21_X1 U18503 ( .B1(n22212), .B2(n22386), .A(n16347), .ZN(P1_U2991) );
  OAI21_X1 U18504 ( .B1(n16299), .B2(n16349), .A(n16348), .ZN(n16971) );
  NAND2_X1 U18505 ( .A1(n16303), .A2(n16350), .ZN(n16351) );
  NAND2_X1 U18506 ( .A1(n16707), .A2(n16351), .ZN(n22244) );
  INV_X1 U18507 ( .A(n22244), .ZN(n16359) );
  NOR3_X1 U18508 ( .A1(n20735), .A2(n20734), .A3(n16352), .ZN(n22313) );
  OAI21_X1 U18509 ( .B1(n22373), .B2(n22313), .A(n16584), .ZN(n22330) );
  NAND2_X1 U18510 ( .A1(n22330), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16355) );
  OAI21_X1 U18511 ( .B1(n22370), .B2(n16965), .A(n16666), .ZN(n16353) );
  AOI21_X1 U18512 ( .B1(n22376), .B2(P1_EBX_REG_10__SCAN_IN), .A(n16353), .ZN(
        n16354) );
  OAI211_X1 U18513 ( .C1(n16964), .C2(n22384), .A(n16355), .B(n16354), .ZN(
        n16358) );
  NOR3_X1 U18514 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20734), .A3(n16356), 
        .ZN(n16357) );
  AOI211_X1 U18515 ( .C1(n16359), .C2(n22359), .A(n16358), .B(n16357), .ZN(
        n16360) );
  OAI21_X1 U18516 ( .B1(n16971), .B2(n22379), .A(n16360), .ZN(P1_U2830) );
  INV_X1 U18517 ( .A(n16718), .ZN(n16362) );
  OAI222_X1 U18518 ( .A1(n16971), .A2(n16782), .B1(n16794), .B2(n16362), .C1(
        n16361), .C2(n16791), .ZN(P1_U2894) );
  OAI222_X1 U18519 ( .A1(n22244), .A2(n20820), .B1(n16363), .B2(n20830), .C1(
        n20805), .C2(n16971), .ZN(P1_U2862) );
  OR2_X1 U18520 ( .A1(n16255), .A2(n16364), .ZN(n16365) );
  AND2_X1 U18521 ( .A1(n14534), .A2(n16365), .ZN(n19336) );
  INV_X1 U18522 ( .A(n19336), .ZN(n16366) );
  NOR2_X1 U18523 ( .A1(n16366), .A2(n17432), .ZN(n16371) );
  AOI211_X1 U18524 ( .C1(n16369), .C2(n16368), .A(n17452), .B(n16367), .ZN(
        n16370) );
  AOI211_X1 U18525 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n17432), .A(n16371), .B(
        n16370), .ZN(n16372) );
  INV_X1 U18526 ( .A(n16372), .ZN(P2_U2873) );
  INV_X1 U18527 ( .A(n17416), .ZN(n16373) );
  OAI211_X1 U18528 ( .C1(n16367), .C2(n16374), .A(n16373), .B(n17419), .ZN(
        n16377) );
  INV_X1 U18529 ( .A(n17911), .ZN(n16375) );
  NAND2_X1 U18530 ( .A1(n16375), .A2(n17411), .ZN(n16376) );
  OAI211_X1 U18531 ( .C1(n17411), .C2(n14530), .A(n16377), .B(n16376), .ZN(
        P2_U2872) );
  OAI21_X1 U18532 ( .B1(n16380), .B2(n16379), .A(n16378), .ZN(n22227) );
  INV_X1 U18533 ( .A(n16381), .ZN(n16386) );
  INV_X1 U18534 ( .A(n16382), .ZN(n16384) );
  NOR2_X1 U18535 ( .A1(n16939), .A2(n20734), .ZN(n22229) );
  AOI21_X1 U18536 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n22229), .ZN(n16383) );
  OAI21_X1 U18537 ( .B1(n20856), .B2(n16384), .A(n16383), .ZN(n16385) );
  AOI21_X1 U18538 ( .B1(n16386), .B2(n20860), .A(n16385), .ZN(n16387) );
  OAI21_X1 U18539 ( .B1(n22227), .B2(n22386), .A(n16387), .ZN(P1_U2990) );
  OAI21_X1 U18540 ( .B1(n17416), .B2(n16388), .A(n17427), .ZN(n16402) );
  NOR2_X1 U18541 ( .A1(n16389), .A2(n14537), .ZN(n16390) );
  OR2_X1 U18542 ( .A1(n16391), .A2(n16390), .ZN(n16392) );
  NAND2_X1 U18543 ( .A1(n17546), .A2(n16392), .ZN(n19347) );
  OAI22_X1 U18544 ( .A1(n20515), .A2(n19347), .B1(n16393), .B2(n20513), .ZN(
        n16395) );
  NOR2_X1 U18545 ( .A1(n20009), .A2(n20526), .ZN(n16394) );
  NOR2_X1 U18546 ( .A1(n16395), .A2(n16394), .ZN(n16397) );
  AOI22_X1 U18547 ( .A1(n20003), .A2(BUF2_REG_16__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n16396) );
  OAI211_X1 U18548 ( .C1(n16402), .C2(n20517), .A(n16397), .B(n16396), .ZN(
        P2_U2903) );
  NAND2_X1 U18549 ( .A1(n17432), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16401) );
  OR2_X1 U18550 ( .A1(n11382), .A2(n16398), .ZN(n17448) );
  NAND2_X1 U18551 ( .A1(n11382), .A2(n16398), .ZN(n16399) );
  NAND2_X1 U18552 ( .A1(n19346), .A2(n17411), .ZN(n16400) );
  OAI211_X1 U18553 ( .C1(n16402), .C2(n17452), .A(n16401), .B(n16400), .ZN(
        P2_U2871) );
  INV_X1 U18554 ( .A(n19455), .ZN(n17465) );
  NOR3_X1 U18555 ( .A1(n16404), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17557), .ZN(n16405) );
  NOR2_X1 U18556 ( .A1(n16409), .A2(n19508), .ZN(n16410) );
  XNOR2_X1 U18557 ( .A(n16413), .B(n16412), .ZN(n16435) );
  INV_X1 U18558 ( .A(n16435), .ZN(n16429) );
  INV_X1 U18559 ( .A(n20408), .ZN(n16414) );
  OAI22_X1 U18560 ( .A1(n16416), .A2(n16415), .B1(n16414), .B2(n18066), .ZN(
        n16428) );
  AOI21_X1 U18561 ( .B1(n16419), .B2(n16418), .A(n16417), .ZN(n16431) );
  NAND2_X1 U18562 ( .A1(n12603), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n16432) );
  INV_X1 U18563 ( .A(n16432), .ZN(n16423) );
  AOI21_X1 U18564 ( .B1(n16421), .B2(n16420), .A(n17877), .ZN(n16422) );
  AOI211_X1 U18565 ( .C1(n16431), .C2(n18055), .A(n16423), .B(n16422), .ZN(
        n16424) );
  OAI21_X1 U18566 ( .B1(n16426), .B2(n16425), .A(n16424), .ZN(n16427) );
  AOI211_X1 U18567 ( .C1(n14175), .C2(n16429), .A(n16428), .B(n16427), .ZN(
        n16430) );
  OAI21_X1 U18568 ( .B1(n16440), .B2(n18061), .A(n16430), .ZN(P2_U3044) );
  INV_X1 U18569 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16434) );
  NAND2_X1 U18570 ( .A1(n16431), .A2(n18198), .ZN(n16433) );
  OAI211_X1 U18571 ( .C1(n18204), .C2(n16434), .A(n16433), .B(n16432), .ZN(
        n16437) );
  NOR2_X1 U18572 ( .A1(n16435), .A2(n18184), .ZN(n16436) );
  AOI211_X1 U18573 ( .C1(n18196), .C2(n16438), .A(n16437), .B(n16436), .ZN(
        n16439) );
  OAI21_X1 U18574 ( .B1(n16440), .B2(n18190), .A(n16439), .ZN(P2_U3012) );
  NAND2_X1 U18575 ( .A1(n17432), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n16441) );
  OAI21_X1 U18576 ( .B1(n16442), .B2(n17432), .A(n16441), .ZN(P2_U2856) );
  NAND2_X1 U18577 ( .A1(n11196), .A2(n17411), .ZN(n16444) );
  NAND2_X1 U18578 ( .A1(n17432), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n16443) );
  OAI211_X1 U18579 ( .C1(n20262), .C2(n17452), .A(n16444), .B(n16443), .ZN(
        P2_U2884) );
  NAND2_X1 U18580 ( .A1(n11186), .A2(n16445), .ZN(n16446) );
  XNOR2_X1 U18581 ( .A(n17750), .B(n16446), .ZN(n16447) );
  NAND2_X1 U18582 ( .A1(n16447), .A2(n19481), .ZN(n16453) );
  AOI22_X1 U18583 ( .A1(n19471), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n19459), 
        .B2(n20358), .ZN(n16449) );
  AOI22_X1 U18584 ( .A1(n19470), .A2(P2_EBX_REG_3__SCAN_IN), .B1(n19472), .B2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16448) );
  OAI211_X1 U18585 ( .C1(n16450), .C2(n19441), .A(n16449), .B(n16448), .ZN(
        n16451) );
  AOI21_X1 U18586 ( .B1(n11196), .B2(n19461), .A(n16451), .ZN(n16452) );
  OAI211_X1 U18587 ( .C1(n19276), .C2(n20262), .A(n16453), .B(n16452), .ZN(
        P2_U2852) );
  INV_X1 U18588 ( .A(n16454), .ZN(n16455) );
  OAI211_X1 U18589 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11223), .A(n22482), 
        .B(n16455), .ZN(n16458) );
  INV_X1 U18590 ( .A(n18165), .ZN(n16456) );
  NAND2_X1 U18591 ( .A1(n16456), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n16457) );
  OAI211_X1 U18592 ( .C1(n16459), .C2(n11222), .A(n16458), .B(n16457), .ZN(
        P1_U3477) );
  INV_X1 U18593 ( .A(n16474), .ZN(n16460) );
  OAI21_X1 U18594 ( .B1(n16460), .B2(n22406), .A(P1_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n16464) );
  INV_X1 U18595 ( .A(n16461), .ZN(n16462) );
  NAND3_X1 U18596 ( .A1(n16464), .A2(n16463), .A3(n16462), .ZN(P1_U2801) );
  INV_X1 U18597 ( .A(n16465), .ZN(n16473) );
  OAI21_X1 U18598 ( .B1(n16467), .B2(n16473), .A(n16466), .ZN(n16470) );
  NAND2_X1 U18599 ( .A1(n16468), .A2(n16472), .ZN(n16469) );
  OAI211_X1 U18600 ( .C1(n14238), .C2(n16471), .A(n16470), .B(n16469), .ZN(
        n18147) );
  OAI22_X1 U18601 ( .A1(n16474), .A2(n16473), .B1(n13166), .B2(n16472), .ZN(
        n20866) );
  NOR2_X1 U18602 ( .A1(n16475), .A2(n13211), .ZN(n17200) );
  INV_X1 U18603 ( .A(n17200), .ZN(n16476) );
  AOI21_X1 U18604 ( .B1(n16476), .B2(n18155), .A(n22389), .ZN(n22131) );
  NOR2_X1 U18605 ( .A1(n20866), .A2(n22131), .ZN(n18140) );
  NOR2_X1 U18606 ( .A1(n18140), .A2(n22406), .ZN(n22388) );
  MUX2_X1 U18607 ( .A(P1_MORE_REG_SCAN_IN), .B(n18147), .S(n22388), .Z(
        P1_U3484) );
  INV_X1 U18608 ( .A(n16477), .ZN(n16486) );
  INV_X1 U18609 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20754) );
  INV_X1 U18610 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20744) );
  INV_X1 U18611 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20740) );
  AND2_X1 U18612 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22313), .ZN(n22332) );
  NAND2_X1 U18613 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n22332), .ZN(n16613) );
  NAND3_X1 U18614 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .ZN(n22352) );
  NOR4_X1 U18615 ( .A1(n20744), .A2(n20740), .A3(n16613), .A4(n22352), .ZN(
        n16478) );
  NAND3_X1 U18616 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(n16478), .ZN(n16596) );
  NOR2_X1 U18617 ( .A1(n20754), .A2(n16596), .ZN(n22371) );
  NAND2_X1 U18618 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22371), .ZN(n16571) );
  INV_X1 U18619 ( .A(n16571), .ZN(n16479) );
  AND3_X1 U18620 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(n16479), .ZN(n16546) );
  NAND2_X1 U18621 ( .A1(n22333), .A2(n16546), .ZN(n16559) );
  INV_X1 U18622 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20761) );
  NAND2_X1 U18623 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n16480) );
  NOR2_X1 U18624 ( .A1(n16549), .A2(n16480), .ZN(n16537) );
  NAND2_X1 U18625 ( .A1(n16523), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16509) );
  INV_X1 U18626 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20771) );
  NOR2_X1 U18627 ( .A1(n16509), .A2(n20771), .ZN(n16499) );
  NAND2_X1 U18628 ( .A1(n16499), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16483) );
  NAND3_X1 U18629 ( .A1(n16483), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n22339), 
        .ZN(n16482) );
  AOI22_X1 U18630 ( .A1(n22376), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n22355), .ZN(n16481) );
  OAI211_X1 U18631 ( .C1(n16483), .C2(P1_REIP_REG_31__SCAN_IN), .A(n16482), 
        .B(n16481), .ZN(n16484) );
  AOI21_X1 U18632 ( .B1(n16677), .B2(n22359), .A(n16484), .ZN(n16485) );
  OAI21_X1 U18633 ( .B1(n16486), .B2(n22379), .A(n16485), .ZN(P1_U2809) );
  XNOR2_X1 U18634 ( .A(n16489), .B(n16488), .ZN(n16979) );
  XNOR2_X1 U18635 ( .A(n16499), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n16492) );
  INV_X1 U18636 ( .A(n22339), .ZN(n16671) );
  AOI22_X1 U18637 ( .A1(n22376), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n22355), .ZN(n16491) );
  NAND2_X1 U18638 ( .A1(n22357), .A2(n16799), .ZN(n16490) );
  OAI211_X1 U18639 ( .C1(n16492), .C2(n16671), .A(n16491), .B(n16490), .ZN(
        n16493) );
  AOI21_X1 U18640 ( .B1(n16979), .B2(n22359), .A(n16493), .ZN(n16494) );
  OAI21_X1 U18641 ( .B1(n16681), .B2(n22379), .A(n16494), .ZN(P1_U2810) );
  AOI21_X1 U18642 ( .B1(n16496), .B2(n14210), .A(n16495), .ZN(n16810) );
  INV_X1 U18643 ( .A(n16810), .ZN(n16712) );
  AOI21_X1 U18644 ( .B1(n11243), .B2(n16498), .A(n16497), .ZN(n16986) );
  NAND2_X1 U18645 ( .A1(n22339), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16500) );
  AOI21_X1 U18646 ( .B1(n16509), .B2(n16500), .A(n16499), .ZN(n16503) );
  AOI22_X1 U18647 ( .A1(n22376), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22355), .ZN(n16501) );
  OAI21_X1 U18648 ( .B1(n22384), .B2(n16808), .A(n16501), .ZN(n16502) );
  AOI211_X1 U18649 ( .C1(n16986), .C2(n22359), .A(n16503), .B(n16502), .ZN(
        n16504) );
  OAI21_X1 U18650 ( .B1(n16712), .B2(n22379), .A(n16504), .ZN(P1_U2811) );
  OAI21_X1 U18651 ( .B1(n16522), .B2(n16505), .A(n11243), .ZN(n16990) );
  INV_X1 U18652 ( .A(n16506), .ZN(n16507) );
  NAND2_X1 U18653 ( .A1(n16507), .A2(n22360), .ZN(n16516) );
  INV_X1 U18654 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16683) );
  OAI22_X1 U18655 ( .A1(n22342), .A2(n16683), .B1(n16508), .B2(n22370), .ZN(
        n16513) );
  AOI21_X1 U18656 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n22339), .A(n16523), 
        .ZN(n16511) );
  INV_X1 U18657 ( .A(n16509), .ZN(n16510) );
  NOR2_X1 U18658 ( .A1(n16511), .A2(n16510), .ZN(n16512) );
  AOI211_X1 U18659 ( .C1(n22357), .C2(n16514), .A(n16513), .B(n16512), .ZN(
        n16515) );
  OAI211_X1 U18660 ( .C1(n22377), .C2(n16990), .A(n16516), .B(n16515), .ZN(
        P1_U2812) );
  AOI21_X1 U18661 ( .B1(n16519), .B2(n16518), .A(n14209), .ZN(n16817) );
  INV_X1 U18662 ( .A(n16817), .ZN(n16717) );
  AND2_X1 U18663 ( .A1(n16531), .A2(n16520), .ZN(n16521) );
  NOR2_X1 U18664 ( .A1(n16522), .A2(n16521), .ZN(n17008) );
  AOI21_X1 U18665 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n22339), .A(n16537), 
        .ZN(n16524) );
  NOR2_X1 U18666 ( .A1(n16524), .A2(n16523), .ZN(n16527) );
  AOI22_X1 U18667 ( .A1(n22376), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n22355), .ZN(n16525) );
  OAI21_X1 U18668 ( .B1(n22384), .B2(n16815), .A(n16525), .ZN(n16526) );
  AOI211_X1 U18669 ( .C1(n17008), .C2(n22359), .A(n16527), .B(n16526), .ZN(
        n16528) );
  OAI21_X1 U18670 ( .B1(n16717), .B2(n22379), .A(n16528), .ZN(P1_U2813) );
  OAI21_X1 U18671 ( .B1(n16529), .B2(n16530), .A(n16518), .ZN(n16823) );
  INV_X1 U18672 ( .A(n16531), .ZN(n16532) );
  AOI21_X1 U18673 ( .B1(n16533), .B2(n16541), .A(n16532), .ZN(n17019) );
  INV_X1 U18674 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20762) );
  NOR3_X1 U18675 ( .A1(n16559), .A2(n20762), .A3(n20761), .ZN(n16534) );
  AOI21_X1 U18676 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n22339), .A(n16534), 
        .ZN(n16538) );
  AOI22_X1 U18677 ( .A1(n22376), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n22355), .ZN(n16536) );
  NAND2_X1 U18678 ( .A1(n22357), .A2(n16824), .ZN(n16535) );
  OAI211_X1 U18679 ( .C1(n16538), .C2(n16537), .A(n16536), .B(n16535), .ZN(
        n16539) );
  AOI21_X1 U18680 ( .B1(n17019), .B2(n22359), .A(n16539), .ZN(n16540) );
  OAI21_X1 U18681 ( .B1(n16823), .B2(n22379), .A(n16540), .ZN(P1_U2814) );
  OAI21_X1 U18682 ( .B1(n16560), .B2(n16542), .A(n16541), .ZN(n17027) );
  AOI21_X1 U18683 ( .B1(n16545), .B2(n16544), .A(n16529), .ZN(n16837) );
  NAND2_X1 U18684 ( .A1(n16837), .A2(n22360), .ZN(n16554) );
  INV_X1 U18685 ( .A(n16546), .ZN(n16547) );
  OAI21_X1 U18686 ( .B1(n22279), .B2(n16547), .A(n22339), .ZN(n16573) );
  OAI21_X1 U18687 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n22373), .A(n16573), 
        .ZN(n16552) );
  AOI22_X1 U18688 ( .A1(n22376), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n22355), .ZN(n16548) );
  OAI21_X1 U18689 ( .B1(n22384), .B2(n16835), .A(n16548), .ZN(n16551) );
  NOR2_X1 U18690 ( .A1(n16549), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16550) );
  AOI211_X1 U18691 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n16552), .A(n16551), 
        .B(n16550), .ZN(n16553) );
  OAI211_X1 U18692 ( .C1(n22377), .C2(n17027), .A(n16554), .B(n16553), .ZN(
        P1_U2815) );
  OAI21_X1 U18693 ( .B1(n16555), .B2(n16556), .A(n16544), .ZN(n16843) );
  INV_X1 U18694 ( .A(n16573), .ZN(n16565) );
  AOI22_X1 U18695 ( .A1(n22376), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n22355), .ZN(n16558) );
  NAND2_X1 U18696 ( .A1(n22357), .A2(n16844), .ZN(n16557) );
  OAI211_X1 U18697 ( .C1(n16559), .C2(P1_REIP_REG_24__SCAN_IN), .A(n16558), 
        .B(n16557), .ZN(n16564) );
  INV_X1 U18698 ( .A(n16560), .ZN(n16561) );
  OAI21_X1 U18699 ( .B1(n16569), .B2(n16562), .A(n16561), .ZN(n17037) );
  NOR2_X1 U18700 ( .A1(n17037), .A2(n22377), .ZN(n16563) );
  AOI211_X1 U18701 ( .C1(n16565), .C2(P1_REIP_REG_24__SCAN_IN), .A(n16564), 
        .B(n16563), .ZN(n16566) );
  OAI21_X1 U18702 ( .B1(n16843), .B2(n22379), .A(n16566), .ZN(P1_U2816) );
  AOI21_X1 U18703 ( .B1(n16568), .B2(n16567), .A(n16555), .ZN(n16855) );
  INV_X1 U18704 ( .A(n16855), .ZN(n16734) );
  AOI21_X1 U18705 ( .B1(n16570), .B2(n16580), .A(n16569), .ZN(n17047) );
  NOR2_X1 U18706 ( .A1(n22373), .A2(n16571), .ZN(n16586) );
  AOI21_X1 U18707 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n16586), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n16572) );
  NOR2_X1 U18708 ( .A1(n16573), .A2(n16572), .ZN(n16576) );
  AOI22_X1 U18709 ( .A1(n22376), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n22355), .ZN(n16574) );
  OAI21_X1 U18710 ( .B1(n22384), .B2(n16853), .A(n16574), .ZN(n16575) );
  AOI211_X1 U18711 ( .C1(n17047), .C2(n22359), .A(n16576), .B(n16575), .ZN(
        n16577) );
  OAI21_X1 U18712 ( .B1(n16734), .B2(n22379), .A(n16577), .ZN(P1_U2817) );
  OAI21_X1 U18713 ( .B1(n16578), .B2(n16579), .A(n16567), .ZN(n16863) );
  INV_X1 U18714 ( .A(n16580), .ZN(n16581) );
  AOI21_X1 U18715 ( .B1(n16582), .B2(n17071), .A(n16581), .ZN(n17062) );
  INV_X1 U18716 ( .A(n16583), .ZN(n16865) );
  OAI21_X1 U18717 ( .B1(n22373), .B2(n22371), .A(n16584), .ZN(n16604) );
  INV_X1 U18718 ( .A(n16604), .ZN(n22368) );
  OAI21_X1 U18719 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n22373), .A(n22368), 
        .ZN(n16585) );
  MUX2_X1 U18720 ( .A(n16586), .B(n16585), .S(P1_REIP_REG_22__SCAN_IN), .Z(
        n16587) );
  AOI21_X1 U18721 ( .B1(n22355), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16587), .ZN(n16589) );
  NAND2_X1 U18722 ( .A1(n22376), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n16588) );
  OAI211_X1 U18723 ( .C1(n22384), .C2(n16865), .A(n16589), .B(n16588), .ZN(
        n16590) );
  AOI21_X1 U18724 ( .B1(n17062), .B2(n22359), .A(n16590), .ZN(n16591) );
  OAI21_X1 U18725 ( .B1(n16863), .B2(n22379), .A(n16591), .ZN(P1_U2818) );
  INV_X1 U18726 ( .A(n16594), .ZN(n16741) );
  AOI21_X1 U18727 ( .B1(n16595), .B2(n16592), .A(n16594), .ZN(n16882) );
  INV_X1 U18728 ( .A(n16882), .ZN(n16749) );
  OAI21_X1 U18729 ( .B1(n22373), .B2(n16596), .A(n20754), .ZN(n16603) );
  INV_X1 U18730 ( .A(n16881), .ZN(n16598) );
  AOI22_X1 U18731 ( .A1(n22376), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n22355), .ZN(n16597) );
  OAI21_X1 U18732 ( .B1(n22384), .B2(n16598), .A(n16597), .ZN(n16602) );
  OAI21_X1 U18733 ( .B1(n17100), .B2(n16600), .A(n16599), .ZN(n17076) );
  NOR2_X1 U18734 ( .A1(n17076), .A2(n22377), .ZN(n16601) );
  AOI211_X1 U18735 ( .C1(n16604), .C2(n16603), .A(n16602), .B(n16601), .ZN(
        n16605) );
  OAI21_X1 U18736 ( .B1(n16749), .B2(n22379), .A(n16605), .ZN(P1_U2820) );
  OR2_X1 U18737 ( .A1(n11180), .A2(n16607), .ZN(n16623) );
  AND2_X1 U18738 ( .A1(n16606), .A2(n16608), .ZN(n16751) );
  AOI21_X1 U18739 ( .B1(n16609), .B2(n16623), .A(n16751), .ZN(n16891) );
  INV_X1 U18740 ( .A(n16891), .ZN(n16760) );
  INV_X1 U18741 ( .A(n17098), .ZN(n16611) );
  AOI21_X1 U18742 ( .B1(n16612), .B2(n16610), .A(n16611), .ZN(n17104) );
  INV_X1 U18743 ( .A(n16893), .ZN(n16620) );
  INV_X1 U18744 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20747) );
  INV_X1 U18745 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20742) );
  NOR2_X1 U18746 ( .A1(n22373), .A2(n16613), .ZN(n16674) );
  NAND2_X1 U18747 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16674), .ZN(n16672) );
  NOR2_X1 U18748 ( .A1(n20742), .A2(n16672), .ZN(n22338) );
  NAND2_X1 U18749 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22338), .ZN(n22351) );
  INV_X1 U18750 ( .A(n22351), .ZN(n22350) );
  NAND2_X1 U18751 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22350), .ZN(n16643) );
  NOR2_X1 U18752 ( .A1(n20747), .A2(n16643), .ZN(n16614) );
  NOR2_X1 U18753 ( .A1(n16671), .A2(n16614), .ZN(n22363) );
  NAND2_X1 U18754 ( .A1(n22363), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16619) );
  INV_X1 U18755 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20750) );
  AND2_X1 U18756 ( .A1(n20750), .A2(n16614), .ZN(n22362) );
  INV_X1 U18757 ( .A(n22362), .ZN(n16615) );
  OAI211_X1 U18758 ( .C1(n22370), .C2(n16616), .A(n16615), .B(n16666), .ZN(
        n16617) );
  AOI21_X1 U18759 ( .B1(n22376), .B2(P1_EBX_REG_18__SCAN_IN), .A(n16617), .ZN(
        n16618) );
  OAI211_X1 U18760 ( .C1(n22384), .C2(n16620), .A(n16619), .B(n16618), .ZN(
        n16621) );
  AOI21_X1 U18761 ( .B1(n17104), .B2(n22359), .A(n16621), .ZN(n16622) );
  OAI21_X1 U18762 ( .B1(n16760), .B2(n22379), .A(n16622), .ZN(P1_U2822) );
  OR2_X1 U18763 ( .A1(n11180), .A2(n16634), .ZN(n16635) );
  INV_X1 U18764 ( .A(n16623), .ZN(n16624) );
  AOI21_X1 U18765 ( .B1(n16625), .B2(n16635), .A(n16624), .ZN(n20861) );
  INV_X1 U18766 ( .A(n20861), .ZN(n16769) );
  NAND2_X1 U18767 ( .A1(n20747), .A2(n16643), .ZN(n16629) );
  INV_X1 U18768 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20808) );
  AOI21_X1 U18769 ( .B1(n22355), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n22353), .ZN(n16627) );
  NAND2_X1 U18770 ( .A1(n22357), .A2(n20858), .ZN(n16626) );
  OAI211_X1 U18771 ( .C1(n22342), .C2(n20808), .A(n16627), .B(n16626), .ZN(
        n16628) );
  AOI21_X1 U18772 ( .B1(n22363), .B2(n16629), .A(n16628), .ZN(n16633) );
  INV_X1 U18773 ( .A(n16610), .ZN(n16630) );
  AOI21_X1 U18774 ( .B1(n16631), .B2(n11256), .A(n16630), .ZN(n20806) );
  NAND2_X1 U18775 ( .A1(n20806), .A2(n22359), .ZN(n16632) );
  OAI211_X1 U18776 ( .C1(n16769), .C2(n22379), .A(n16633), .B(n16632), .ZN(
        P1_U2823) );
  INV_X1 U18777 ( .A(n16634), .ZN(n16636) );
  INV_X1 U18778 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20746) );
  OAI21_X1 U18779 ( .B1(n16671), .B2(n20746), .A(n22351), .ZN(n16642) );
  OAI21_X1 U18780 ( .B1(n11495), .B2(n16637), .A(n11256), .ZN(n17147) );
  AOI21_X1 U18781 ( .B1(n22355), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n22353), .ZN(n16638) );
  OAI21_X1 U18782 ( .B1(n22342), .B2(n16692), .A(n16638), .ZN(n16639) );
  AOI21_X1 U18783 ( .B1(n16908), .B2(n22357), .A(n16639), .ZN(n16640) );
  OAI21_X1 U18784 ( .B1(n17147), .B2(n22377), .A(n16640), .ZN(n16641) );
  AOI21_X1 U18785 ( .B1(n16643), .B2(n16642), .A(n16641), .ZN(n16644) );
  OAI21_X1 U18786 ( .B1(n16911), .B2(n22379), .A(n16644), .ZN(P1_U2824) );
  NOR2_X1 U18787 ( .A1(n11229), .A2(n16646), .ZN(n16647) );
  OR2_X1 U18788 ( .A1(n16645), .A2(n16647), .ZN(n16931) );
  NAND2_X1 U18789 ( .A1(n16665), .A2(n16649), .ZN(n16650) );
  NAND2_X1 U18790 ( .A1(n17148), .A2(n16650), .ZN(n22146) );
  INV_X1 U18791 ( .A(n22146), .ZN(n16655) );
  OAI21_X1 U18792 ( .B1(n22370), .B2(n16926), .A(n16666), .ZN(n16651) );
  AOI21_X1 U18793 ( .B1(n22376), .B2(P1_EBX_REG_14__SCAN_IN), .A(n16651), .ZN(
        n16652) );
  OAI21_X1 U18794 ( .B1(n22384), .B2(n16925), .A(n16652), .ZN(n16654) );
  AOI211_X1 U18795 ( .C1(n20742), .C2(n16672), .A(n22338), .B(n16671), .ZN(
        n16653) );
  AOI211_X1 U18796 ( .C1(n16655), .C2(n22359), .A(n16654), .B(n16653), .ZN(
        n16656) );
  OAI21_X1 U18797 ( .B1(n16931), .B2(n22379), .A(n16656), .ZN(P1_U2826) );
  NAND2_X1 U18798 ( .A1(n16348), .A2(n16658), .ZN(n16659) );
  NAND2_X1 U18799 ( .A1(n16657), .A2(n16659), .ZN(n16703) );
  OR2_X1 U18800 ( .A1(n16703), .A2(n16704), .ZN(n16660) );
  NAND2_X1 U18801 ( .A1(n16660), .A2(n16657), .ZN(n16697) );
  NAND2_X1 U18802 ( .A1(n16697), .A2(n16696), .ZN(n16695) );
  INV_X1 U18803 ( .A(n16661), .ZN(n16662) );
  AOI21_X1 U18804 ( .B1(n16695), .B2(n16662), .A(n11229), .ZN(n16943) );
  INV_X1 U18805 ( .A(n16943), .ZN(n16786) );
  OR2_X1 U18806 ( .A1(n16699), .A2(n16663), .ZN(n16664) );
  AND2_X1 U18807 ( .A1(n16665), .A2(n16664), .ZN(n17170) );
  OAI21_X1 U18808 ( .B1(n22370), .B2(n16667), .A(n16666), .ZN(n16668) );
  AOI21_X1 U18809 ( .B1(n22376), .B2(P1_EBX_REG_13__SCAN_IN), .A(n16668), .ZN(
        n16669) );
  OAI21_X1 U18810 ( .B1(n22384), .B2(n16941), .A(n16669), .ZN(n16670) );
  AOI21_X1 U18811 ( .B1(n17170), .B2(n22359), .A(n16670), .ZN(n16676) );
  NOR2_X1 U18812 ( .A1(n16671), .A2(n20740), .ZN(n16673) );
  OAI21_X1 U18813 ( .B1(n16674), .B2(n16673), .A(n16672), .ZN(n16675) );
  OAI211_X1 U18814 ( .C1(n16786), .C2(n22379), .A(n16676), .B(n16675), .ZN(
        P1_U2827) );
  INV_X1 U18815 ( .A(n16677), .ZN(n16679) );
  OAI22_X1 U18816 ( .A1(n16679), .A2(n20820), .B1(n16678), .B2(n20830), .ZN(
        P1_U2841) );
  AOI22_X1 U18817 ( .A1(n16979), .A2(n20826), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n16708), .ZN(n16680) );
  OAI21_X1 U18818 ( .B1(n16681), .B2(n20805), .A(n16680), .ZN(P1_U2842) );
  AOI22_X1 U18819 ( .A1(n16986), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n16682) );
  OAI21_X1 U18820 ( .B1(n16712), .B2(n20805), .A(n16682), .ZN(P1_U2843) );
  OAI222_X1 U18821 ( .A1(n16683), .A2(n20830), .B1(n20820), .B2(n16990), .C1(
        n16506), .C2(n20805), .ZN(P1_U2844) );
  AOI22_X1 U18822 ( .A1(n17008), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n16684) );
  OAI21_X1 U18823 ( .B1(n16717), .B2(n20805), .A(n16684), .ZN(P1_U2845) );
  AOI22_X1 U18824 ( .A1(n17019), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n16685) );
  OAI21_X1 U18825 ( .B1(n16823), .B2(n20805), .A(n16685), .ZN(P1_U2846) );
  INV_X1 U18826 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16686) );
  INV_X1 U18827 ( .A(n16837), .ZN(n16727) );
  OAI222_X1 U18828 ( .A1(n16686), .A2(n20830), .B1(n20820), .B2(n17027), .C1(
        n16727), .C2(n20805), .ZN(P1_U2847) );
  OAI222_X1 U18829 ( .A1(n16687), .A2(n20830), .B1(n20820), .B2(n17037), .C1(
        n16843), .C2(n20805), .ZN(P1_U2848) );
  AOI22_X1 U18830 ( .A1(n17047), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n16688) );
  OAI21_X1 U18831 ( .B1(n16734), .B2(n20805), .A(n16688), .ZN(P1_U2849) );
  AOI22_X1 U18832 ( .A1(n17062), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n16689) );
  OAI21_X1 U18833 ( .B1(n16863), .B2(n20805), .A(n16689), .ZN(P1_U2850) );
  OAI222_X1 U18834 ( .A1(n16690), .A2(n20830), .B1(n20820), .B2(n17076), .C1(
        n16749), .C2(n20805), .ZN(P1_U2852) );
  AOI22_X1 U18835 ( .A1(n17104), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n16691) );
  OAI21_X1 U18836 ( .B1(n16760), .B2(n20805), .A(n16691), .ZN(P1_U2854) );
  OAI222_X1 U18837 ( .A1(n17147), .A2(n20820), .B1(n16692), .B2(n20830), .C1(
        n16911), .C2(n20805), .ZN(P1_U2856) );
  OAI222_X1 U18838 ( .A1(n22146), .A2(n20820), .B1(n16693), .B2(n20830), .C1(
        n20805), .C2(n16931), .ZN(P1_U2858) );
  AOI22_X1 U18839 ( .A1(n17170), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n16694) );
  OAI21_X1 U18840 ( .B1(n16786), .B2(n20805), .A(n16694), .ZN(P1_U2859) );
  OAI21_X1 U18841 ( .B1(n16697), .B2(n16696), .A(n16695), .ZN(n16949) );
  INV_X1 U18842 ( .A(n16698), .ZN(n16701) );
  INV_X1 U18843 ( .A(n16705), .ZN(n16700) );
  AOI21_X1 U18844 ( .B1(n16701), .B2(n16700), .A(n16699), .ZN(n22324) );
  AOI22_X1 U18845 ( .A1(n22324), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n16702) );
  OAI21_X1 U18846 ( .B1(n16949), .B2(n20805), .A(n16702), .ZN(P1_U2860) );
  XOR2_X1 U18847 ( .A(n16704), .B(n16703), .Z(n22320) );
  INV_X1 U18848 ( .A(n22320), .ZN(n16795) );
  AOI21_X1 U18849 ( .B1(n16707), .B2(n16706), .A(n16705), .ZN(n22314) );
  AOI22_X1 U18850 ( .A1(n22314), .A2(n20826), .B1(n16708), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16709) );
  OAI21_X1 U18851 ( .B1(n16795), .B2(n20805), .A(n16709), .ZN(P1_U2861) );
  AOI22_X1 U18852 ( .A1(n16771), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16770), .ZN(n16711) );
  AOI22_X1 U18853 ( .A1(n16774), .A2(BUF1_REG_29__SCAN_IN), .B1(n16773), .B2(
        n16783), .ZN(n16710) );
  OAI211_X1 U18854 ( .C1(n16712), .C2(n16782), .A(n16711), .B(n16710), .ZN(
        P1_U2875) );
  AOI22_X1 U18855 ( .A1(n16771), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16770), .ZN(n16714) );
  AOI22_X1 U18856 ( .A1(n16774), .A2(BUF1_REG_28__SCAN_IN), .B1(n16773), .B2(
        n16787), .ZN(n16713) );
  OAI211_X1 U18857 ( .C1(n16506), .C2(n16782), .A(n16714), .B(n16713), .ZN(
        P1_U2876) );
  AOI22_X1 U18858 ( .A1(n16771), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16770), .ZN(n16716) );
  AOI22_X1 U18859 ( .A1(n16774), .A2(BUF1_REG_27__SCAN_IN), .B1(n16773), .B2(
        n16790), .ZN(n16715) );
  OAI211_X1 U18860 ( .C1(n16717), .C2(n16782), .A(n16716), .B(n16715), .ZN(
        P1_U2877) );
  AOI22_X1 U18861 ( .A1(n16771), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16770), .ZN(n16720) );
  AOI22_X1 U18862 ( .A1(n16774), .A2(BUF1_REG_26__SCAN_IN), .B1(n16773), .B2(
        n16718), .ZN(n16719) );
  OAI211_X1 U18863 ( .C1(n16823), .C2(n16782), .A(n16720), .B(n16719), .ZN(
        P1_U2878) );
  OAI22_X1 U18864 ( .A1(n16763), .A2(n16722), .B1(n16721), .B2(n16791), .ZN(
        n16723) );
  INV_X1 U18865 ( .A(n16723), .ZN(n16726) );
  AOI22_X1 U18866 ( .A1(n16774), .A2(BUF1_REG_25__SCAN_IN), .B1(n16773), .B2(
        n16724), .ZN(n16725) );
  OAI211_X1 U18867 ( .C1(n16727), .C2(n16782), .A(n16726), .B(n16725), .ZN(
        P1_U2879) );
  AOI22_X1 U18868 ( .A1(n16771), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16770), .ZN(n16730) );
  AOI22_X1 U18869 ( .A1(n16774), .A2(BUF1_REG_24__SCAN_IN), .B1(n16773), .B2(
        n16728), .ZN(n16729) );
  OAI211_X1 U18870 ( .C1(n16843), .C2(n16782), .A(n16730), .B(n16729), .ZN(
        P1_U2880) );
  AOI22_X1 U18871 ( .A1(n16771), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16770), .ZN(n16733) );
  AOI22_X1 U18872 ( .A1(n16774), .A2(BUF1_REG_23__SCAN_IN), .B1(n16773), .B2(
        n16731), .ZN(n16732) );
  OAI211_X1 U18873 ( .C1(n16734), .C2(n16782), .A(n16733), .B(n16732), .ZN(
        P1_U2881) );
  OAI22_X1 U18874 ( .A1(n16763), .A2(n14975), .B1(n16735), .B2(n16791), .ZN(
        n16738) );
  INV_X1 U18875 ( .A(n16773), .ZN(n16765) );
  NOR2_X1 U18876 ( .A1(n16765), .A2(n16736), .ZN(n16737) );
  AOI211_X1 U18877 ( .C1(n16774), .C2(BUF1_REG_22__SCAN_IN), .A(n16738), .B(
        n16737), .ZN(n16739) );
  OAI21_X1 U18878 ( .B1(n16863), .B2(n16782), .A(n16739), .ZN(P1_U2882) );
  AND2_X1 U18879 ( .A1(n16741), .A2(n16740), .ZN(n16742) );
  OR2_X1 U18880 ( .A1(n16742), .A2(n16578), .ZN(n22380) );
  AOI22_X1 U18881 ( .A1(n16771), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16770), .ZN(n16745) );
  AOI22_X1 U18882 ( .A1(n16774), .A2(BUF1_REG_21__SCAN_IN), .B1(n16773), .B2(
        n16743), .ZN(n16744) );
  OAI211_X1 U18883 ( .C1(n22380), .C2(n16782), .A(n16745), .B(n16744), .ZN(
        P1_U2883) );
  AOI22_X1 U18884 ( .A1(n16771), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16770), .ZN(n16748) );
  AOI22_X1 U18885 ( .A1(n16774), .A2(BUF1_REG_20__SCAN_IN), .B1(n16773), .B2(
        n16746), .ZN(n16747) );
  OAI211_X1 U18886 ( .C1(n16749), .C2(n16782), .A(n16748), .B(n16747), .ZN(
        P1_U2884) );
  OR2_X1 U18887 ( .A1(n16751), .A2(n16750), .ZN(n16752) );
  AND2_X1 U18888 ( .A1(n16592), .A2(n16752), .ZN(n22361) );
  INV_X1 U18889 ( .A(n22361), .ZN(n16756) );
  AOI22_X1 U18890 ( .A1(n16771), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16770), .ZN(n16755) );
  AOI22_X1 U18891 ( .A1(n16774), .A2(BUF1_REG_19__SCAN_IN), .B1(n16773), .B2(
        n16753), .ZN(n16754) );
  OAI211_X1 U18892 ( .C1(n16756), .C2(n16782), .A(n16755), .B(n16754), .ZN(
        P1_U2885) );
  AOI22_X1 U18893 ( .A1(n16771), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16770), .ZN(n16759) );
  AOI22_X1 U18894 ( .A1(n16774), .A2(BUF1_REG_18__SCAN_IN), .B1(n16773), .B2(
        n16757), .ZN(n16758) );
  OAI211_X1 U18895 ( .C1(n16760), .C2(n16782), .A(n16759), .B(n16758), .ZN(
        P1_U2886) );
  OAI22_X1 U18896 ( .A1(n16763), .A2(n16762), .B1(n16761), .B2(n16791), .ZN(
        n16767) );
  NOR2_X1 U18897 ( .A1(n16765), .A2(n16764), .ZN(n16766) );
  AOI211_X1 U18898 ( .C1(n16774), .C2(BUF1_REG_17__SCAN_IN), .A(n16767), .B(
        n16766), .ZN(n16768) );
  OAI21_X1 U18899 ( .B1(n16769), .B2(n16782), .A(n16768), .ZN(P1_U2887) );
  AOI22_X1 U18900 ( .A1(n16771), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16770), .ZN(n16776) );
  AOI22_X1 U18901 ( .A1(n16774), .A2(BUF1_REG_16__SCAN_IN), .B1(n16773), .B2(
        n16772), .ZN(n16775) );
  OAI211_X1 U18902 ( .C1(n16911), .C2(n16782), .A(n16776), .B(n16775), .ZN(
        P1_U2888) );
  OAI21_X1 U18903 ( .B1(n16645), .B2(n16777), .A(n11180), .ZN(n20809) );
  OAI222_X1 U18904 ( .A1(n20809), .A2(n16782), .B1(n16794), .B2(n16778), .C1(
        n16791), .C2(n20719), .ZN(P1_U2889) );
  INV_X1 U18905 ( .A(n16779), .ZN(n16781) );
  OAI222_X1 U18906 ( .A1(n16931), .A2(n16782), .B1(n16794), .B2(n16781), .C1(
        n16780), .C2(n16791), .ZN(P1_U2890) );
  INV_X1 U18907 ( .A(n16783), .ZN(n16785) );
  OAI222_X1 U18908 ( .A1(n16786), .A2(n16782), .B1(n16794), .B2(n16785), .C1(
        n16784), .C2(n16791), .ZN(P1_U2891) );
  INV_X1 U18909 ( .A(n16787), .ZN(n16789) );
  OAI222_X1 U18910 ( .A1(n16949), .A2(n16782), .B1(n16794), .B2(n16789), .C1(
        n16788), .C2(n16791), .ZN(P1_U2892) );
  INV_X1 U18911 ( .A(n16790), .ZN(n16793) );
  OAI222_X1 U18912 ( .A1(n16782), .A2(n16795), .B1(n16794), .B2(n16793), .C1(
        n16792), .C2(n16791), .ZN(P1_U2893) );
  XNOR2_X1 U18913 ( .A(n16955), .B(n16797), .ZN(n16805) );
  XNOR2_X1 U18914 ( .A(n11249), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16981) );
  NAND2_X1 U18915 ( .A1(n16799), .A2(n20859), .ZN(n16800) );
  NAND2_X1 U18916 ( .A1(n22241), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16975) );
  OAI211_X1 U18917 ( .C1(n16966), .C2(n16801), .A(n16800), .B(n16975), .ZN(
        n16802) );
  AOI21_X1 U18918 ( .B1(n16803), .B2(n20860), .A(n16802), .ZN(n16804) );
  OAI21_X1 U18919 ( .B1(n16981), .B2(n22386), .A(n16804), .ZN(P1_U2969) );
  XNOR2_X1 U18920 ( .A(n16806), .B(n16805), .ZN(n16989) );
  NOR2_X1 U18921 ( .A1(n16939), .A2(n20771), .ZN(n16984) );
  AOI21_X1 U18922 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16984), .ZN(n16807) );
  OAI21_X1 U18923 ( .B1(n16808), .B2(n20856), .A(n16807), .ZN(n16809) );
  AOI21_X1 U18924 ( .B1(n16810), .B2(n20860), .A(n16809), .ZN(n16811) );
  OAI21_X1 U18925 ( .B1(n22386), .B2(n16989), .A(n16811), .ZN(P1_U2970) );
  XNOR2_X1 U18926 ( .A(n16956), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16813) );
  XNOR2_X1 U18927 ( .A(n16812), .B(n16813), .ZN(n17011) );
  INV_X1 U18928 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20767) );
  NOR2_X1 U18929 ( .A1(n16939), .A2(n20767), .ZN(n17005) );
  AOI21_X1 U18930 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17005), .ZN(n16814) );
  OAI21_X1 U18931 ( .B1(n20856), .B2(n16815), .A(n16814), .ZN(n16816) );
  AOI21_X1 U18932 ( .B1(n16817), .B2(n20860), .A(n16816), .ZN(n16818) );
  OAI21_X1 U18933 ( .B1(n17011), .B2(n22386), .A(n16818), .ZN(P1_U2972) );
  INV_X1 U18934 ( .A(n16819), .ZN(n16821) );
  NAND3_X1 U18935 ( .A1(n16821), .A2(n16831), .A3(n16820), .ZN(n16822) );
  XNOR2_X1 U18936 ( .A(n16822), .B(n17014), .ZN(n17022) );
  INV_X1 U18937 ( .A(n16823), .ZN(n16828) );
  INV_X1 U18938 ( .A(n16824), .ZN(n16826) );
  INV_X1 U18939 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20765) );
  NOR2_X1 U18940 ( .A1(n16939), .A2(n20765), .ZN(n17017) );
  AOI21_X1 U18941 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17017), .ZN(n16825) );
  OAI21_X1 U18942 ( .B1(n20856), .B2(n16826), .A(n16825), .ZN(n16827) );
  AOI21_X1 U18943 ( .B1(n16828), .B2(n20860), .A(n16827), .ZN(n16829) );
  OAI21_X1 U18944 ( .B1(n22386), .B2(n17022), .A(n16829), .ZN(P1_U2973) );
  INV_X1 U18945 ( .A(n16830), .ZN(n16832) );
  OAI211_X1 U18946 ( .C1(n16832), .C2(n17034), .A(n16850), .B(n16831), .ZN(
        n16833) );
  XOR2_X1 U18947 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n16833), .Z(
        n17031) );
  NOR2_X1 U18948 ( .A1(n16939), .A2(n20762), .ZN(n17025) );
  AOI21_X1 U18949 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17025), .ZN(n16834) );
  OAI21_X1 U18950 ( .B1(n20856), .B2(n16835), .A(n16834), .ZN(n16836) );
  AOI21_X1 U18951 ( .B1(n16837), .B2(n20860), .A(n16836), .ZN(n16838) );
  OAI21_X1 U18952 ( .B1(n22386), .B2(n17031), .A(n16838), .ZN(P1_U2974) );
  NAND3_X1 U18953 ( .A1(n13431), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n13412), .ZN(n16841) );
  INV_X1 U18954 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16839) );
  NAND3_X1 U18955 ( .A1(n16861), .A2(n16956), .A3(n16839), .ZN(n16840) );
  NAND2_X1 U18956 ( .A1(n16841), .A2(n16840), .ZN(n16842) );
  XNOR2_X1 U18957 ( .A(n16842), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17041) );
  INV_X1 U18958 ( .A(n16843), .ZN(n16848) );
  INV_X1 U18959 ( .A(n16844), .ZN(n16846) );
  NOR2_X1 U18960 ( .A1(n16939), .A2(n20761), .ZN(n17036) );
  AOI21_X1 U18961 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n17036), .ZN(n16845) );
  OAI21_X1 U18962 ( .B1(n20856), .B2(n16846), .A(n16845), .ZN(n16847) );
  AOI21_X1 U18963 ( .B1(n16848), .B2(n20860), .A(n16847), .ZN(n16849) );
  OAI21_X1 U18964 ( .B1(n17041), .B2(n22386), .A(n16849), .ZN(P1_U2975) );
  OAI21_X1 U18965 ( .B1(n16956), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16850), .ZN(n16851) );
  XNOR2_X1 U18966 ( .A(n16861), .B(n16851), .ZN(n17049) );
  INV_X1 U18967 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20759) );
  NOR2_X1 U18968 ( .A1(n16939), .A2(n20759), .ZN(n17042) );
  AOI21_X1 U18969 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17042), .ZN(n16852) );
  OAI21_X1 U18970 ( .B1(n20856), .B2(n16853), .A(n16852), .ZN(n16854) );
  AOI21_X1 U18971 ( .B1(n16855), .B2(n20860), .A(n16854), .ZN(n16856) );
  OAI21_X1 U18972 ( .B1(n17049), .B2(n22386), .A(n16856), .ZN(P1_U2976) );
  INV_X1 U18973 ( .A(n16857), .ZN(n16859) );
  NAND2_X1 U18974 ( .A1(n16859), .A2(n16858), .ZN(n16862) );
  AOI22_X1 U18975 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16862), .B1(
        n16861), .B2(n16860), .ZN(n17065) );
  INV_X1 U18976 ( .A(n16863), .ZN(n16867) );
  INV_X1 U18977 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20756) );
  NOR2_X1 U18978 ( .A1(n16939), .A2(n20756), .ZN(n17060) );
  AOI21_X1 U18979 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17060), .ZN(n16864) );
  OAI21_X1 U18980 ( .B1(n20856), .B2(n16865), .A(n16864), .ZN(n16866) );
  AOI21_X1 U18981 ( .B1(n16867), .B2(n20860), .A(n16866), .ZN(n16868) );
  OAI21_X1 U18982 ( .B1(n17065), .B2(n22386), .A(n16868), .ZN(P1_U2977) );
  XNOR2_X1 U18983 ( .A(n16955), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16892) );
  NAND2_X1 U18984 ( .A1(n16869), .A2(n16892), .ZN(n17105) );
  OAI21_X1 U18985 ( .B1(n16870), .B2(n16955), .A(n17105), .ZN(n16886) );
  AOI22_X1 U18986 ( .A1(n16886), .A2(n17095), .B1(n16955), .B2(n17105), .ZN(
        n16877) );
  NAND2_X1 U18987 ( .A1(n16956), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16871) );
  OAI211_X1 U18988 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n17095), .A(
        n16877), .B(n16871), .ZN(n16872) );
  XOR2_X1 U18989 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n16872), .Z(
        n17075) );
  INV_X1 U18990 ( .A(n22380), .ZN(n16875) );
  INV_X1 U18991 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n22369) );
  NOR2_X1 U18992 ( .A1(n16939), .A2(n22369), .ZN(n17067) );
  AOI21_X1 U18993 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17067), .ZN(n16873) );
  OAI21_X1 U18994 ( .B1(n20856), .B2(n22385), .A(n16873), .ZN(n16874) );
  AOI21_X1 U18995 ( .B1(n16875), .B2(n20860), .A(n16874), .ZN(n16876) );
  OAI21_X1 U18996 ( .B1(n17075), .B2(n22386), .A(n16876), .ZN(P1_U2978) );
  OAI21_X1 U18997 ( .B1(n13412), .B2(n17095), .A(n16877), .ZN(n16878) );
  XOR2_X1 U18998 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n16878), .Z(
        n17090) );
  NOR2_X1 U18999 ( .A1(n16939), .A2(n20754), .ZN(n17086) );
  NOR2_X1 U19000 ( .A1(n16966), .A2(n16879), .ZN(n16880) );
  AOI211_X1 U19001 ( .C1(n20859), .C2(n16881), .A(n17086), .B(n16880), .ZN(
        n16884) );
  NAND2_X1 U19002 ( .A1(n16882), .A2(n20860), .ZN(n16883) );
  OAI211_X1 U19003 ( .C1(n17090), .C2(n22386), .A(n16884), .B(n16883), .ZN(
        P1_U2979) );
  XNOR2_X1 U19004 ( .A(n16955), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16885) );
  XNOR2_X1 U19005 ( .A(n16886), .B(n16885), .ZN(n17103) );
  INV_X1 U19006 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20751) );
  NOR2_X1 U19007 ( .A1(n16939), .A2(n20751), .ZN(n17093) );
  AOI21_X1 U19008 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17093), .ZN(n16887) );
  OAI21_X1 U19009 ( .B1(n20856), .B2(n16888), .A(n16887), .ZN(n16889) );
  AOI21_X1 U19010 ( .B1(n22361), .B2(n20860), .A(n16889), .ZN(n16890) );
  OAI21_X1 U19011 ( .B1(n17103), .B2(n22386), .A(n16890), .ZN(P1_U2980) );
  NAND2_X1 U19012 ( .A1(n16891), .A2(n20860), .ZN(n16897) );
  NOR2_X1 U19013 ( .A1(n16939), .A2(n20750), .ZN(n17121) );
  AOI21_X1 U19014 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17121), .ZN(n16896) );
  OR2_X1 U19015 ( .A1(n16869), .A2(n16892), .ZN(n17106) );
  NAND3_X1 U19016 ( .A1(n17106), .A2(n17105), .A3(n20853), .ZN(n16895) );
  NAND2_X1 U19017 ( .A1(n20859), .A2(n16893), .ZN(n16894) );
  NAND4_X1 U19018 ( .A1(n16897), .A2(n16896), .A3(n16895), .A4(n16894), .ZN(
        P1_U2981) );
  INV_X1 U19019 ( .A(n16898), .ZN(n16919) );
  OAI211_X1 U19020 ( .C1(n16919), .C2(n17125), .A(n16899), .B(n16918), .ZN(
        n16914) );
  INV_X1 U19021 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17152) );
  NAND2_X1 U19022 ( .A1(n16955), .A2(n17152), .ZN(n16901) );
  NAND2_X1 U19023 ( .A1(n16900), .A2(n16901), .ZN(n16913) );
  NOR2_X1 U19024 ( .A1(n16914), .A2(n16913), .ZN(n16912) );
  INV_X1 U19025 ( .A(n16901), .ZN(n16902) );
  NOR2_X1 U19026 ( .A1(n16912), .A2(n16902), .ZN(n16905) );
  INV_X1 U19027 ( .A(n17130), .ZN(n16903) );
  AOI21_X1 U19028 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16955), .A(
        n16903), .ZN(n16904) );
  XNOR2_X1 U19029 ( .A(n16905), .B(n16904), .ZN(n17139) );
  NAND2_X1 U19030 ( .A1(n17139), .A2(n20853), .ZN(n16910) );
  NOR2_X1 U19031 ( .A1(n16939), .A2(n20746), .ZN(n17143) );
  NOR2_X1 U19032 ( .A1(n16966), .A2(n16906), .ZN(n16907) );
  AOI211_X1 U19033 ( .C1(n20859), .C2(n16908), .A(n17143), .B(n16907), .ZN(
        n16909) );
  OAI211_X1 U19034 ( .C1(n16972), .C2(n16911), .A(n16910), .B(n16909), .ZN(
        P1_U2983) );
  AOI21_X1 U19035 ( .B1(n16914), .B2(n16913), .A(n16912), .ZN(n17156) );
  OAI22_X1 U19036 ( .A1(n16966), .A2(n22340), .B1(n16939), .B2(n20744), .ZN(
        n16916) );
  NOR2_X1 U19037 ( .A1(n20809), .A2(n16972), .ZN(n16915) );
  AOI211_X1 U19038 ( .C1(n20859), .C2(n22344), .A(n16916), .B(n16915), .ZN(
        n16917) );
  OAI21_X1 U19039 ( .B1(n17156), .B2(n22386), .A(n16917), .ZN(P1_U2984) );
  NAND2_X1 U19040 ( .A1(n16919), .A2(n16918), .ZN(n17128) );
  INV_X1 U19041 ( .A(n16920), .ZN(n16921) );
  AOI21_X1 U19042 ( .B1(n17128), .B2(n16922), .A(n16921), .ZN(n16924) );
  XNOR2_X1 U19043 ( .A(n16955), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16923) );
  XNOR2_X1 U19044 ( .A(n16924), .B(n16923), .ZN(n22143) );
  NAND2_X1 U19045 ( .A1(n22143), .A2(n20853), .ZN(n16930) );
  INV_X1 U19046 ( .A(n16925), .ZN(n16928) );
  OAI22_X1 U19047 ( .A1(n16966), .A2(n16926), .B1(n16939), .B2(n20742), .ZN(
        n16927) );
  AOI21_X1 U19048 ( .B1(n16928), .B2(n20859), .A(n16927), .ZN(n16929) );
  OAI211_X1 U19049 ( .C1(n16972), .C2(n16931), .A(n16930), .B(n16929), .ZN(
        P1_U2985) );
  INV_X1 U19050 ( .A(n16932), .ZN(n16933) );
  AOI21_X1 U19051 ( .B1(n16898), .B2(n16934), .A(n16933), .ZN(n16947) );
  AND2_X1 U19052 ( .A1(n16935), .A2(n16936), .ZN(n16946) );
  NAND2_X1 U19053 ( .A1(n16947), .A2(n16946), .ZN(n16945) );
  NAND2_X1 U19054 ( .A1(n16945), .A2(n16936), .ZN(n16938) );
  XNOR2_X1 U19055 ( .A(n16938), .B(n16937), .ZN(n17172) );
  OR2_X1 U19056 ( .A1(n16939), .A2(n20740), .ZN(n17166) );
  NAND2_X1 U19057 ( .A1(n20857), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16940) );
  OAI211_X1 U19058 ( .C1(n20856), .C2(n16941), .A(n17166), .B(n16940), .ZN(
        n16942) );
  AOI21_X1 U19059 ( .B1(n16943), .B2(n20860), .A(n16942), .ZN(n16944) );
  OAI21_X1 U19060 ( .B1(n17172), .B2(n22386), .A(n16944), .ZN(P1_U2986) );
  OAI21_X1 U19061 ( .B1(n16947), .B2(n16946), .A(n16945), .ZN(n16948) );
  INV_X1 U19062 ( .A(n16948), .ZN(n17186) );
  INV_X1 U19063 ( .A(n16949), .ZN(n22328) );
  NAND2_X1 U19064 ( .A1(n20859), .A2(n22329), .ZN(n16951) );
  INV_X1 U19065 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n16950) );
  OR2_X1 U19066 ( .A1(n16939), .A2(n16950), .ZN(n17180) );
  OAI211_X1 U19067 ( .C1(n16966), .C2(n16952), .A(n16951), .B(n17180), .ZN(
        n16953) );
  AOI21_X1 U19068 ( .B1(n22328), .B2(n20860), .A(n16953), .ZN(n16954) );
  OAI21_X1 U19069 ( .B1(n17186), .B2(n22386), .A(n16954), .ZN(P1_U2987) );
  NOR2_X1 U19070 ( .A1(n16898), .A2(n16955), .ZN(n16957) );
  MUX2_X1 U19071 ( .A(n16378), .B(n16898), .S(n16956), .Z(n16963) );
  NOR2_X1 U19072 ( .A1(n16963), .A2(n22235), .ZN(n16962) );
  MUX2_X1 U19073 ( .A(n16957), .B(n13412), .S(n16962), .Z(n16958) );
  XNOR2_X1 U19074 ( .A(n16958), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17192) );
  NOR2_X1 U19075 ( .A1(n16939), .A2(n22317), .ZN(n17187) );
  AOI21_X1 U19076 ( .B1(n20857), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17187), .ZN(n16959) );
  OAI21_X1 U19077 ( .B1(n20856), .B2(n22323), .A(n16959), .ZN(n16960) );
  AOI21_X1 U19078 ( .B1(n22320), .B2(n20860), .A(n16960), .ZN(n16961) );
  OAI21_X1 U19079 ( .B1(n17192), .B2(n22386), .A(n16961), .ZN(P1_U2988) );
  AOI21_X1 U19080 ( .B1(n22235), .B2(n16963), .A(n16962), .ZN(n22240) );
  NAND2_X1 U19081 ( .A1(n22240), .A2(n20853), .ZN(n16970) );
  INV_X1 U19082 ( .A(n16964), .ZN(n16968) );
  OAI22_X1 U19083 ( .A1(n16966), .A2(n16965), .B1(n16939), .B2(n20735), .ZN(
        n16967) );
  AOI21_X1 U19084 ( .B1(n20859), .B2(n16968), .A(n16967), .ZN(n16969) );
  OAI211_X1 U19085 ( .C1(n16972), .C2(n16971), .A(n16970), .B(n16969), .ZN(
        P1_U2989) );
  NOR2_X1 U19086 ( .A1(n16974), .A2(n16973), .ZN(n16978) );
  OAI21_X1 U19087 ( .B1(n16976), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16975), .ZN(n16977) );
  AOI211_X1 U19088 ( .C1(n16979), .C2(n22231), .A(n16978), .B(n16977), .ZN(
        n16980) );
  OAI21_X1 U19089 ( .B1(n16981), .B2(n22226), .A(n16980), .ZN(P1_U3001) );
  NOR3_X1 U19090 ( .A1(n17001), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16982), .ZN(n16983) );
  AOI211_X1 U19091 ( .C1(n16985), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16984), .B(n16983), .ZN(n16988) );
  NAND2_X1 U19092 ( .A1(n16986), .A2(n22231), .ZN(n16987) );
  OAI211_X1 U19093 ( .C1(n16989), .C2(n22226), .A(n16988), .B(n16987), .ZN(
        P1_U3002) );
  NOR2_X1 U19094 ( .A1(n16990), .A2(n22245), .ZN(n16998) );
  INV_X1 U19095 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16991) );
  NOR3_X1 U19096 ( .A1(n17003), .A2(n17002), .A3(n16991), .ZN(n16997) );
  INV_X1 U19097 ( .A(n16992), .ZN(n16996) );
  NOR3_X1 U19098 ( .A1(n17001), .A2(n16994), .A3(n16993), .ZN(n16995) );
  NOR4_X1 U19099 ( .A1(n16998), .A2(n16997), .A3(n16996), .A4(n16995), .ZN(
        n16999) );
  OAI21_X1 U19100 ( .B1(n17000), .B2(n22226), .A(n16999), .ZN(P1_U3003) );
  INV_X1 U19101 ( .A(n17001), .ZN(n17007) );
  INV_X1 U19102 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17006) );
  NOR3_X1 U19103 ( .A1(n17003), .A2(n17002), .A3(n17006), .ZN(n17004) );
  AOI211_X1 U19104 ( .C1(n17007), .C2(n17006), .A(n17005), .B(n17004), .ZN(
        n17010) );
  NAND2_X1 U19105 ( .A1(n17008), .A2(n22231), .ZN(n17009) );
  OAI211_X1 U19106 ( .C1(n17011), .C2(n22226), .A(n17010), .B(n17009), .ZN(
        P1_U3004) );
  NOR2_X1 U19107 ( .A1(n17012), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17018) );
  INV_X1 U19108 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17013) );
  NAND3_X1 U19109 ( .A1(n17032), .A2(n17034), .A3(n17013), .ZN(n17023) );
  INV_X1 U19110 ( .A(n17026), .ZN(n17015) );
  AOI21_X1 U19111 ( .B1(n17023), .B2(n17015), .A(n17014), .ZN(n17016) );
  AOI211_X1 U19112 ( .C1(n17018), .C2(n17032), .A(n17017), .B(n17016), .ZN(
        n17021) );
  NAND2_X1 U19113 ( .A1(n17019), .A2(n22231), .ZN(n17020) );
  OAI211_X1 U19114 ( .C1(n17022), .C2(n22226), .A(n17021), .B(n17020), .ZN(
        P1_U3005) );
  INV_X1 U19115 ( .A(n17023), .ZN(n17024) );
  AOI211_X1 U19116 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n17026), .A(
        n17025), .B(n17024), .ZN(n17030) );
  INV_X1 U19117 ( .A(n17027), .ZN(n17028) );
  NAND2_X1 U19118 ( .A1(n17028), .A2(n22231), .ZN(n17029) );
  OAI211_X1 U19119 ( .C1(n17031), .C2(n22226), .A(n17030), .B(n17029), .ZN(
        P1_U3006) );
  INV_X1 U19120 ( .A(n17032), .ZN(n17045) );
  NOR3_X1 U19121 ( .A1(n17045), .A2(n17034), .A3(n17033), .ZN(n17035) );
  AOI211_X1 U19122 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n17043), .A(
        n17036), .B(n17035), .ZN(n17040) );
  INV_X1 U19123 ( .A(n17037), .ZN(n17038) );
  NAND2_X1 U19124 ( .A1(n17038), .A2(n22231), .ZN(n17039) );
  OAI211_X1 U19125 ( .C1(n17041), .C2(n22226), .A(n17040), .B(n17039), .ZN(
        P1_U3007) );
  AOI21_X1 U19126 ( .B1(n17043), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17042), .ZN(n17044) );
  OAI21_X1 U19127 ( .B1(n17045), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17044), .ZN(n17046) );
  AOI21_X1 U19128 ( .B1(n17047), .B2(n22231), .A(n17046), .ZN(n17048) );
  OAI21_X1 U19129 ( .B1(n17049), .B2(n22226), .A(n17048), .ZN(P1_U3008) );
  INV_X1 U19130 ( .A(n22160), .ZN(n22184) );
  NOR2_X1 U19131 ( .A1(n22184), .A2(n17173), .ZN(n17178) );
  NOR2_X1 U19132 ( .A1(n22151), .A2(n17050), .ZN(n17080) );
  NOR2_X1 U19133 ( .A1(n17178), .A2(n17080), .ZN(n22139) );
  NAND3_X1 U19134 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n17057), .ZN(n17053) );
  NOR3_X1 U19135 ( .A1(n22139), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17053), .ZN(n17066) );
  AOI21_X1 U19136 ( .B1(n17164), .B2(n17051), .A(n22221), .ZN(n17052) );
  OR2_X1 U19137 ( .A1(n17052), .A2(n22163), .ZN(n17077) );
  INV_X1 U19138 ( .A(n17077), .ZN(n17056) );
  INV_X1 U19139 ( .A(n17053), .ZN(n17055) );
  NOR2_X1 U19140 ( .A1(n17054), .A2(n22163), .ZN(n22199) );
  AOI21_X1 U19141 ( .B1(n17056), .B2(n17055), .A(n22199), .ZN(n17068) );
  OR2_X1 U19142 ( .A1(n17066), .A2(n17068), .ZN(n17061) );
  INV_X1 U19143 ( .A(n22139), .ZN(n17179) );
  NAND2_X1 U19144 ( .A1(n17179), .A2(n17057), .ZN(n17091) );
  NOR3_X1 U19145 ( .A1(n17091), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17058), .ZN(n17059) );
  AOI211_X1 U19146 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17061), .A(
        n17060), .B(n17059), .ZN(n17064) );
  NAND2_X1 U19147 ( .A1(n17062), .A2(n22231), .ZN(n17063) );
  OAI211_X1 U19148 ( .C1(n17065), .C2(n22226), .A(n17064), .B(n17063), .ZN(
        P1_U3009) );
  AOI211_X1 U19149 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n17068), .A(
        n17067), .B(n17066), .ZN(n17074) );
  NAND2_X1 U19150 ( .A1(n16599), .A2(n17069), .ZN(n17070) );
  NAND2_X1 U19151 ( .A1(n17071), .A2(n17070), .ZN(n22378) );
  INV_X1 U19152 ( .A(n22378), .ZN(n17072) );
  NAND2_X1 U19153 ( .A1(n17072), .A2(n22231), .ZN(n17073) );
  OAI211_X1 U19154 ( .C1(n17075), .C2(n22226), .A(n17074), .B(n17073), .ZN(
        P1_U3010) );
  NOR2_X1 U19155 ( .A1(n17076), .A2(n22245), .ZN(n17088) );
  NOR3_X1 U19156 ( .A1(n17091), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n17095), .ZN(n17087) );
  AOI21_X1 U19157 ( .B1(n22225), .B2(n17078), .A(n17077), .ZN(n17092) );
  INV_X1 U19158 ( .A(n22137), .ZN(n17079) );
  NAND2_X1 U19159 ( .A1(n17080), .A2(n17079), .ZN(n17083) );
  NAND3_X1 U19160 ( .A1(n17081), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n17164), .ZN(n17082) );
  NAND2_X1 U19161 ( .A1(n17083), .A2(n17082), .ZN(n17163) );
  OAI21_X1 U19162 ( .B1(n17163), .B2(n17165), .A(n17095), .ZN(n17084) );
  AOI21_X1 U19163 ( .B1(n17092), .B2(n17084), .A(n13428), .ZN(n17085) );
  NOR4_X1 U19164 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17089) );
  OAI21_X1 U19165 ( .B1(n17090), .B2(n22226), .A(n17089), .ZN(P1_U3011) );
  INV_X1 U19166 ( .A(n17091), .ZN(n17096) );
  NOR2_X1 U19167 ( .A1(n17092), .A2(n17095), .ZN(n17094) );
  AOI211_X1 U19168 ( .C1(n17096), .C2(n17095), .A(n17094), .B(n17093), .ZN(
        n17102) );
  AND2_X1 U19169 ( .A1(n17098), .A2(n17097), .ZN(n17099) );
  NOR2_X1 U19170 ( .A1(n17100), .A2(n17099), .ZN(n22358) );
  NAND2_X1 U19171 ( .A1(n22358), .A2(n22231), .ZN(n17101) );
  OAI211_X1 U19172 ( .C1(n17103), .C2(n22226), .A(n17102), .B(n17101), .ZN(
        P1_U3012) );
  INV_X1 U19173 ( .A(n17104), .ZN(n17124) );
  NAND3_X1 U19174 ( .A1(n17106), .A2(n17105), .A3(n22239), .ZN(n17123) );
  INV_X1 U19175 ( .A(n17119), .ZN(n17115) );
  INV_X1 U19176 ( .A(n22221), .ZN(n22166) );
  INV_X1 U19177 ( .A(n17109), .ZN(n17107) );
  NAND2_X1 U19178 ( .A1(n17164), .A2(n17107), .ZN(n17116) );
  NAND2_X1 U19179 ( .A1(n22166), .A2(n17116), .ZN(n17113) );
  INV_X1 U19180 ( .A(n17108), .ZN(n17159) );
  NOR2_X1 U19181 ( .A1(n17109), .A2(n17159), .ZN(n17117) );
  INV_X1 U19182 ( .A(n17117), .ZN(n17110) );
  NAND2_X1 U19183 ( .A1(n22225), .A2(n17110), .ZN(n17111) );
  AND2_X1 U19184 ( .A1(n22182), .A2(n17111), .ZN(n17112) );
  AND2_X1 U19185 ( .A1(n17113), .A2(n17112), .ZN(n17151) );
  OAI21_X1 U19186 ( .B1(n17115), .B2(n17114), .A(n17151), .ZN(n17136) );
  INV_X1 U19187 ( .A(n17116), .ZN(n17118) );
  AOI22_X1 U19188 ( .A1(n22160), .A2(n17118), .B1(n22225), .B2(n17117), .ZN(
        n17153) );
  NOR3_X1 U19189 ( .A1(n17153), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17119), .ZN(n17120) );
  AOI211_X1 U19190 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n17136), .A(
        n17121), .B(n17120), .ZN(n17122) );
  OAI211_X1 U19191 ( .C1(n22245), .C2(n17124), .A(n17123), .B(n17122), .ZN(
        P1_U3013) );
  NAND2_X1 U19192 ( .A1(n13412), .A2(n17140), .ZN(n17131) );
  INV_X1 U19193 ( .A(n17125), .ZN(n17127) );
  AOI21_X1 U19194 ( .B1(n17128), .B2(n17127), .A(n17126), .ZN(n17129) );
  MUX2_X1 U19195 ( .A(n17131), .B(n17130), .S(n17129), .Z(n17132) );
  XOR2_X1 U19196 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n17132), .Z(
        n20864) );
  INV_X1 U19197 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17133) );
  OAI21_X1 U19198 ( .B1(n17153), .B2(n17134), .A(n17133), .ZN(n17135) );
  AOI22_X1 U19199 ( .A1(n17136), .A2(n17135), .B1(n22241), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n17138) );
  NAND2_X1 U19200 ( .A1(n20806), .A2(n22231), .ZN(n17137) );
  OAI211_X1 U19201 ( .C1(n20864), .C2(n22226), .A(n17138), .B(n17137), .ZN(
        P1_U3014) );
  NAND2_X1 U19202 ( .A1(n17139), .A2(n22239), .ZN(n17146) );
  INV_X1 U19203 ( .A(n17151), .ZN(n17144) );
  AOI211_X1 U19204 ( .C1(n17141), .C2(n17152), .A(n17140), .B(n17153), .ZN(
        n17142) );
  AOI211_X1 U19205 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17144), .A(
        n17143), .B(n17142), .ZN(n17145) );
  OAI211_X1 U19206 ( .C1(n22245), .C2(n17147), .A(n17146), .B(n17145), .ZN(
        P1_U3015) );
  AOI21_X1 U19207 ( .B1(n17149), .B2(n17148), .A(n11495), .ZN(n22345) );
  NAND2_X1 U19208 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22241), .ZN(n17150) );
  OAI221_X1 U19209 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17153), 
        .C1(n17152), .C2(n17151), .A(n17150), .ZN(n17154) );
  AOI21_X1 U19210 ( .B1(n22345), .B2(n22231), .A(n17154), .ZN(n17155) );
  OAI21_X1 U19211 ( .B1(n17156), .B2(n22226), .A(n17155), .ZN(P1_U3016) );
  AOI21_X1 U19212 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17164), .A(
        n17157), .ZN(n17158) );
  AOI21_X1 U19213 ( .B1(n22225), .B2(n17159), .A(n17158), .ZN(n17160) );
  OAI211_X1 U19214 ( .C1(n17164), .C2(n17161), .A(n22182), .B(n17160), .ZN(
        n17162) );
  AOI21_X1 U19215 ( .B1(n22138), .B2(n17163), .A(n17162), .ZN(n22141) );
  NOR2_X1 U19216 ( .A1(n17163), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17168) );
  NAND3_X1 U19217 ( .A1(n17165), .A2(n17164), .A3(n22138), .ZN(n17167) );
  OAI211_X1 U19218 ( .C1(n22141), .C2(n17168), .A(n17167), .B(n17166), .ZN(
        n17169) );
  AOI21_X1 U19219 ( .B1(n17170), .B2(n22231), .A(n17169), .ZN(n17171) );
  OAI21_X1 U19220 ( .B1(n17172), .B2(n22226), .A(n17171), .ZN(P1_U3018) );
  INV_X1 U19221 ( .A(n17173), .ZN(n17176) );
  NAND2_X1 U19222 ( .A1(n22225), .A2(n17174), .ZN(n17175) );
  OAI211_X1 U19223 ( .C1(n22221), .C2(n17176), .A(n22182), .B(n17175), .ZN(
        n17188) );
  AOI21_X1 U19224 ( .B1(n17178), .B2(n17177), .A(n17188), .ZN(n17183) );
  NAND3_X1 U19225 ( .A1(n17179), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17182), .ZN(n17181) );
  OAI211_X1 U19226 ( .C1(n17183), .C2(n17182), .A(n17181), .B(n17180), .ZN(
        n17184) );
  AOI21_X1 U19227 ( .B1(n22231), .B2(n22324), .A(n17184), .ZN(n17185) );
  OAI21_X1 U19228 ( .B1(n17186), .B2(n22226), .A(n17185), .ZN(P1_U3019) );
  AOI21_X1 U19229 ( .B1(n17188), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17187), .ZN(n17189) );
  OAI21_X1 U19230 ( .B1(n22139), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17189), .ZN(n17190) );
  AOI21_X1 U19231 ( .B1(n22231), .B2(n22314), .A(n17190), .ZN(n17191) );
  OAI21_X1 U19232 ( .B1(n17192), .B2(n22226), .A(n17191), .ZN(P1_U3020) );
  INV_X1 U19233 ( .A(n17193), .ZN(n17194) );
  NOR2_X1 U19234 ( .A1(n17194), .A2(n22395), .ZN(n22404) );
  AOI21_X1 U19235 ( .B1(n11176), .B2(n17195), .A(n22404), .ZN(n17196) );
  OAI21_X1 U19236 ( .B1(n11212), .B2(n22534), .A(n17196), .ZN(n17197) );
  MUX2_X1 U19237 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17197), .S(
        n18165), .Z(P1_U3478) );
  XNOR2_X1 U19238 ( .A(n14713), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17214) );
  NAND2_X1 U19239 ( .A1(n17199), .A2(n17198), .ZN(n17225) );
  NAND2_X1 U19240 ( .A1(n17201), .A2(n17200), .ZN(n17216) );
  MUX2_X1 U19241 ( .A(n17225), .B(n17216), .S(n17214), .Z(n17206) );
  NAND2_X1 U19242 ( .A1(n17202), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17204) );
  MUX2_X1 U19243 ( .A(n17204), .B(n17203), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17205) );
  OAI211_X1 U19244 ( .C1(n17208), .C2(n17207), .A(n17206), .B(n17205), .ZN(
        n18125) );
  NAND2_X1 U19245 ( .A1(n18125), .A2(n20865), .ZN(n17213) );
  INV_X1 U19246 ( .A(n17209), .ZN(n17210) );
  NAND2_X1 U19247 ( .A1(n17211), .A2(n17210), .ZN(n17212) );
  OAI211_X1 U19248 ( .C1(n17230), .C2(n17214), .A(n17213), .B(n17212), .ZN(
        n17215) );
  MUX2_X1 U19249 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17215), .S(
        n17233), .Z(P1_U3472) );
  NAND2_X1 U19250 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17218) );
  NOR2_X1 U19251 ( .A1(n14713), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17217) );
  OAI22_X1 U19252 ( .A1(n18127), .A2(n17218), .B1(n17217), .B2(n17216), .ZN(
        n17220) );
  MUX2_X1 U19253 ( .A(n17220), .B(n17219), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n17227) );
  AOI21_X1 U19254 ( .B1(n14713), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13027), .ZN(n17221) );
  NOR2_X1 U19255 ( .A1(n13985), .A2(n17221), .ZN(n17231) );
  NAND2_X1 U19256 ( .A1(n18127), .A2(n14713), .ZN(n17223) );
  NAND2_X1 U19257 ( .A1(n17223), .A2(n17222), .ZN(n17224) );
  OAI21_X1 U19258 ( .B1(n17231), .B2(n17225), .A(n17224), .ZN(n17226) );
  AOI211_X1 U19259 ( .C1(n17229), .C2(n17228), .A(n17227), .B(n17226), .ZN(
        n18123) );
  INV_X1 U19260 ( .A(n20865), .ZN(n17232) );
  OAI22_X1 U19261 ( .A1(n18123), .A2(n17232), .B1(n17231), .B2(n17230), .ZN(
        n17234) );
  MUX2_X1 U19262 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17234), .S(
        n17233), .Z(P1_U3469) );
  INV_X1 U19263 ( .A(n17235), .ZN(n17241) );
  NAND2_X1 U19264 ( .A1(n17241), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n17240) );
  AOI22_X1 U19265 ( .A1(n17236), .A2(n17243), .B1(n17242), .B2(n22595), .ZN(
        n17239) );
  NAND2_X1 U19266 ( .A1(n22728), .A2(n22602), .ZN(n17238) );
  NAND2_X1 U19267 ( .A1(n17252), .A2(n22596), .ZN(n17237) );
  NAND4_X1 U19268 ( .A1(n17240), .A2(n17239), .A3(n17238), .A4(n17237), .ZN(
        P1_U3067) );
  NAND2_X1 U19269 ( .A1(n17241), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n17248) );
  AOI22_X1 U19270 ( .A1(n17244), .A2(n17243), .B1(n17242), .B2(n22617), .ZN(
        n17247) );
  NAND2_X1 U19271 ( .A1(n22728), .A2(n22624), .ZN(n17246) );
  NAND2_X1 U19272 ( .A1(n17252), .A2(n22618), .ZN(n17245) );
  NAND4_X1 U19273 ( .A1(n17248), .A2(n17247), .A3(n17246), .A4(n17245), .ZN(
        P1_U3068) );
  NAND2_X1 U19274 ( .A1(n17249), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n17256) );
  AOI22_X1 U19275 ( .A1(n17251), .A2(n22691), .B1(n22697), .B2(n17250), .ZN(
        n17255) );
  NAND2_X1 U19276 ( .A1(n17252), .A2(n22709), .ZN(n17254) );
  NAND2_X1 U19277 ( .A1(n22737), .A2(n22698), .ZN(n17253) );
  NAND4_X1 U19278 ( .A1(n17256), .A2(n17255), .A3(n17254), .A4(n17253), .ZN(
        P1_U3079) );
  NAND2_X1 U19279 ( .A1(n17257), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n17263) );
  AOI22_X1 U19280 ( .A1(n17259), .A2(n22691), .B1(n22697), .B2(n17258), .ZN(
        n17262) );
  INV_X1 U19281 ( .A(n22735), .ZN(n22614) );
  NAND2_X1 U19282 ( .A1(n22614), .A2(n22709), .ZN(n17261) );
  NAND2_X1 U19283 ( .A1(n22693), .A2(n22698), .ZN(n17260) );
  NAND4_X1 U19284 ( .A1(n17263), .A2(n17262), .A3(n17261), .A4(n17260), .ZN(
        P1_U3095) );
  INV_X1 U19285 ( .A(n17264), .ZN(n17277) );
  OAI211_X1 U19286 ( .C1(n17266), .C2(n17558), .A(n19481), .B(n17265), .ZN(
        n17276) );
  AOI21_X1 U19287 ( .B1(n17268), .B2(n11238), .A(n17267), .ZN(n17758) );
  INV_X1 U19288 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18305) );
  AOI22_X1 U19289 ( .A1(n19470), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19472), .ZN(n17269) );
  OAI21_X1 U19290 ( .B1(n18305), .B2(n19371), .A(n17269), .ZN(n17274) );
  AND2_X1 U19291 ( .A1(n17270), .A2(n17271), .ZN(n17272) );
  OR2_X1 U19292 ( .A1(n17272), .A2(n14201), .ZN(n17762) );
  NOR2_X1 U19293 ( .A1(n17762), .A2(n19477), .ZN(n17273) );
  AOI211_X1 U19294 ( .C1(n17758), .C2(n19459), .A(n17274), .B(n17273), .ZN(
        n17275) );
  OAI211_X1 U19295 ( .C1(n17277), .C2(n19441), .A(n17276), .B(n17275), .ZN(
        P2_U2828) );
  NOR2_X1 U19296 ( .A1(n17279), .A2(n17280), .ZN(n17281) );
  OR2_X1 U19297 ( .A1(n17278), .A2(n17281), .ZN(n17793) );
  NAND2_X1 U19298 ( .A1(n17282), .A2(n19473), .ZN(n17292) );
  XNOR2_X1 U19299 ( .A(n17283), .B(n17284), .ZN(n17798) );
  INV_X1 U19300 ( .A(n17798), .ZN(n17493) );
  OAI211_X1 U19301 ( .C1(n17593), .C2(n17286), .A(n19481), .B(n17285), .ZN(
        n17287) );
  OAI21_X1 U19302 ( .B1(n19443), .B2(n14473), .A(n17287), .ZN(n17288) );
  AOI21_X1 U19303 ( .B1(n19470), .B2(P2_EBX_REG_24__SCAN_IN), .A(n17288), .ZN(
        n17289) );
  OAI21_X1 U19304 ( .B1(n18302), .B2(n19371), .A(n17289), .ZN(n17290) );
  AOI21_X1 U19305 ( .B1(n17493), .B2(n19459), .A(n17290), .ZN(n17291) );
  OAI211_X1 U19306 ( .C1(n19477), .C2(n17793), .A(n17292), .B(n17291), .ZN(
        P2_U2831) );
  OAI211_X1 U19307 ( .C1(n17294), .C2(n17603), .A(n19481), .B(n17293), .ZN(
        n17306) );
  INV_X1 U19308 ( .A(n17279), .ZN(n17295) );
  OAI21_X1 U19309 ( .B1(n17406), .B2(n17296), .A(n17295), .ZN(n17811) );
  NOR2_X1 U19310 ( .A1(n17297), .A2(n17298), .ZN(n17299) );
  OR2_X1 U19311 ( .A1(n17283), .A2(n17299), .ZN(n17808) );
  INV_X1 U19312 ( .A(n17808), .ZN(n17499) );
  INV_X1 U19313 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18301) );
  NOR2_X1 U19314 ( .A1(n19371), .A2(n18301), .ZN(n17301) );
  OAI22_X1 U19315 ( .A1(n19409), .A2(n12275), .B1(n19443), .B2(n11336), .ZN(
        n17300) );
  AOI211_X1 U19316 ( .C1(n17499), .C2(n19459), .A(n17301), .B(n17300), .ZN(
        n17302) );
  OAI21_X1 U19317 ( .B1(n17811), .B2(n19477), .A(n17302), .ZN(n17303) );
  AOI21_X1 U19318 ( .B1(n17304), .B2(n19473), .A(n17303), .ZN(n17305) );
  NAND2_X1 U19319 ( .A1(n17306), .A2(n17305), .ZN(P2_U2832) );
  NAND2_X1 U19320 ( .A1(n11185), .A2(n17307), .ZN(n17308) );
  XOR2_X1 U19321 ( .A(n17634), .B(n17308), .Z(n17309) );
  NAND2_X1 U19322 ( .A1(n17309), .A2(n19481), .ZN(n17325) );
  INV_X1 U19323 ( .A(n17310), .ZN(n17323) );
  OR2_X1 U19324 ( .A1(n17311), .A2(n17312), .ZN(n17313) );
  NAND2_X1 U19325 ( .A1(n12658), .A2(n17313), .ZN(n17861) );
  INV_X1 U19326 ( .A(n17521), .ZN(n17316) );
  NAND2_X1 U19327 ( .A1(n17537), .A2(n17314), .ZN(n17315) );
  NAND2_X1 U19328 ( .A1(n17316), .A2(n17315), .ZN(n17857) );
  INV_X1 U19329 ( .A(n17857), .ZN(n17320) );
  NAND2_X1 U19330 ( .A1(n19470), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U19331 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19472), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19471), .ZN(n17317) );
  NAND3_X1 U19332 ( .A1(n17318), .A2(n17317), .A3(n14452), .ZN(n17319) );
  AOI21_X1 U19333 ( .B1(n17320), .B2(n19459), .A(n17319), .ZN(n17321) );
  OAI21_X1 U19334 ( .B1(n17861), .B2(n19477), .A(n17321), .ZN(n17322) );
  AOI21_X1 U19335 ( .B1(n17323), .B2(n19473), .A(n17322), .ZN(n17324) );
  NAND2_X1 U19336 ( .A1(n17325), .A2(n17324), .ZN(P2_U2836) );
  OAI21_X1 U19337 ( .B1(n17326), .B2(n17328), .A(n17327), .ZN(n17943) );
  INV_X1 U19338 ( .A(n17943), .ZN(n20017) );
  AOI22_X1 U19339 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19472), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19471), .ZN(n17329) );
  OAI211_X1 U19340 ( .C1(n17330), .C2(n17686), .A(n14452), .B(n17329), .ZN(
        n17332) );
  NOR2_X1 U19341 ( .A1(n19409), .A2(n12234), .ZN(n17331) );
  AOI211_X1 U19342 ( .C1(n19459), .C2(n20017), .A(n17332), .B(n17331), .ZN(
        n17333) );
  OAI21_X1 U19343 ( .B1(n17937), .B2(n19477), .A(n17333), .ZN(n17338) );
  OR2_X1 U19344 ( .A1(n11184), .A2(n17334), .ZN(n19335) );
  AOI211_X1 U19345 ( .C1(n17336), .C2(n17335), .A(n19518), .B(n19335), .ZN(
        n17337) );
  AOI211_X1 U19346 ( .C1(n19473), .C2(n17339), .A(n17338), .B(n17337), .ZN(
        n17340) );
  INV_X1 U19347 ( .A(n17340), .ZN(P2_U2842) );
  NOR2_X1 U19348 ( .A1(n11184), .A2(n17341), .ZN(n19326) );
  OAI211_X1 U19349 ( .C1(n17342), .C2(n17716), .A(n19481), .B(n19326), .ZN(
        n17351) );
  XNOR2_X1 U19350 ( .A(n17343), .B(n17991), .ZN(n20025) );
  INV_X1 U19351 ( .A(n20025), .ZN(n17968) );
  INV_X1 U19352 ( .A(n17716), .ZN(n17346) );
  AOI22_X1 U19353 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19472), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19471), .ZN(n17344) );
  INV_X1 U19354 ( .A(n17344), .ZN(n17345) );
  AOI211_X1 U19355 ( .C1(n17346), .C2(n17354), .A(n17345), .B(n12603), .ZN(
        n17347) );
  OAI21_X1 U19356 ( .B1(n19409), .B2(n12227), .A(n17347), .ZN(n17349) );
  NOR2_X1 U19357 ( .A1(n17971), .A2(n19477), .ZN(n17348) );
  AOI211_X1 U19358 ( .C1(n19459), .C2(n17968), .A(n17349), .B(n17348), .ZN(
        n17350) );
  OAI211_X1 U19359 ( .C1(n17352), .C2(n19441), .A(n17351), .B(n17350), .ZN(
        P2_U2844) );
  NAND2_X1 U19360 ( .A1(n17353), .A2(n19481), .ZN(n17362) );
  AOI22_X1 U19361 ( .A1(n19471), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n19459), 
        .B2(n20458), .ZN(n17357) );
  MUX2_X1 U19362 ( .A(n17354), .B(n19472), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n17355) );
  AOI21_X1 U19363 ( .B1(n19470), .B2(P2_EBX_REG_1__SCAN_IN), .A(n17355), .ZN(
        n17356) );
  OAI211_X1 U19364 ( .C1(n19441), .C2(n17358), .A(n17357), .B(n17356), .ZN(
        n17359) );
  AOI21_X1 U19365 ( .B1(n17360), .B2(n19461), .A(n17359), .ZN(n17361) );
  OAI211_X1 U19366 ( .C1(n18214), .C2(n19276), .A(n17362), .B(n17361), .ZN(
        P2_U2854) );
  AOI21_X1 U19367 ( .B1(n17365), .B2(n17364), .A(n17363), .ZN(n17453) );
  NAND2_X1 U19368 ( .A1(n17453), .A2(n17419), .ZN(n17367) );
  NAND2_X1 U19369 ( .A1(n17432), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n17366) );
  OAI211_X1 U19370 ( .C1(n19457), .C2(n17432), .A(n17367), .B(n17366), .ZN(
        P2_U2858) );
  INV_X1 U19371 ( .A(n17368), .ZN(n17375) );
  NOR2_X1 U19372 ( .A1(n17375), .A2(n17369), .ZN(n17371) );
  XNOR2_X1 U19373 ( .A(n17371), .B(n17370), .ZN(n17468) );
  NAND2_X1 U19374 ( .A1(n17432), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n17373) );
  NAND2_X1 U19375 ( .A1(n19445), .A2(n17411), .ZN(n17372) );
  OAI211_X1 U19376 ( .C1(n17468), .C2(n17452), .A(n17373), .B(n17372), .ZN(
        P2_U2859) );
  NOR2_X1 U19377 ( .A1(n17376), .A2(n17375), .ZN(n17378) );
  XNOR2_X1 U19378 ( .A(n17378), .B(n17377), .ZN(n17469) );
  NAND2_X1 U19379 ( .A1(n17469), .A2(n17419), .ZN(n17380) );
  NAND2_X1 U19380 ( .A1(n17432), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n17379) );
  OAI211_X1 U19381 ( .C1(n17432), .C2(n17762), .A(n17380), .B(n17379), .ZN(
        P2_U2860) );
  OAI21_X1 U19382 ( .B1(n17383), .B2(n17382), .A(n17381), .ZN(n17480) );
  NAND2_X1 U19383 ( .A1(n17432), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n17388) );
  NAND2_X1 U19384 ( .A1(n17384), .A2(n17385), .ZN(n17386) );
  AND2_X1 U19385 ( .A1(n17270), .A2(n17386), .ZN(n19433) );
  NAND2_X1 U19386 ( .A1(n19433), .A2(n17411), .ZN(n17387) );
  OAI211_X1 U19387 ( .C1(n17480), .C2(n17452), .A(n17388), .B(n17387), .ZN(
        P2_U2861) );
  OAI21_X1 U19388 ( .B1(n17391), .B2(n17390), .A(n17389), .ZN(n17490) );
  OAI21_X1 U19389 ( .B1(n17278), .B2(n17392), .A(n17384), .ZN(n17781) );
  NOR2_X1 U19390 ( .A1(n17781), .A2(n17432), .ZN(n17393) );
  AOI21_X1 U19391 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n17432), .A(n17393), .ZN(
        n17394) );
  OAI21_X1 U19392 ( .B1(n17490), .B2(n17452), .A(n17394), .ZN(P2_U2862) );
  OAI21_X1 U19393 ( .B1(n17397), .B2(n17396), .A(n17395), .ZN(n17496) );
  NOR2_X1 U19394 ( .A1(n17793), .A2(n17432), .ZN(n17398) );
  AOI21_X1 U19395 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n17432), .A(n17398), .ZN(
        n17399) );
  OAI21_X1 U19396 ( .B1(n17496), .B2(n17452), .A(n17399), .ZN(P2_U2863) );
  XNOR2_X1 U19397 ( .A(n17400), .B(n17401), .ZN(n17502) );
  NOR2_X1 U19398 ( .A1(n17811), .A2(n17432), .ZN(n17402) );
  AOI21_X1 U19399 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n17432), .A(n17402), .ZN(
        n17403) );
  OAI21_X1 U19400 ( .B1(n17502), .B2(n17452), .A(n17403), .ZN(P2_U2864) );
  AND2_X1 U19401 ( .A1(n17416), .A2(n17404), .ZN(n17417) );
  OAI21_X1 U19402 ( .B1(n17417), .B2(n17405), .A(n17400), .ZN(n17511) );
  INV_X1 U19403 ( .A(n17406), .ZN(n17410) );
  NAND2_X1 U19404 ( .A1(n17408), .A2(n17407), .ZN(n17409) );
  NAND2_X1 U19405 ( .A1(n17410), .A2(n17409), .ZN(n19412) );
  MUX2_X1 U19406 ( .A(n12271), .B(n19412), .S(n17411), .Z(n17412) );
  OAI21_X1 U19407 ( .B1(n17511), .B2(n17452), .A(n17412), .ZN(P2_U2865) );
  XNOR2_X1 U19408 ( .A(n17414), .B(n17413), .ZN(n19398) );
  NAND2_X1 U19409 ( .A1(n17416), .A2(n17415), .ZN(n17423) );
  AOI21_X1 U19410 ( .B1(n17418), .B2(n17423), .A(n17417), .ZN(n17518) );
  NAND2_X1 U19411 ( .A1(n17518), .A2(n17419), .ZN(n17421) );
  NAND2_X1 U19412 ( .A1(n17432), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n17420) );
  OAI211_X1 U19413 ( .C1(n19398), .C2(n17432), .A(n17421), .B(n17420), .ZN(
        P2_U2866) );
  INV_X1 U19414 ( .A(n17427), .ZN(n17446) );
  OAI21_X1 U19415 ( .B1(n17428), .B2(n17424), .A(n17423), .ZN(n17528) );
  NOR2_X1 U19416 ( .A1(n19384), .A2(n17432), .ZN(n17425) );
  AOI21_X1 U19417 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n17432), .A(n17425), .ZN(
        n17426) );
  OAI21_X1 U19418 ( .B1(n17528), .B2(n17452), .A(n17426), .ZN(P2_U2867) );
  AOI21_X1 U19419 ( .B1(n17429), .B2(n17435), .A(n17428), .ZN(n17430) );
  INV_X1 U19420 ( .A(n17430), .ZN(n17534) );
  NOR2_X1 U19421 ( .A1(n17861), .A2(n17432), .ZN(n17431) );
  AOI21_X1 U19422 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n17432), .A(n17431), .ZN(
        n17433) );
  OAI21_X1 U19423 ( .B1(n17534), .B2(n17452), .A(n17433), .ZN(P2_U2868) );
  INV_X1 U19424 ( .A(n17444), .ZN(n17437) );
  INV_X1 U19425 ( .A(n17434), .ZN(n17436) );
  OAI21_X1 U19426 ( .B1(n17437), .B2(n17436), .A(n17435), .ZN(n17544) );
  INV_X1 U19427 ( .A(n17311), .ZN(n17439) );
  OAI21_X1 U19428 ( .B1(n17438), .B2(n17440), .A(n17439), .ZN(n19377) );
  NOR2_X1 U19429 ( .A1(n19377), .A2(n17432), .ZN(n17441) );
  AOI21_X1 U19430 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n17432), .A(n17441), .ZN(
        n17442) );
  OAI21_X1 U19431 ( .B1(n17544), .B2(n17452), .A(n17442), .ZN(P2_U2869) );
  INV_X1 U19432 ( .A(n17443), .ZN(n17445) );
  OAI21_X1 U19433 ( .B1(n17446), .B2(n17445), .A(n17444), .ZN(n17554) );
  AND2_X1 U19434 ( .A1(n17448), .A2(n17447), .ZN(n17449) );
  OR2_X1 U19435 ( .A1(n17449), .A2(n17438), .ZN(n19362) );
  NOR2_X1 U19436 ( .A1(n19362), .A2(n17432), .ZN(n17450) );
  AOI21_X1 U19437 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n17432), .A(n17450), .ZN(
        n17451) );
  OAI21_X1 U19438 ( .B1(n17554), .B2(n17452), .A(n17451), .ZN(P2_U2870) );
  NAND2_X1 U19439 ( .A1(n17453), .A2(n20461), .ZN(n17459) );
  OAI22_X1 U19440 ( .A1(n20009), .A2(n20019), .B1(n17454), .B2(n20513), .ZN(
        n17457) );
  INV_X1 U19441 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17455) );
  NOR2_X1 U19442 ( .A1(n17462), .A2(n17455), .ZN(n17456) );
  AOI211_X1 U19443 ( .C1(BUF1_REG_29__SCAN_IN), .C2(n20005), .A(n17457), .B(
        n17456), .ZN(n17458) );
  OAI211_X1 U19444 ( .C1(n19458), .C2(n20515), .A(n17459), .B(n17458), .ZN(
        P2_U2890) );
  OAI22_X1 U19445 ( .A1(n20009), .A2(n20020), .B1(n17460), .B2(n20513), .ZN(
        n17464) );
  INV_X1 U19446 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17461) );
  NOR2_X1 U19447 ( .A1(n17462), .A2(n17461), .ZN(n17463) );
  AOI211_X1 U19448 ( .C1(BUF1_REG_28__SCAN_IN), .C2(n20005), .A(n17464), .B(
        n17463), .ZN(n17467) );
  NAND2_X1 U19449 ( .A1(n17465), .A2(n20459), .ZN(n17466) );
  OAI211_X1 U19450 ( .C1(n17468), .C2(n20517), .A(n17467), .B(n17466), .ZN(
        P2_U2891) );
  NAND2_X1 U19451 ( .A1(n17469), .A2(n20461), .ZN(n17473) );
  INV_X1 U19452 ( .A(n20009), .ZN(n17541) );
  INV_X1 U19453 ( .A(n20513), .ZN(n20457) );
  AOI22_X1 U19454 ( .A1(n17541), .A2(n20023), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20457), .ZN(n17472) );
  AOI22_X1 U19455 ( .A1(n17758), .A2(n20459), .B1(n20005), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n17471) );
  NAND2_X1 U19456 ( .A1(n20003), .A2(BUF2_REG_27__SCAN_IN), .ZN(n17470) );
  NAND4_X1 U19457 ( .A1(n17473), .A2(n17472), .A3(n17471), .A4(n17470), .ZN(
        P2_U2892) );
  NAND2_X1 U19458 ( .A1(n17484), .A2(n17474), .ZN(n17475) );
  NAND2_X1 U19459 ( .A1(n11238), .A2(n17475), .ZN(n17771) );
  INV_X1 U19460 ( .A(n17771), .ZN(n19432) );
  OAI22_X1 U19461 ( .A1(n20009), .A2(n20026), .B1(n17476), .B2(n20513), .ZN(
        n17477) );
  AOI21_X1 U19462 ( .B1(n19432), .B2(n20459), .A(n17477), .ZN(n17479) );
  AOI22_X1 U19463 ( .A1(n20003), .A2(BUF2_REG_26__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n17478) );
  OAI211_X1 U19464 ( .C1(n17480), .C2(n20517), .A(n17479), .B(n17478), .ZN(
        P2_U2893) );
  NAND2_X1 U19465 ( .A1(n17482), .A2(n17481), .ZN(n17483) );
  NAND2_X1 U19466 ( .A1(n17484), .A2(n17483), .ZN(n19422) );
  OAI22_X1 U19467 ( .A1(n19422), .A2(n20515), .B1(n17485), .B2(n20513), .ZN(
        n17487) );
  NOR2_X1 U19468 ( .A1(n20009), .A2(n20031), .ZN(n17486) );
  NOR2_X1 U19469 ( .A1(n17487), .A2(n17486), .ZN(n17489) );
  AOI22_X1 U19470 ( .A1(n20003), .A2(BUF2_REG_25__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n17488) );
  OAI211_X1 U19471 ( .C1(n17490), .C2(n20517), .A(n17489), .B(n17488), .ZN(
        P2_U2894) );
  OAI22_X1 U19472 ( .A1(n20009), .A2(n20032), .B1(n17491), .B2(n20513), .ZN(
        n17492) );
  AOI21_X1 U19473 ( .B1(n17493), .B2(n20459), .A(n17492), .ZN(n17495) );
  AOI22_X1 U19474 ( .A1(n20003), .A2(BUF2_REG_24__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n17494) );
  OAI211_X1 U19475 ( .C1(n17496), .C2(n20517), .A(n17495), .B(n17494), .ZN(
        P2_U2895) );
  OAI22_X1 U19476 ( .A1(n20009), .A2(n20037), .B1(n17497), .B2(n20513), .ZN(
        n17498) );
  AOI21_X1 U19477 ( .B1(n17499), .B2(n20459), .A(n17498), .ZN(n17501) );
  AOI22_X1 U19478 ( .A1(n20003), .A2(BUF2_REG_23__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n17500) );
  OAI211_X1 U19479 ( .C1(n17502), .C2(n20517), .A(n17501), .B(n17500), .ZN(
        P2_U2896) );
  OR2_X1 U19480 ( .A1(n17503), .A2(n17512), .ZN(n17514) );
  AND2_X1 U19481 ( .A1(n17514), .A2(n17504), .ZN(n17505) );
  OR2_X1 U19482 ( .A1(n17505), .A2(n17297), .ZN(n19420) );
  OAI22_X1 U19483 ( .A1(n19420), .A2(n20515), .B1(n17506), .B2(n20513), .ZN(
        n17508) );
  NOR2_X1 U19484 ( .A1(n20009), .A2(n20213), .ZN(n17507) );
  NOR2_X1 U19485 ( .A1(n17508), .A2(n17507), .ZN(n17510) );
  AOI22_X1 U19486 ( .A1(n20003), .A2(BUF2_REG_22__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n17509) );
  OAI211_X1 U19487 ( .C1(n17511), .C2(n20517), .A(n17510), .B(n17509), .ZN(
        P2_U2897) );
  AOI22_X1 U19488 ( .A1(n20003), .A2(BUF2_REG_21__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n17516) );
  NAND2_X1 U19489 ( .A1(n17503), .A2(n17512), .ZN(n17513) );
  AOI22_X1 U19490 ( .A1(n20459), .A2(n19396), .B1(n20457), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n17515) );
  OAI211_X1 U19491 ( .C1(n20268), .C2(n20009), .A(n17516), .B(n17515), .ZN(
        n17517) );
  AOI21_X1 U19492 ( .B1(n17518), .B2(n20461), .A(n17517), .ZN(n17519) );
  INV_X1 U19493 ( .A(n17519), .ZN(P2_U2898) );
  OR2_X1 U19494 ( .A1(n17521), .A2(n17520), .ZN(n17522) );
  NAND2_X1 U19495 ( .A1(n17503), .A2(n17522), .ZN(n19394) );
  OAI22_X1 U19496 ( .A1(n20515), .A2(n19394), .B1(n17523), .B2(n20513), .ZN(
        n17525) );
  NOR2_X1 U19497 ( .A1(n20009), .A2(n20317), .ZN(n17524) );
  NOR2_X1 U19498 ( .A1(n17525), .A2(n17524), .ZN(n17527) );
  AOI22_X1 U19499 ( .A1(n20003), .A2(BUF2_REG_20__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n17526) );
  OAI211_X1 U19500 ( .C1(n17528), .C2(n20517), .A(n17527), .B(n17526), .ZN(
        P2_U2899) );
  OAI22_X1 U19501 ( .A1(n20009), .A2(n20365), .B1(n17529), .B2(n20513), .ZN(
        n17531) );
  NOR2_X1 U19502 ( .A1(n20515), .A2(n17857), .ZN(n17530) );
  NOR2_X1 U19503 ( .A1(n17531), .A2(n17530), .ZN(n17533) );
  AOI22_X1 U19504 ( .A1(n20003), .A2(BUF2_REG_19__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n17532) );
  OAI211_X1 U19505 ( .C1(n17534), .C2(n20517), .A(n17533), .B(n17532), .ZN(
        P2_U2900) );
  INV_X1 U19506 ( .A(n20414), .ZN(n17540) );
  NAND2_X1 U19507 ( .A1(n17548), .A2(n17535), .ZN(n17536) );
  NAND2_X1 U19508 ( .A1(n17537), .A2(n17536), .ZN(n19373) );
  OAI22_X1 U19509 ( .A1(n20515), .A2(n19373), .B1(n17538), .B2(n20513), .ZN(
        n17539) );
  AOI21_X1 U19510 ( .B1(n17541), .B2(n17540), .A(n17539), .ZN(n17543) );
  AOI22_X1 U19511 ( .A1(n20003), .A2(BUF2_REG_18__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n17542) );
  OAI211_X1 U19512 ( .C1(n17544), .C2(n20517), .A(n17543), .B(n17542), .ZN(
        P2_U2901) );
  NAND2_X1 U19513 ( .A1(n17546), .A2(n17545), .ZN(n17547) );
  AND2_X1 U19514 ( .A1(n17548), .A2(n17547), .ZN(n17882) );
  INV_X1 U19515 ( .A(n17882), .ZN(n19361) );
  OAI22_X1 U19516 ( .A1(n20515), .A2(n19361), .B1(n17549), .B2(n20513), .ZN(
        n17551) );
  NOR2_X1 U19517 ( .A1(n20009), .A2(n20466), .ZN(n17550) );
  NOR2_X1 U19518 ( .A1(n17551), .A2(n17550), .ZN(n17553) );
  AOI22_X1 U19519 ( .A1(n20003), .A2(BUF2_REG_17__SCAN_IN), .B1(n20005), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n17552) );
  OAI211_X1 U19520 ( .C1(n17554), .C2(n20517), .A(n17553), .B(n17552), .ZN(
        P2_U2902) );
  XNOR2_X1 U19521 ( .A(n17555), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17766) );
  AOI21_X1 U19522 ( .B1(n17557), .B2(n17565), .A(n17556), .ZN(n17764) );
  NOR2_X1 U19523 ( .A1(n14452), .A2(n18305), .ZN(n17756) );
  NOR2_X1 U19524 ( .A1(n18181), .A2(n17558), .ZN(n17559) );
  AOI211_X1 U19525 ( .C1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18174), .A(
        n17756), .B(n17559), .ZN(n17560) );
  OAI21_X1 U19526 ( .B1(n17762), .B2(n18190), .A(n17560), .ZN(n17561) );
  AOI21_X1 U19527 ( .B1(n17764), .B2(n18198), .A(n17561), .ZN(n17562) );
  OAI21_X1 U19528 ( .B1(n17766), .B2(n18184), .A(n17562), .ZN(P2_U2987) );
  NAND2_X1 U19529 ( .A1(n17563), .A2(n17768), .ZN(n17564) );
  NAND2_X1 U19530 ( .A1(n17565), .A2(n17564), .ZN(n17776) );
  INV_X1 U19531 ( .A(n17566), .ZN(n17567) );
  OAI21_X1 U19532 ( .B1(n17567), .B2(n17580), .A(n12084), .ZN(n17569) );
  MUX2_X1 U19533 ( .A(n17580), .B(n17569), .S(n17568), .Z(n17571) );
  NOR2_X1 U19534 ( .A1(n17571), .A2(n17570), .ZN(n17778) );
  NAND2_X1 U19535 ( .A1(n17778), .A2(n18200), .ZN(n17577) );
  INV_X1 U19536 ( .A(n19436), .ZN(n17572) );
  NAND2_X1 U19537 ( .A1(n18196), .A2(n17572), .ZN(n17573) );
  NAND2_X1 U19538 ( .A1(n19360), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n17769) );
  OAI211_X1 U19539 ( .C1(n17574), .C2(n18204), .A(n17573), .B(n17769), .ZN(
        n17575) );
  AOI21_X1 U19540 ( .B1(n19433), .B2(n18199), .A(n17575), .ZN(n17576) );
  OAI211_X1 U19541 ( .C1(n18185), .C2(n17776), .A(n17577), .B(n17576), .ZN(
        P2_U2988) );
  OAI21_X1 U19542 ( .B1(n17578), .B2(n17794), .A(n17784), .ZN(n17579) );
  NAND2_X1 U19543 ( .A1(n17579), .A2(n17563), .ZN(n17791) );
  NOR2_X1 U19544 ( .A1(n17581), .A2(n17580), .ZN(n17582) );
  XNOR2_X1 U19545 ( .A(n17566), .B(n17582), .ZN(n17780) );
  NAND2_X1 U19546 ( .A1(n17780), .A2(n18200), .ZN(n17588) );
  NAND2_X1 U19547 ( .A1(n19360), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17786) );
  OAI21_X1 U19548 ( .B1(n18204), .B2(n17583), .A(n17786), .ZN(n17585) );
  NOR2_X1 U19549 ( .A1(n17781), .A2(n18190), .ZN(n17584) );
  AOI211_X1 U19550 ( .C1(n18196), .C2(n17586), .A(n17585), .B(n17584), .ZN(
        n17587) );
  OAI211_X1 U19551 ( .C1(n18185), .C2(n17791), .A(n17588), .B(n17587), .ZN(
        P2_U2989) );
  XNOR2_X1 U19552 ( .A(n17578), .B(n17794), .ZN(n17804) );
  OAI21_X1 U19553 ( .B1(n17591), .B2(n17590), .A(n17589), .ZN(n17792) );
  NOR2_X1 U19554 ( .A1(n17793), .A2(n18190), .ZN(n17595) );
  NAND2_X1 U19555 ( .A1(n12603), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n17796) );
  NAND2_X1 U19556 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17592) );
  OAI211_X1 U19557 ( .C1(n18181), .C2(n17593), .A(n17796), .B(n17592), .ZN(
        n17594) );
  AOI211_X1 U19558 ( .C1(n17792), .C2(n18200), .A(n17595), .B(n17594), .ZN(
        n17596) );
  OAI21_X1 U19559 ( .B1(n18185), .B2(n17804), .A(n17596), .ZN(P2_U2990) );
  AND2_X1 U19560 ( .A1(n17598), .A2(n17597), .ZN(n17608) );
  OAI21_X1 U19561 ( .B1(n17608), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17578), .ZN(n17815) );
  OAI21_X1 U19562 ( .B1(n17601), .B2(n17600), .A(n17599), .ZN(n17813) );
  NOR2_X1 U19563 ( .A1(n17811), .A2(n18190), .ZN(n17605) );
  NAND2_X1 U19564 ( .A1(n19360), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17806) );
  NAND2_X1 U19565 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17602) );
  OAI211_X1 U19566 ( .C1(n18181), .C2(n17603), .A(n17806), .B(n17602), .ZN(
        n17604) );
  AOI211_X1 U19567 ( .C1(n17813), .C2(n18200), .A(n17605), .B(n17604), .ZN(
        n17606) );
  OAI21_X1 U19568 ( .B1(n18185), .B2(n17815), .A(n17606), .ZN(P2_U2991) );
  AOI21_X1 U19569 ( .B1(n17624), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17607) );
  OAI21_X1 U19570 ( .B1(n17609), .B2(n17611), .A(n11167), .ZN(n17823) );
  INV_X1 U19571 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n18300) );
  NOR2_X1 U19572 ( .A1(n14452), .A2(n18300), .ZN(n17817) );
  NOR2_X1 U19573 ( .A1(n18181), .A2(n19417), .ZN(n17612) );
  AOI211_X1 U19574 ( .C1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n18174), .A(
        n17817), .B(n17612), .ZN(n17613) );
  OAI21_X1 U19575 ( .B1(n19412), .B2(n18190), .A(n17613), .ZN(n17614) );
  AOI21_X1 U19576 ( .B1(n17823), .B2(n18200), .A(n17614), .ZN(n17615) );
  OAI21_X1 U19577 ( .B1(n18185), .B2(n17825), .A(n17615), .ZN(P2_U2992) );
  INV_X1 U19578 ( .A(n17616), .ZN(n17618) );
  AOI22_X1 U19579 ( .A1(n17619), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17618), .B2(n17617), .ZN(n17622) );
  XNOR2_X1 U19580 ( .A(n17620), .B(n17623), .ZN(n17621) );
  XNOR2_X1 U19581 ( .A(n17622), .B(n17621), .ZN(n17836) );
  XNOR2_X1 U19582 ( .A(n17624), .B(n17623), .ZN(n17834) );
  NOR2_X1 U19583 ( .A1(n19398), .A2(n18190), .ZN(n17627) );
  NAND2_X1 U19584 ( .A1(n19360), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n17828) );
  NAND2_X1 U19585 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17625) );
  OAI211_X1 U19586 ( .C1(n18181), .C2(n19403), .A(n17828), .B(n17625), .ZN(
        n17626) );
  AOI211_X1 U19587 ( .C1(n17834), .C2(n18198), .A(n17627), .B(n17626), .ZN(
        n17628) );
  OAI21_X1 U19588 ( .B1(n17836), .B2(n18184), .A(n17628), .ZN(P2_U2993) );
  NAND2_X1 U19589 ( .A1(n17638), .A2(n17639), .ZN(n17637) );
  NAND2_X1 U19590 ( .A1(n17637), .A2(n17641), .ZN(n17632) );
  NAND2_X1 U19591 ( .A1(n17630), .A2(n17629), .ZN(n17631) );
  XNOR2_X1 U19592 ( .A(n17632), .B(n17631), .ZN(n17865) );
  NOR2_X1 U19593 ( .A1(n17861), .A2(n18190), .ZN(n17636) );
  NAND2_X1 U19594 ( .A1(n19360), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17855) );
  NAND2_X1 U19595 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17633) );
  OAI211_X1 U19596 ( .C1(n18181), .C2(n17634), .A(n17855), .B(n17633), .ZN(
        n17635) );
  INV_X1 U19597 ( .A(n17637), .ZN(n17642) );
  AOI21_X1 U19598 ( .B1(n17641), .B2(n17639), .A(n17638), .ZN(n17640) );
  AOI21_X1 U19599 ( .B1(n17642), .B2(n17641), .A(n17640), .ZN(n17876) );
  INV_X1 U19600 ( .A(n17878), .ZN(n17643) );
  AOI21_X1 U19601 ( .B1(n17643), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17644) );
  NOR2_X1 U19602 ( .A1(n11195), .A2(n17644), .ZN(n17873) );
  NAND2_X1 U19603 ( .A1(n19360), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n17868) );
  OAI21_X1 U19604 ( .B1(n18204), .B2(n19370), .A(n17868), .ZN(n17646) );
  AOI21_X1 U19605 ( .B1(n18196), .B2(n17647), .A(n17646), .ZN(n17648) );
  OAI21_X1 U19606 ( .B1(n19377), .B2(n18190), .A(n17648), .ZN(n17649) );
  OAI21_X1 U19607 ( .B1(n17876), .B2(n18184), .A(n17650), .ZN(P2_U2996) );
  INV_X1 U19608 ( .A(n17651), .ZN(n17653) );
  NOR2_X1 U19609 ( .A1(n17653), .A2(n17652), .ZN(n17654) );
  XNOR2_X1 U19610 ( .A(n17655), .B(n17654), .ZN(n17892) );
  XNOR2_X1 U19611 ( .A(n17878), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17659) );
  NAND2_X1 U19612 ( .A1(n19360), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17884) );
  OAI21_X1 U19613 ( .B1(n18204), .B2(n19358), .A(n17884), .ZN(n17656) );
  AOI21_X1 U19614 ( .B1(n18196), .B2(n19355), .A(n17656), .ZN(n17657) );
  OAI21_X1 U19615 ( .B1(n19362), .B2(n18190), .A(n17657), .ZN(n17658) );
  AOI21_X1 U19616 ( .B1(n17659), .B2(n18198), .A(n17658), .ZN(n17660) );
  OAI21_X1 U19617 ( .B1(n17892), .B2(n18184), .A(n17660), .ZN(P2_U2997) );
  OAI21_X1 U19618 ( .B1(n17663), .B2(n17662), .A(n17661), .ZN(n17893) );
  NAND2_X1 U19619 ( .A1(n12603), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17899) );
  NAND2_X1 U19620 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17664) );
  OAI211_X1 U19621 ( .C1(n18181), .C2(n19342), .A(n17899), .B(n17664), .ZN(
        n17665) );
  AOI21_X1 U19622 ( .B1(n19346), .B2(n18199), .A(n17665), .ZN(n17667) );
  OAI211_X1 U19623 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17896), .A(
        n17878), .B(n18198), .ZN(n17666) );
  OAI211_X1 U19624 ( .C1(n17893), .C2(n18184), .A(n17667), .B(n17666), .ZN(
        P2_U2998) );
  NAND2_X1 U19625 ( .A1(n17668), .A2(n17682), .ZN(n17918) );
  NAND2_X1 U19626 ( .A1(n17918), .A2(n17916), .ZN(n17921) );
  NAND2_X1 U19627 ( .A1(n17921), .A2(n17917), .ZN(n17672) );
  NAND2_X1 U19628 ( .A1(n17670), .A2(n17669), .ZN(n17671) );
  XNOR2_X1 U19629 ( .A(n17672), .B(n17671), .ZN(n17915) );
  AOI21_X1 U19630 ( .B1(n17908), .B2(n17930), .A(n17896), .ZN(n17913) );
  NAND2_X1 U19631 ( .A1(n12603), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17904) );
  OAI21_X1 U19632 ( .B1(n18204), .B2(n17673), .A(n17904), .ZN(n17674) );
  AOI21_X1 U19633 ( .B1(n18196), .B2(n17675), .A(n17674), .ZN(n17676) );
  OAI21_X1 U19634 ( .B1(n17911), .B2(n18190), .A(n17676), .ZN(n17677) );
  AOI21_X1 U19635 ( .B1(n17913), .B2(n18198), .A(n17677), .ZN(n17678) );
  OAI21_X1 U19636 ( .B1(n17915), .B2(n18184), .A(n17678), .ZN(P2_U2999) );
  NAND2_X1 U19637 ( .A1(n17679), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18001) );
  NOR2_X2 U19638 ( .A1(n18001), .A2(n17979), .ZN(n17978) );
  NAND2_X1 U19639 ( .A1(n17978), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17701) );
  OAI21_X1 U19640 ( .B1(n17701), .B2(n17691), .A(n17680), .ZN(n17681) );
  NAND2_X1 U19641 ( .A1(n17681), .A2(n12655), .ZN(n17948) );
  NAND2_X1 U19642 ( .A1(n17683), .A2(n17682), .ZN(n17685) );
  XOR2_X1 U19643 ( .A(n17685), .B(n17684), .Z(n17946) );
  INV_X1 U19644 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n18294) );
  NOR2_X1 U19645 ( .A1(n14452), .A2(n18294), .ZN(n17940) );
  NOR2_X1 U19646 ( .A1(n18181), .A2(n17686), .ZN(n17687) );
  AOI211_X1 U19647 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18174), .A(
        n17940), .B(n17687), .ZN(n17688) );
  OAI21_X1 U19648 ( .B1(n18190), .B2(n17937), .A(n17688), .ZN(n17689) );
  AOI21_X1 U19649 ( .B1(n17946), .B2(n18200), .A(n17689), .ZN(n17690) );
  OAI21_X1 U19650 ( .B1(n18185), .B2(n17948), .A(n17690), .ZN(P2_U3001) );
  XNOR2_X1 U19651 ( .A(n17701), .B(n17691), .ZN(n17962) );
  NAND2_X1 U19652 ( .A1(n12603), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17955) );
  NAND2_X1 U19653 ( .A1(n18174), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17692) );
  OAI211_X1 U19654 ( .C1(n18181), .C2(n19325), .A(n17955), .B(n17692), .ZN(
        n17699) );
  AOI21_X1 U19655 ( .B1(n17694), .B2(n17696), .A(n17693), .ZN(n17695) );
  AOI21_X1 U19656 ( .B1(n17697), .B2(n17696), .A(n17695), .ZN(n17959) );
  NOR2_X1 U19657 ( .A1(n17959), .A2(n18184), .ZN(n17698) );
  AOI211_X1 U19658 ( .C1(n18199), .C2(n19327), .A(n17699), .B(n17698), .ZN(
        n17700) );
  OAI21_X1 U19659 ( .B1(n18185), .B2(n17962), .A(n17700), .ZN(P2_U3002) );
  OAI21_X1 U19660 ( .B1(n17978), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17701), .ZN(n17977) );
  NAND2_X1 U19661 ( .A1(n17702), .A2(n17703), .ZN(n17705) );
  NAND2_X1 U19662 ( .A1(n17705), .A2(n17704), .ZN(n17737) );
  OR2_X1 U19663 ( .A1(n17737), .A2(n17706), .ZN(n17708) );
  NAND2_X1 U19664 ( .A1(n17708), .A2(n17707), .ZN(n17710) );
  NAND2_X1 U19665 ( .A1(n11501), .A2(n17711), .ZN(n17715) );
  NAND2_X1 U19666 ( .A1(n17713), .A2(n17712), .ZN(n17714) );
  XNOR2_X1 U19667 ( .A(n17715), .B(n17714), .ZN(n17974) );
  INV_X1 U19668 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n18292) );
  NOR2_X1 U19669 ( .A1(n14452), .A2(n18292), .ZN(n17967) );
  NOR2_X1 U19670 ( .A1(n18181), .A2(n17716), .ZN(n17717) );
  AOI211_X1 U19671 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18174), .A(
        n17967), .B(n17717), .ZN(n17718) );
  OAI21_X1 U19672 ( .B1(n18190), .B2(n17971), .A(n17718), .ZN(n17719) );
  AOI21_X1 U19673 ( .B1(n17974), .B2(n18200), .A(n17719), .ZN(n17720) );
  OAI21_X1 U19674 ( .B1(n17977), .B2(n18185), .A(n17720), .ZN(P2_U3003) );
  NAND2_X1 U19675 ( .A1(n18018), .A2(n17721), .ZN(n17722) );
  INV_X1 U19676 ( .A(n17980), .ZN(n17726) );
  OAI21_X1 U19677 ( .B1(n17724), .B2(n17726), .A(n17723), .ZN(n17725) );
  OAI21_X1 U19678 ( .B1(n17981), .B2(n17726), .A(n17725), .ZN(n18013) );
  INV_X1 U19679 ( .A(n17679), .ZN(n17728) );
  NAND2_X1 U19680 ( .A1(n17728), .A2(n17727), .ZN(n18002) );
  NAND3_X1 U19681 ( .A1(n18002), .A2(n18198), .A3(n18001), .ZN(n17733) );
  NOR2_X1 U19682 ( .A1(n18190), .A2(n18006), .ZN(n17731) );
  INV_X1 U19683 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n18288) );
  OAI22_X1 U19684 ( .A1(n18288), .A2(n14452), .B1(n18181), .B2(n17729), .ZN(
        n17730) );
  AOI211_X1 U19685 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18174), .A(
        n17731), .B(n17730), .ZN(n17732) );
  OAI211_X1 U19686 ( .C1(n18013), .C2(n18184), .A(n17733), .B(n17732), .ZN(
        P2_U3005) );
  INV_X1 U19687 ( .A(n18017), .ZN(n17735) );
  NOR2_X1 U19688 ( .A1(n17735), .A2(n17734), .ZN(n17736) );
  XNOR2_X1 U19689 ( .A(n17737), .B(n17736), .ZN(n18052) );
  OR2_X1 U19690 ( .A1(n17739), .A2(n17738), .ZN(n18042) );
  NAND3_X1 U19691 ( .A1(n18042), .A2(n18198), .A3(n17740), .ZN(n17746) );
  NOR2_X1 U19692 ( .A1(n18190), .A2(n18043), .ZN(n17743) );
  INV_X1 U19693 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18285) );
  OAI22_X1 U19694 ( .A1(n17741), .A2(n18204), .B1(n18285), .B2(n14452), .ZN(
        n17742) );
  AOI211_X1 U19695 ( .C1(n18196), .C2(n17744), .A(n17743), .B(n17742), .ZN(
        n17745) );
  OAI211_X1 U19696 ( .C1(n18052), .C2(n18184), .A(n17746), .B(n17745), .ZN(
        P2_U3007) );
  OR2_X1 U19697 ( .A1(n17747), .A2(n18184), .ZN(n17755) );
  OAI22_X1 U19698 ( .A1(n17748), .A2(n18204), .B1(n18277), .B2(n14452), .ZN(
        n17749) );
  AOI21_X1 U19699 ( .B1(n18196), .B2(n17750), .A(n17749), .ZN(n17754) );
  NAND3_X1 U19700 ( .A1(n15563), .A2(n17751), .A3(n18198), .ZN(n17753) );
  NAND2_X1 U19701 ( .A1(n11196), .A2(n18199), .ZN(n17752) );
  NAND4_X1 U19702 ( .A1(n17755), .A2(n17754), .A3(n17753), .A4(n17752), .ZN(
        P2_U3011) );
  AOI211_X1 U19703 ( .C1(n17758), .C2(n19500), .A(n17757), .B(n17756), .ZN(
        n17761) );
  NAND2_X1 U19704 ( .A1(n17759), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17760) );
  OAI211_X1 U19705 ( .C1(n17762), .C2(n18061), .A(n17761), .B(n17760), .ZN(
        n17763) );
  AOI21_X1 U19706 ( .B1(n17764), .B2(n18055), .A(n17763), .ZN(n17765) );
  OAI21_X1 U19707 ( .B1(n17766), .B2(n19495), .A(n17765), .ZN(P2_U3019) );
  OAI21_X1 U19708 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17767), .A(
        n17782), .ZN(n17773) );
  NAND3_X1 U19709 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17783), .A3(
        n17768), .ZN(n17770) );
  OAI211_X1 U19710 ( .C1(n17771), .C2(n18066), .A(n17770), .B(n17769), .ZN(
        n17772) );
  AOI21_X1 U19711 ( .B1(n17773), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17772), .ZN(n17775) );
  NAND2_X1 U19712 ( .A1(n19433), .A2(n19504), .ZN(n17774) );
  OAI211_X1 U19713 ( .C1(n17776), .C2(n19508), .A(n17775), .B(n17774), .ZN(
        n17777) );
  AOI21_X1 U19714 ( .B1(n17778), .B2(n14175), .A(n17777), .ZN(n17779) );
  INV_X1 U19715 ( .A(n17779), .ZN(P2_U3020) );
  NAND2_X1 U19716 ( .A1(n17780), .A2(n14175), .ZN(n17790) );
  INV_X1 U19717 ( .A(n17781), .ZN(n19424) );
  NOR2_X1 U19718 ( .A1(n17782), .A2(n17784), .ZN(n17788) );
  NAND2_X1 U19719 ( .A1(n17784), .A2(n17783), .ZN(n17785) );
  OAI211_X1 U19720 ( .C1(n19422), .C2(n18066), .A(n17786), .B(n17785), .ZN(
        n17787) );
  AOI211_X1 U19721 ( .C1(n19424), .C2(n19504), .A(n17788), .B(n17787), .ZN(
        n17789) );
  OAI211_X1 U19722 ( .C1(n17791), .C2(n19508), .A(n17790), .B(n17789), .ZN(
        P2_U3021) );
  NAND2_X1 U19723 ( .A1(n17792), .A2(n14175), .ZN(n17803) );
  INV_X1 U19724 ( .A(n17793), .ZN(n17801) );
  NOR2_X1 U19725 ( .A1(n17795), .A2(n17794), .ZN(n17800) );
  OAI211_X1 U19726 ( .C1(n17798), .C2(n18066), .A(n17797), .B(n17796), .ZN(
        n17799) );
  AOI211_X1 U19727 ( .C1(n17801), .C2(n19504), .A(n17800), .B(n17799), .ZN(
        n17802) );
  OAI211_X1 U19728 ( .C1(n17804), .C2(n19508), .A(n17803), .B(n17802), .ZN(
        P2_U3022) );
  XOR2_X1 U19729 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17805) );
  NAND2_X1 U19730 ( .A1(n17819), .A2(n17805), .ZN(n17807) );
  OAI211_X1 U19731 ( .C1(n18066), .C2(n17808), .A(n17807), .B(n17806), .ZN(
        n17809) );
  AOI21_X1 U19732 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17826), .A(
        n17809), .ZN(n17810) );
  OAI21_X1 U19733 ( .B1(n17811), .B2(n18061), .A(n17810), .ZN(n17812) );
  AOI21_X1 U19734 ( .B1(n17813), .B2(n14175), .A(n17812), .ZN(n17814) );
  OAI21_X1 U19735 ( .B1(n19508), .B2(n17815), .A(n17814), .ZN(P2_U3023) );
  INV_X1 U19736 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17818) );
  NOR2_X1 U19737 ( .A1(n19420), .A2(n18066), .ZN(n17816) );
  AOI211_X1 U19738 ( .C1(n17819), .C2(n17818), .A(n17817), .B(n17816), .ZN(
        n17821) );
  NAND2_X1 U19739 ( .A1(n17826), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17820) );
  OAI211_X1 U19740 ( .C1(n19412), .C2(n18061), .A(n17821), .B(n17820), .ZN(
        n17822) );
  AOI21_X1 U19741 ( .B1(n17823), .B2(n14175), .A(n17822), .ZN(n17824) );
  OAI21_X1 U19742 ( .B1(n19508), .B2(n17825), .A(n17824), .ZN(P2_U3024) );
  NOR2_X1 U19743 ( .A1(n19398), .A2(n18061), .ZN(n17833) );
  INV_X1 U19744 ( .A(n17826), .ZN(n17831) );
  AOI21_X1 U19745 ( .B1(n17964), .B2(n17827), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17830) );
  NAND2_X1 U19746 ( .A1(n19500), .A2(n19396), .ZN(n17829) );
  OAI211_X1 U19747 ( .C1(n17831), .C2(n17830), .A(n17829), .B(n17828), .ZN(
        n17832) );
  AOI211_X1 U19748 ( .C1(n17834), .C2(n18055), .A(n17833), .B(n17832), .ZN(
        n17835) );
  OAI21_X1 U19749 ( .B1(n17836), .B2(n19495), .A(n17835), .ZN(P2_U3025) );
  INV_X1 U19750 ( .A(n17841), .ZN(n17839) );
  INV_X1 U19751 ( .A(n17837), .ZN(n17840) );
  OAI21_X1 U19752 ( .B1(n19502), .B2(n17840), .A(n18003), .ZN(n17879) );
  AOI21_X1 U19753 ( .B1(n17839), .B2(n17838), .A(n17879), .ZN(n17867) );
  AND2_X1 U19754 ( .A1(n17964), .A2(n17840), .ZN(n17909) );
  NAND2_X1 U19755 ( .A1(n17909), .A2(n17841), .ZN(n17843) );
  INV_X1 U19756 ( .A(n17843), .ZN(n17854) );
  NAND2_X1 U19757 ( .A1(n17854), .A2(n17866), .ZN(n17869) );
  NAND2_X1 U19758 ( .A1(n17867), .A2(n17869), .ZN(n17859) );
  OAI21_X1 U19759 ( .B1(n18066), .B2(n19394), .A(n17842), .ZN(n17847) );
  AOI21_X1 U19760 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17845), .A(
        n17853), .ZN(n17844) );
  AOI211_X1 U19761 ( .C1(n17853), .C2(n17845), .A(n17844), .B(n17843), .ZN(
        n17846) );
  AOI211_X1 U19762 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n17859), .A(
        n17847), .B(n17846), .ZN(n17848) );
  OAI21_X1 U19763 ( .B1(n19384), .B2(n18061), .A(n17848), .ZN(n17849) );
  AOI21_X1 U19764 ( .B1(n17850), .B2(n18055), .A(n17849), .ZN(n17851) );
  OAI21_X1 U19765 ( .B1(n17852), .B2(n19495), .A(n17851), .ZN(P2_U3026) );
  NAND3_X1 U19766 ( .A1(n17854), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17853), .ZN(n17856) );
  OAI211_X1 U19767 ( .C1(n18066), .C2(n17857), .A(n17856), .B(n17855), .ZN(
        n17858) );
  AOI21_X1 U19768 ( .B1(n17859), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n17858), .ZN(n17860) );
  OAI21_X1 U19769 ( .B1(n17861), .B2(n18061), .A(n17860), .ZN(n17862) );
  AOI21_X1 U19770 ( .B1(n17863), .B2(n18055), .A(n17862), .ZN(n17864) );
  OAI21_X1 U19771 ( .B1(n17865), .B2(n19495), .A(n17864), .ZN(P2_U3027) );
  INV_X1 U19772 ( .A(n19377), .ZN(n17872) );
  NOR2_X1 U19773 ( .A1(n17867), .A2(n17866), .ZN(n17871) );
  OAI211_X1 U19774 ( .C1(n18066), .C2(n19373), .A(n17869), .B(n17868), .ZN(
        n17870) );
  AOI211_X1 U19775 ( .C1(n17872), .C2(n19504), .A(n17871), .B(n17870), .ZN(
        n17875) );
  NAND2_X1 U19776 ( .A1(n17873), .A2(n18055), .ZN(n17874) );
  OAI211_X1 U19777 ( .C1(n17876), .C2(n19495), .A(n17875), .B(n17874), .ZN(
        P2_U3028) );
  NAND2_X1 U19778 ( .A1(n19508), .A2(n17877), .ZN(n17894) );
  NAND2_X1 U19779 ( .A1(n17878), .A2(n17894), .ZN(n17881) );
  AOI21_X1 U19780 ( .B1(n17880), .B2(n17908), .A(n17879), .ZN(n17905) );
  OAI211_X1 U19781 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n19502), .A(
        n17881), .B(n17905), .ZN(n17890) );
  NAND2_X1 U19782 ( .A1(n19500), .A2(n17882), .ZN(n17883) );
  OAI211_X1 U19783 ( .C1(n19362), .C2(n18061), .A(n17884), .B(n17883), .ZN(
        n17889) );
  INV_X1 U19784 ( .A(n17909), .ZN(n17885) );
  OAI21_X1 U19785 ( .B1(n17930), .B2(n19508), .A(n17885), .ZN(n17886) );
  NAND2_X1 U19786 ( .A1(n17886), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17903) );
  INV_X1 U19787 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17887) );
  NOR3_X1 U19788 ( .A1(n17903), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n17887), .ZN(n17888) );
  OAI21_X1 U19789 ( .B1(n17892), .B2(n19495), .A(n17891), .ZN(P2_U3029) );
  INV_X1 U19790 ( .A(n17893), .ZN(n17898) );
  INV_X1 U19791 ( .A(n17894), .ZN(n17895) );
  OAI21_X1 U19792 ( .B1(n17896), .B2(n17895), .A(n17905), .ZN(n17897) );
  AOI22_X1 U19793 ( .A1(n17898), .A2(n14175), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17897), .ZN(n17902) );
  OAI21_X1 U19794 ( .B1(n18066), .B2(n19347), .A(n17899), .ZN(n17900) );
  AOI21_X1 U19795 ( .B1(n19346), .B2(n19504), .A(n17900), .ZN(n17901) );
  OAI211_X1 U19796 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17903), .A(
        n17902), .B(n17901), .ZN(P2_U3030) );
  OAI21_X1 U19797 ( .B1(n18066), .B2(n20013), .A(n17904), .ZN(n17907) );
  NOR2_X1 U19798 ( .A1(n17905), .A2(n17908), .ZN(n17906) );
  AOI211_X1 U19799 ( .C1(n17909), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        n17910) );
  OAI21_X1 U19800 ( .B1(n18061), .B2(n17911), .A(n17910), .ZN(n17912) );
  AOI21_X1 U19801 ( .B1(n17913), .B2(n18055), .A(n17912), .ZN(n17914) );
  OAI21_X1 U19802 ( .B1(n17915), .B2(n19495), .A(n17914), .ZN(P2_U3031) );
  INV_X1 U19803 ( .A(n17917), .ZN(n17920) );
  AND2_X1 U19804 ( .A1(n17917), .A2(n17916), .ZN(n17919) );
  OAI22_X1 U19805 ( .A1(n17921), .A2(n17920), .B1(n17919), .B2(n17918), .ZN(
        n18201) );
  NAND2_X1 U19806 ( .A1(n18201), .A2(n14175), .ZN(n17936) );
  NAND2_X1 U19807 ( .A1(n17327), .A2(n17922), .ZN(n17923) );
  NAND2_X1 U19808 ( .A1(n14537), .A2(n17923), .ZN(n20016) );
  OAI22_X1 U19809 ( .A1(n18066), .A2(n20016), .B1(n17924), .B2(n14452), .ZN(
        n17927) );
  INV_X1 U19810 ( .A(n17964), .ZN(n18007) );
  NOR3_X1 U19811 ( .A1(n18007), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n11446), .ZN(n17926) );
  AOI211_X1 U19812 ( .C1(n19336), .C2(n19504), .A(n17927), .B(n17926), .ZN(
        n17935) );
  NAND2_X1 U19813 ( .A1(n12655), .A2(n17928), .ZN(n17929) );
  AND2_X1 U19814 ( .A1(n17930), .A2(n17929), .ZN(n18197) );
  NAND2_X1 U19815 ( .A1(n18197), .A2(n18055), .ZN(n17934) );
  AND2_X1 U19816 ( .A1(n17964), .A2(n17931), .ZN(n17966) );
  NAND2_X1 U19817 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17966), .ZN(
        n17932) );
  NOR2_X1 U19818 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17932), .ZN(
        n17938) );
  OR2_X1 U19819 ( .A1(n17932), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17956) );
  OAI211_X1 U19820 ( .C1(n17952), .C2(n19502), .A(n18003), .B(n17956), .ZN(
        n17939) );
  OAI21_X1 U19821 ( .B1(n17938), .B2(n17939), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17933) );
  NAND4_X1 U19822 ( .A1(n17936), .A2(n17935), .A3(n17934), .A4(n17933), .ZN(
        P2_U3032) );
  NOR2_X1 U19823 ( .A1(n17937), .A2(n18061), .ZN(n17945) );
  AOI22_X1 U19824 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17939), .B1(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17938), .ZN(n17942) );
  INV_X1 U19825 ( .A(n17940), .ZN(n17941) );
  OAI211_X1 U19826 ( .C1(n18066), .C2(n17943), .A(n17942), .B(n17941), .ZN(
        n17944) );
  AOI211_X1 U19827 ( .C1(n17946), .C2(n14175), .A(n17945), .B(n17944), .ZN(
        n17947) );
  OAI21_X1 U19828 ( .B1(n19508), .B2(n17948), .A(n17947), .ZN(P2_U3033) );
  INV_X1 U19829 ( .A(n17326), .ZN(n17949) );
  OAI21_X1 U19830 ( .B1(n17951), .B2(n17950), .A(n17949), .ZN(n20022) );
  OAI21_X1 U19831 ( .B1(n17952), .B2(n19502), .A(n18003), .ZN(n17953) );
  NAND2_X1 U19832 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17953), .ZN(
        n17954) );
  OAI211_X1 U19833 ( .C1(n18066), .C2(n20022), .A(n17955), .B(n17954), .ZN(
        n17958) );
  INV_X1 U19834 ( .A(n17956), .ZN(n17957) );
  AOI211_X1 U19835 ( .C1(n19504), .C2(n19327), .A(n17958), .B(n17957), .ZN(
        n17961) );
  OR2_X1 U19836 ( .A1(n17959), .A2(n19495), .ZN(n17960) );
  OAI211_X1 U19837 ( .C1(n17962), .C2(n19508), .A(n17961), .B(n17960), .ZN(
        P2_U3034) );
  AND2_X1 U19838 ( .A1(n17979), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17963) );
  NAND2_X1 U19839 ( .A1(n17964), .A2(n17963), .ZN(n17996) );
  OAI211_X1 U19840 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n19502), .A(
        n18003), .B(n17996), .ZN(n17973) );
  NAND2_X1 U19841 ( .A1(n17966), .A2(n17965), .ZN(n17970) );
  AOI21_X1 U19842 ( .B1(n19500), .B2(n17968), .A(n17967), .ZN(n17969) );
  OAI211_X1 U19843 ( .C1(n17971), .C2(n18061), .A(n17970), .B(n17969), .ZN(
        n17972) );
  AOI21_X1 U19844 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n17973), .A(
        n17972), .ZN(n17976) );
  NAND2_X1 U19845 ( .A1(n17974), .A2(n14175), .ZN(n17975) );
  OAI211_X1 U19846 ( .C1(n17977), .C2(n19508), .A(n17976), .B(n17975), .ZN(
        P2_U3035) );
  AOI21_X1 U19847 ( .B1(n17979), .B2(n18001), .A(n17978), .ZN(n18191) );
  INV_X1 U19848 ( .A(n18191), .ZN(n18000) );
  NAND2_X1 U19849 ( .A1(n17981), .A2(n17980), .ZN(n17986) );
  INV_X1 U19850 ( .A(n17982), .ZN(n17984) );
  OR2_X1 U19851 ( .A1(n17984), .A2(n17983), .ZN(n17985) );
  XNOR2_X1 U19852 ( .A(n17986), .B(n17985), .ZN(n18192) );
  INV_X1 U19853 ( .A(n17987), .ZN(n19318) );
  NAND2_X1 U19854 ( .A1(n19318), .A2(n19504), .ZN(n17997) );
  OAI21_X1 U19855 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19502), .A(
        n18003), .ZN(n17988) );
  AOI22_X1 U19856 ( .A1(n12603), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17988), .ZN(n17995) );
  OR2_X1 U19857 ( .A1(n17990), .A2(n17989), .ZN(n17992) );
  NAND2_X1 U19858 ( .A1(n17992), .A2(n17991), .ZN(n20028) );
  INV_X1 U19859 ( .A(n20028), .ZN(n17993) );
  NAND2_X1 U19860 ( .A1(n19500), .A2(n17993), .ZN(n17994) );
  NAND4_X1 U19861 ( .A1(n17997), .A2(n17996), .A3(n17995), .A4(n17994), .ZN(
        n17998) );
  AOI21_X1 U19862 ( .B1(n18192), .B2(n14175), .A(n17998), .ZN(n17999) );
  OAI21_X1 U19863 ( .B1(n18000), .B2(n19508), .A(n17999), .ZN(P2_U3036) );
  NAND3_X1 U19864 ( .A1(n18002), .A2(n18055), .A3(n18001), .ZN(n18012) );
  INV_X1 U19865 ( .A(n18003), .ZN(n18010) );
  NAND2_X1 U19866 ( .A1(n19500), .A2(n20029), .ZN(n18005) );
  NAND2_X1 U19867 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19360), .ZN(n18004) );
  OAI211_X1 U19868 ( .C1(n18006), .C2(n18061), .A(n18005), .B(n18004), .ZN(
        n18009) );
  NOR2_X1 U19869 ( .A1(n18007), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18008) );
  AOI211_X1 U19870 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18010), .A(
        n18009), .B(n18008), .ZN(n18011) );
  OAI211_X1 U19871 ( .C1(n19495), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        P2_U3037) );
  OAI21_X1 U19872 ( .B1(n18016), .B2(n18015), .A(n18014), .ZN(n18186) );
  NAND2_X1 U19873 ( .A1(n18018), .A2(n18017), .ZN(n18022) );
  NAND2_X1 U19874 ( .A1(n18020), .A2(n18019), .ZN(n18021) );
  XNOR2_X1 U19875 ( .A(n18022), .B(n18021), .ZN(n18183) );
  INV_X1 U19876 ( .A(n18183), .ZN(n18040) );
  NOR2_X1 U19877 ( .A1(n18026), .A2(n18023), .ZN(n18069) );
  NAND2_X1 U19878 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18069), .ZN(
        n18047) );
  AOI211_X1 U19879 ( .C1(n18037), .C2(n18046), .A(n18024), .B(n18047), .ZN(
        n18039) );
  OAI21_X1 U19880 ( .B1(n18026), .B2(n18025), .A(n18030), .ZN(n18027) );
  OAI211_X1 U19881 ( .C1(n18029), .C2(n18028), .A(n18027), .B(n19497), .ZN(
        n18064) );
  AOI21_X1 U19882 ( .B1(n18030), .B2(n18068), .A(n18064), .ZN(n18045) );
  INV_X1 U19883 ( .A(n19305), .ZN(n18031) );
  AOI22_X1 U19884 ( .A1(n19504), .A2(n18031), .B1(P2_REIP_REG_8__SCAN_IN), 
        .B2(n12603), .ZN(n18036) );
  OAI21_X1 U19885 ( .B1(n18033), .B2(n15197), .A(n18032), .ZN(n20034) );
  INV_X1 U19886 ( .A(n20034), .ZN(n18034) );
  NAND2_X1 U19887 ( .A1(n19500), .A2(n18034), .ZN(n18035) );
  OAI211_X1 U19888 ( .C1(n18045), .C2(n18037), .A(n18036), .B(n18035), .ZN(
        n18038) );
  AOI211_X1 U19889 ( .C1(n18040), .C2(n14175), .A(n18039), .B(n18038), .ZN(
        n18041) );
  OAI21_X1 U19890 ( .B1(n18186), .B2(n19508), .A(n18041), .ZN(P2_U3038) );
  NAND3_X1 U19891 ( .A1(n18042), .A2(n18055), .A3(n17740), .ZN(n18051) );
  NOR2_X1 U19892 ( .A1(n18043), .A2(n18061), .ZN(n18049) );
  NAND2_X1 U19893 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19360), .ZN(n18044) );
  OAI221_X1 U19894 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18047), .C1(
        n18046), .C2(n18045), .A(n18044), .ZN(n18048) );
  AOI211_X1 U19895 ( .C1(n20035), .C2(n19500), .A(n18049), .B(n18048), .ZN(
        n18050) );
  OAI211_X1 U19896 ( .C1(n18052), .C2(n19495), .A(n18051), .B(n18050), .ZN(
        P2_U3039) );
  XNOR2_X1 U19897 ( .A(n17702), .B(n17703), .ZN(n18176) );
  NOR2_X1 U19898 ( .A1(n18053), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18175) );
  INV_X1 U19899 ( .A(n18175), .ZN(n18056) );
  NAND3_X1 U19900 ( .A1(n18056), .A2(n18055), .A3(n18054), .ZN(n18071) );
  AOI21_X1 U19901 ( .B1(n18059), .B2(n18058), .A(n18057), .ZN(n18060) );
  INV_X1 U19902 ( .A(n18060), .ZN(n20210) );
  INV_X1 U19903 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n18283) );
  NOR2_X1 U19904 ( .A1(n18283), .A2(n14452), .ZN(n18063) );
  NOR2_X1 U19905 ( .A1(n18061), .A2(n19292), .ZN(n18062) );
  AOI211_X1 U19906 ( .C1(n18064), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n18063), .B(n18062), .ZN(n18065) );
  OAI21_X1 U19907 ( .B1(n20210), .B2(n18066), .A(n18065), .ZN(n18067) );
  AOI21_X1 U19908 ( .B1(n18069), .B2(n18068), .A(n18067), .ZN(n18070) );
  OAI211_X1 U19909 ( .C1(n18176), .C2(n19495), .A(n18071), .B(n18070), .ZN(
        P2_U3040) );
  AOI222_X1 U19910 ( .A1(n18074), .A2(n18078), .B1(n18073), .B2(n18072), .C1(
        n19529), .C2(n20255), .ZN(n18077) );
  NAND2_X1 U19911 ( .A1(n18076), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n18075) );
  OAI21_X1 U19912 ( .B1(n18077), .B2(n18076), .A(n18075), .ZN(P2_U3600) );
  INV_X1 U19913 ( .A(n19529), .ZN(n18080) );
  INV_X1 U19914 ( .A(n18078), .ZN(n19512) );
  OAI22_X1 U19915 ( .A1(n20262), .A2(n18080), .B1(n18079), .B2(n19512), .ZN(
        n18081) );
  MUX2_X1 U19916 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n18081), .S(
        n19493), .Z(P2_U3596) );
  NAND2_X1 U19917 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19594) );
  NAND2_X1 U19918 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19098) );
  NAND2_X1 U19919 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18082) );
  INV_X1 U19920 ( .A(n18082), .ZN(n18700) );
  NOR2_X1 U19921 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18700), .ZN(n20944) );
  AND2_X1 U19922 ( .A1(n19098), .A2(n20944), .ZN(n18084) );
  NAND2_X1 U19923 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19617), .ZN(n19570) );
  NOR2_X1 U19924 ( .A1(n22113), .A2(n18082), .ZN(n22098) );
  INV_X1 U19925 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21044) );
  OAI21_X1 U19926 ( .B1(n21622), .B2(n21640), .A(n21044), .ZN(n18091) );
  NOR2_X1 U19927 ( .A1(n18548), .A2(n18091), .ZN(n18701) );
  INV_X1 U19928 ( .A(n18701), .ZN(n18083) );
  AOI21_X1 U19929 ( .B1(n22102), .B2(n18082), .A(n22105), .ZN(n19568) );
  AOI221_X1 U19930 ( .B1(n22098), .B2(n18083), .C1(n22098), .C2(
        P3_FLUSH_REG_SCAN_IN), .A(n19854), .ZN(n18703) );
  INV_X1 U19931 ( .A(n18703), .ZN(n18096) );
  NAND2_X1 U19932 ( .A1(n19570), .A2(n18096), .ZN(n19149) );
  AOI221_X1 U19933 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19594), .C1(n18084), 
        .C2(n19594), .A(n19149), .ZN(n19148) );
  NOR2_X1 U19934 ( .A1(n22100), .A2(n19617), .ZN(n19584) );
  OAI21_X1 U19935 ( .B1(n18084), .B2(n19584), .A(n18096), .ZN(n19151) );
  INV_X1 U19936 ( .A(n19151), .ZN(n18085) );
  NAND3_X1 U19937 ( .A1(n22091), .A2(n22100), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19596) );
  INV_X1 U19938 ( .A(n19596), .ZN(n19613) );
  AOI22_X1 U19939 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18085), .B1(
        n19613), .B2(n18096), .ZN(n19147) );
  AOI22_X1 U19940 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19148), .B1(
        n19147), .B2(n22076), .ZN(P3_U2865) );
  NAND2_X1 U19941 ( .A1(n22063), .A2(n20941), .ZN(n21426) );
  NAND2_X1 U19942 ( .A1(n20936), .A2(n18087), .ZN(n18097) );
  OAI221_X1 U19943 ( .B1(n21426), .B2(n21427), .C1(n21426), .C2(n18097), .A(
        n18088), .ZN(n18089) );
  NOR2_X1 U19944 ( .A1(n18319), .A2(n18089), .ZN(n22074) );
  NAND2_X1 U19945 ( .A1(n22113), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19567) );
  NAND2_X1 U19946 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n22098), .ZN(n18090) );
  OAI211_X1 U19947 ( .C1(n22088), .C2(n22074), .A(n19567), .B(n18090), .ZN(
        n21654) );
  NOR2_X1 U19948 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21652) );
  AND2_X1 U19949 ( .A1(n18091), .A2(n21616), .ZN(n22064) );
  NAND3_X1 U19950 ( .A1(n21654), .A2(n21652), .A3(n22064), .ZN(n18092) );
  OAI21_X1 U19951 ( .B1(n21654), .B2(n21044), .A(n18092), .ZN(P3_U3284) );
  OAI21_X1 U19952 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n22419), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n19217) );
  NAND2_X1 U19953 ( .A1(n19239), .A2(n19217), .ZN(n18094) );
  INV_X1 U19954 ( .A(n18094), .ZN(n22418) );
  NOR2_X1 U19955 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n19177) );
  OAI21_X1 U19956 ( .B1(BS16), .B2(n19177), .A(n22418), .ZN(n22416) );
  OAI21_X1 U19957 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n22418), .A(n22416), 
        .ZN(n18093) );
  INV_X1 U19958 ( .A(n18093), .ZN(P3_U3280) );
  AND2_X1 U19959 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18094), .ZN(P3_U3028) );
  AND2_X1 U19960 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18094), .ZN(P3_U3027) );
  AND2_X1 U19961 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18094), .ZN(P3_U3026) );
  AND2_X1 U19962 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18094), .ZN(P3_U3025) );
  AND2_X1 U19963 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18094), .ZN(P3_U3024) );
  AND2_X1 U19964 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18094), .ZN(P3_U3023) );
  AND2_X1 U19965 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18094), .ZN(P3_U3022) );
  AND2_X1 U19966 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18094), .ZN(P3_U3021) );
  AND2_X1 U19967 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18094), .ZN(
        P3_U3020) );
  AND2_X1 U19968 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18094), .ZN(
        P3_U3019) );
  AND2_X1 U19969 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18094), .ZN(
        P3_U3018) );
  AND2_X1 U19970 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18094), .ZN(
        P3_U3017) );
  AND2_X1 U19971 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18094), .ZN(
        P3_U3016) );
  AND2_X1 U19972 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18094), .ZN(
        P3_U3015) );
  AND2_X1 U19973 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18094), .ZN(
        P3_U3014) );
  AND2_X1 U19974 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18094), .ZN(
        P3_U3013) );
  AND2_X1 U19975 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18094), .ZN(
        P3_U3012) );
  AND2_X1 U19976 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18094), .ZN(
        P3_U3011) );
  AND2_X1 U19977 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18094), .ZN(
        P3_U3010) );
  AND2_X1 U19978 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18094), .ZN(
        P3_U3009) );
  AND2_X1 U19979 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18094), .ZN(
        P3_U3008) );
  AND2_X1 U19980 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18094), .ZN(
        P3_U3007) );
  AND2_X1 U19981 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18094), .ZN(
        P3_U3006) );
  AND2_X1 U19982 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18094), .ZN(
        P3_U3005) );
  AND2_X1 U19983 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18094), .ZN(
        P3_U3004) );
  AND2_X1 U19984 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18094), .ZN(
        P3_U3003) );
  AND2_X1 U19985 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18094), .ZN(
        P3_U3002) );
  AND2_X1 U19986 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18094), .ZN(
        P3_U3001) );
  AND2_X1 U19987 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18094), .ZN(
        P3_U3000) );
  AND2_X1 U19988 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18094), .ZN(
        P3_U2999) );
  AOI21_X1 U19989 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18095)
         );
  NOR4_X1 U19990 ( .A1(n21612), .A2(n22113), .A3(n20941), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n22058) );
  AOI211_X1 U19991 ( .C1(n19098), .C2(n18095), .A(n22098), .B(n22058), .ZN(
        P3_U2998) );
  NOR2_X1 U19992 ( .A1(n22080), .A2(n18096), .ZN(P3_U2867) );
  NAND2_X1 U19993 ( .A1(n22113), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18899) );
  NOR2_X1 U19994 ( .A1(n21612), .A2(n18899), .ZN(n19206) );
  AND2_X1 U19995 ( .A1(n19208), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NOR2_X1 U19996 ( .A1(n18696), .A2(n20942), .ZN(n18098) );
  INV_X1 U19997 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19175) );
  AOI22_X1 U19998 ( .A1(n18098), .A2(n19175), .B1(n20942), .B2(n20939), .ZN(
        P3_U3298) );
  INV_X1 U19999 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19174) );
  NAND2_X1 U20000 ( .A1(n19905), .A2(n20942), .ZN(n21423) );
  INV_X1 U20001 ( .A(n21423), .ZN(n21021) );
  AOI21_X1 U20002 ( .B1(n18098), .B2(n19174), .A(n21021), .ZN(P3_U3299) );
  AOI21_X1 U20003 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n18100), .A(n18099), 
        .ZN(n18102) );
  INV_X1 U20004 ( .A(n18102), .ZN(n22414) );
  NOR2_X1 U20005 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n22429) );
  OAI21_X1 U20006 ( .B1(BS16), .B2(n22429), .A(n22414), .ZN(n22412) );
  OAI21_X1 U20007 ( .B1(n22414), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n22412), 
        .ZN(n18101) );
  INV_X1 U20008 ( .A(n18101), .ZN(P2_U3591) );
  AND2_X1 U20009 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n18102), .ZN(P2_U3208) );
  AND2_X1 U20010 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n18102), .ZN(P2_U3207) );
  INV_X1 U20011 ( .A(n22414), .ZN(n18103) );
  AND2_X1 U20012 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n18103), .ZN(P2_U3206) );
  AND2_X1 U20013 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n18102), .ZN(P2_U3205) );
  AND2_X1 U20014 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n18103), .ZN(P2_U3204) );
  AND2_X1 U20015 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n18102), .ZN(P2_U3203) );
  AND2_X1 U20016 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n18103), .ZN(P2_U3202) );
  AND2_X1 U20017 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n18103), .ZN(P2_U3201) );
  AND2_X1 U20018 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n18103), .ZN(
        P2_U3200) );
  AND2_X1 U20019 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n18103), .ZN(
        P2_U3199) );
  AND2_X1 U20020 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n18103), .ZN(
        P2_U3198) );
  AND2_X1 U20021 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n18103), .ZN(
        P2_U3197) );
  AND2_X1 U20022 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n18103), .ZN(
        P2_U3196) );
  AND2_X1 U20023 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n18102), .ZN(
        P2_U3195) );
  AND2_X1 U20024 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n18102), .ZN(
        P2_U3194) );
  AND2_X1 U20025 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n18102), .ZN(
        P2_U3193) );
  AND2_X1 U20026 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n18102), .ZN(
        P2_U3192) );
  AND2_X1 U20027 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n18102), .ZN(
        P2_U3191) );
  AND2_X1 U20028 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n18102), .ZN(
        P2_U3190) );
  AND2_X1 U20029 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n18102), .ZN(
        P2_U3189) );
  AND2_X1 U20030 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n18102), .ZN(
        P2_U3188) );
  AND2_X1 U20031 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n18102), .ZN(
        P2_U3187) );
  AND2_X1 U20032 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n18103), .ZN(
        P2_U3186) );
  AND2_X1 U20033 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n18103), .ZN(
        P2_U3185) );
  AND2_X1 U20034 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n18103), .ZN(
        P2_U3184) );
  AND2_X1 U20035 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n18103), .ZN(
        P2_U3183) );
  AND2_X1 U20036 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n18103), .ZN(
        P2_U3182) );
  AND2_X1 U20037 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n18103), .ZN(
        P2_U3181) );
  AND2_X1 U20038 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n18103), .ZN(
        P2_U3180) );
  AND2_X1 U20039 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n18103), .ZN(
        P2_U3179) );
  NAND2_X1 U20040 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19531), .ZN(n19513) );
  AOI21_X1 U20041 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19247), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18106) );
  AOI221_X1 U20042 ( .B1(n19513), .B2(n18106), .C1(n18105), .C2(n18106), .A(
        n18104), .ZN(P2_U3178) );
  INV_X1 U20043 ( .A(n19523), .ZN(n18107) );
  OAI221_X1 U20044 ( .B1(n19540), .B2(n19522), .C1(n18107), .C2(n19522), .A(
        n20525), .ZN(n18217) );
  NOR2_X1 U20045 ( .A1(n18108), .A2(n18217), .ZN(P2_U3047) );
  AND2_X1 U20046 ( .A1(n18251), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U20047 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18112) );
  NOR4_X1 U20048 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18111) );
  NOR4_X1 U20049 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18110) );
  NOR4_X1 U20050 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18109) );
  NAND4_X1 U20051 ( .A1(n18112), .A2(n18111), .A3(n18110), .A4(n18109), .ZN(
        n18118) );
  NOR4_X1 U20052 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18116) );
  AOI211_X1 U20053 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18115) );
  NOR4_X1 U20054 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18114) );
  NOR4_X1 U20055 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18113) );
  NAND4_X1 U20056 ( .A1(n18116), .A2(n18115), .A3(n18114), .A4(n18113), .ZN(
        n18117) );
  NOR2_X1 U20057 ( .A1(n18118), .A2(n18117), .ZN(n18234) );
  INV_X1 U20058 ( .A(n18234), .ZN(n18232) );
  NOR2_X1 U20059 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18232), .ZN(n18226) );
  OR3_X1 U20060 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18231) );
  INV_X1 U20061 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U20062 ( .A1(n18226), .A2(n18231), .B1(n18232), .B2(n18119), .ZN(
        P2_U2821) );
  INV_X1 U20063 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18227) );
  INV_X1 U20064 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U20065 ( .A1(n18226), .A2(n18227), .B1(n18232), .B2(n18120), .ZN(
        P2_U2820) );
  INV_X1 U20066 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20792) );
  INV_X1 U20067 ( .A(n22410), .ZN(n18122) );
  INV_X1 U20068 ( .A(n22408), .ZN(n18121) );
  AOI21_X1 U20069 ( .B1(n20792), .B2(n18122), .A(n18121), .ZN(P1_U3464) );
  AND2_X1 U20070 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n18122), .ZN(P1_U3193) );
  AND2_X1 U20071 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n18122), .ZN(P1_U3192) );
  AND2_X1 U20072 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n18122), .ZN(P1_U3191) );
  AND2_X1 U20073 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n18122), .ZN(P1_U3190) );
  AND2_X1 U20074 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n18122), .ZN(P1_U3189) );
  AND2_X1 U20075 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n18122), .ZN(P1_U3188) );
  AND2_X1 U20076 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n18122), .ZN(P1_U3187) );
  AND2_X1 U20077 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n18122), .ZN(P1_U3186) );
  AND2_X1 U20078 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n18122), .ZN(
        P1_U3185) );
  AND2_X1 U20079 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n18122), .ZN(
        P1_U3184) );
  AND2_X1 U20080 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n18122), .ZN(
        P1_U3183) );
  AND2_X1 U20081 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n18122), .ZN(
        P1_U3182) );
  AND2_X1 U20082 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n18122), .ZN(
        P1_U3181) );
  AND2_X1 U20083 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n18122), .ZN(
        P1_U3180) );
  AND2_X1 U20084 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n18122), .ZN(
        P1_U3179) );
  AND2_X1 U20085 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n18122), .ZN(
        P1_U3178) );
  AND2_X1 U20086 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n18122), .ZN(
        P1_U3177) );
  AND2_X1 U20087 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n18122), .ZN(
        P1_U3176) );
  AND2_X1 U20088 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n18122), .ZN(
        P1_U3175) );
  AND2_X1 U20089 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n18122), .ZN(
        P1_U3174) );
  AND2_X1 U20090 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n18122), .ZN(
        P1_U3173) );
  AND2_X1 U20091 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n18122), .ZN(
        P1_U3172) );
  AND2_X1 U20092 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n18122), .ZN(
        P1_U3171) );
  AND2_X1 U20093 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n18122), .ZN(
        P1_U3170) );
  AND2_X1 U20094 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n18122), .ZN(
        P1_U3169) );
  AND2_X1 U20095 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n18122), .ZN(
        P1_U3168) );
  AND2_X1 U20096 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n18122), .ZN(
        P1_U3167) );
  AND2_X1 U20097 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n18122), .ZN(
        P1_U3166) );
  AND2_X1 U20098 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n18122), .ZN(
        P1_U3165) );
  AND2_X1 U20099 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n18122), .ZN(
        P1_U3164) );
  INV_X1 U20100 ( .A(n18151), .ZN(n18133) );
  INV_X1 U20101 ( .A(n18123), .ZN(n18124) );
  AOI22_X1 U20102 ( .A1(n18133), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18124), .B2(n18151), .ZN(n18142) );
  MUX2_X1 U20103 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18125), .S(
        n18151), .Z(n18139) );
  OAI211_X1 U20104 ( .C1(n18128), .C2(n18127), .A(n18126), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18130) );
  OAI21_X1 U20105 ( .B1(n18130), .B2(n22475), .A(n18129), .ZN(n18132) );
  NAND2_X1 U20106 ( .A1(n18130), .A2(n22475), .ZN(n18131) );
  OAI21_X1 U20107 ( .B1(n18133), .B2(n18132), .A(n18131), .ZN(n18134) );
  AOI222_X1 U20108 ( .A1(n18139), .A2(n18135), .B1(n18139), .B2(n18134), .C1(
        n18135), .C2(n18134), .ZN(n18136) );
  OR2_X1 U20109 ( .A1(n18136), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18137) );
  AOI221_X1 U20110 ( .B1(n18142), .B2(n18137), .C1(n18136), .C2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18153) );
  NAND2_X1 U20111 ( .A1(n18138), .A2(n22251), .ZN(n18149) );
  INV_X1 U20112 ( .A(n18139), .ZN(n18143) );
  OAI21_X1 U20113 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n18140), .ZN(n18141) );
  OAI21_X1 U20114 ( .B1(n18143), .B2(n18142), .A(n18141), .ZN(n18144) );
  OR2_X1 U20115 ( .A1(n18145), .A2(n18144), .ZN(n18146) );
  NOR2_X1 U20116 ( .A1(n18147), .A2(n18146), .ZN(n18148) );
  OAI211_X1 U20117 ( .C1(n18151), .C2(n18150), .A(n18149), .B(n18148), .ZN(
        n18152) );
  NOR2_X1 U20118 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22489), .ZN(n18157) );
  INV_X1 U20119 ( .A(n13211), .ZN(n22132) );
  OAI221_X1 U20120 ( .B1(n22390), .B2(n18157), .C1(n22390), .C2(n22389), .A(
        n11491), .ZN(n18163) );
  AOI221_X1 U20121 ( .B1(n22396), .B2(n18164), .C1(n22398), .C2(n18164), .A(
        n18163), .ZN(n22399) );
  NOR2_X1 U20122 ( .A1(n22399), .A2(n22396), .ZN(n22397) );
  NOR2_X1 U20123 ( .A1(n22129), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n18161) );
  INV_X1 U20124 ( .A(n18161), .ZN(n18158) );
  OAI211_X1 U20125 ( .C1(n18159), .C2(n15600), .A(n22397), .B(n18158), .ZN(
        n22403) );
  NOR2_X1 U20126 ( .A1(n22396), .A2(n18164), .ZN(n22391) );
  AOI21_X1 U20127 ( .B1(n18161), .B2(n22391), .A(n18160), .ZN(n18162) );
  OAI221_X1 U20128 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n22403), .C1(n18164), 
        .C2(n18163), .A(n18162), .ZN(P1_U3162) );
  NOR2_X1 U20129 ( .A1(n18166), .A2(n18165), .ZN(P1_U3032) );
  AND2_X1 U20130 ( .A1(n20711), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U20131 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18167) );
  OAI22_X1 U20132 ( .A1(n18168), .A2(n18167), .B1(n19512), .B2(n19521), .ZN(
        P2_U2816) );
  AOI22_X1 U20133 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18174), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19360), .ZN(n18173) );
  AOI222_X1 U20134 ( .A1(n18171), .A2(n18200), .B1(n18199), .B2(n18170), .C1(
        n18169), .C2(n18198), .ZN(n18172) );
  OAI211_X1 U20135 ( .C1(n18181), .C2(n19278), .A(n18173), .B(n18172), .ZN(
        P2_U3010) );
  AOI22_X1 U20136 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18174), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19360), .ZN(n18180) );
  NOR2_X1 U20137 ( .A1(n18175), .A2(n18185), .ZN(n18178) );
  OAI22_X1 U20138 ( .A1(n18176), .A2(n18184), .B1(n18190), .B2(n19292), .ZN(
        n18177) );
  AOI21_X1 U20139 ( .B1(n18178), .B2(n18054), .A(n18177), .ZN(n18179) );
  OAI211_X1 U20140 ( .C1(n18181), .C2(n19291), .A(n18180), .B(n18179), .ZN(
        P2_U3008) );
  INV_X1 U20141 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19310) );
  OAI22_X1 U20142 ( .A1(n19310), .A2(n18204), .B1(n18181), .B2(n19304), .ZN(
        n18182) );
  AOI21_X1 U20143 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(n19360), .A(n18182), .ZN(
        n18189) );
  OAI22_X1 U20144 ( .A1(n18186), .A2(n18185), .B1(n18184), .B2(n18183), .ZN(
        n18187) );
  INV_X1 U20145 ( .A(n18187), .ZN(n18188) );
  OAI211_X1 U20146 ( .C1(n18190), .C2(n19305), .A(n18189), .B(n18188), .ZN(
        P2_U3006) );
  AOI22_X1 U20147 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19360), .B1(n18196), 
        .B2(n19316), .ZN(n18194) );
  AOI222_X1 U20148 ( .A1(n18192), .A2(n18200), .B1(n18199), .B2(n19318), .C1(
        n18198), .C2(n18191), .ZN(n18193) );
  OAI211_X1 U20149 ( .C1(n19313), .C2(n18204), .A(n18194), .B(n18193), .ZN(
        P2_U3004) );
  AOI22_X1 U20150 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19360), .B1(n18196), 
        .B2(n18195), .ZN(n18203) );
  AOI222_X1 U20151 ( .A1(n18201), .A2(n18200), .B1(n18199), .B2(n19336), .C1(
        n18198), .C2(n18197), .ZN(n18202) );
  OAI211_X1 U20152 ( .C1(n11338), .C2(n18204), .A(n18203), .B(n18202), .ZN(
        P2_U3000) );
  INV_X1 U20153 ( .A(n18217), .ZN(n18225) );
  OAI22_X1 U20154 ( .A1(n20519), .A2(n19245), .B1(n18206), .B2(n18205), .ZN(
        n18207) );
  AOI21_X1 U20155 ( .B1(n20122), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n18207), 
        .ZN(n18208) );
  OAI22_X1 U20156 ( .A1(n20122), .A2(n18217), .B1(n18225), .B2(n18208), .ZN(
        P2_U3605) );
  NAND2_X1 U20157 ( .A1(n18209), .A2(n20167), .ZN(n18213) );
  NAND2_X1 U20158 ( .A1(n19512), .A2(n18213), .ZN(n18219) );
  INV_X1 U20159 ( .A(n18209), .ZN(n18210) );
  NAND2_X1 U20160 ( .A1(n20409), .A2(n18210), .ZN(n20148) );
  INV_X1 U20161 ( .A(n20148), .ZN(n18211) );
  AOI222_X1 U20162 ( .A1(n20408), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n18220), 
        .B2(n18219), .C1(n20167), .C2(n18211), .ZN(n18212) );
  AOI22_X1 U20163 ( .A1(n18225), .A2(n20146), .B1(n18212), .B2(n18217), .ZN(
        P2_U3603) );
  AND2_X1 U20164 ( .A1(n18213), .A2(n19512), .ZN(n18215) );
  OAI22_X1 U20165 ( .A1(n18215), .A2(n18214), .B1(n22411), .B2(n18213), .ZN(
        n18216) );
  AOI21_X1 U20166 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20458), .A(n18216), 
        .ZN(n18218) );
  AOI22_X1 U20167 ( .A1(n18225), .A2(n20150), .B1(n18218), .B2(n18217), .ZN(
        P2_U3604) );
  INV_X1 U20168 ( .A(n20262), .ZN(n20149) );
  AOI22_X1 U20169 ( .A1(n20149), .A2(n18219), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20358), .ZN(n18224) );
  INV_X1 U20170 ( .A(n20133), .ZN(n18221) );
  NAND2_X1 U20171 ( .A1(n18221), .A2(n20255), .ZN(n20115) );
  AOI211_X1 U20172 ( .C1(n20092), .C2(n20115), .A(n20192), .B(n22411), .ZN(
        n18222) );
  NOR2_X1 U20173 ( .A1(n18225), .A2(n18222), .ZN(n18223) );
  AOI22_X1 U20174 ( .A1(n20145), .A2(n18225), .B1(n18224), .B2(n18223), .ZN(
        P2_U3602) );
  INV_X1 U20175 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22413) );
  NAND2_X1 U20176 ( .A1(n18226), .A2(n22413), .ZN(n18230) );
  INV_X1 U20177 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n18273) );
  OAI21_X1 U20178 ( .B1(n18273), .B2(n18227), .A(n18234), .ZN(n18228) );
  OAI21_X1 U20179 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18234), .A(n18228), 
        .ZN(n18229) );
  OAI221_X1 U20180 ( .B1(n18230), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18230), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18229), .ZN(P2_U2822) );
  INV_X1 U20181 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18233) );
  OAI221_X1 U20182 ( .B1(n18234), .B2(n18233), .C1(n18232), .C2(n18231), .A(
        n18230), .ZN(P2_U2823) );
  OAI22_X1 U20183 ( .A1(n18316), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n18311), .ZN(n18235) );
  INV_X1 U20184 ( .A(n18235), .ZN(P2_U3611) );
  INV_X1 U20185 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n18236) );
  AOI22_X1 U20186 ( .A1(n18311), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n18236), 
        .B2(n18316), .ZN(P2_U3608) );
  AOI21_X1 U20187 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n22414), .ZN(n18237) );
  INV_X1 U20188 ( .A(n18237), .ZN(P2_U2815) );
  INV_X1 U20189 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n20514) );
  AOI22_X1 U20190 ( .A1(n18266), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18239) );
  OAI21_X1 U20191 ( .B1(n20514), .B2(n18268), .A(n18239), .ZN(P2_U2951) );
  INV_X1 U20192 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U20193 ( .A1(n18266), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18240) );
  OAI21_X1 U20194 ( .B1(n18241), .B2(n18268), .A(n18240), .ZN(P2_U2950) );
  INV_X1 U20195 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18243) );
  AOI22_X1 U20196 ( .A1(n18266), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18242) );
  OAI21_X1 U20197 ( .B1(n18243), .B2(n18268), .A(n18242), .ZN(P2_U2949) );
  INV_X1 U20198 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18245) );
  AOI22_X1 U20199 ( .A1(n18257), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18244) );
  OAI21_X1 U20200 ( .B1(n18245), .B2(n18268), .A(n18244), .ZN(P2_U2948) );
  INV_X1 U20201 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U20202 ( .A1(n18266), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18246) );
  OAI21_X1 U20203 ( .B1(n18247), .B2(n18268), .A(n18246), .ZN(P2_U2947) );
  INV_X1 U20204 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18249) );
  AOI22_X1 U20205 ( .A1(n18257), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18248) );
  OAI21_X1 U20206 ( .B1(n18249), .B2(n18268), .A(n18248), .ZN(P2_U2946) );
  INV_X1 U20207 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U20208 ( .A1(n18257), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18250) );
  OAI21_X1 U20209 ( .B1(n20208), .B2(n18268), .A(n18250), .ZN(P2_U2945) );
  INV_X1 U20210 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U20211 ( .A1(n18257), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18251), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18252) );
  OAI21_X1 U20212 ( .B1(n18253), .B2(n18268), .A(n18252), .ZN(P2_U2944) );
  INV_X1 U20213 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20033) );
  AOI22_X1 U20214 ( .A1(n18257), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18254) );
  OAI21_X1 U20215 ( .B1(n20033), .B2(n18268), .A(n18254), .ZN(P2_U2943) );
  INV_X1 U20216 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U20217 ( .A1(n18266), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18255) );
  OAI21_X1 U20218 ( .B1(n18256), .B2(n18268), .A(n18255), .ZN(P2_U2942) );
  INV_X1 U20219 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20027) );
  AOI22_X1 U20220 ( .A1(n18257), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18258) );
  OAI21_X1 U20221 ( .B1(n20027), .B2(n18268), .A(n18258), .ZN(P2_U2941) );
  AOI22_X1 U20222 ( .A1(n18266), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18259) );
  OAI21_X1 U20223 ( .B1(n18260), .B2(n18268), .A(n18259), .ZN(P2_U2940) );
  INV_X1 U20224 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U20225 ( .A1(n18266), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18261) );
  OAI21_X1 U20226 ( .B1(n20021), .B2(n18268), .A(n18261), .ZN(P2_U2939) );
  INV_X1 U20227 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18263) );
  AOI22_X1 U20228 ( .A1(n18266), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18262) );
  OAI21_X1 U20229 ( .B1(n18263), .B2(n18268), .A(n18262), .ZN(P2_U2938) );
  INV_X1 U20230 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U20231 ( .A1(n18266), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18264) );
  OAI21_X1 U20232 ( .B1(n20015), .B2(n18268), .A(n18264), .ZN(P2_U2937) );
  AOI22_X1 U20233 ( .A1(n18266), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18265), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18267) );
  OAI21_X1 U20234 ( .B1(n20012), .B2(n18268), .A(n18267), .ZN(P2_U2936) );
  AOI21_X1 U20235 ( .B1(n18270), .B2(n18269), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18271) );
  AOI21_X1 U20236 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n18311), .A(n18271), 
        .ZN(P2_U2817) );
  INV_X1 U20237 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n18275) );
  NOR2_X1 U20238 ( .A1(n18272), .A2(n18316), .ZN(n22435) );
  OAI222_X1 U20239 ( .A1(n18313), .A2(n18275), .B1(n18274), .B2(n18311), .C1(
        n18273), .C2(n18306), .ZN(P2_U3212) );
  INV_X1 U20240 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n18276) );
  OAI222_X1 U20241 ( .A1(n18308), .A2(n18277), .B1(n18276), .B2(n18311), .C1(
        n18275), .C2(n18306), .ZN(P2_U3213) );
  INV_X1 U20242 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n18279) );
  INV_X1 U20243 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n18278) );
  OAI222_X1 U20244 ( .A1(n18308), .A2(n18279), .B1(n18278), .B2(n18311), .C1(
        n18277), .C2(n18306), .ZN(P2_U3214) );
  INV_X1 U20245 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n18280) );
  OAI222_X1 U20246 ( .A1(n18308), .A2(n18281), .B1(n18280), .B2(n18311), .C1(
        n18279), .C2(n18306), .ZN(P2_U3215) );
  INV_X1 U20247 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n18282) );
  OAI222_X1 U20248 ( .A1(n18308), .A2(n18283), .B1(n18282), .B2(n18311), .C1(
        n18281), .C2(n18306), .ZN(P2_U3216) );
  INV_X1 U20249 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n18284) );
  OAI222_X1 U20250 ( .A1(n18308), .A2(n18285), .B1(n18284), .B2(n18311), .C1(
        n18283), .C2(n18306), .ZN(P2_U3217) );
  INV_X1 U20251 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n18287) );
  INV_X1 U20252 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n18286) );
  OAI222_X1 U20253 ( .A1(n18308), .A2(n18287), .B1(n18286), .B2(n18311), .C1(
        n18285), .C2(n18306), .ZN(P2_U3218) );
  INV_X1 U20254 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20651) );
  OAI222_X1 U20255 ( .A1(n18313), .A2(n18288), .B1(n20651), .B2(n18311), .C1(
        n18287), .C2(n18306), .ZN(P2_U3219) );
  INV_X1 U20256 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20653) );
  INV_X1 U20257 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n18290) );
  OAI222_X1 U20258 ( .A1(n18306), .A2(n18288), .B1(n20653), .B2(n18311), .C1(
        n18290), .C2(n18308), .ZN(P2_U3220) );
  INV_X1 U20259 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n18289) );
  OAI222_X1 U20260 ( .A1(n18306), .A2(n18290), .B1(n18289), .B2(n18311), .C1(
        n18292), .C2(n18308), .ZN(P2_U3221) );
  INV_X1 U20261 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n18291) );
  INV_X1 U20262 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n18293) );
  OAI222_X1 U20263 ( .A1(n18306), .A2(n18292), .B1(n18291), .B2(n18311), .C1(
        n18293), .C2(n18308), .ZN(P2_U3222) );
  INV_X1 U20264 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20657) );
  OAI222_X1 U20265 ( .A1(n18306), .A2(n18293), .B1(n20657), .B2(n18311), .C1(
        n18294), .C2(n18308), .ZN(P2_U3223) );
  INV_X1 U20266 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20659) );
  OAI222_X1 U20267 ( .A1(n18306), .A2(n18294), .B1(n20659), .B2(n18311), .C1(
        n17924), .C2(n18308), .ZN(P2_U3224) );
  INV_X1 U20268 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20661) );
  OAI222_X1 U20269 ( .A1(n18306), .A2(n17924), .B1(n20661), .B2(n18311), .C1(
        n18295), .C2(n18308), .ZN(P2_U3225) );
  INV_X1 U20270 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20663) );
  INV_X1 U20271 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19345) );
  OAI222_X1 U20272 ( .A1(n18306), .A2(n18295), .B1(n20663), .B2(n18311), .C1(
        n19345), .C2(n18308), .ZN(P2_U3226) );
  INV_X1 U20273 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20665) );
  INV_X1 U20274 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n18296) );
  OAI222_X1 U20275 ( .A1(n18306), .A2(n19345), .B1(n20665), .B2(n18311), .C1(
        n18296), .C2(n18308), .ZN(P2_U3227) );
  INV_X1 U20276 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20667) );
  OAI222_X1 U20277 ( .A1(n18306), .A2(n18296), .B1(n20667), .B2(n18311), .C1(
        n19372), .C2(n18308), .ZN(P2_U3228) );
  INV_X1 U20278 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18297) );
  INV_X1 U20279 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20669) );
  OAI222_X1 U20280 ( .A1(n18313), .A2(n18297), .B1(n20669), .B2(n18311), .C1(
        n19372), .C2(n18306), .ZN(P2_U3229) );
  INV_X1 U20281 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20671) );
  OAI222_X1 U20282 ( .A1(n18306), .A2(n18297), .B1(n20671), .B2(n18311), .C1(
        n18298), .C2(n18308), .ZN(P2_U3230) );
  INV_X1 U20283 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n18299) );
  INV_X1 U20284 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20673) );
  OAI222_X1 U20285 ( .A1(n18313), .A2(n18299), .B1(n20673), .B2(n18311), .C1(
        n18298), .C2(n18306), .ZN(P2_U3231) );
  INV_X1 U20286 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20675) );
  OAI222_X1 U20287 ( .A1(n18313), .A2(n18300), .B1(n20675), .B2(n18311), .C1(
        n18299), .C2(n18306), .ZN(P2_U3232) );
  INV_X1 U20288 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20677) );
  OAI222_X1 U20289 ( .A1(n18313), .A2(n18301), .B1(n20677), .B2(n18311), .C1(
        n18300), .C2(n18306), .ZN(P2_U3233) );
  INV_X1 U20290 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20679) );
  OAI222_X1 U20291 ( .A1(n18313), .A2(n18302), .B1(n20679), .B2(n18311), .C1(
        n18301), .C2(n18306), .ZN(P2_U3234) );
  INV_X1 U20292 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20681) );
  OAI222_X1 U20293 ( .A1(n18313), .A2(n18303), .B1(n20681), .B2(n18311), .C1(
        n18302), .C2(n18306), .ZN(P2_U3235) );
  INV_X1 U20294 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20683) );
  INV_X1 U20295 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n18304) );
  OAI222_X1 U20296 ( .A1(n18306), .A2(n18303), .B1(n20683), .B2(n18311), .C1(
        n18304), .C2(n18308), .ZN(P2_U3236) );
  INV_X1 U20297 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20685) );
  OAI222_X1 U20298 ( .A1(n18313), .A2(n18305), .B1(n20685), .B2(n18311), .C1(
        n18304), .C2(n18306), .ZN(P2_U3237) );
  INV_X1 U20299 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20687) );
  OAI222_X1 U20300 ( .A1(n18306), .A2(n18305), .B1(n20687), .B2(n18311), .C1(
        n18307), .C2(n18308), .ZN(P2_U3238) );
  INV_X1 U20301 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20689) );
  OAI222_X1 U20302 ( .A1(n18313), .A2(n18309), .B1(n20689), .B2(n18311), .C1(
        n18307), .C2(n18306), .ZN(P2_U3239) );
  INV_X1 U20303 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20691) );
  INV_X1 U20304 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n18310) );
  OAI222_X1 U20305 ( .A1(n18306), .A2(n18309), .B1(n20691), .B2(n18311), .C1(
        n18310), .C2(n18308), .ZN(P2_U3240) );
  INV_X1 U20306 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18312) );
  INV_X1 U20307 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20694) );
  OAI222_X1 U20308 ( .A1(n18313), .A2(n18312), .B1(n20694), .B2(n18311), .C1(
        n18310), .C2(n18306), .ZN(P2_U3241) );
  OAI22_X1 U20309 ( .A1(n18316), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n18311), .ZN(n18314) );
  INV_X1 U20310 ( .A(n18314), .ZN(P2_U3588) );
  OAI22_X1 U20311 ( .A1(n18316), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n18311), .ZN(n18315) );
  INV_X1 U20312 ( .A(n18315), .ZN(P2_U3587) );
  MUX2_X1 U20313 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n18316), .Z(P2_U3586) );
  OAI22_X1 U20314 ( .A1(n18316), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n18311), .ZN(n18317) );
  INV_X1 U20315 ( .A(n18317), .ZN(P2_U3585) );
  NOR2_X1 U20316 ( .A1(n21521), .A2(n18318), .ZN(n18320) );
  NAND2_X1 U20317 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18688) );
  INV_X1 U20318 ( .A(n18688), .ZN(n18328) );
  AND2_X1 U20319 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n18328), .ZN(n18322) );
  INV_X1 U20320 ( .A(n11217), .ZN(n18692) );
  INV_X1 U20321 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n21035) );
  NAND3_X1 U20322 ( .A1(n18687), .A2(n11217), .A3(n18322), .ZN(n18325) );
  NOR2_X1 U20323 ( .A1(n21035), .A2(n18325), .ZN(n18327) );
  AOI21_X1 U20324 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18689), .A(n18327), .ZN(
        n18324) );
  OAI22_X1 U20325 ( .A1(n18351), .A2(n18324), .B1(n18323), .B2(n18689), .ZN(
        P3_U2699) );
  INV_X1 U20326 ( .A(n18325), .ZN(n18329) );
  AOI21_X1 U20327 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18689), .A(n18329), .ZN(
        n18326) );
  OAI22_X1 U20328 ( .A1(n18327), .A2(n18326), .B1(n18535), .B2(n18689), .ZN(
        P3_U2700) );
  INV_X1 U20329 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18331) );
  AOI221_X1 U20330 ( .B1(n18328), .B2(n11217), .C1(n21521), .C2(n11217), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18330) );
  AOI211_X1 U20331 ( .C1(n18693), .C2(n18331), .A(n18330), .B(n18329), .ZN(
        P3_U2701) );
  AOI22_X1 U20332 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U20333 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18334) );
  AOI22_X1 U20334 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18333) );
  AOI22_X1 U20335 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18332) );
  NAND4_X1 U20336 ( .A1(n18335), .A2(n18334), .A3(n18333), .A4(n18332), .ZN(
        n18341) );
  AOI22_X1 U20337 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U20338 ( .A1(n16134), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U20339 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18337) );
  AOI22_X1 U20340 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18336) );
  NAND4_X1 U20341 ( .A1(n18339), .A2(n18338), .A3(n18337), .A4(n18336), .ZN(
        n18340) );
  NOR2_X1 U20342 ( .A1(n18341), .A2(n18340), .ZN(n21591) );
  NAND4_X1 U20343 ( .A1(n18687), .A2(P3_EBX_REG_7__SCAN_IN), .A3(
        P3_EBX_REG_6__SCAN_IN), .A4(n18353), .ZN(n18342) );
  NOR2_X1 U20344 ( .A1(n21110), .A2(n18342), .ZN(n18450) );
  INV_X1 U20345 ( .A(n18342), .ZN(n18346) );
  AOI21_X1 U20346 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n18689), .A(n18346), .ZN(
        n18343) );
  OAI22_X1 U20347 ( .A1(n21591), .A2(n18689), .B1(n18450), .B2(n18343), .ZN(
        P3_U2695) );
  NAND2_X1 U20348 ( .A1(n18687), .A2(n18353), .ZN(n18347) );
  NOR2_X1 U20349 ( .A1(n21080), .A2(n18347), .ZN(n18344) );
  AOI21_X1 U20350 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18689), .A(n18344), .ZN(
        n18345) );
  OAI22_X1 U20351 ( .A1(n18346), .A2(n18345), .B1(n18710), .B2(n18689), .ZN(
        P3_U2696) );
  AOI21_X1 U20352 ( .B1(n21080), .B2(n18347), .A(n18364), .ZN(n18348) );
  INV_X1 U20353 ( .A(n18348), .ZN(n18349) );
  AOI22_X1 U20354 ( .A1(n18693), .A2(n18350), .B1(n18349), .B2(n18689), .ZN(
        P3_U2697) );
  OAI21_X1 U20355 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18351), .A(n18689), .ZN(
        n18352) );
  OAI22_X1 U20356 ( .A1(n18353), .A2(n18352), .B1(n18546), .B2(n18689), .ZN(
        P3_U2698) );
  AOI22_X1 U20357 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18357) );
  AOI22_X1 U20358 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18524), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U20359 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18355) );
  AOI22_X1 U20360 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18354) );
  NAND4_X1 U20361 ( .A1(n18357), .A2(n18356), .A3(n18355), .A4(n18354), .ZN(
        n18363) );
  AOI22_X1 U20362 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18475), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18361) );
  AOI22_X1 U20363 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18360) );
  AOI22_X1 U20364 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U20365 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18358) );
  NAND4_X1 U20366 ( .A1(n18361), .A2(n18360), .A3(n18359), .A4(n18358), .ZN(
        n18362) );
  NOR2_X1 U20367 ( .A1(n18363), .A2(n18362), .ZN(n21574) );
  INV_X1 U20368 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21207) );
  INV_X1 U20369 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n21152) );
  NAND4_X1 U20370 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(n18420), .ZN(n18377) );
  NOR2_X2 U20371 ( .A1(n21207), .A2(n18377), .ZN(n18464) );
  NOR2_X1 U20372 ( .A1(n18693), .A2(n18464), .ZN(n18378) );
  OAI222_X1 U20373 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18687), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n18464), .C1(n18378), .C2(n21218), .ZN(
        n18365) );
  OAI21_X1 U20374 ( .B1(n21574), .B2(n18689), .A(n18365), .ZN(P3_U2687) );
  AOI22_X1 U20375 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18370) );
  AOI22_X1 U20376 ( .A1(n18366), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U20377 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18368) );
  AOI22_X1 U20378 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18367) );
  NAND4_X1 U20379 ( .A1(n18370), .A2(n18369), .A3(n18368), .A4(n18367), .ZN(
        n18376) );
  AOI22_X1 U20380 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14067), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18374) );
  AOI22_X1 U20381 ( .A1(n18621), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U20382 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n21034), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18372) );
  AOI22_X1 U20383 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18371) );
  NAND4_X1 U20384 ( .A1(n18374), .A2(n18373), .A3(n18372), .A4(n18371), .ZN(
        n18375) );
  NOR2_X1 U20385 ( .A1(n18376), .A2(n18375), .ZN(n21584) );
  INV_X1 U20386 ( .A(n18377), .ZN(n18379) );
  OAI21_X1 U20387 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18379), .A(n18378), .ZN(
        n18380) );
  OAI21_X1 U20388 ( .B1(n21584), .B2(n18689), .A(n18380), .ZN(P3_U2688) );
  AOI22_X1 U20389 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18384) );
  AOI22_X1 U20390 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18383) );
  AOI22_X1 U20391 ( .A1(n21034), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18382) );
  AOI22_X1 U20392 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18381) );
  NAND4_X1 U20393 ( .A1(n18384), .A2(n18383), .A3(n18382), .A4(n18381), .ZN(
        n18390) );
  AOI22_X1 U20394 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18388) );
  AOI22_X1 U20395 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18387) );
  AOI22_X1 U20396 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18386) );
  AOI22_X1 U20397 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18385) );
  NAND4_X1 U20398 ( .A1(n18388), .A2(n18387), .A3(n18386), .A4(n18385), .ZN(
        n18389) );
  NOR2_X1 U20399 ( .A1(n18390), .A2(n18389), .ZN(n21434) );
  NAND2_X1 U20400 ( .A1(n18687), .A2(n18420), .ZN(n18421) );
  NOR2_X1 U20401 ( .A1(n21162), .A2(n18421), .ZN(n18391) );
  NAND2_X1 U20402 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18391), .ZN(n18404) );
  OAI211_X1 U20403 ( .C1(n18391), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18689), .B(
        n18404), .ZN(n18392) );
  OAI21_X1 U20404 ( .B1(n21434), .B2(n18689), .A(n18392), .ZN(P3_U2690) );
  AOI22_X1 U20405 ( .A1(n16134), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14067), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18396) );
  AOI22_X1 U20406 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18395) );
  AOI22_X1 U20407 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U20408 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18393) );
  NAND4_X1 U20409 ( .A1(n18396), .A2(n18395), .A3(n18394), .A4(n18393), .ZN(
        n18403) );
  AOI22_X1 U20410 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18401) );
  AOI22_X1 U20411 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18397), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18400) );
  AOI22_X1 U20412 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18399) );
  AOI22_X1 U20413 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18398) );
  NAND4_X1 U20414 ( .A1(n18401), .A2(n18400), .A3(n18399), .A4(n18398), .ZN(
        n18402) );
  NOR2_X1 U20415 ( .A1(n18403), .A2(n18402), .ZN(n21578) );
  NAND3_X1 U20416 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n18406) );
  OAI21_X1 U20417 ( .B1(n18693), .B2(n21192), .A(n18404), .ZN(n18405) );
  OAI21_X1 U20418 ( .B1(n18421), .B2(n18406), .A(n18405), .ZN(n18407) );
  OAI21_X1 U20419 ( .B1(n21578), .B2(n18689), .A(n18407), .ZN(P3_U2689) );
  AOI22_X1 U20420 ( .A1(n18713), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18413) );
  AOI22_X1 U20421 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U20422 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18409), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18411) );
  AOI22_X1 U20423 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18410) );
  NAND4_X1 U20424 ( .A1(n18413), .A2(n18412), .A3(n18411), .A4(n18410), .ZN(
        n18419) );
  AOI22_X1 U20425 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18417) );
  AOI22_X1 U20426 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18416) );
  AOI22_X1 U20427 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18415) );
  AOI22_X1 U20428 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18414) );
  NAND4_X1 U20429 ( .A1(n18417), .A2(n18416), .A3(n18415), .A4(n18414), .ZN(
        n18418) );
  NOR2_X1 U20430 ( .A1(n18419), .A2(n18418), .ZN(n21439) );
  NOR2_X1 U20431 ( .A1(n18693), .A2(n18420), .ZN(n18435) );
  INV_X1 U20432 ( .A(n18421), .ZN(n18422) );
  AOI22_X1 U20433 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18435), .B1(n18422), 
        .B2(n21162), .ZN(n18423) );
  OAI21_X1 U20434 ( .B1(n21439), .B2(n18689), .A(n18423), .ZN(P3_U2691) );
  AOI22_X1 U20435 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18428) );
  AOI22_X1 U20436 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18427) );
  AOI22_X1 U20437 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18426) );
  AOI22_X1 U20438 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18425) );
  NAND4_X1 U20439 ( .A1(n18428), .A2(n18427), .A3(n18426), .A4(n18425), .ZN(
        n18434) );
  AOI22_X1 U20440 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18432) );
  AOI22_X1 U20441 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18431) );
  AOI22_X1 U20442 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U20443 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18429) );
  NAND4_X1 U20444 ( .A1(n18432), .A2(n18431), .A3(n18430), .A4(n18429), .ZN(
        n18433) );
  NOR2_X1 U20445 ( .A1(n18434), .A2(n18433), .ZN(n21444) );
  INV_X1 U20446 ( .A(n18448), .ZN(n18436) );
  OAI21_X1 U20447 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18436), .A(n18435), .ZN(
        n18437) );
  OAI21_X1 U20448 ( .B1(n21444), .B2(n18689), .A(n18437), .ZN(P3_U2692) );
  AOI22_X1 U20449 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18441) );
  AOI22_X1 U20450 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18440) );
  AOI22_X1 U20451 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18439) );
  AOI22_X1 U20452 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18438) );
  NAND4_X1 U20453 ( .A1(n18441), .A2(n18440), .A3(n18439), .A4(n18438), .ZN(
        n18447) );
  AOI22_X1 U20454 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18445) );
  AOI22_X1 U20455 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18408), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18444) );
  AOI22_X1 U20456 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18443) );
  AOI22_X1 U20457 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18442) );
  NAND4_X1 U20458 ( .A1(n18445), .A2(n18444), .A3(n18443), .A4(n18442), .ZN(
        n18446) );
  NOR2_X1 U20459 ( .A1(n18447), .A2(n18446), .ZN(n21451) );
  OAI21_X1 U20460 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18463), .A(n18448), .ZN(
        n18449) );
  AOI22_X1 U20461 ( .A1(n18693), .A2(n21451), .B1(n18449), .B2(n18689), .ZN(
        P3_U2693) );
  AOI21_X1 U20462 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18689), .A(n18450), .ZN(
        n18462) );
  AOI22_X1 U20463 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18524), .B1(
        n18548), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U20464 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11165), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18453) );
  AOI22_X1 U20465 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18673), .ZN(n18452) );
  AOI22_X1 U20466 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18674), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n21637), .ZN(n18451) );
  NAND4_X1 U20467 ( .A1(n18454), .A2(n18453), .A3(n18452), .A4(n18451), .ZN(
        n18461) );
  AOI22_X1 U20468 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11159), .ZN(n18459) );
  AOI22_X1 U20469 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18714), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U20470 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18457) );
  AOI22_X1 U20471 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18716), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18456) );
  NAND4_X1 U20472 ( .A1(n18459), .A2(n18458), .A3(n18457), .A4(n18456), .ZN(
        n18460) );
  NOR2_X1 U20473 ( .A1(n18461), .A2(n18460), .ZN(n21452) );
  OAI22_X1 U20474 ( .A1(n18463), .A2(n18462), .B1(n21452), .B2(n18689), .ZN(
        P3_U2694) );
  INV_X1 U20475 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21403) );
  INV_X1 U20476 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n21309) );
  INV_X1 U20477 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21256) );
  INV_X1 U20478 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21237) );
  NAND2_X1 U20479 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18584), .ZN(n18583) );
  NAND4_X1 U20480 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n18465)
         );
  NOR4_X1 U20481 ( .A1(n21309), .A2(n21297), .A3(n18583), .A4(n18465), .ZN(
        n18466) );
  NAND4_X1 U20482 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n18466), .ZN(n18469) );
  NOR2_X1 U20483 ( .A1(n21403), .A2(n18469), .ZN(n18572) );
  NAND2_X1 U20484 ( .A1(n18689), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18468) );
  NAND2_X1 U20485 ( .A1(n18572), .A2(n18687), .ZN(n18467) );
  OAI22_X1 U20486 ( .A1(n18572), .A2(n18468), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18467), .ZN(P3_U2672) );
  NAND2_X1 U20487 ( .A1(n21403), .A2(n18469), .ZN(n18470) );
  NAND2_X1 U20488 ( .A1(n18470), .A2(n18689), .ZN(n18571) );
  AOI22_X1 U20489 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18474) );
  AOI22_X1 U20490 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18473) );
  AOI22_X1 U20491 ( .A1(n18713), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18472) );
  AOI22_X1 U20492 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18471) );
  NAND4_X1 U20493 ( .A1(n18474), .A2(n18473), .A3(n18472), .A4(n18471), .ZN(
        n18481) );
  AOI22_X1 U20494 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18479) );
  AOI22_X1 U20495 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18478) );
  INV_X1 U20496 ( .A(n18547), .ZN(n18715) );
  AOI22_X1 U20497 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18477) );
  BUF_X1 U20498 ( .A(n18475), .Z(n18706) );
  AOI22_X1 U20499 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18476) );
  NAND4_X1 U20500 ( .A1(n18479), .A2(n18478), .A3(n18477), .A4(n18476), .ZN(
        n18480) );
  NOR2_X1 U20501 ( .A1(n18481), .A2(n18480), .ZN(n18590) );
  AOI22_X1 U20502 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18485) );
  AOI22_X1 U20503 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18484) );
  AOI22_X1 U20504 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18483) );
  AOI22_X1 U20505 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18482) );
  NAND4_X1 U20506 ( .A1(n18485), .A2(n18484), .A3(n18483), .A4(n18482), .ZN(
        n18491) );
  AOI22_X1 U20507 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18707), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18489) );
  AOI22_X1 U20508 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U20509 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U20510 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18486) );
  NAND4_X1 U20511 ( .A1(n18489), .A2(n18488), .A3(n18487), .A4(n18486), .ZN(
        n18490) );
  NOR2_X1 U20512 ( .A1(n18491), .A2(n18490), .ZN(n18587) );
  AOI22_X1 U20513 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18495) );
  AOI22_X1 U20514 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18494) );
  AOI22_X1 U20515 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18493) );
  AOI22_X1 U20516 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18492) );
  NAND4_X1 U20517 ( .A1(n18495), .A2(n18494), .A3(n18493), .A4(n18492), .ZN(
        n18501) );
  AOI22_X1 U20518 ( .A1(n18621), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18499) );
  AOI22_X1 U20519 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18498) );
  AOI22_X1 U20520 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18497) );
  AOI22_X1 U20521 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18496) );
  NAND4_X1 U20522 ( .A1(n18499), .A2(n18498), .A3(n18497), .A4(n18496), .ZN(
        n18500) );
  NOR2_X1 U20523 ( .A1(n18501), .A2(n18500), .ZN(n18603) );
  AOI22_X1 U20524 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18505) );
  AOI22_X1 U20525 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18504) );
  AOI22_X1 U20526 ( .A1(n18621), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18503) );
  AOI22_X1 U20527 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18502) );
  NAND4_X1 U20528 ( .A1(n18505), .A2(n18504), .A3(n18503), .A4(n18502), .ZN(
        n18511) );
  AOI22_X1 U20529 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U20530 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18622), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18508) );
  AOI22_X1 U20531 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18507) );
  AOI22_X1 U20532 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18506) );
  NAND4_X1 U20533 ( .A1(n18509), .A2(n18508), .A3(n18507), .A4(n18506), .ZN(
        n18510) );
  NOR2_X1 U20534 ( .A1(n18511), .A2(n18510), .ZN(n18614) );
  AOI22_X1 U20535 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18515) );
  AOI22_X1 U20536 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18714), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18514) );
  AOI22_X1 U20537 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U20538 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18512) );
  NAND4_X1 U20539 ( .A1(n18515), .A2(n18514), .A3(n18513), .A4(n18512), .ZN(
        n18521) );
  AOI22_X1 U20540 ( .A1(n18713), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18519) );
  AOI22_X1 U20541 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U20542 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U20543 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18516) );
  NAND4_X1 U20544 ( .A1(n18519), .A2(n18518), .A3(n18517), .A4(n18516), .ZN(
        n18520) );
  NOR2_X1 U20545 ( .A1(n18521), .A2(n18520), .ZN(n18613) );
  NOR2_X1 U20546 ( .A1(n18614), .A2(n18613), .ZN(n18609) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18622), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18716), .ZN(n18533) );
  AOI22_X1 U20548 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18522), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11158), .ZN(n18532) );
  AOI22_X1 U20549 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18713), .ZN(n18523) );
  OAI21_X1 U20550 ( .B1(n18547), .B2(n18690), .A(n18523), .ZN(n18530) );
  AOI22_X1 U20551 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18528) );
  AOI22_X1 U20552 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11165), .B1(
        n18524), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U20553 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n21637), .ZN(n18526) );
  AOI22_X1 U20554 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18673), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18525) );
  NAND4_X1 U20555 ( .A1(n18528), .A2(n18527), .A3(n18526), .A4(n18525), .ZN(
        n18529) );
  AOI211_X1 U20556 ( .C1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .C2(n18475), .A(
        n18530), .B(n18529), .ZN(n18531) );
  NAND3_X1 U20557 ( .A1(n18533), .A2(n18532), .A3(n18531), .ZN(n18608) );
  NAND2_X1 U20558 ( .A1(n18609), .A2(n18608), .ZN(n18607) );
  NOR2_X1 U20559 ( .A1(n18603), .A2(n18607), .ZN(n18600) );
  AOI22_X1 U20560 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18544) );
  AOI22_X1 U20561 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18543) );
  AOI22_X1 U20562 ( .A1(n18713), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18534) );
  OAI21_X1 U20563 ( .B1(n18547), .B2(n18535), .A(n18534), .ZN(n18541) );
  AOI22_X1 U20564 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18539) );
  AOI22_X1 U20565 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18672), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18538) );
  AOI22_X1 U20566 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18537) );
  AOI22_X1 U20567 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18536) );
  NAND4_X1 U20568 ( .A1(n18539), .A2(n18538), .A3(n18537), .A4(n18536), .ZN(
        n18540) );
  AOI211_X1 U20569 ( .C1(n18712), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n18541), .B(n18540), .ZN(n18542) );
  NAND3_X1 U20570 ( .A1(n18544), .A2(n18543), .A3(n18542), .ZN(n18599) );
  NAND2_X1 U20571 ( .A1(n18600), .A2(n18599), .ZN(n18598) );
  NOR2_X1 U20572 ( .A1(n18587), .A2(n18598), .ZN(n18594) );
  AOI22_X1 U20573 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18557) );
  AOI22_X1 U20574 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18660), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18556) );
  AOI22_X1 U20575 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18545) );
  OAI21_X1 U20576 ( .B1(n18547), .B2(n18546), .A(n18545), .ZN(n18554) );
  AOI22_X1 U20577 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18552) );
  AOI22_X1 U20578 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18551) );
  AOI22_X1 U20579 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18550) );
  AOI22_X1 U20580 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18549) );
  NAND4_X1 U20581 ( .A1(n18552), .A2(n18551), .A3(n18550), .A4(n18549), .ZN(
        n18553) );
  AOI211_X1 U20582 ( .C1(n18711), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n18554), .B(n18553), .ZN(n18555) );
  NAND3_X1 U20583 ( .A1(n18557), .A2(n18556), .A3(n18555), .ZN(n18593) );
  NAND2_X1 U20584 ( .A1(n18594), .A2(n18593), .ZN(n18592) );
  NOR2_X1 U20585 ( .A1(n18590), .A2(n18592), .ZN(n18570) );
  AOI22_X1 U20586 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18562) );
  AOI22_X1 U20587 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18561) );
  AOI22_X1 U20588 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n21637), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18560) );
  AOI22_X1 U20589 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18558), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18559) );
  NAND4_X1 U20590 ( .A1(n18562), .A2(n18561), .A3(n18560), .A4(n18559), .ZN(
        n18568) );
  AOI22_X1 U20591 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18566) );
  AOI22_X1 U20592 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18565) );
  AOI22_X1 U20593 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18564) );
  AOI22_X1 U20594 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18563) );
  NAND4_X1 U20595 ( .A1(n18566), .A2(n18565), .A3(n18564), .A4(n18563), .ZN(
        n18567) );
  NOR2_X1 U20596 ( .A1(n18568), .A2(n18567), .ZN(n18569) );
  XOR2_X1 U20597 ( .A(n18570), .B(n18569), .Z(n21536) );
  OAI22_X1 U20598 ( .A1(n18572), .A2(n18571), .B1(n21536), .B2(n18689), .ZN(
        P3_U2673) );
  AOI22_X1 U20599 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18576) );
  AOI22_X1 U20600 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18714), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18575) );
  AOI22_X1 U20601 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18574) );
  AOI22_X1 U20602 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n21637), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18573) );
  NAND4_X1 U20603 ( .A1(n18576), .A2(n18575), .A3(n18574), .A4(n18573), .ZN(
        n18582) );
  AOI22_X1 U20604 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18580) );
  AOI22_X1 U20605 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18579) );
  AOI22_X1 U20606 ( .A1(n16155), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18578) );
  AOI22_X1 U20607 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18577) );
  NAND4_X1 U20608 ( .A1(n18580), .A2(n18579), .A3(n18578), .A4(n18577), .ZN(
        n18581) );
  NOR2_X1 U20609 ( .A1(n18582), .A2(n18581), .ZN(n21491) );
  AND2_X1 U20610 ( .A1(n18689), .A2(n18583), .ZN(n18642) );
  NAND2_X1 U20611 ( .A1(n18687), .A2(n18584), .ZN(n18641) );
  INV_X1 U20612 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21283) );
  AOI22_X1 U20613 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18642), .B1(n18586), 
        .B2(n21283), .ZN(n18585) );
  OAI21_X1 U20614 ( .B1(n21491), .B2(n18689), .A(n18585), .ZN(P3_U2682) );
  NAND2_X1 U20615 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18612), .ZN(n18606) );
  XNOR2_X1 U20616 ( .A(n18587), .B(n18598), .ZN(n21557) );
  NAND3_X1 U20617 ( .A1(n18589), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18689), 
        .ZN(n18588) );
  NAND3_X1 U20618 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n18602), .ZN(n18595) );
  XNOR2_X1 U20619 ( .A(n18590), .B(n18592), .ZN(n21545) );
  NAND3_X1 U20620 ( .A1(n18595), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n18689), 
        .ZN(n18591) );
  OAI221_X1 U20621 ( .B1(n18595), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18689), 
        .C2(n21545), .A(n18591), .ZN(P3_U2674) );
  OAI21_X1 U20622 ( .B1(n18594), .B2(n18593), .A(n18592), .ZN(n21552) );
  NAND3_X1 U20623 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18602), .A3(n21376), 
        .ZN(n18597) );
  NAND3_X1 U20624 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18689), .A3(n18595), 
        .ZN(n18596) );
  OAI211_X1 U20625 ( .C1(n18689), .C2(n21552), .A(n18597), .B(n18596), .ZN(
        P3_U2675) );
  AOI21_X1 U20626 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18689), .A(n18605), .ZN(
        n18601) );
  OAI21_X1 U20627 ( .B1(n18600), .B2(n18599), .A(n18598), .ZN(n21531) );
  OAI22_X1 U20628 ( .A1(n18602), .A2(n18601), .B1(n18689), .B2(n21531), .ZN(
        P3_U2677) );
  AOI21_X1 U20629 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18689), .A(n18611), .ZN(
        n18604) );
  XNOR2_X1 U20630 ( .A(n18603), .B(n18607), .ZN(n21525) );
  OAI22_X1 U20631 ( .A1(n18605), .A2(n18604), .B1(n18689), .B2(n21525), .ZN(
        P3_U2678) );
  INV_X1 U20632 ( .A(n18606), .ZN(n18616) );
  AOI21_X1 U20633 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18689), .A(n18616), .ZN(
        n18610) );
  OAI21_X1 U20634 ( .B1(n18609), .B2(n18608), .A(n18607), .ZN(n21563) );
  OAI22_X1 U20635 ( .A1(n18611), .A2(n18610), .B1(n18689), .B2(n21563), .ZN(
        P3_U2679) );
  AOI21_X1 U20636 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18689), .A(n18612), .ZN(
        n18615) );
  XNOR2_X1 U20637 ( .A(n18614), .B(n18613), .ZN(n21568) );
  OAI22_X1 U20638 ( .A1(n18616), .A2(n18615), .B1(n18689), .B2(n21568), .ZN(
        P3_U2680) );
  AOI22_X1 U20639 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18620) );
  AOI22_X1 U20640 ( .A1(n18672), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18619) );
  AOI22_X1 U20641 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18618) );
  AOI22_X1 U20642 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n21637), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18617) );
  NAND4_X1 U20643 ( .A1(n18620), .A2(n18619), .A3(n18618), .A4(n18617), .ZN(
        n18628) );
  AOI22_X1 U20644 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18626) );
  AOI22_X1 U20645 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18625) );
  AOI22_X1 U20646 ( .A1(n16134), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18621), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18624) );
  AOI22_X1 U20647 ( .A1(n18622), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18623) );
  NAND4_X1 U20648 ( .A1(n18626), .A2(n18625), .A3(n18624), .A4(n18623), .ZN(
        n18627) );
  NOR2_X1 U20649 ( .A1(n18628), .A2(n18627), .ZN(n21497) );
  NAND3_X1 U20650 ( .A1(n18630), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18689), 
        .ZN(n18629) );
  OAI221_X1 U20651 ( .B1(n18630), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18689), 
        .C2(n21497), .A(n18629), .ZN(P3_U2681) );
  AOI22_X1 U20652 ( .A1(n16155), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18634) );
  AOI22_X1 U20653 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18633) );
  AOI22_X1 U20654 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n21637), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18632) );
  AOI22_X1 U20655 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18631) );
  NAND4_X1 U20656 ( .A1(n18634), .A2(n18633), .A3(n18632), .A4(n18631), .ZN(
        n18640) );
  AOI22_X1 U20657 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18705), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18638) );
  AOI22_X1 U20658 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18637) );
  AOI22_X1 U20659 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18714), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18636) );
  AOI22_X1 U20660 ( .A1(n18711), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18635) );
  NAND4_X1 U20661 ( .A1(n18638), .A2(n18637), .A3(n18636), .A4(n18635), .ZN(
        n18639) );
  NOR2_X1 U20662 ( .A1(n18640), .A2(n18639), .ZN(n21495) );
  INV_X1 U20663 ( .A(n18641), .ZN(n18643) );
  OAI21_X1 U20664 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18643), .A(n18642), .ZN(
        n18644) );
  OAI21_X1 U20665 ( .B1(n21495), .B2(n18689), .A(n18644), .ZN(P3_U2683) );
  AOI22_X1 U20666 ( .A1(n16155), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18707), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18648) );
  AOI22_X1 U20667 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18647) );
  AOI22_X1 U20668 ( .A1(n21637), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18646) );
  AOI22_X1 U20669 ( .A1(n18674), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18673), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18645) );
  NAND4_X1 U20670 ( .A1(n18648), .A2(n18647), .A3(n18646), .A4(n18645), .ZN(
        n18654) );
  AOI22_X1 U20671 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14079), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18652) );
  AOI22_X1 U20672 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18714), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18651) );
  AOI22_X1 U20673 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18650) );
  AOI22_X1 U20674 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18649) );
  NAND4_X1 U20675 ( .A1(n18652), .A2(n18651), .A3(n18650), .A4(n18649), .ZN(
        n18653) );
  NOR2_X1 U20676 ( .A1(n18654), .A2(n18653), .ZN(n21512) );
  OAI211_X1 U20677 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18686), .A(n18667), .B(
        n18689), .ZN(n18655) );
  OAI21_X1 U20678 ( .B1(n21512), .B2(n18689), .A(n18655), .ZN(P3_U2685) );
  AOI22_X1 U20679 ( .A1(n18713), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18659) );
  AOI22_X1 U20680 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18711), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18658) );
  AOI22_X1 U20681 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18674), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18657) );
  AOI22_X1 U20682 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14127), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18656) );
  NAND4_X1 U20683 ( .A1(n18659), .A2(n18658), .A3(n18657), .A4(n18656), .ZN(
        n18666) );
  AOI22_X1 U20684 ( .A1(n11165), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18664) );
  AOI22_X1 U20685 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18707), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18663) );
  AOI22_X1 U20686 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18397), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18662) );
  AOI22_X1 U20687 ( .A1(n18660), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18661) );
  NAND4_X1 U20688 ( .A1(n18664), .A2(n18663), .A3(n18662), .A4(n18661), .ZN(
        n18665) );
  NOR2_X1 U20689 ( .A1(n18666), .A2(n18665), .ZN(n21507) );
  NAND3_X1 U20690 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18689), .A3(n18667), 
        .ZN(n18669) );
  OR3_X1 U20691 ( .A1(n21521), .A2(n18667), .A3(P3_EBX_REG_19__SCAN_IN), .ZN(
        n18668) );
  OAI211_X1 U20692 ( .C1(n21507), .C2(n18689), .A(n18669), .B(n18668), .ZN(
        P3_U2684) );
  AOI21_X1 U20693 ( .B1(n21237), .B2(n18670), .A(n18693), .ZN(n18671) );
  INV_X1 U20694 ( .A(n18671), .ZN(n18685) );
  AOI22_X1 U20695 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18711), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18678) );
  AOI22_X1 U20696 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18672), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18677) );
  AOI22_X1 U20697 ( .A1(n16155), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18673), .ZN(n18676) );
  AOI22_X1 U20698 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21637), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18674), .ZN(n18675) );
  NAND4_X1 U20699 ( .A1(n18678), .A2(n18677), .A3(n18676), .A4(n18675), .ZN(
        n18684) );
  AOI22_X1 U20700 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18682) );
  AOI22_X1 U20701 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11159), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n14090), .ZN(n18681) );
  AOI22_X1 U20702 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18621), .B1(
        n18717), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18680) );
  AOI22_X1 U20703 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18716), .ZN(n18679) );
  NAND4_X1 U20704 ( .A1(n18682), .A2(n18681), .A3(n18680), .A4(n18679), .ZN(
        n18683) );
  NOR2_X1 U20705 ( .A1(n18684), .A2(n18683), .ZN(n21517) );
  OAI22_X1 U20706 ( .A1(n18686), .A2(n18685), .B1(n21517), .B2(n18689), .ZN(
        P3_U2686) );
  NAND2_X1 U20707 ( .A1(n18687), .A2(n11217), .ZN(n18695) );
  NAND2_X1 U20708 ( .A1(n21025), .A2(n18688), .ZN(n21006) );
  INV_X1 U20709 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n21009) );
  OAI222_X1 U20710 ( .A1(n18695), .A2(n21006), .B1(n21009), .B2(n11217), .C1(
        n18690), .C2(n18689), .ZN(P3_U2702) );
  AOI22_X1 U20711 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18693), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18692), .ZN(n18694) );
  OAI21_X1 U20712 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18695), .A(n18694), .ZN(
        P3_U2703) );
  INV_X1 U20713 ( .A(n18696), .ZN(n18699) );
  OAI21_X1 U20714 ( .B1(n18697), .B2(n20949), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18698) );
  OAI21_X1 U20715 ( .B1(n18699), .B2(n22113), .A(n18698), .ZN(P3_U2634) );
  OAI21_X1 U20716 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18701), .A(n18700), .ZN(
        n22111) );
  OAI21_X1 U20717 ( .B1(n20944), .B2(n18703), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18702) );
  OAI221_X1 U20718 ( .B1(n18703), .B2(n22111), .C1(n18703), .C2(n19570), .A(
        n18702), .ZN(P3_U2863) );
  INV_X2 U20719 ( .A(n22117), .ZN(n21930) );
  OAI22_X2 U20720 ( .A1(n22116), .A2(n21930), .B1(n22118), .B2(n21745), .ZN(
        n18733) );
  NOR2_X1 U20721 ( .A1(n19855), .A2(n22088), .ZN(n18704) );
  AOI22_X1 U20722 ( .A1(n18705), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18726) );
  AOI22_X1 U20723 ( .A1(n18707), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18706), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18725) );
  AOI22_X1 U20724 ( .A1(n18708), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n21637), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18709) );
  OAI21_X1 U20725 ( .B1(n11234), .B2(n18710), .A(n18709), .ZN(n18723) );
  AOI22_X1 U20726 ( .A1(n18712), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18711), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18721) );
  AOI22_X1 U20727 ( .A1(n18714), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18713), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18720) );
  AOI22_X1 U20728 ( .A1(n18715), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11165), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18719) );
  AOI22_X1 U20729 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18716), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18718) );
  NAND4_X1 U20730 ( .A1(n18721), .A2(n18720), .A3(n18719), .A4(n18718), .ZN(
        n18722) );
  AOI211_X1 U20731 ( .C1(n18621), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n18723), .B(n18722), .ZN(n18724) );
  INV_X1 U20732 ( .A(n21673), .ZN(n21459) );
  INV_X1 U20733 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21752) );
  OAI221_X1 U20734 ( .B1(n21673), .B2(n21934), .C1(n21673), .C2(n21932), .A(
        n19044), .ZN(n18731) );
  NOR2_X1 U20735 ( .A1(n18769), .A2(n18731), .ZN(n18732) );
  INV_X1 U20736 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19063) );
  XNOR2_X1 U20737 ( .A(n18769), .B(n18731), .ZN(n19059) );
  NOR2_X1 U20738 ( .A1(n19063), .A2(n19059), .ZN(n19058) );
  NAND2_X1 U20739 ( .A1(n19046), .A2(n19044), .ZN(n19010) );
  INV_X1 U20740 ( .A(n21769), .ZN(n19013) );
  NAND2_X2 U20741 ( .A1(n19855), .A2(n22124), .ZN(n19140) );
  AOI222_X1 U20742 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18735), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18734), .C1(n18735), .C2(
        n18734), .ZN(n19062) );
  NAND3_X1 U20743 ( .A1(n18736), .A2(n21932), .A3(n21673), .ZN(n18739) );
  NOR3_X1 U20744 ( .A1(n19062), .A2(n19063), .A3(n18739), .ZN(n18742) );
  NAND2_X1 U20745 ( .A1(n21932), .A2(n18736), .ZN(n18737) );
  XOR2_X1 U20746 ( .A(n18737), .B(n21459), .Z(n19064) );
  NAND2_X1 U20747 ( .A1(n19062), .A2(n19063), .ZN(n18741) );
  NOR2_X1 U20748 ( .A1(n19062), .A2(n19063), .ZN(n18738) );
  XNOR2_X1 U20749 ( .A(n18739), .B(n18738), .ZN(n18740) );
  AOI21_X1 U20750 ( .B1(n19064), .B2(n18741), .A(n18740), .ZN(n19049) );
  OAI22_X1 U20751 ( .A1(n18965), .A2(n19013), .B1(n19140), .B2(n21990), .ZN(
        n18812) );
  INV_X1 U20752 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21818) );
  INV_X1 U20753 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n22024) );
  INV_X1 U20754 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n22023) );
  NAND2_X1 U20755 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19011) );
  NOR3_X1 U20756 ( .A1(n22024), .A2(n22023), .A3(n19011), .ZN(n21778) );
  NAND2_X1 U20757 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21778), .ZN(
        n21819) );
  NOR2_X1 U20758 ( .A1(n21818), .A2(n21819), .ZN(n21807) );
  NAND2_X1 U20759 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21807), .ZN(
        n21661) );
  INV_X1 U20760 ( .A(n21661), .ZN(n21985) );
  NAND2_X1 U20761 ( .A1(n18812), .A2(n21985), .ZN(n18822) );
  INV_X1 U20762 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n22004) );
  INV_X1 U20763 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n22012) );
  NOR2_X1 U20764 ( .A1(n22004), .A2(n22012), .ZN(n21665) );
  INV_X1 U20765 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21997) );
  NAND2_X1 U20766 ( .A1(n21665), .A2(n21997), .ZN(n22003) );
  INV_X1 U20767 ( .A(n19098), .ZN(n18901) );
  INV_X1 U20768 ( .A(n18743), .ZN(n18745) );
  AOI21_X1 U20769 ( .B1(n18901), .B2(n18745), .A(n19141), .ZN(n18981) );
  OAI21_X1 U20770 ( .B1(n18744), .B2(n18899), .A(n18981), .ZN(n18761) );
  INV_X1 U20771 ( .A(n18899), .ZN(n19142) );
  NOR3_X1 U20772 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18898), .A3(
        n18745), .ZN(n18762) );
  INV_X1 U20773 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21252) );
  OAI22_X1 U20774 ( .A1(n18767), .A2(n21252), .B1(n21245), .B2(n18979), .ZN(
        n18746) );
  AOI211_X1 U20775 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18761), .A(
        n18762), .B(n18746), .ZN(n18757) );
  NAND2_X1 U20776 ( .A1(n21778), .A2(n21769), .ZN(n18790) );
  INV_X1 U20777 ( .A(n18790), .ZN(n21782) );
  NAND2_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21782), .ZN(
        n18998) );
  INV_X1 U20779 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21813) );
  NOR2_X1 U20780 ( .A1(n21990), .A2(n21819), .ZN(n18991) );
  NAND2_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18991), .ZN(
        n18990) );
  NOR2_X2 U20782 ( .A1(n21813), .A2(n18990), .ZN(n21811) );
  OAI22_X1 U20783 ( .A1(n18965), .A2(n21810), .B1(n19140), .B2(n21811), .ZN(
        n18747) );
  INV_X1 U20784 ( .A(n18747), .ZN(n18789) );
  OAI21_X1 U20785 ( .B1(n21665), .B2(n18822), .A(n18789), .ZN(n18987) );
  NAND2_X1 U20786 ( .A1(n19044), .A2(n21997), .ZN(n18845) );
  OAI21_X1 U20787 ( .B1(n19044), .B2(n21997), .A(n18845), .ZN(n18755) );
  NOR2_X1 U20788 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19022) );
  NOR3_X2 U20789 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n18791), .ZN(n18772) );
  NAND3_X1 U20790 ( .A1(n18772), .A2(n21813), .A3(n21818), .ZN(n18750) );
  NAND2_X1 U20791 ( .A1(n18750), .A2(n19044), .ZN(n18754) );
  NOR2_X1 U20792 ( .A1(n19020), .A2(n21661), .ZN(n18752) );
  INV_X1 U20793 ( .A(n18752), .ZN(n18753) );
  NAND2_X1 U20794 ( .A1(n18754), .A2(n18753), .ZN(n18873) );
  XNOR2_X1 U20795 ( .A(n18755), .B(n18816), .ZN(n22000) );
  AOI22_X1 U20796 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18987), .B1(
        n19040), .B2(n22000), .ZN(n18756) );
  OAI211_X1 U20797 ( .C1(n18822), .C2(n22003), .A(n18757), .B(n18756), .ZN(
        P3_U2812) );
  NAND2_X1 U20798 ( .A1(n21665), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21662) );
  INV_X1 U20799 ( .A(n21662), .ZN(n21675) );
  NAND2_X1 U20800 ( .A1(n21675), .A2(n18986), .ZN(n18834) );
  INV_X1 U20801 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21976) );
  NOR2_X1 U20802 ( .A1(n21662), .A2(n21976), .ZN(n21663) );
  NAND2_X1 U20803 ( .A1(n21811), .A2(n21663), .ZN(n21968) );
  NAND2_X1 U20804 ( .A1(n21810), .A2(n21663), .ZN(n21966) );
  AOI22_X1 U20805 ( .A1(n19074), .A2(n21968), .B1(n19047), .B2(n21966), .ZN(
        n18852) );
  INV_X1 U20806 ( .A(n18845), .ZN(n18815) );
  NAND2_X1 U20807 ( .A1(n18815), .A2(n18816), .ZN(n18832) );
  NAND3_X1 U20808 ( .A1(n18749), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18758), .ZN(n18846) );
  NAND2_X1 U20809 ( .A1(n18832), .A2(n18846), .ZN(n18759) );
  XOR2_X1 U20810 ( .A(n18759), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n21972) );
  NOR3_X1 U20811 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18898), .A3(
        n18760), .ZN(n18765) );
  INV_X2 U20812 ( .A(n18767), .ZN(n22043) );
  NAND2_X1 U20813 ( .A1(n22043), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21973) );
  OAI21_X1 U20814 ( .B1(n18762), .B2(n18761), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18763) );
  OAI211_X1 U20815 ( .C1(n18979), .C2(n21259), .A(n21973), .B(n18763), .ZN(
        n18764) );
  AOI211_X1 U20816 ( .C1(n19040), .C2(n21972), .A(n18765), .B(n18764), .ZN(
        n18766) );
  OAI221_X1 U20817 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18834), 
        .C1(n21976), .C2(n18852), .A(n18766), .ZN(P3_U2811) );
  NAND2_X1 U20818 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18993), .ZN(
        n18781) );
  OAI21_X1 U20819 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18993), .A(
        n18781), .ZN(n21202) );
  NOR2_X1 U20820 ( .A1(n18898), .A2(n21201), .ZN(n18784) );
  AOI21_X1 U20821 ( .B1(n18901), .B2(n21201), .A(n19141), .ZN(n18994) );
  OAI21_X1 U20822 ( .B1(n18993), .B2(n18899), .A(n18994), .ZN(n18782) );
  INV_X1 U20823 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n21212) );
  NOR2_X1 U20824 ( .A1(n18767), .A2(n21212), .ZN(n21815) );
  AOI221_X1 U20825 ( .B1(n18784), .B2(n21206), .C1(n18782), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n21815), .ZN(n18777) );
  NOR2_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18990), .ZN(
        n21816) );
  NOR2_X1 U20827 ( .A1(n19013), .A2(n18965), .ZN(n18768) );
  AOI21_X1 U20828 ( .B1(n21807), .B2(n18768), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18774) );
  INV_X1 U20829 ( .A(n21819), .ZN(n18770) );
  NAND2_X1 U20830 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21660) );
  NOR3_X1 U20831 ( .A1(n18769), .A2(n19044), .A3(n21660), .ZN(n19031) );
  NAND2_X1 U20832 ( .A1(n18770), .A2(n19031), .ZN(n18999) );
  NAND2_X1 U20833 ( .A1(n18772), .A2(n18771), .ZN(n19000) );
  AOI22_X1 U20834 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18999), .B1(
        n19000), .B2(n21818), .ZN(n18773) );
  XOR2_X1 U20835 ( .A(n21813), .B(n18773), .Z(n21824) );
  OAI22_X1 U20836 ( .A1(n18789), .A2(n18774), .B1(n21824), .B2(n19057), .ZN(
        n18775) );
  AOI21_X1 U20837 ( .B1(n19074), .B2(n21816), .A(n18775), .ZN(n18776) );
  OAI211_X1 U20838 ( .C1(n18979), .C2(n21202), .A(n18777), .B(n18776), .ZN(
        P3_U2815) );
  AOI22_X1 U20839 ( .A1(n18749), .A2(n22012), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19044), .ZN(n18778) );
  XOR2_X1 U20840 ( .A(n18873), .B(n18778), .Z(n22017) );
  INV_X1 U20841 ( .A(n18979), .ZN(n18971) );
  INV_X1 U20842 ( .A(n18779), .ZN(n18780) );
  AOI21_X1 U20843 ( .B1(n21221), .B2(n18781), .A(n18780), .ZN(n21217) );
  AOI22_X1 U20844 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18782), .B1(
        n18971), .B2(n21217), .ZN(n18786) );
  NAND2_X1 U20845 ( .A1(n22043), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n22018) );
  NAND2_X1 U20846 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18783) );
  OAI211_X1 U20847 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18784), .B(n18783), .ZN(n18785) );
  NAND3_X1 U20848 ( .A1(n18786), .A2(n22018), .A3(n18785), .ZN(n18787) );
  AOI21_X1 U20849 ( .B1(n19040), .B2(n22017), .A(n18787), .ZN(n18788) );
  OAI221_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18822), 
        .C1(n22012), .C2(n18789), .A(n18788), .ZN(P3_U2814) );
  INV_X1 U20851 ( .A(n21990), .ZN(n21674) );
  NAND2_X1 U20852 ( .A1(n21778), .A2(n21674), .ZN(n21780) );
  AOI22_X1 U20853 ( .A1(n19074), .A2(n21780), .B1(n19047), .B2(n18790), .ZN(
        n18810) );
  NOR2_X1 U20854 ( .A1(n22024), .A2(n19011), .ZN(n21784) );
  NAND2_X1 U20855 ( .A1(n19044), .A2(n18791), .ZN(n18807) );
  OAI221_X1 U20856 ( .B1(n19044), .B2(n18792), .C1(n19044), .C2(n21784), .A(
        n18807), .ZN(n18793) );
  XOR2_X1 U20857 ( .A(n22023), .B(n18793), .Z(n21785) );
  INV_X1 U20858 ( .A(n18812), .ZN(n19043) );
  INV_X1 U20859 ( .A(n21784), .ZN(n21765) );
  NOR3_X1 U20860 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19043), .A3(
        n21765), .ZN(n18800) );
  NAND2_X1 U20861 ( .A1(n18794), .A2(n18935), .ZN(n18802) );
  NOR2_X1 U20862 ( .A1(n21115), .A2(n21012), .ZN(n19023) );
  INV_X1 U20863 ( .A(n19023), .ZN(n19035) );
  NOR2_X1 U20864 ( .A1(n18795), .A2(n19035), .ZN(n18797) );
  AOI21_X1 U20865 ( .B1(n18901), .B2(n21147), .A(n19142), .ZN(n18796) );
  OAI21_X1 U20866 ( .B1(n18797), .B2(n18796), .A(n19097), .ZN(n18805) );
  INV_X1 U20867 ( .A(n18797), .ZN(n19004) );
  NOR2_X1 U20868 ( .A1(n21165), .A2(n19004), .ZN(n21170) );
  AOI21_X1 U20869 ( .B1(n21165), .B2(n19004), .A(n21170), .ZN(n21161) );
  AOI22_X1 U20870 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18805), .B1(
        n18971), .B2(n21161), .ZN(n18798) );
  NAND2_X1 U20871 ( .A1(n22043), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21786) );
  OAI211_X1 U20872 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18802), .A(
        n18798), .B(n21786), .ZN(n18799) );
  AOI211_X1 U20873 ( .C1(n21785), .C2(n19040), .A(n18800), .B(n18799), .ZN(
        n18801) );
  OAI21_X1 U20874 ( .B1(n18810), .B2(n22023), .A(n18801), .ZN(P3_U2818) );
  INV_X1 U20875 ( .A(n18992), .ZN(n18995) );
  OAI22_X1 U20876 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n21170), .B1(
        n21012), .B2(n18995), .ZN(n21183) );
  INV_X1 U20877 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21180) );
  NOR2_X1 U20878 ( .A1(n18767), .A2(n21180), .ZN(n18804) );
  AOI221_X1 U20879 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C1(n21165), .C2(n21177), .A(
        n18802), .ZN(n18803) );
  AOI211_X1 U20880 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18805), .A(
        n18804), .B(n18803), .ZN(n18814) );
  INV_X1 U20881 ( .A(n21778), .ZN(n18806) );
  NOR2_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18806), .ZN(
        n22021) );
  INV_X1 U20883 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21792) );
  OAI22_X1 U20884 ( .A1(n19020), .A2(n18806), .B1(n18749), .B2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18808) );
  NAND2_X1 U20885 ( .A1(n18808), .A2(n18807), .ZN(n18809) );
  XOR2_X1 U20886 ( .A(n18809), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n22032) );
  OAI22_X1 U20887 ( .A1(n18810), .A2(n21792), .B1(n19057), .B2(n22032), .ZN(
        n18811) );
  AOI21_X1 U20888 ( .B1(n22021), .B2(n18812), .A(n18811), .ZN(n18813) );
  OAI211_X1 U20889 ( .C1(n18979), .C2(n21183), .A(n18814), .B(n18813), .ZN(
        P3_U2817) );
  INV_X1 U20890 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21836) );
  INV_X1 U20891 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21670) );
  INV_X1 U20892 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18837) );
  NAND4_X1 U20893 ( .A1(n18815), .A2(n21670), .A3(n21976), .A4(n18837), .ZN(
        n18863) );
  NOR2_X1 U20894 ( .A1(n21670), .A2(n21976), .ZN(n21668) );
  NAND2_X1 U20895 ( .A1(n21668), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21835) );
  NOR3_X1 U20896 ( .A1(n18816), .A2(n21835), .A3(n21997), .ZN(n18876) );
  INV_X1 U20897 ( .A(n18876), .ZN(n18817) );
  AOI21_X1 U20898 ( .B1(n18863), .B2(n18817), .A(n18875), .ZN(n18864) );
  XOR2_X1 U20899 ( .A(n21836), .B(n18864), .Z(n21828) );
  OAI21_X1 U20900 ( .B1(n18818), .B2(n18899), .A(n19097), .ZN(n18819) );
  AOI21_X1 U20901 ( .B1(n18901), .B2(n11269), .A(n18819), .ZN(n18841) );
  OAI21_X1 U20902 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18980), .A(
        n18841), .ZN(n18830) );
  NAND2_X1 U20903 ( .A1(n22043), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21830) );
  NOR2_X1 U20904 ( .A1(n18898), .A2(n11269), .ZN(n18831) );
  OAI211_X1 U20905 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18831), .B(n18820), .ZN(n18821) );
  OAI211_X1 U20906 ( .C1(n18979), .C2(n21296), .A(n21830), .B(n18821), .ZN(
        n18827) );
  NOR2_X1 U20907 ( .A1(n21662), .A2(n21835), .ZN(n18823) );
  INV_X1 U20908 ( .A(n18823), .ZN(n18853) );
  NOR2_X1 U20909 ( .A1(n18853), .A2(n18822), .ZN(n18825) );
  NAND2_X1 U20910 ( .A1(n18823), .A2(n21811), .ZN(n21659) );
  NAND2_X1 U20911 ( .A1(n18823), .A2(n21810), .ZN(n21658) );
  AOI22_X1 U20912 ( .A1(n19074), .A2(n21659), .B1(n19047), .B2(n21658), .ZN(
        n18838) );
  INV_X1 U20913 ( .A(n18838), .ZN(n18824) );
  MUX2_X1 U20914 ( .A(n18825), .B(n18824), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18826) );
  AOI211_X1 U20915 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n18830), .A(
        n18827), .B(n18826), .ZN(n18828) );
  OAI21_X1 U20916 ( .B1(n19057), .B2(n21828), .A(n18828), .ZN(P3_U2808) );
  OAI22_X1 U20917 ( .A1(n18767), .A2(n21680), .B1(n21288), .B2(n18979), .ZN(
        n18829) );
  AOI221_X1 U20918 ( .B1(n18831), .B2(n21282), .C1(n18830), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18829), .ZN(n18836) );
  OAI33_X1 U20919 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n18832), .B1(n21976), .B2(
        n18846), .B3(n21670), .ZN(n18833) );
  XOR2_X1 U20920 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18833), .Z(
        n21678) );
  AND2_X1 U20921 ( .A1(n18837), .A2(n21668), .ZN(n21677) );
  INV_X1 U20922 ( .A(n18834), .ZN(n18848) );
  AOI22_X1 U20923 ( .A1(n19040), .A2(n21678), .B1(n21677), .B2(n18848), .ZN(
        n18835) );
  OAI211_X1 U20924 ( .C1(n18838), .C2(n18837), .A(n18836), .B(n18835), .ZN(
        P3_U2809) );
  INV_X1 U20925 ( .A(n21272), .ZN(n18844) );
  INV_X1 U20926 ( .A(n18980), .ZN(n18843) );
  INV_X2 U20927 ( .A(n19653), .ZN(n19901) );
  AOI21_X1 U20928 ( .B1(n18839), .B2(n19901), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18840) );
  NAND2_X1 U20929 ( .A1(n22043), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21982) );
  OAI21_X1 U20930 ( .B1(n18841), .B2(n18840), .A(n21982), .ZN(n18842) );
  AOI221_X1 U20931 ( .B1(n18971), .B2(n18844), .C1(n18843), .C2(n18844), .A(
        n18842), .ZN(n18851) );
  AOI221_X1 U20932 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18846), 
        .C1(n21976), .C2(n18845), .A(n18875), .ZN(n18847) );
  XOR2_X1 U20933 ( .A(n21670), .B(n18847), .Z(n21984) );
  INV_X1 U20934 ( .A(n21984), .ZN(n18849) );
  NOR2_X1 U20935 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21976), .ZN(
        n21979) );
  AOI22_X1 U20936 ( .A1(n19040), .A2(n18849), .B1(n18848), .B2(n21979), .ZN(
        n18850) );
  OAI211_X1 U20937 ( .C1(n18852), .C2(n21670), .A(n18851), .B(n18850), .ZN(
        P3_U2810) );
  NAND2_X1 U20938 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18871) );
  NOR2_X1 U20939 ( .A1(n18871), .A2(n18853), .ZN(n18880) );
  NAND2_X1 U20940 ( .A1(n18880), .A2(n21811), .ZN(n21942) );
  AOI22_X1 U20941 ( .A1(n19047), .A2(n21946), .B1(n19074), .B2(n21942), .ZN(
        n18890) );
  INV_X1 U20942 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21956) );
  INV_X1 U20943 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21308) );
  OAI21_X1 U20944 ( .B1(n18854), .B2(n18980), .A(n21308), .ZN(n18860) );
  NAND2_X1 U20945 ( .A1(n18856), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18896) );
  AOI22_X1 U20946 ( .A1(n19901), .A2(n18896), .B1(n19142), .B2(n18854), .ZN(
        n18855) );
  OAI211_X1 U20947 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18899), .A(
        n18855), .B(n19097), .ZN(n18884) );
  INV_X1 U20948 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21303) );
  NOR2_X1 U20949 ( .A1(n18767), .A2(n21303), .ZN(n21952) );
  INV_X1 U20950 ( .A(n18856), .ZN(n18858) );
  NAND2_X1 U20951 ( .A1(n19901), .A2(n18896), .ZN(n18857) );
  OAI22_X1 U20952 ( .A1(n18858), .A2(n18857), .B1(n21314), .B2(n18979), .ZN(
        n18859) );
  AOI211_X1 U20953 ( .C1(n18860), .C2(n18884), .A(n21952), .B(n18859), .ZN(
        n18868) );
  NAND2_X1 U20954 ( .A1(n19047), .A2(n21946), .ZN(n18862) );
  NAND2_X1 U20955 ( .A1(n19074), .A2(n21942), .ZN(n18861) );
  OAI22_X1 U20956 ( .A1(n21658), .A2(n18862), .B1(n21659), .B2(n18861), .ZN(
        n18866) );
  NOR2_X1 U20957 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18863), .ZN(
        n18872) );
  OAI221_X1 U20958 ( .B1(n18872), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n18872), .C2(n18749), .A(n18864), .ZN(n18865) );
  XOR2_X1 U20959 ( .A(n21956), .B(n18865), .Z(n21953) );
  AOI22_X1 U20960 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18866), .B1(
        n19040), .B2(n21953), .ZN(n18867) );
  OAI211_X1 U20961 ( .C1(n18890), .C2(n21956), .A(n18868), .B(n18867), .ZN(
        P3_U2807) );
  INV_X1 U20962 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21840) );
  INV_X1 U20963 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21959) );
  NOR2_X1 U20964 ( .A1(n21959), .A2(n21946), .ZN(n18908) );
  XOR2_X1 U20965 ( .A(n21840), .B(n18908), .Z(n21839) );
  NAND2_X1 U20966 ( .A1(n22043), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21845) );
  NOR2_X1 U20967 ( .A1(n18898), .A2(n18896), .ZN(n18886) );
  OAI211_X1 U20968 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18886), .B(n18897), .ZN(n18869) );
  OAI211_X1 U20969 ( .C1(n18979), .C2(n21336), .A(n21845), .B(n18869), .ZN(
        n18870) );
  AOI21_X1 U20970 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18884), .A(
        n18870), .ZN(n18879) );
  NAND2_X1 U20971 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21857) );
  NOR2_X1 U20972 ( .A1(n21857), .A2(n21942), .ZN(n18909) );
  AOI221_X1 U20973 ( .B1(n21959), .B2(n21840), .C1(n21942), .C2(n21840), .A(
        n18909), .ZN(n21834) );
  INV_X1 U20974 ( .A(n18871), .ZN(n21856) );
  AOI22_X1 U20975 ( .A1(n18880), .A2(n18873), .B1(n18872), .B2(n21956), .ZN(
        n18874) );
  NAND2_X1 U20976 ( .A1(n18882), .A2(n21959), .ZN(n18881) );
  NAND3_X1 U20977 ( .A1(n21856), .A2(n18876), .A3(n18881), .ZN(n18893) );
  INV_X1 U20978 ( .A(n18893), .ZN(n18923) );
  NAND2_X1 U20979 ( .A1(n19044), .A2(n18881), .ZN(n18922) );
  OAI21_X1 U20980 ( .B1(n19044), .B2(n18923), .A(n18922), .ZN(n18877) );
  XOR2_X1 U20981 ( .A(n18877), .B(n21840), .Z(n21833) );
  AOI22_X1 U20982 ( .A1(n19074), .A2(n21834), .B1(n19040), .B2(n21833), .ZN(
        n18878) );
  OAI211_X1 U20983 ( .C1(n18965), .C2(n21839), .A(n18879), .B(n18878), .ZN(
        P3_U2805) );
  NAND2_X1 U20984 ( .A1(n18880), .A2(n18986), .ZN(n18891) );
  OAI21_X1 U20985 ( .B1(n18882), .B2(n21959), .A(n18881), .ZN(n21963) );
  NOR2_X1 U20986 ( .A1(n18767), .A2(n21965), .ZN(n18883) );
  AOI221_X1 U20987 ( .B1(n18886), .B2(n18885), .C1(n18884), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18883), .ZN(n18887) );
  OAI21_X1 U20988 ( .B1(n21323), .B2(n18979), .A(n18887), .ZN(n18888) );
  AOI21_X1 U20989 ( .B1(n19040), .B2(n21963), .A(n18888), .ZN(n18889) );
  OAI221_X1 U20990 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18891), 
        .C1(n21959), .C2(n18890), .A(n18889), .ZN(P3_U2806) );
  INV_X1 U20991 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21850) );
  INV_X1 U20992 ( .A(n18919), .ZN(n18952) );
  INV_X1 U20993 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21925) );
  NAND2_X1 U20994 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21925), .ZN(
        n18912) );
  NAND2_X1 U20995 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21865) );
  OAI21_X1 U20996 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n19044), .ZN(n18892) );
  OAI211_X1 U20997 ( .C1(n18893), .C2(n21865), .A(n18892), .B(n18922), .ZN(
        n18894) );
  AND2_X1 U20998 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18894), .ZN(
        n18945) );
  AOI22_X1 U20999 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n19044), .B1(
        n18749), .B2(n21925), .ZN(n21938) );
  AOI211_X1 U21000 ( .C1(n18895), .C2(n21938), .A(n21923), .B(n19057), .ZN(
        n18907) );
  NOR2_X1 U21001 ( .A1(n18897), .A2(n18896), .ZN(n18925) );
  NAND2_X1 U21002 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18925), .ZN(
        n18902) );
  NOR3_X1 U21003 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18898), .A3(
        n18902), .ZN(n18916) );
  OAI21_X1 U21004 ( .B1(n14034), .B2(n18899), .A(n19097), .ZN(n18900) );
  AOI21_X1 U21005 ( .B1(n18901), .B2(n18902), .A(n18900), .ZN(n18927) );
  OAI21_X1 U21006 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18980), .A(
        n18927), .ZN(n18917) );
  OAI21_X1 U21007 ( .B1(n18916), .B2(n18917), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18905) );
  NOR2_X1 U21008 ( .A1(n18903), .A2(n18902), .ZN(n18934) );
  NAND3_X1 U21009 ( .A1(n18934), .A2(n11349), .A3(n18935), .ZN(n18904) );
  OAI211_X1 U21010 ( .C1(n18979), .C2(n21382), .A(n18905), .B(n18904), .ZN(
        n18906) );
  AOI211_X1 U21011 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n22043), .A(n18907), 
        .B(n18906), .ZN(n18911) );
  NAND3_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n18908), .ZN(n21848) );
  NAND2_X1 U21013 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18909), .ZN(
        n21852) );
  AOI22_X1 U21014 ( .A1(n19047), .A2(n21848), .B1(n19074), .B2(n21852), .ZN(
        n18931) );
  NAND2_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18931), .ZN(
        n18918) );
  OAI211_X1 U21016 ( .C1(n19074), .C2(n19047), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18918), .ZN(n18910) );
  OAI211_X1 U21017 ( .C1(n18952), .C2(n18912), .A(n18911), .B(n18910), .ZN(
        P3_U2802) );
  AOI21_X1 U21018 ( .B1(n19044), .B2(n18914), .A(n18913), .ZN(n21877) );
  OAI22_X1 U21019 ( .A1(n18767), .A2(n21862), .B1(n21367), .B2(n18979), .ZN(
        n18915) );
  AOI211_X1 U21020 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18917), .A(
        n18916), .B(n18915), .ZN(n18921) );
  OAI21_X1 U21021 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18919), .A(
        n18918), .ZN(n18920) );
  OAI211_X1 U21022 ( .C1(n21877), .C2(n19057), .A(n18921), .B(n18920), .ZN(
        P3_U2803) );
  OAI221_X1 U21023 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n19044), 
        .C1(n21840), .C2(n18923), .A(n18922), .ZN(n18924) );
  XOR2_X1 U21024 ( .A(n21850), .B(n18924), .Z(n21847) );
  AOI21_X1 U21025 ( .B1(n18979), .B2(n18980), .A(n21356), .ZN(n18929) );
  AOI21_X1 U21026 ( .B1(n18925), .B2(n19901), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18926) );
  OAI22_X1 U21027 ( .A1(n18927), .A2(n18926), .B1(n18767), .B2(n21359), .ZN(
        n18928) );
  AOI211_X1 U21028 ( .C1(n21847), .C2(n19040), .A(n18929), .B(n18928), .ZN(
        n18930) );
  OAI221_X1 U21029 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18932), 
        .C1(n21850), .C2(n18931), .A(n18930), .ZN(P3_U2804) );
  INV_X1 U21030 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21913) );
  NAND2_X1 U21031 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21881) );
  INV_X1 U21032 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21908) );
  NOR2_X1 U21033 ( .A1(n21881), .A2(n21908), .ZN(n21899) );
  INV_X1 U21034 ( .A(n21899), .ZN(n18953) );
  NOR2_X1 U21035 ( .A1(n21852), .A2(n18953), .ZN(n21892) );
  NAND2_X1 U21036 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21892), .ZN(
        n18933) );
  XNOR2_X1 U21037 ( .A(n21913), .B(n18933), .ZN(n21912) );
  NAND2_X1 U21038 ( .A1(n22043), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n21919) );
  INV_X1 U21039 ( .A(n21919), .ZN(n18943) );
  NAND2_X1 U21040 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18934), .ZN(
        n18962) );
  NOR2_X1 U21041 ( .A1(n18961), .A2(n18962), .ZN(n18936) );
  NAND2_X1 U21042 ( .A1(n18936), .A2(n18935), .ZN(n18957) );
  XNOR2_X1 U21043 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18941) );
  NOR2_X1 U21044 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18980), .ZN(
        n18972) );
  INV_X1 U21045 ( .A(n18936), .ZN(n18938) );
  AOI22_X1 U21046 ( .A1(n19901), .A2(n18938), .B1(n19142), .B2(n18937), .ZN(
        n18939) );
  NAND2_X1 U21047 ( .A1(n18939), .A2(n19097), .ZN(n18964) );
  NOR2_X1 U21048 ( .A1(n18972), .A2(n18964), .ZN(n18956) );
  OAI22_X1 U21049 ( .A1(n18957), .A2(n18941), .B1(n18956), .B2(n18940), .ZN(
        n18942) );
  AOI211_X1 U21050 ( .C1(n14024), .C2(n18971), .A(n18943), .B(n18942), .ZN(
        n18948) );
  NOR2_X1 U21051 ( .A1(n21848), .A2(n18953), .ZN(n21891) );
  NAND2_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21891), .ZN(
        n18944) );
  XOR2_X1 U21053 ( .A(n21913), .B(n18944), .Z(n21917) );
  NAND3_X1 U21054 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18749), .A3(
        n18945), .ZN(n21924) );
  NOR2_X1 U21055 ( .A1(n21924), .A2(n21908), .ZN(n18949) );
  NAND3_X1 U21056 ( .A1(n21939), .A2(n21925), .A3(n19044), .ZN(n18966) );
  NOR2_X1 U21057 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n18966), .ZN(
        n18950) );
  INV_X1 U21058 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21910) );
  AOI22_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18949), .B1(
        n18950), .B2(n21910), .ZN(n18946) );
  XOR2_X1 U21060 ( .A(n21913), .B(n18946), .Z(n21918) );
  AOI22_X1 U21061 ( .A1(n21917), .A2(n19047), .B1(n19040), .B2(n21918), .ZN(
        n18947) );
  OAI211_X1 U21062 ( .C1(n21912), .C2(n19140), .A(n18948), .B(n18947), .ZN(
        P3_U2799) );
  NOR2_X1 U21063 ( .A1(n18950), .A2(n18949), .ZN(n18951) );
  XOR2_X1 U21064 ( .A(n18951), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n21906) );
  NOR2_X1 U21065 ( .A1(n18953), .A2(n18952), .ZN(n18959) );
  OAI22_X1 U21066 ( .A1(n21891), .A2(n18965), .B1(n21892), .B2(n19140), .ZN(
        n18969) );
  OAI22_X1 U21067 ( .A1(n18767), .A2(n19235), .B1(n21407), .B2(n18979), .ZN(
        n18954) );
  INV_X1 U21068 ( .A(n18954), .ZN(n18955) );
  OAI221_X1 U21069 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18957), .C1(
        n11351), .C2(n18956), .A(n18955), .ZN(n18958) );
  AOI221_X1 U21070 ( .B1(n18959), .B2(n21910), .C1(n18969), .C2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n18958), .ZN(n18960) );
  OAI21_X1 U21071 ( .B1(n21906), .B2(n19057), .A(n18960), .ZN(P3_U2800) );
  OAI21_X1 U21072 ( .B1(n18962), .B2(n19653), .A(n18961), .ZN(n18963) );
  AOI22_X1 U21073 ( .A1(n22043), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18964), 
        .B2(n18963), .ZN(n18976) );
  NOR2_X1 U21074 ( .A1(n21881), .A2(n21848), .ZN(n21929) );
  NOR2_X1 U21075 ( .A1(n21891), .A2(n18965), .ZN(n18968) );
  NAND2_X1 U21076 ( .A1(n18966), .A2(n21924), .ZN(n18967) );
  XOR2_X1 U21077 ( .A(n18967), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21878) );
  AOI22_X1 U21078 ( .A1(n21929), .A2(n18968), .B1(n19040), .B2(n21878), .ZN(
        n18975) );
  NOR2_X1 U21079 ( .A1(n21881), .A2(n21852), .ZN(n21931) );
  OAI221_X1 U21080 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21931), 
        .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n19074), .A(n18969), .ZN(
        n18974) );
  OAI21_X1 U21081 ( .B1(n18972), .B2(n18971), .A(n18970), .ZN(n18973) );
  NAND4_X1 U21082 ( .A1(n18976), .A2(n18975), .A3(n18974), .A4(n18973), .ZN(
        P3_U2801) );
  AOI21_X1 U21083 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18978), .A(
        n18977), .ZN(n22011) );
  NOR2_X1 U21084 ( .A1(n18767), .A2(n21242), .ZN(n22007) );
  AOI221_X1 U21085 ( .B1(n18983), .B2(n18982), .C1(n19653), .C2(n18982), .A(
        n18981), .ZN(n18984) );
  AOI211_X1 U21086 ( .C1(n18985), .C2(n19137), .A(n22007), .B(n18984), .ZN(
        n18989) );
  NOR2_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n22012), .ZN(
        n22009) );
  AOI22_X1 U21088 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18987), .B1(
        n18986), .B2(n22009), .ZN(n18988) );
  OAI211_X1 U21089 ( .C1(n22011), .C2(n19057), .A(n18989), .B(n18988), .ZN(
        P3_U2813) );
  OAI21_X1 U21090 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18991), .A(
        n18990), .ZN(n21804) );
  INV_X1 U21091 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21196) );
  NAND2_X1 U21092 ( .A1(n18992), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21186) );
  AOI21_X1 U21093 ( .B1(n21196), .B2(n21186), .A(n18993), .ZN(n21188) );
  AOI221_X1 U21094 ( .B1(n18995), .B2(n21196), .C1(n19653), .C2(n21196), .A(
        n18994), .ZN(n18997) );
  INV_X1 U21095 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19231) );
  NOR2_X1 U21096 ( .A1(n18767), .A2(n19231), .ZN(n18996) );
  AOI211_X1 U21097 ( .C1(n21188), .C2(n19137), .A(n18997), .B(n18996), .ZN(
        n19003) );
  AOI21_X1 U21098 ( .B1(n21818), .B2(n18998), .A(n21820), .ZN(n21797) );
  NAND2_X1 U21099 ( .A1(n19000), .A2(n18999), .ZN(n19001) );
  XOR2_X1 U21100 ( .A(n19001), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n21800) );
  AOI22_X1 U21101 ( .A1(n19047), .A2(n21797), .B1(n19040), .B2(n21800), .ZN(
        n19002) );
  OAI211_X1 U21102 ( .C1(n19140), .C2(n21804), .A(n19003), .B(n19002), .ZN(
        P3_U2816) );
  NOR2_X1 U21103 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19011), .ZN(
        n21764) );
  AOI21_X1 U21104 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n19011), .A(
        n21764), .ZN(n19017) );
  NAND2_X1 U21105 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19023), .ZN(
        n21133) );
  INV_X1 U21106 ( .A(n21133), .ZN(n19005) );
  OAI21_X1 U21107 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19005), .A(
        n19004), .ZN(n21149) );
  INV_X1 U21108 ( .A(n21149), .ZN(n21150) );
  INV_X1 U21109 ( .A(n19006), .ZN(n19076) );
  NOR2_X1 U21110 ( .A1(n19076), .A2(n19653), .ZN(n19072) );
  NAND2_X1 U21111 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19072), .ZN(
        n19070) );
  NOR2_X1 U21112 ( .A1(n19007), .A2(n19070), .ZN(n19037) );
  NAND2_X1 U21113 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19037), .ZN(
        n19024) );
  NAND2_X1 U21114 ( .A1(n19024), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19009) );
  NAND2_X1 U21115 ( .A1(n19097), .A2(n19098), .ZN(n19138) );
  INV_X1 U21116 ( .A(n19138), .ZN(n19073) );
  NAND2_X1 U21117 ( .A1(n22043), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n19008) );
  OAI221_X1 U21118 ( .B1(n19024), .B2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C1(
        n19009), .C2(n19073), .A(n19008), .ZN(n19015) );
  NOR2_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19010), .ZN(
        n19032) );
  INV_X1 U21120 ( .A(n19011), .ZN(n21771) );
  AOI22_X1 U21121 ( .A1(n19022), .A2(n19032), .B1(n21771), .B2(n19031), .ZN(
        n19012) );
  XOR2_X1 U21122 ( .A(n19012), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n21776) );
  AOI22_X1 U21123 ( .A1(n21990), .A2(n19074), .B1(n19047), .B2(n19013), .ZN(
        n19042) );
  OAI22_X1 U21124 ( .A1(n21776), .A2(n19057), .B1(n19042), .B2(n22024), .ZN(
        n19014) );
  AOI211_X1 U21125 ( .C1(n21150), .C2(n19137), .A(n19015), .B(n19014), .ZN(
        n19016) );
  OAI21_X1 U21126 ( .B1(n19043), .B2(n19017), .A(n19016), .ZN(P3_U2819) );
  INV_X1 U21127 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19030) );
  INV_X1 U21128 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n22049) );
  OAI221_X1 U21129 ( .B1(n19044), .B2(n19031), .C1(n22049), .C2(n19031), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19018) );
  INV_X1 U21130 ( .A(n19018), .ZN(n19021) );
  AOI221_X1 U21131 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19031), .C1(
        n22049), .C2(n19032), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19019) );
  AOI221_X1 U21132 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19021), .C1(
        n19020), .C2(n19021), .A(n19019), .ZN(n22038) );
  NOR3_X1 U21133 ( .A1(n19022), .A2(n21771), .A3(n19043), .ZN(n19028) );
  OAI21_X1 U21134 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19023), .A(
        n21133), .ZN(n21137) );
  OAI211_X1 U21135 ( .C1(n19037), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19138), .B(n19024), .ZN(n19026) );
  NAND2_X1 U21136 ( .A1(n22043), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n19025) );
  OAI211_X1 U21137 ( .C1(n19128), .C2(n21137), .A(n19026), .B(n19025), .ZN(
        n19027) );
  AOI211_X1 U21138 ( .C1(n22038), .C2(n19040), .A(n19028), .B(n19027), .ZN(
        n19029) );
  OAI21_X1 U21139 ( .B1(n19042), .B2(n19030), .A(n19029), .ZN(P3_U2820) );
  NOR2_X1 U21140 ( .A1(n19032), .A2(n19031), .ZN(n19033) );
  XOR2_X1 U21141 ( .A(n19033), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n22056) );
  INV_X1 U21142 ( .A(n22056), .ZN(n19039) );
  INV_X1 U21143 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21130) );
  NOR2_X1 U21144 ( .A1(n18767), .A2(n21130), .ZN(n22052) );
  INV_X1 U21145 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21114) );
  INV_X1 U21146 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21104) );
  NOR2_X1 U21147 ( .A1(n21114), .A2(n21104), .ZN(n19050) );
  INV_X1 U21148 ( .A(n19070), .ZN(n19034) );
  AOI22_X1 U21149 ( .A1(n19050), .A2(n19034), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19138), .ZN(n19036) );
  NAND3_X1 U21150 ( .A1(n19060), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19061) );
  NOR2_X1 U21151 ( .A1(n21114), .A2(n19061), .ZN(n21119) );
  OAI21_X1 U21152 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n21119), .A(
        n19035), .ZN(n21121) );
  OAI22_X1 U21153 ( .A1(n19037), .A2(n19036), .B1(n19128), .B2(n21121), .ZN(
        n19038) );
  AOI211_X1 U21154 ( .C1(n19040), .C2(n19039), .A(n22052), .B(n19038), .ZN(
        n19041) );
  OAI221_X1 U21155 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19043), .C1(
        n22049), .C2(n19042), .A(n19041), .ZN(P3_U2821) );
  AOI22_X1 U21156 ( .A1(n18749), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n21752), .B2(n19044), .ZN(n19045) );
  XOR2_X1 U21157 ( .A(n19046), .B(n19045), .Z(n21755) );
  INV_X1 U21158 ( .A(n21755), .ZN(n21760) );
  AOI21_X1 U21159 ( .B1(n19060), .B2(n19097), .A(n19073), .ZN(n19067) );
  AOI22_X1 U21160 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19067), .B1(
        n19047), .B2(n21760), .ZN(n19056) );
  AOI21_X1 U21161 ( .B1(n19049), .B2(n21752), .A(n19048), .ZN(n21756) );
  NAND2_X1 U21162 ( .A1(n19060), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19051) );
  AOI211_X1 U21163 ( .C1(n21114), .C2(n19051), .A(n19050), .B(n19653), .ZN(
        n19054) );
  AOI21_X1 U21164 ( .B1(n21114), .B2(n19061), .A(n21119), .ZN(n21106) );
  INV_X1 U21165 ( .A(n21106), .ZN(n19052) );
  OAI22_X1 U21166 ( .A1(n19128), .A2(n19052), .B1(n18767), .B2(n21126), .ZN(
        n19053) );
  AOI211_X1 U21167 ( .C1(n21756), .C2(n19074), .A(n19054), .B(n19053), .ZN(
        n19055) );
  OAI211_X1 U21168 ( .C1(n21760), .C2(n19057), .A(n19056), .B(n19055), .ZN(
        P3_U2822) );
  AOI21_X1 U21169 ( .B1(n19063), .B2(n19059), .A(n19058), .ZN(n21737) );
  AOI22_X1 U21170 ( .A1(n22043), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n19082), 
        .B2(n21737), .ZN(n19069) );
  NOR2_X1 U21171 ( .A1(n21074), .A2(n21012), .ZN(n19077) );
  OAI21_X1 U21172 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19077), .A(
        n19061), .ZN(n21095) );
  XOR2_X1 U21173 ( .A(n19063), .B(n19062), .Z(n19065) );
  XNOR2_X1 U21174 ( .A(n19065), .B(n19064), .ZN(n21750) );
  OAI22_X1 U21175 ( .A1(n19128), .A2(n21095), .B1(n19140), .B2(n21750), .ZN(
        n19066) );
  AOI21_X1 U21176 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19067), .A(
        n19066), .ZN(n19068) );
  OAI211_X1 U21177 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19070), .A(
        n19069), .B(n19068), .ZN(P3_U2823) );
  INV_X1 U21178 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U21179 ( .A1(n19071), .A2(n19082), .B1(n19072), .B2(n21075), .ZN(
        n19081) );
  NOR2_X1 U21180 ( .A1(n19073), .A2(n19072), .ZN(n19093) );
  AOI22_X1 U21181 ( .A1(n19075), .A2(n19074), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19093), .ZN(n19080) );
  NOR2_X1 U21182 ( .A1(n19076), .A2(n21012), .ZN(n21079) );
  INV_X1 U21183 ( .A(n21079), .ZN(n19087) );
  AOI21_X1 U21184 ( .B1(n21075), .B2(n19087), .A(n19077), .ZN(n21078) );
  NAND2_X1 U21185 ( .A1(n21078), .A2(n19137), .ZN(n19078) );
  NAND4_X1 U21186 ( .A1(n19081), .A2(n19080), .A3(n19079), .A4(n19078), .ZN(
        P3_U2824) );
  OAI21_X1 U21187 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n19084), .A(
        n19083), .ZN(n21731) );
  OAI21_X1 U21188 ( .B1(n19141), .B2(n19086), .A(n19085), .ZN(n19092) );
  NOR2_X1 U21189 ( .A1(n19086), .A2(n21012), .ZN(n21047) );
  OAI21_X1 U21190 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n21047), .A(
        n19087), .ZN(n21066) );
  OAI21_X1 U21191 ( .B1(n19090), .B2(n19089), .A(n19088), .ZN(n21730) );
  OAI22_X1 U21192 ( .A1(n19128), .A2(n21066), .B1(n19140), .B2(n21730), .ZN(
        n19091) );
  AOI21_X1 U21193 ( .B1(n19093), .B2(n19092), .A(n19091), .ZN(n19094) );
  NAND2_X1 U21194 ( .A1(n22043), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21735) );
  OAI211_X1 U21195 ( .C1(n19135), .C2(n21731), .A(n19094), .B(n21735), .ZN(
        P3_U2825) );
  INV_X1 U21196 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21057) );
  NAND2_X1 U21197 ( .A1(n19099), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19095) );
  AOI21_X1 U21198 ( .B1(n21057), .B2(n19095), .A(n21047), .ZN(n21056) );
  INV_X1 U21199 ( .A(n21056), .ZN(n21048) );
  NOR3_X1 U21200 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19113), .A3(
        n19653), .ZN(n19096) );
  AOI21_X1 U21201 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n22043), .A(n19096), .ZN(
        n19109) );
  OAI21_X1 U21202 ( .B1(n19099), .B2(n19098), .A(n19097), .ZN(n19119) );
  OAI211_X1 U21203 ( .C1(n19102), .C2(n19101), .A(n22119), .B(n19100), .ZN(
        n19107) );
  OAI211_X1 U21204 ( .C1(n19105), .C2(n19104), .A(n22117), .B(n19103), .ZN(
        n19106) );
  NAND2_X1 U21205 ( .A1(n19107), .A2(n19106), .ZN(n21722) );
  AOI22_X1 U21206 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19119), .B1(
        n22124), .B2(n21722), .ZN(n19108) );
  OAI211_X1 U21207 ( .C1(n19128), .C2(n21048), .A(n19109), .B(n19108), .ZN(
        P3_U2826) );
  OAI21_X1 U21208 ( .B1(n19112), .B2(n19111), .A(n19110), .ZN(n21712) );
  INV_X1 U21209 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21018) );
  NOR2_X1 U21210 ( .A1(n19141), .A2(n21018), .ZN(n19118) );
  NOR2_X1 U21211 ( .A1(n21018), .A2(n21012), .ZN(n19124) );
  OAI22_X1 U21212 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n19124), .B1(
        n21012), .B2(n19113), .ZN(n21040) );
  OAI21_X1 U21213 ( .B1(n19116), .B2(n19115), .A(n19114), .ZN(n21716) );
  OAI22_X1 U21214 ( .A1(n19128), .A2(n21040), .B1(n19140), .B2(n21716), .ZN(
        n19117) );
  AOI221_X1 U21215 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19119), .C1(
        n19118), .C2(n19119), .A(n19117), .ZN(n19120) );
  NAND2_X1 U21216 ( .A1(n22043), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21714) );
  OAI211_X1 U21217 ( .C1(n19135), .C2(n21712), .A(n19120), .B(n21714), .ZN(
        P3_U2827) );
  OAI21_X1 U21218 ( .B1(n19123), .B2(n19122), .A(n19121), .ZN(n21702) );
  INV_X1 U21219 ( .A(n19124), .ZN(n21022) );
  OAI21_X1 U21220 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n21022), .ZN(n21030) );
  OAI21_X1 U21221 ( .B1(n19127), .B2(n19126), .A(n19125), .ZN(n21706) );
  OAI22_X1 U21222 ( .A1(n19128), .A2(n21030), .B1(n19140), .B2(n21706), .ZN(
        n19129) );
  AOI221_X1 U21223 ( .B1(n19141), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19901), .C2(n21018), .A(n19129), .ZN(n19130) );
  NAND2_X1 U21224 ( .A1(n22043), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21704) );
  OAI211_X1 U21225 ( .C1(n19135), .C2(n21702), .A(n19130), .B(n21704), .ZN(
        P3_U2828) );
  NOR2_X1 U21226 ( .A1(n19131), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19132) );
  XNOR2_X1 U21227 ( .A(n19132), .B(n19134), .ZN(n21689) );
  INV_X1 U21228 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n21016) );
  OAI22_X1 U21229 ( .A1(n18767), .A2(n21016), .B1(n19135), .B2(n21688), .ZN(
        n19136) );
  AOI221_X1 U21230 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19138), .C1(
        n21012), .C2(n19137), .A(n19136), .ZN(n19139) );
  OAI21_X1 U21231 ( .B1(n21689), .B2(n19140), .A(n19139), .ZN(P3_U2829) );
  NOR3_X1 U21232 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19142), .A3(n19141), 
        .ZN(n19145) );
  MUX2_X1 U21233 ( .A(n22117), .B(n22119), .S(n19143), .Z(n21682) );
  AOI22_X1 U21234 ( .A1(n22043), .A2(P3_REIP_REG_0__SCAN_IN), .B1(n22124), 
        .B2(n21682), .ZN(n19144) );
  OAI21_X1 U21235 ( .B1(n19145), .B2(n21415), .A(n19144), .ZN(P3_U2830) );
  NAND2_X1 U21236 ( .A1(n22079), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19618) );
  INV_X1 U21237 ( .A(n19618), .ZN(n19619) );
  NAND2_X1 U21238 ( .A1(n22076), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19600) );
  INV_X1 U21239 ( .A(n19600), .ZN(n19601) );
  NOR2_X1 U21240 ( .A1(n19619), .A2(n19601), .ZN(n19146) );
  OAI22_X1 U21241 ( .A1(n19148), .A2(n22079), .B1(n19147), .B2(n19146), .ZN(
        P3_U2866) );
  OAI21_X1 U21242 ( .B1(n19149), .B2(n19613), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U21243 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19151), .A(
        n19150), .ZN(P3_U2864) );
  NOR4_X1 U21244 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19155) );
  NOR4_X1 U21245 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19154) );
  NOR4_X1 U21246 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19153) );
  NOR4_X1 U21247 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19152) );
  NAND4_X1 U21248 ( .A1(n19155), .A2(n19154), .A3(n19153), .A4(n19152), .ZN(
        n19161) );
  NOR4_X1 U21249 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19159) );
  AOI211_X1 U21250 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19158) );
  NOR4_X1 U21251 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19157) );
  NOR4_X1 U21252 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19156) );
  NAND4_X1 U21253 ( .A1(n19159), .A2(n19158), .A3(n19157), .A4(n19156), .ZN(
        n19160) );
  NOR2_X1 U21254 ( .A1(n19161), .A2(n19160), .ZN(n19173) );
  INV_X1 U21255 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19163) );
  OAI21_X1 U21256 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19173), .ZN(n19162) );
  OAI21_X1 U21257 ( .B1(n19173), .B2(n19163), .A(n19162), .ZN(P3_U3293) );
  INV_X1 U21258 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19166) );
  AOI21_X1 U21259 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19164) );
  OAI221_X1 U21260 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n19164), .C1(n21016), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n19173), .ZN(n19165) );
  OAI21_X1 U21261 ( .B1(n19173), .B2(n19166), .A(n19165), .ZN(P3_U3292) );
  INV_X1 U21262 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19168) );
  NOR3_X1 U21263 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19169) );
  OAI21_X1 U21264 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n19169), .A(n19173), .ZN(
        n19167) );
  OAI21_X1 U21265 ( .B1(n19173), .B2(n19168), .A(n19167), .ZN(P3_U2638) );
  INV_X1 U21266 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22417) );
  AOI21_X1 U21267 ( .B1(n21016), .B2(n22417), .A(n19169), .ZN(n19172) );
  INV_X1 U21268 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19171) );
  INV_X1 U21269 ( .A(n19173), .ZN(n19170) );
  AOI22_X1 U21270 ( .A1(n19173), .A2(n19172), .B1(n19171), .B2(n19170), .ZN(
        P3_U2639) );
  INV_X1 U21271 ( .A(n19239), .ZN(n22439) );
  INV_X1 U21272 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19241) );
  AOI22_X1 U21273 ( .A1(n22439), .A2(n19174), .B1(n19241), .B2(n19239), .ZN(
        P3_U3297) );
  OAI22_X1 U21274 ( .A1(n19239), .A2(n19175), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n22439), .ZN(n19176) );
  INV_X1 U21275 ( .A(n19176), .ZN(P3_U3294) );
  OAI21_X1 U21276 ( .B1(n19177), .B2(P3_D_C_N_REG_SCAN_IN), .A(n19239), .ZN(
        n19178) );
  OAI21_X1 U21277 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n19239), .A(n19178), 
        .ZN(P3_U2635) );
  INV_X1 U21278 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21605) );
  AOI22_X1 U21279 ( .A1(n22057), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U21280 ( .B1(n21605), .B2(n19195), .A(n19179), .ZN(P3_U2767) );
  INV_X1 U21281 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20978) );
  AOI22_X1 U21282 ( .A1(n22057), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n19180) );
  OAI21_X1 U21283 ( .B1(n20978), .B2(n19195), .A(n19180), .ZN(P3_U2766) );
  INV_X1 U21284 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21476) );
  AOI22_X1 U21285 ( .A1(n22057), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U21286 ( .B1(n21476), .B2(n19195), .A(n19181), .ZN(P3_U2765) );
  INV_X1 U21287 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20981) );
  AOI22_X1 U21288 ( .A1(n22057), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n19182) );
  OAI21_X1 U21289 ( .B1(n20981), .B2(n19195), .A(n19182), .ZN(P3_U2764) );
  INV_X1 U21290 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21431) );
  AOI22_X1 U21291 ( .A1(n22057), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U21292 ( .B1(n21431), .B2(n19195), .A(n19183), .ZN(P3_U2763) );
  INV_X1 U21293 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21430) );
  AOI22_X1 U21294 ( .A1(n22057), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U21295 ( .B1(n21430), .B2(n19195), .A(n19184), .ZN(P3_U2762) );
  INV_X1 U21296 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21458) );
  AOI22_X1 U21297 ( .A1(n22057), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U21298 ( .B1(n21458), .B2(n19195), .A(n19185), .ZN(P3_U2761) );
  INV_X1 U21299 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20986) );
  AOI22_X1 U21300 ( .A1(n22057), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U21301 ( .B1(n20986), .B2(n19195), .A(n19186), .ZN(P3_U2760) );
  INV_X1 U21302 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21585) );
  AOI22_X1 U21303 ( .A1(n22057), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U21304 ( .B1(n21585), .B2(n19195), .A(n19187), .ZN(P3_U2759) );
  INV_X1 U21305 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20989) );
  AOI22_X1 U21306 ( .A1(n19206), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U21307 ( .B1(n20989), .B2(n19195), .A(n19188), .ZN(P3_U2758) );
  INV_X1 U21308 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U21309 ( .A1(n19206), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n19189) );
  OAI21_X1 U21310 ( .B1(n20992), .B2(n19195), .A(n19189), .ZN(P3_U2757) );
  INV_X1 U21311 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21438) );
  AOI22_X1 U21312 ( .A1(n19206), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U21313 ( .B1(n21438), .B2(n19195), .A(n19190), .ZN(P3_U2756) );
  INV_X1 U21314 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U21315 ( .A1(n19206), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U21316 ( .B1(n20995), .B2(n19195), .A(n19191), .ZN(P3_U2755) );
  INV_X1 U21317 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20997) );
  AOI22_X1 U21318 ( .A1(n19206), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U21319 ( .B1(n20997), .B2(n19195), .A(n19192), .ZN(P3_U2754) );
  INV_X1 U21320 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21000) );
  AOI22_X1 U21321 ( .A1(n19206), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U21322 ( .B1(n21000), .B2(n19195), .A(n19193), .ZN(P3_U2753) );
  INV_X1 U21323 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21580) );
  AOI22_X1 U21324 ( .A1(n19206), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U21325 ( .B1(n21580), .B2(n19195), .A(n19194), .ZN(P3_U2752) );
  INV_X1 U21326 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20953) );
  NAND2_X1 U21327 ( .A1(n19197), .A2(n19196), .ZN(n19216) );
  AOI22_X1 U21328 ( .A1(n19206), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U21329 ( .B1(n20953), .B2(n19216), .A(n19198), .ZN(P3_U2751) );
  INV_X1 U21330 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20955) );
  AOI22_X1 U21331 ( .A1(n19206), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U21332 ( .B1(n20955), .B2(n19216), .A(n19199), .ZN(P3_U2750) );
  INV_X1 U21333 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20957) );
  AOI22_X1 U21334 ( .A1(n19206), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U21335 ( .B1(n20957), .B2(n19216), .A(n19200), .ZN(P3_U2749) );
  INV_X1 U21336 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21503) );
  AOI22_X1 U21337 ( .A1(n22057), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U21338 ( .B1(n21503), .B2(n19216), .A(n19201), .ZN(P3_U2748) );
  INV_X1 U21339 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20960) );
  AOI22_X1 U21340 ( .A1(n22057), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U21341 ( .B1(n20960), .B2(n19216), .A(n19202), .ZN(P3_U2747) );
  INV_X1 U21342 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21519) );
  AOI22_X1 U21343 ( .A1(n22057), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U21344 ( .B1(n21519), .B2(n19216), .A(n19203), .ZN(P3_U2746) );
  INV_X1 U21345 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n21520) );
  AOI22_X1 U21346 ( .A1(n22057), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U21347 ( .B1(n21520), .B2(n19216), .A(n19204), .ZN(P3_U2745) );
  INV_X1 U21348 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20964) );
  AOI22_X1 U21349 ( .A1(n22057), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U21350 ( .B1(n20964), .B2(n19216), .A(n19205), .ZN(P3_U2744) );
  INV_X1 U21351 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U21352 ( .A1(n19206), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U21353 ( .B1(n20966), .B2(n19216), .A(n19207), .ZN(P3_U2743) );
  INV_X1 U21354 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20968) );
  AOI22_X1 U21355 ( .A1(n22057), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n19208), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U21356 ( .B1(n20968), .B2(n19216), .A(n19209), .ZN(P3_U2742) );
  INV_X1 U21357 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21527) );
  AOI22_X1 U21358 ( .A1(n22057), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n19210) );
  OAI21_X1 U21359 ( .B1(n21527), .B2(n19216), .A(n19210), .ZN(P3_U2741) );
  INV_X1 U21360 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U21361 ( .A1(n22057), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U21362 ( .B1(n20971), .B2(n19216), .A(n19211), .ZN(P3_U2740) );
  INV_X1 U21363 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21548) );
  AOI22_X1 U21364 ( .A1(n22057), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n19212) );
  OAI21_X1 U21365 ( .B1(n21548), .B2(n19216), .A(n19212), .ZN(P3_U2739) );
  INV_X1 U21366 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U21367 ( .A1(n22057), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U21368 ( .B1(n20974), .B2(n19216), .A(n19213), .ZN(P3_U2738) );
  INV_X1 U21369 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n21540) );
  AOI22_X1 U21370 ( .A1(n22057), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n19214), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U21371 ( .B1(n21540), .B2(n19216), .A(n19215), .ZN(P3_U2737) );
  NOR2_X1 U21372 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n19217), .ZN(n19218) );
  NOR2_X1 U21373 ( .A1(n22421), .A2(n19218), .ZN(P3_U2633) );
  INV_X1 U21374 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n21017) );
  NOR2_X1 U21375 ( .A1(n19239), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19227) );
  AOI22_X1 U21376 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n19229), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n19239), .ZN(n19219) );
  OAI21_X1 U21377 ( .B1(n21017), .B2(n19233), .A(n19219), .ZN(P3_U3032) );
  INV_X1 U21378 ( .A(n19229), .ZN(n19234) );
  AOI22_X1 U21379 ( .A1(n19227), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n19239), .ZN(n19220) );
  OAI21_X1 U21380 ( .B1(n19234), .B2(n21017), .A(n19220), .ZN(P3_U3033) );
  AOI22_X1 U21381 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n19229), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n19239), .ZN(n19221) );
  OAI21_X1 U21382 ( .B1(n21060), .B2(n19233), .A(n19221), .ZN(P3_U3034) );
  AOI22_X1 U21383 ( .A1(n19227), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n19239), .ZN(n19222) );
  OAI21_X1 U21384 ( .B1(n19234), .B2(n21060), .A(n19222), .ZN(P3_U3035) );
  AOI22_X1 U21385 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n19229), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n19239), .ZN(n19223) );
  OAI21_X1 U21386 ( .B1(n19225), .B2(n19233), .A(n19223), .ZN(P3_U3036) );
  AOI22_X1 U21387 ( .A1(n19227), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n19239), .ZN(n19224) );
  OAI21_X1 U21388 ( .B1(n19225), .B2(n19234), .A(n19224), .ZN(P3_U3037) );
  AOI22_X1 U21389 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n19229), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n19239), .ZN(n19226) );
  OAI21_X1 U21390 ( .B1(n21126), .B2(n19233), .A(n19226), .ZN(P3_U3038) );
  INV_X1 U21391 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20652) );
  OAI222_X1 U21392 ( .A1(n19233), .A2(n21130), .B1(n20652), .B2(n22439), .C1(
        n21126), .C2(n19234), .ZN(P3_U3039) );
  INV_X1 U21393 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20654) );
  INV_X1 U21394 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n22041) );
  OAI222_X1 U21395 ( .A1(n21130), .A2(n19234), .B1(n20654), .B2(n22439), .C1(
        n22041), .C2(n19233), .ZN(P3_U3040) );
  AOI22_X1 U21396 ( .A1(n19227), .A2(P3_REIP_REG_11__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n19239), .ZN(n19228) );
  OAI21_X1 U21397 ( .B1(n19234), .B2(n22041), .A(n19228), .ZN(P3_U3041) );
  INV_X1 U21398 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n21171) );
  AOI22_X1 U21399 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n19229), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n19239), .ZN(n19230) );
  OAI21_X1 U21400 ( .B1(n21171), .B2(n19233), .A(n19230), .ZN(P3_U3042) );
  INV_X1 U21401 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20658) );
  OAI222_X1 U21402 ( .A1(n19233), .A2(n21180), .B1(n20658), .B2(n22439), .C1(
        n21171), .C2(n19234), .ZN(P3_U3043) );
  INV_X1 U21403 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20660) );
  OAI222_X1 U21404 ( .A1(n21180), .A2(n19234), .B1(n20660), .B2(n22439), .C1(
        n19231), .C2(n19233), .ZN(P3_U3044) );
  INV_X1 U21405 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20662) );
  OAI222_X1 U21406 ( .A1(n19231), .A2(n19234), .B1(n20662), .B2(n22439), .C1(
        n21212), .C2(n19233), .ZN(P3_U3045) );
  INV_X1 U21407 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21227) );
  INV_X1 U21408 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20664) );
  OAI222_X1 U21409 ( .A1(n19233), .A2(n21227), .B1(n20664), .B2(n22439), .C1(
        n21212), .C2(n19234), .ZN(P3_U3046) );
  INV_X1 U21410 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20666) );
  OAI222_X1 U21411 ( .A1(n19233), .A2(n21242), .B1(n20666), .B2(n22439), .C1(
        n21227), .C2(n19234), .ZN(P3_U3047) );
  INV_X1 U21412 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20668) );
  OAI222_X1 U21413 ( .A1(n21242), .A2(n19234), .B1(n20668), .B2(n22439), .C1(
        n21252), .C2(n19233), .ZN(P3_U3048) );
  INV_X1 U21414 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20670) );
  INV_X1 U21415 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n21263) );
  OAI222_X1 U21416 ( .A1(n21252), .A2(n19234), .B1(n20670), .B2(n22439), .C1(
        n21263), .C2(n19233), .ZN(P3_U3049) );
  INV_X1 U21417 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20672) );
  OAI222_X1 U21418 ( .A1(n19233), .A2(n19232), .B1(n20672), .B2(n22439), .C1(
        n21263), .C2(n19234), .ZN(P3_U3050) );
  INV_X1 U21419 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20674) );
  OAI222_X1 U21420 ( .A1(n19232), .A2(n19234), .B1(n20674), .B2(n22439), .C1(
        n21680), .C2(n19233), .ZN(P3_U3051) );
  INV_X1 U21421 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20676) );
  OAI222_X1 U21422 ( .A1(n19233), .A2(n21291), .B1(n20676), .B2(n22439), .C1(
        n21680), .C2(n19234), .ZN(P3_U3052) );
  INV_X1 U21423 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20678) );
  OAI222_X1 U21424 ( .A1(n19233), .A2(n21303), .B1(n20678), .B2(n22439), .C1(
        n21291), .C2(n19234), .ZN(P3_U3053) );
  INV_X1 U21425 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20680) );
  OAI222_X1 U21426 ( .A1(n19233), .A2(n21965), .B1(n20680), .B2(n22439), .C1(
        n21303), .C2(n19234), .ZN(P3_U3054) );
  INV_X1 U21427 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21337) );
  INV_X1 U21428 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20682) );
  OAI222_X1 U21429 ( .A1(n19233), .A2(n21337), .B1(n20682), .B2(n22439), .C1(
        n21965), .C2(n19234), .ZN(P3_U3055) );
  INV_X1 U21430 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20684) );
  OAI222_X1 U21431 ( .A1(n19233), .A2(n21359), .B1(n20684), .B2(n22439), .C1(
        n21337), .C2(n19234), .ZN(P3_U3056) );
  INV_X1 U21432 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20686) );
  OAI222_X1 U21433 ( .A1(n19233), .A2(n21862), .B1(n20686), .B2(n22439), .C1(
        n21359), .C2(n19234), .ZN(P3_U3057) );
  INV_X1 U21434 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20688) );
  OAI222_X1 U21435 ( .A1(n19233), .A2(n21940), .B1(n20688), .B2(n22439), .C1(
        n21862), .C2(n19234), .ZN(P3_U3058) );
  INV_X1 U21436 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20690) );
  OAI222_X1 U21437 ( .A1(n21940), .A2(n19234), .B1(n20690), .B2(n22439), .C1(
        n21898), .C2(n19233), .ZN(P3_U3059) );
  INV_X1 U21438 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20692) );
  OAI222_X1 U21439 ( .A1(n19233), .A2(n19235), .B1(n20692), .B2(n22439), .C1(
        n21898), .C2(n19234), .ZN(P3_U3060) );
  INV_X1 U21440 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20695) );
  INV_X1 U21441 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21409) );
  OAI222_X1 U21442 ( .A1(n19235), .A2(n19234), .B1(n20695), .B2(n22439), .C1(
        n21409), .C2(n19233), .ZN(P3_U3061) );
  OAI22_X1 U21443 ( .A1(n19239), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n22421), .ZN(n19236) );
  INV_X1 U21444 ( .A(n19236), .ZN(P3_U3277) );
  OAI22_X1 U21445 ( .A1(n19239), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n22421), .ZN(n19237) );
  INV_X1 U21446 ( .A(n19237), .ZN(P3_U3276) );
  OAI22_X1 U21447 ( .A1(n19239), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n22421), .ZN(n19238) );
  INV_X1 U21448 ( .A(n19238), .ZN(P3_U3275) );
  OAI22_X1 U21449 ( .A1(n19239), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n22421), .ZN(n19240) );
  INV_X1 U21450 ( .A(n19240), .ZN(P3_U3274) );
  NOR4_X1 U21451 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n19243)
         );
  NOR4_X1 U21452 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n19241), .ZN(n19242) );
  INV_X2 U21453 ( .A(n19897), .ZN(U215) );
  NAND3_X1 U21454 ( .A1(n19243), .A2(n19242), .A3(U215), .ZN(U213) );
  NOR2_X1 U21455 ( .A1(n20103), .A2(n19514), .ZN(n19248) );
  OAI21_X1 U21456 ( .B1(n19511), .B2(n19245), .A(n19244), .ZN(n19246) );
  AOI21_X1 U21457 ( .B1(n19247), .B2(n19248), .A(n19246), .ZN(n19258) );
  INV_X1 U21458 ( .A(n19248), .ZN(n19255) );
  NOR4_X1 U21459 ( .A1(n19249), .A2(n19252), .A3(n12819), .A4(n19251), .ZN(
        n19254) );
  AOI211_X1 U21460 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19252), .A(n19251), 
        .B(n19250), .ZN(n19253) );
  AOI211_X1 U21461 ( .C1(n19528), .C2(n19255), .A(n19254), .B(n19253), .ZN(
        n19257) );
  NAND2_X1 U21462 ( .A1(n19258), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19256) );
  OAI21_X1 U21463 ( .B1(n19258), .B2(n19257), .A(n19256), .ZN(P2_U3610) );
  NAND2_X1 U21464 ( .A1(n19505), .A2(n19461), .ZN(n19266) );
  AOI22_X1 U21465 ( .A1(n19471), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19470), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n19265) );
  NAND2_X1 U21466 ( .A1(n19473), .A2(n19260), .ZN(n19264) );
  OAI21_X1 U21467 ( .B1(n19262), .B2(n19261), .A(n12395), .ZN(n20518) );
  INV_X1 U21468 ( .A(n20518), .ZN(n19499) );
  NAND2_X1 U21469 ( .A1(n19459), .A2(n19499), .ZN(n19263) );
  NAND4_X1 U21470 ( .A1(n19266), .A2(n19265), .A3(n19264), .A4(n19263), .ZN(
        n19267) );
  AOI21_X1 U21471 ( .B1(n19269), .B2(n19268), .A(n19267), .ZN(n19271) );
  NAND2_X1 U21472 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19472), .ZN(
        n19270) );
  OAI211_X1 U21473 ( .C1(n14486), .C2(n19518), .A(n19271), .B(n19270), .ZN(
        P2_U2855) );
  AOI22_X1 U21474 ( .A1(n19272), .A2(n19473), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19470), .ZN(n19286) );
  INV_X1 U21475 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19273) );
  OAI22_X1 U21476 ( .A1(n19273), .A2(n19443), .B1(n19475), .B2(n20310), .ZN(
        n19274) );
  AOI211_X1 U21477 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19471), .A(n19360), .B(
        n19274), .ZN(n19285) );
  OAI22_X1 U21478 ( .A1(n20313), .A2(n19276), .B1(n19275), .B2(n19477), .ZN(
        n19277) );
  INV_X1 U21479 ( .A(n19277), .ZN(n19284) );
  INV_X1 U21480 ( .A(n19278), .ZN(n19282) );
  NOR2_X1 U21481 ( .A1(n11184), .A2(n19279), .ZN(n19281) );
  AOI21_X1 U21482 ( .B1(n19282), .B2(n19281), .A(n19518), .ZN(n19280) );
  OAI21_X1 U21483 ( .B1(n19282), .B2(n19281), .A(n19280), .ZN(n19283) );
  NAND4_X1 U21484 ( .A1(n19286), .A2(n19285), .A3(n19284), .A4(n19283), .ZN(
        P2_U2851) );
  INV_X1 U21485 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19297) );
  OAI22_X1 U21486 ( .A1(n19287), .A2(n19441), .B1(n12209), .B2(n19409), .ZN(
        n19288) );
  AOI211_X1 U21487 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19471), .A(n19360), .B(
        n19288), .ZN(n19296) );
  NOR2_X1 U21488 ( .A1(n11184), .A2(n19289), .ZN(n19290) );
  XNOR2_X1 U21489 ( .A(n19291), .B(n19290), .ZN(n19294) );
  OAI22_X1 U21490 ( .A1(n20210), .A2(n19475), .B1(n19292), .B2(n19477), .ZN(
        n19293) );
  AOI21_X1 U21491 ( .B1(n19294), .B2(n19481), .A(n19293), .ZN(n19295) );
  OAI211_X1 U21492 ( .C1(n19297), .C2(n19443), .A(n19296), .B(n19295), .ZN(
        P2_U2849) );
  OAI21_X1 U21493 ( .B1(n19409), .B2(n19298), .A(n14452), .ZN(n19301) );
  NOR2_X1 U21494 ( .A1(n19299), .A2(n19441), .ZN(n19300) );
  AOI211_X1 U21495 ( .C1(n19471), .C2(P2_REIP_REG_8__SCAN_IN), .A(n19301), .B(
        n19300), .ZN(n19309) );
  NOR2_X1 U21496 ( .A1(n11184), .A2(n19302), .ZN(n19303) );
  XNOR2_X1 U21497 ( .A(n19304), .B(n19303), .ZN(n19307) );
  OAI22_X1 U21498 ( .A1(n19305), .A2(n19477), .B1(n20034), .B2(n19475), .ZN(
        n19306) );
  AOI21_X1 U21499 ( .B1(n19307), .B2(n19481), .A(n19306), .ZN(n19308) );
  OAI211_X1 U21500 ( .C1(n19310), .C2(n19443), .A(n19309), .B(n19308), .ZN(
        P2_U2847) );
  AOI22_X1 U21501 ( .A1(n19311), .A2(n19473), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19470), .ZN(n19312) );
  OAI21_X1 U21502 ( .B1(n19313), .B2(n19443), .A(n19312), .ZN(n19314) );
  AOI211_X1 U21503 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19471), .A(n19360), 
        .B(n19314), .ZN(n19321) );
  AND2_X1 U21504 ( .A1(n11185), .A2(n19315), .ZN(n19317) );
  XOR2_X1 U21505 ( .A(n19317), .B(n19316), .Z(n19319) );
  AOI22_X1 U21506 ( .A1(n19319), .A2(n19481), .B1(n19318), .B2(n19461), .ZN(
        n19320) );
  OAI211_X1 U21507 ( .C1(n20028), .C2(n19475), .A(n19321), .B(n19320), .ZN(
        P2_U2845) );
  AOI22_X1 U21508 ( .A1(n19470), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19472), .ZN(n19322) );
  OAI21_X1 U21509 ( .B1(n19323), .B2(n19441), .A(n19322), .ZN(n19324) );
  AOI211_X1 U21510 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19471), .A(n19360), 
        .B(n19324), .ZN(n19330) );
  XNOR2_X1 U21511 ( .A(n19326), .B(n19325), .ZN(n19328) );
  AOI22_X1 U21512 ( .A1(n19328), .A2(n19481), .B1(n19327), .B2(n19461), .ZN(
        n19329) );
  OAI211_X1 U21513 ( .C1(n20022), .C2(n19475), .A(n19330), .B(n19329), .ZN(
        P2_U2843) );
  AOI22_X1 U21514 ( .A1(n19331), .A2(n19473), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19470), .ZN(n19332) );
  OAI21_X1 U21515 ( .B1(n11338), .B2(n19443), .A(n19332), .ZN(n19333) );
  AOI211_X1 U21516 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19471), .A(n19360), 
        .B(n19333), .ZN(n19339) );
  XOR2_X1 U21517 ( .A(n19335), .B(n19334), .Z(n19337) );
  AOI22_X1 U21518 ( .A1(n19337), .A2(n19481), .B1(n19336), .B2(n19461), .ZN(
        n19338) );
  OAI211_X1 U21519 ( .C1(n20016), .C2(n19475), .A(n19339), .B(n19338), .ZN(
        P2_U2841) );
  NOR2_X1 U21520 ( .A1(n11184), .A2(n19340), .ZN(n19341) );
  XOR2_X1 U21521 ( .A(n19342), .B(n19341), .Z(n19352) );
  AOI22_X1 U21522 ( .A1(n19343), .A2(n19473), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19470), .ZN(n19344) );
  OAI211_X1 U21523 ( .C1(n19345), .C2(n19371), .A(n19344), .B(n14452), .ZN(
        n19350) );
  INV_X1 U21524 ( .A(n19346), .ZN(n19348) );
  OAI22_X1 U21525 ( .A1(n19348), .A2(n19477), .B1(n19347), .B2(n19475), .ZN(
        n19349) );
  AOI211_X1 U21526 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19472), .A(
        n19350), .B(n19349), .ZN(n19351) );
  OAI21_X1 U21527 ( .B1(n19518), .B2(n19352), .A(n19351), .ZN(P2_U2839) );
  NAND2_X1 U21528 ( .A1(n11186), .A2(n19353), .ZN(n19354) );
  XOR2_X1 U21529 ( .A(n19355), .B(n19354), .Z(n19366) );
  AOI22_X1 U21530 ( .A1(n19356), .A2(n19473), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n19470), .ZN(n19357) );
  OAI21_X1 U21531 ( .B1(n19358), .B2(n19443), .A(n19357), .ZN(n19359) );
  AOI211_X1 U21532 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19471), .A(n19360), 
        .B(n19359), .ZN(n19365) );
  OAI22_X1 U21533 ( .A1(n19362), .A2(n19477), .B1(n19361), .B2(n19475), .ZN(
        n19363) );
  INV_X1 U21534 ( .A(n19363), .ZN(n19364) );
  OAI211_X1 U21535 ( .C1(n19518), .C2(n19366), .A(n19365), .B(n19364), .ZN(
        P2_U2838) );
  NOR2_X1 U21536 ( .A1(n11184), .A2(n19367), .ZN(n19369) );
  XOR2_X1 U21537 ( .A(n19369), .B(n19368), .Z(n19381) );
  OAI21_X1 U21538 ( .B1(n19443), .B2(n19370), .A(n14452), .ZN(n19375) );
  OAI22_X1 U21539 ( .A1(n19475), .A2(n19373), .B1(n19372), .B2(n19371), .ZN(
        n19374) );
  AOI211_X1 U21540 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19470), .A(n19375), .B(
        n19374), .ZN(n19376) );
  OAI21_X1 U21541 ( .B1(n19377), .B2(n19477), .A(n19376), .ZN(n19378) );
  AOI21_X1 U21542 ( .B1(n19379), .B2(n19473), .A(n19378), .ZN(n19380) );
  OAI21_X1 U21543 ( .B1(n19518), .B2(n19381), .A(n19380), .ZN(P2_U2837) );
  AOI22_X1 U21544 ( .A1(n19470), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19472), .ZN(n19383) );
  NAND2_X1 U21545 ( .A1(n19471), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n19382) );
  OAI211_X1 U21546 ( .C1(n19384), .C2(n19477), .A(n19383), .B(n19382), .ZN(
        n19385) );
  AOI21_X1 U21547 ( .B1(n19386), .B2(n19473), .A(n19385), .ZN(n19393) );
  INV_X1 U21548 ( .A(n19387), .ZN(n19391) );
  NOR2_X1 U21549 ( .A1(n11184), .A2(n19388), .ZN(n19390) );
  NAND2_X1 U21550 ( .A1(n19391), .A2(n19390), .ZN(n19389) );
  OAI211_X1 U21551 ( .C1(n19391), .C2(n19390), .A(n19481), .B(n19389), .ZN(
        n19392) );
  OAI211_X1 U21552 ( .C1(n19475), .C2(n19394), .A(n19393), .B(n19392), .ZN(
        P2_U2835) );
  AOI22_X1 U21553 ( .A1(n19471), .A2(P2_REIP_REG_21__SCAN_IN), .B1(n19470), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n19407) );
  AOI22_X1 U21554 ( .A1(n19395), .A2(n19473), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19472), .ZN(n19406) );
  INV_X1 U21555 ( .A(n19396), .ZN(n19397) );
  OAI22_X1 U21556 ( .A1(n19398), .A2(n19477), .B1(n19475), .B2(n19397), .ZN(
        n19399) );
  INV_X1 U21557 ( .A(n19399), .ZN(n19405) );
  NAND2_X1 U21558 ( .A1(n11185), .A2(n19400), .ZN(n19402) );
  NAND2_X1 U21559 ( .A1(n19403), .A2(n19402), .ZN(n19401) );
  OAI211_X1 U21560 ( .C1(n19403), .C2(n19402), .A(n19481), .B(n19401), .ZN(
        n19404) );
  NAND4_X1 U21561 ( .A1(n19407), .A2(n19406), .A3(n19405), .A4(n19404), .ZN(
        P2_U2834) );
  INV_X1 U21562 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n19408) );
  OAI22_X1 U21563 ( .A1(n19409), .A2(n12271), .B1(n19443), .B2(n19408), .ZN(
        n19410) );
  AOI21_X1 U21564 ( .B1(P2_REIP_REG_22__SCAN_IN), .B2(n19471), .A(n19410), 
        .ZN(n19411) );
  OAI21_X1 U21565 ( .B1(n19412), .B2(n19477), .A(n19411), .ZN(n19413) );
  AOI21_X1 U21566 ( .B1(n19414), .B2(n19473), .A(n19413), .ZN(n19419) );
  OAI211_X1 U21567 ( .C1(n19417), .C2(n19416), .A(n19481), .B(n19415), .ZN(
        n19418) );
  OAI211_X1 U21568 ( .C1(n19475), .C2(n19420), .A(n19419), .B(n19418), .ZN(
        P2_U2833) );
  AOI22_X1 U21569 ( .A1(n19471), .A2(P2_REIP_REG_25__SCAN_IN), .B1(n19470), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n19431) );
  AOI22_X1 U21570 ( .A1(n19421), .A2(n19473), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19472), .ZN(n19430) );
  INV_X1 U21571 ( .A(n19422), .ZN(n19423) );
  AOI22_X1 U21572 ( .A1(n19424), .A2(n19461), .B1(n19423), .B2(n19459), .ZN(
        n19429) );
  OAI211_X1 U21573 ( .C1(n19427), .C2(n19426), .A(n19481), .B(n19425), .ZN(
        n19428) );
  NAND4_X1 U21574 ( .A1(n19431), .A2(n19430), .A3(n19429), .A4(n19428), .ZN(
        P2_U2830) );
  AOI22_X1 U21575 ( .A1(n19471), .A2(P2_REIP_REG_26__SCAN_IN), .B1(n19470), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n19440) );
  AOI22_X1 U21576 ( .A1(n12100), .A2(n19473), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19472), .ZN(n19439) );
  AOI22_X1 U21577 ( .A1(n19433), .A2(n19461), .B1(n19432), .B2(n19459), .ZN(
        n19438) );
  OAI211_X1 U21578 ( .C1(n19436), .C2(n19435), .A(n19481), .B(n19434), .ZN(
        n19437) );
  NAND4_X1 U21579 ( .A1(n19440), .A2(n19439), .A3(n19438), .A4(n19437), .ZN(
        P2_U2829) );
  OR2_X1 U21580 ( .A1(n19442), .A2(n19441), .ZN(n19449) );
  NOR2_X1 U21581 ( .A1(n19443), .A2(n14204), .ZN(n19444) );
  AOI21_X1 U21582 ( .B1(n19470), .B2(P2_EBX_REG_28__SCAN_IN), .A(n19444), .ZN(
        n19448) );
  NAND2_X1 U21583 ( .A1(n19445), .A2(n19461), .ZN(n19447) );
  NAND2_X1 U21584 ( .A1(n19471), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n19446) );
  OAI211_X1 U21585 ( .C1(n19452), .C2(n19451), .A(n19481), .B(n19450), .ZN(
        n19453) );
  OAI211_X1 U21586 ( .C1(n19475), .C2(n19455), .A(n19454), .B(n19453), .ZN(
        P2_U2827) );
  AOI22_X1 U21587 ( .A1(n19471), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n19470), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n19469) );
  AOI22_X1 U21588 ( .A1(n19456), .A2(n19473), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19472), .ZN(n19468) );
  INV_X1 U21589 ( .A(n19457), .ZN(n19462) );
  INV_X1 U21590 ( .A(n19458), .ZN(n19460) );
  AOI22_X1 U21591 ( .A1(n19462), .A2(n19461), .B1(n19460), .B2(n19459), .ZN(
        n19467) );
  OAI211_X1 U21592 ( .C1(n19465), .C2(n19464), .A(n19481), .B(n19463), .ZN(
        n19466) );
  NAND4_X1 U21593 ( .A1(n19469), .A2(n19468), .A3(n19467), .A4(n19466), .ZN(
        P2_U2826) );
  AOI22_X1 U21594 ( .A1(n19471), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n19470), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n19487) );
  AOI22_X1 U21595 ( .A1(n19474), .A2(n19473), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19472), .ZN(n19486) );
  OAI22_X1 U21596 ( .A1(n19478), .A2(n19477), .B1(n19476), .B2(n19475), .ZN(
        n19479) );
  INV_X1 U21597 ( .A(n19479), .ZN(n19485) );
  OAI211_X1 U21598 ( .C1(n19483), .C2(n19482), .A(n19481), .B(n19480), .ZN(
        n19484) );
  NAND4_X1 U21599 ( .A1(n19487), .A2(n19486), .A3(n19485), .A4(n19484), .ZN(
        P2_U2825) );
  NOR2_X1 U21600 ( .A1(n19488), .A2(n19512), .ZN(n19489) );
  OAI21_X1 U21601 ( .B1(n19493), .B2(n19492), .A(n19491), .ZN(P2_U3595) );
  OAI22_X1 U21602 ( .A1(n19497), .A2(n19496), .B1(n19495), .B2(n19494), .ZN(
        n19498) );
  AOI21_X1 U21603 ( .B1(n19500), .B2(n19499), .A(n19498), .ZN(n19501) );
  OAI21_X1 U21604 ( .B1(n19502), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19501), .ZN(n19503) );
  AOI21_X1 U21605 ( .B1(n19505), .B2(n19504), .A(n19503), .ZN(n19507) );
  OAI211_X1 U21606 ( .C1(n19509), .C2(n19508), .A(n19507), .B(n19506), .ZN(
        P2_U3046) );
  NAND2_X1 U21607 ( .A1(n19527), .A2(n19510), .ZN(n19532) );
  INV_X1 U21608 ( .A(n19511), .ZN(n19536) );
  OAI21_X1 U21609 ( .B1(n19513), .B2(n19512), .A(n19536), .ZN(n19517) );
  NAND2_X1 U21610 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19514), .ZN(n19515) );
  AOI21_X1 U21611 ( .B1(n19521), .B2(n19532), .A(n19515), .ZN(n19516) );
  AOI21_X1 U21612 ( .B1(n19532), .B2(n19517), .A(n19516), .ZN(n19519) );
  NAND2_X1 U21613 ( .A1(n19519), .A2(n19518), .ZN(P2_U3177) );
  INV_X1 U21614 ( .A(n19520), .ZN(n19535) );
  OAI22_X1 U21615 ( .A1(n19523), .A2(n19522), .B1(n19531), .B2(n19521), .ZN(
        n19525) );
  OR2_X1 U21616 ( .A1(n19525), .A2(n19524), .ZN(n19526) );
  AOI21_X1 U21617 ( .B1(n19527), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19526), 
        .ZN(n19534) );
  OAI21_X1 U21618 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19529), .A(n19528), 
        .ZN(n19530) );
  OAI21_X1 U21619 ( .B1(n19532), .B2(n19531), .A(n19530), .ZN(n19533) );
  OAI211_X1 U21620 ( .C1(n19535), .C2(n19536), .A(n19534), .B(n19533), .ZN(
        P2_U3176) );
  NOR2_X1 U21621 ( .A1(n19537), .A2(n19536), .ZN(n19541) );
  MUX2_X1 U21622 ( .A(P2_MORE_REG_SCAN_IN), .B(n19538), .S(n19541), .Z(
        P2_U3609) );
  OAI21_X1 U21623 ( .B1(n19541), .B2(n19540), .A(n19539), .ZN(P2_U2819) );
  INV_X1 U21624 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20934) );
  AOI22_X1 U21625 ( .A1(n19897), .A2(n20934), .B1(n19569), .B2(U215), .ZN(U282) );
  OAI22_X1 U21626 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19897), .ZN(n19542) );
  INV_X1 U21627 ( .A(n19542), .ZN(U281) );
  OAI22_X1 U21628 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19897), .ZN(n19543) );
  INV_X1 U21629 ( .A(n19543), .ZN(U280) );
  OAI22_X1 U21630 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19897), .ZN(n19544) );
  INV_X1 U21631 ( .A(n19544), .ZN(U279) );
  OAI22_X1 U21632 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19897), .ZN(n19545) );
  INV_X1 U21633 ( .A(n19545), .ZN(U278) );
  OAI22_X1 U21634 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19897), .ZN(n19546) );
  INV_X1 U21635 ( .A(n19546), .ZN(U277) );
  OAI22_X1 U21636 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19897), .ZN(n19547) );
  INV_X1 U21637 ( .A(n19547), .ZN(U276) );
  OAI22_X1 U21638 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19897), .ZN(n19548) );
  INV_X1 U21639 ( .A(n19548), .ZN(U275) );
  OAI22_X1 U21640 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19897), .ZN(n19549) );
  INV_X1 U21641 ( .A(n19549), .ZN(U274) );
  OAI22_X1 U21642 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19897), .ZN(n19550) );
  INV_X1 U21643 ( .A(n19550), .ZN(U273) );
  OAI22_X1 U21644 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19897), .ZN(n19551) );
  INV_X1 U21645 ( .A(n19551), .ZN(U272) );
  OAI22_X1 U21646 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19897), .ZN(n19552) );
  INV_X1 U21647 ( .A(n19552), .ZN(U271) );
  OAI22_X1 U21648 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19565), .ZN(n19553) );
  INV_X1 U21649 ( .A(n19553), .ZN(U270) );
  OAI22_X1 U21650 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19897), .ZN(n19554) );
  INV_X1 U21651 ( .A(n19554), .ZN(U269) );
  OAI22_X1 U21652 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19565), .ZN(n19555) );
  INV_X1 U21653 ( .A(n19555), .ZN(U268) );
  OAI22_X1 U21654 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19897), .ZN(n19556) );
  INV_X1 U21655 ( .A(n19556), .ZN(U267) );
  OAI22_X1 U21656 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19565), .ZN(n19557) );
  INV_X1 U21657 ( .A(n19557), .ZN(U266) );
  OAI22_X1 U21658 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19897), .ZN(n19558) );
  INV_X1 U21659 ( .A(n19558), .ZN(U265) );
  OAI22_X1 U21660 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19565), .ZN(n19559) );
  INV_X1 U21661 ( .A(n19559), .ZN(U264) );
  OAI22_X1 U21662 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19565), .ZN(n19560) );
  INV_X1 U21663 ( .A(n19560), .ZN(U263) );
  OAI22_X1 U21664 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19565), .ZN(n19561) );
  INV_X1 U21665 ( .A(n19561), .ZN(U262) );
  OAI22_X1 U21666 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19565), .ZN(n19562) );
  INV_X1 U21667 ( .A(n19562), .ZN(U261) );
  OAI22_X1 U21668 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19565), .ZN(n19563) );
  INV_X1 U21669 ( .A(n19563), .ZN(U260) );
  OAI22_X1 U21670 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19565), .ZN(n19564) );
  INV_X1 U21671 ( .A(n19564), .ZN(U259) );
  OAI22_X1 U21672 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19565), .ZN(n19566) );
  INV_X1 U21673 ( .A(n19566), .ZN(U258) );
  NOR2_X1 U21674 ( .A1(n22079), .A2(n19594), .ZN(n19639) );
  NAND2_X1 U21675 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19639), .ZN(
        n19991) );
  NOR2_X1 U21676 ( .A1(n19568), .A2(n19567), .ZN(n19691) );
  NAND2_X1 U21677 ( .A1(n19691), .A2(n21521), .ZN(n19650) );
  NOR3_X1 U21678 ( .A1(n22076), .A2(n22079), .A3(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19578) );
  NAND2_X1 U21679 ( .A1(n19617), .A2(n19578), .ZN(n19818) );
  INV_X1 U21680 ( .A(n19818), .ZN(n19921) );
  NOR2_X2 U21681 ( .A1(n19569), .A2(n19653), .ZN(n19647) );
  INV_X1 U21682 ( .A(n19628), .ZN(n22092) );
  AND2_X1 U21683 ( .A1(n22092), .A2(n19639), .ZN(n19903) );
  INV_X1 U21684 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21461) );
  NOR2_X2 U21685 ( .A1(n21461), .A2(n19902), .ZN(n19642) );
  AOI22_X1 U21686 ( .A1(n19921), .A2(n19647), .B1(n19903), .B2(n19642), .ZN(
        n19573) );
  NAND2_X1 U21687 ( .A1(n19570), .A2(n19854), .ZN(n19579) );
  INV_X1 U21688 ( .A(n19579), .ZN(n19591) );
  AOI22_X1 U21689 ( .A1(n19901), .A2(n19578), .B1(n19639), .B2(n19591), .ZN(
        n19907) );
  NAND2_X1 U21690 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19578), .ZN(
        n20002) );
  INV_X1 U21691 ( .A(n20002), .ZN(n19916) );
  INV_X1 U21692 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19571) );
  NOR2_X2 U21693 ( .A1(n19571), .A2(n19653), .ZN(n19643) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19907), .B1(
        n19916), .B2(n19643), .ZN(n19572) );
  OAI211_X1 U21695 ( .C1(n19991), .C2(n19650), .A(n19573), .B(n19572), .ZN(
        P3_U2995) );
  NAND2_X1 U21696 ( .A1(n19639), .A2(n19617), .ZN(n19896) );
  NAND2_X1 U21697 ( .A1(n20002), .A2(n19896), .ZN(n19646) );
  INV_X1 U21698 ( .A(n19646), .ZN(n19574) );
  NOR2_X1 U21699 ( .A1(n19628), .A2(n19574), .ZN(n19910) );
  AOI22_X1 U21700 ( .A1(n19643), .A2(n19921), .B1(n19642), .B2(n19910), .ZN(
        n19577) );
  INV_X1 U21701 ( .A(n19896), .ZN(n19995) );
  NOR2_X1 U21702 ( .A1(n22069), .A2(n19600), .ZN(n19590) );
  NAND2_X1 U21703 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19590), .ZN(
        n19914) );
  NAND2_X1 U21704 ( .A1(n19818), .A2(n19914), .ZN(n19585) );
  INV_X1 U21705 ( .A(n19585), .ZN(n19583) );
  OAI21_X1 U21706 ( .B1(n19583), .B2(n19596), .A(n19574), .ZN(n19575) );
  OAI211_X1 U21707 ( .C1(n19995), .C2(n22100), .A(n19854), .B(n19575), .ZN(
        n19911) );
  INV_X1 U21708 ( .A(n19914), .ZN(n19927) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19911), .B1(
        n19647), .B2(n19927), .ZN(n19576) );
  OAI211_X1 U21710 ( .C1(n19650), .C2(n19896), .A(n19577), .B(n19576), .ZN(
        P3_U2987) );
  NAND2_X1 U21711 ( .A1(n19617), .A2(n19590), .ZN(n19925) );
  AND2_X1 U21712 ( .A1(n22092), .A2(n19578), .ZN(n19915) );
  AOI22_X1 U21713 ( .A1(n19647), .A2(n19933), .B1(n19642), .B2(n19915), .ZN(
        n19582) );
  NOR2_X1 U21714 ( .A1(n22076), .A2(n22079), .ZN(n19580) );
  NOR2_X1 U21715 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19579), .ZN(
        n19638) );
  AOI22_X1 U21716 ( .A1(n19901), .A2(n19590), .B1(n19580), .B2(n19638), .ZN(
        n19917) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19917), .B1(
        n19643), .B2(n19927), .ZN(n19581) );
  OAI211_X1 U21718 ( .C1(n20002), .C2(n19650), .A(n19582), .B(n19581), .ZN(
        P3_U2979) );
  NOR2_X1 U21719 ( .A1(n19628), .A2(n19583), .ZN(n19920) );
  AOI22_X1 U21720 ( .A1(n19643), .A2(n19933), .B1(n19642), .B2(n19920), .ZN(
        n19588) );
  NOR2_X1 U21721 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19617), .ZN(
        n19622) );
  NAND2_X1 U21722 ( .A1(n19601), .A2(n19622), .ZN(n19931) );
  INV_X1 U21723 ( .A(n19931), .ZN(n19939) );
  NOR2_X1 U21724 ( .A1(n19933), .A2(n19939), .ZN(n19595) );
  INV_X1 U21725 ( .A(n19595), .ZN(n19586) );
  NOR2_X1 U21726 ( .A1(n19902), .A2(n19584), .ZN(n19645) );
  AOI22_X1 U21727 ( .A1(n19901), .A2(n19586), .B1(n19645), .B2(n19585), .ZN(
        n19922) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19922), .B1(
        n19647), .B2(n19939), .ZN(n19587) );
  OAI211_X1 U21729 ( .C1(n19650), .C2(n19818), .A(n19588), .B(n19587), .ZN(
        P3_U2971) );
  INV_X1 U21730 ( .A(n19590), .ZN(n19589) );
  NOR2_X1 U21731 ( .A1(n19628), .A2(n19589), .ZN(n19926) );
  AOI22_X1 U21732 ( .A1(n19643), .A2(n19939), .B1(n19642), .B2(n19926), .ZN(
        n19593) );
  AOI22_X1 U21733 ( .A1(n19901), .A2(n19601), .B1(n19591), .B2(n19590), .ZN(
        n19928) );
  NAND2_X1 U21734 ( .A1(n22069), .A2(n19617), .ZN(n22072) );
  NOR2_X2 U21735 ( .A1(n22072), .A2(n19600), .ZN(n19945) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19928), .B1(
        n19647), .B2(n19945), .ZN(n19592) );
  OAI211_X1 U21737 ( .C1(n19650), .C2(n19914), .A(n19593), .B(n19592), .ZN(
        P3_U2963) );
  NOR2_X1 U21738 ( .A1(n19628), .A2(n19595), .ZN(n19932) );
  AOI22_X1 U21739 ( .A1(n19643), .A2(n19945), .B1(n19642), .B2(n19932), .ZN(
        n19599) );
  INV_X1 U21740 ( .A(n19945), .ZN(n19937) );
  NOR2_X1 U21741 ( .A1(n19594), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19608) );
  NAND2_X1 U21742 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19608), .ZN(
        n19943) );
  NAND2_X1 U21743 ( .A1(n19937), .A2(n19943), .ZN(n19605) );
  INV_X1 U21744 ( .A(n19605), .ZN(n19604) );
  OAI21_X1 U21745 ( .B1(n19604), .B2(n19596), .A(n19595), .ZN(n19597) );
  OAI211_X1 U21746 ( .C1(n19933), .C2(n22100), .A(n19854), .B(n19597), .ZN(
        n19934) );
  INV_X1 U21747 ( .A(n19943), .ZN(n19951) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19934), .B1(
        n19647), .B2(n19951), .ZN(n19598) );
  OAI211_X1 U21749 ( .C1(n19650), .C2(n19925), .A(n19599), .B(n19598), .ZN(
        P3_U2955) );
  NAND2_X1 U21750 ( .A1(n22069), .A2(n22092), .ZN(n19636) );
  NOR2_X1 U21751 ( .A1(n19600), .A2(n19636), .ZN(n19938) );
  AOI22_X1 U21752 ( .A1(n19643), .A2(n19951), .B1(n19642), .B2(n19938), .ZN(
        n19603) );
  AOI22_X1 U21753 ( .A1(n19901), .A2(n19608), .B1(n19601), .B2(n19638), .ZN(
        n19940) );
  NAND2_X1 U21754 ( .A1(n19617), .A2(n19608), .ZN(n19949) );
  INV_X1 U21755 ( .A(n19949), .ZN(n19957) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19940), .B1(
        n19647), .B2(n19957), .ZN(n19602) );
  OAI211_X1 U21757 ( .C1(n19650), .C2(n19931), .A(n19603), .B(n19602), .ZN(
        P3_U2947) );
  NOR2_X1 U21758 ( .A1(n19628), .A2(n19604), .ZN(n19944) );
  AOI22_X1 U21759 ( .A1(n19643), .A2(n19957), .B1(n19642), .B2(n19944), .ZN(
        n19607) );
  NAND2_X1 U21760 ( .A1(n19619), .A2(n19622), .ZN(n19874) );
  NAND2_X1 U21761 ( .A1(n19949), .A2(n19874), .ZN(n19614) );
  AOI22_X1 U21762 ( .A1(n19901), .A2(n19614), .B1(n19645), .B2(n19605), .ZN(
        n19946) );
  INV_X1 U21763 ( .A(n19874), .ZN(n19963) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19946), .B1(
        n19647), .B2(n19963), .ZN(n19606) );
  OAI211_X1 U21765 ( .C1(n19650), .C2(n19937), .A(n19607), .B(n19606), .ZN(
        P3_U2939) );
  NOR2_X2 U21766 ( .A1(n22072), .A2(n19618), .ZN(n19968) );
  INV_X1 U21767 ( .A(n19608), .ZN(n19609) );
  NOR2_X1 U21768 ( .A1(n19628), .A2(n19609), .ZN(n19950) );
  AOI22_X1 U21769 ( .A1(n19647), .A2(n19968), .B1(n19642), .B2(n19950), .ZN(
        n19612) );
  NAND2_X1 U21770 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22068) );
  OAI21_X1 U21771 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19613), .A(
        n19854), .ZN(n19610) );
  AOI21_X1 U21772 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n22068), .A(n19610), 
        .ZN(n19629) );
  NAND2_X1 U21773 ( .A1(n19619), .A2(n19629), .ZN(n19952) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19952), .B1(
        n19643), .B2(n19963), .ZN(n19611) );
  OAI211_X1 U21775 ( .C1(n19650), .C2(n19943), .A(n19612), .B(n19611), .ZN(
        P3_U2931) );
  NAND2_X1 U21776 ( .A1(n22076), .A2(n22079), .ZN(n19635) );
  NOR2_X1 U21777 ( .A1(n22069), .A2(n19635), .ZN(n19626) );
  NAND2_X1 U21778 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19626), .ZN(
        n19961) );
  INV_X1 U21779 ( .A(n19961), .ZN(n19974) );
  AND2_X1 U21780 ( .A1(n22092), .A2(n19614), .ZN(n19956) );
  AOI22_X1 U21781 ( .A1(n19647), .A2(n19974), .B1(n19642), .B2(n19956), .ZN(
        n19616) );
  INV_X1 U21782 ( .A(n19968), .ZN(n19955) );
  NAND2_X1 U21783 ( .A1(n19955), .A2(n19961), .ZN(n19623) );
  OAI221_X1 U21784 ( .B1(n19614), .B2(n19613), .C1(n19614), .C2(n19623), .A(
        n19645), .ZN(n19958) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19958), .B1(
        n19643), .B2(n19968), .ZN(n19615) );
  OAI211_X1 U21786 ( .C1(n19650), .C2(n19949), .A(n19616), .B(n19615), .ZN(
        P3_U2923) );
  NAND2_X1 U21787 ( .A1(n19617), .A2(n19626), .ZN(n19972) );
  INV_X1 U21788 ( .A(n19972), .ZN(n19980) );
  NOR2_X1 U21789 ( .A1(n19618), .A2(n19636), .ZN(n19962) );
  AOI22_X1 U21790 ( .A1(n19647), .A2(n19980), .B1(n19642), .B2(n19962), .ZN(
        n19621) );
  AOI22_X1 U21791 ( .A1(n19901), .A2(n19626), .B1(n19619), .B2(n19638), .ZN(
        n19964) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19964), .B1(
        n19643), .B2(n19974), .ZN(n19620) );
  OAI211_X1 U21793 ( .C1(n19650), .C2(n19874), .A(n19621), .B(n19620), .ZN(
        P3_U2915) );
  INV_X1 U21794 ( .A(n19635), .ZN(n19637) );
  NAND2_X1 U21795 ( .A1(n19622), .A2(n19637), .ZN(n19881) );
  INV_X1 U21796 ( .A(n19881), .ZN(n19986) );
  AND2_X1 U21797 ( .A1(n22092), .A2(n19623), .ZN(n19967) );
  AOI22_X1 U21798 ( .A1(n19647), .A2(n19986), .B1(n19642), .B2(n19967), .ZN(
        n19625) );
  NAND2_X1 U21799 ( .A1(n19972), .A2(n19881), .ZN(n19632) );
  AOI22_X1 U21800 ( .A1(n19901), .A2(n19632), .B1(n19645), .B2(n19623), .ZN(
        n19969) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19969), .B1(
        n19643), .B2(n19980), .ZN(n19624) );
  OAI211_X1 U21802 ( .C1(n19650), .C2(n19955), .A(n19625), .B(n19624), .ZN(
        P3_U2907) );
  NOR2_X2 U21803 ( .A1(n22072), .A2(n19635), .ZN(n19997) );
  INV_X1 U21804 ( .A(n19626), .ZN(n19627) );
  NOR2_X1 U21805 ( .A1(n19628), .A2(n19627), .ZN(n19973) );
  AOI22_X1 U21806 ( .A1(n19647), .A2(n19997), .B1(n19642), .B2(n19973), .ZN(
        n19631) );
  NAND2_X1 U21807 ( .A1(n19629), .A2(n19637), .ZN(n19975) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19975), .B1(
        n19643), .B2(n19986), .ZN(n19630) );
  OAI211_X1 U21809 ( .C1(n19650), .C2(n19961), .A(n19631), .B(n19630), .ZN(
        P3_U2899) );
  AND2_X1 U21810 ( .A1(n22092), .A2(n19632), .ZN(n19979) );
  AOI22_X1 U21811 ( .A1(n19643), .A2(n19997), .B1(n19642), .B2(n19979), .ZN(
        n19634) );
  INV_X1 U21812 ( .A(n19997), .ZN(n19978) );
  NAND2_X1 U21813 ( .A1(n19991), .A2(n19978), .ZN(n19644) );
  AOI22_X1 U21814 ( .A1(n19901), .A2(n19644), .B1(n19645), .B2(n19632), .ZN(
        n19981) );
  INV_X1 U21815 ( .A(n19991), .ZN(n19906) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19981), .B1(
        n19906), .B2(n19647), .ZN(n19633) );
  OAI211_X1 U21817 ( .C1(n19650), .C2(n19972), .A(n19634), .B(n19633), .ZN(
        P3_U2891) );
  NOR2_X1 U21818 ( .A1(n19636), .A2(n19635), .ZN(n19984) );
  AOI22_X1 U21819 ( .A1(n19643), .A2(n19906), .B1(n19642), .B2(n19984), .ZN(
        n19641) );
  AOI22_X1 U21820 ( .A1(n19901), .A2(n19639), .B1(n19638), .B2(n19637), .ZN(
        n19987) );
  AOI22_X1 U21821 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19987), .B1(
        n19647), .B2(n19995), .ZN(n19640) );
  OAI211_X1 U21822 ( .C1(n19650), .C2(n19881), .A(n19641), .B(n19640), .ZN(
        P3_U2883) );
  AND2_X1 U21823 ( .A1(n22092), .A2(n19644), .ZN(n19993) );
  AOI22_X1 U21824 ( .A1(n19643), .A2(n19995), .B1(n19642), .B2(n19993), .ZN(
        n19649) );
  AOI22_X1 U21825 ( .A1(n19901), .A2(n19646), .B1(n19645), .B2(n19644), .ZN(
        n19998) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19998), .B1(
        n19916), .B2(n19647), .ZN(n19648) );
  OAI211_X1 U21827 ( .C1(n19650), .C2(n19978), .A(n19649), .B(n19648), .ZN(
        P3_U2875) );
  OAI22_X1 U21828 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19897), .ZN(n19651) );
  INV_X1 U21829 ( .A(n19651), .ZN(U257) );
  NAND2_X1 U21830 ( .A1(n19691), .A2(n19652), .ZN(n19689) );
  NOR2_X2 U21831 ( .A1(n12999), .A2(n19653), .ZN(n19686) );
  INV_X1 U21832 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21466) );
  NOR2_X2 U21833 ( .A1(n21466), .A2(n19902), .ZN(n19684) );
  AOI22_X1 U21834 ( .A1(n19921), .A2(n19686), .B1(n19903), .B2(n19684), .ZN(
        n19655) );
  INV_X1 U21835 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n21496) );
  NOR2_X2 U21836 ( .A1(n21496), .A2(n19653), .ZN(n19685) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19907), .B1(
        n19916), .B2(n19685), .ZN(n19654) );
  OAI211_X1 U21838 ( .C1(n19991), .C2(n19689), .A(n19655), .B(n19654), .ZN(
        P3_U2994) );
  AOI22_X1 U21839 ( .A1(n19927), .A2(n19686), .B1(n19910), .B2(n19684), .ZN(
        n19657) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19911), .B1(
        n19921), .B2(n19685), .ZN(n19656) );
  OAI211_X1 U21841 ( .C1(n19896), .C2(n19689), .A(n19657), .B(n19656), .ZN(
        P3_U2986) );
  AOI22_X1 U21842 ( .A1(n19927), .A2(n19685), .B1(n19915), .B2(n19684), .ZN(
        n19659) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19917), .B1(
        n19933), .B2(n19686), .ZN(n19658) );
  OAI211_X1 U21844 ( .C1(n20002), .C2(n19689), .A(n19659), .B(n19658), .ZN(
        P3_U2978) );
  AOI22_X1 U21845 ( .A1(n19939), .A2(n19686), .B1(n19920), .B2(n19684), .ZN(
        n19661) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19922), .B1(
        n19933), .B2(n19685), .ZN(n19660) );
  OAI211_X1 U21847 ( .C1(n19818), .C2(n19689), .A(n19661), .B(n19660), .ZN(
        P3_U2970) );
  AOI22_X1 U21848 ( .A1(n19945), .A2(n19686), .B1(n19926), .B2(n19684), .ZN(
        n19663) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19928), .B1(
        n19939), .B2(n19685), .ZN(n19662) );
  OAI211_X1 U21850 ( .C1(n19914), .C2(n19689), .A(n19663), .B(n19662), .ZN(
        P3_U2962) );
  AOI22_X1 U21851 ( .A1(n19951), .A2(n19686), .B1(n19932), .B2(n19684), .ZN(
        n19665) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19934), .B1(
        n19945), .B2(n19685), .ZN(n19664) );
  OAI211_X1 U21853 ( .C1(n19925), .C2(n19689), .A(n19665), .B(n19664), .ZN(
        P3_U2954) );
  AOI22_X1 U21854 ( .A1(n19951), .A2(n19685), .B1(n19938), .B2(n19684), .ZN(
        n19667) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19940), .B1(
        n19957), .B2(n19686), .ZN(n19666) );
  OAI211_X1 U21856 ( .C1(n19931), .C2(n19689), .A(n19667), .B(n19666), .ZN(
        P3_U2946) );
  AOI22_X1 U21857 ( .A1(n19963), .A2(n19686), .B1(n19944), .B2(n19684), .ZN(
        n19669) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19946), .B1(
        n19957), .B2(n19685), .ZN(n19668) );
  OAI211_X1 U21859 ( .C1(n19937), .C2(n19689), .A(n19669), .B(n19668), .ZN(
        P3_U2938) );
  AOI22_X1 U21860 ( .A1(n19950), .A2(n19684), .B1(n19968), .B2(n19686), .ZN(
        n19671) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19952), .B1(
        n19963), .B2(n19685), .ZN(n19670) );
  OAI211_X1 U21862 ( .C1(n19943), .C2(n19689), .A(n19671), .B(n19670), .ZN(
        P3_U2930) );
  AOI22_X1 U21863 ( .A1(n19974), .A2(n19686), .B1(n19956), .B2(n19684), .ZN(
        n19673) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19958), .B1(
        n19968), .B2(n19685), .ZN(n19672) );
  OAI211_X1 U21865 ( .C1(n19949), .C2(n19689), .A(n19673), .B(n19672), .ZN(
        P3_U2922) );
  AOI22_X1 U21866 ( .A1(n19980), .A2(n19686), .B1(n19962), .B2(n19684), .ZN(
        n19675) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19964), .B1(
        n19974), .B2(n19685), .ZN(n19674) );
  OAI211_X1 U21868 ( .C1(n19874), .C2(n19689), .A(n19675), .B(n19674), .ZN(
        P3_U2914) );
  AOI22_X1 U21869 ( .A1(n19986), .A2(n19686), .B1(n19967), .B2(n19684), .ZN(
        n19677) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19969), .B1(
        n19980), .B2(n19685), .ZN(n19676) );
  OAI211_X1 U21871 ( .C1(n19955), .C2(n19689), .A(n19677), .B(n19676), .ZN(
        P3_U2906) );
  AOI22_X1 U21872 ( .A1(n19997), .A2(n19686), .B1(n19973), .B2(n19684), .ZN(
        n19679) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19975), .B1(
        n19986), .B2(n19685), .ZN(n19678) );
  OAI211_X1 U21874 ( .C1(n19961), .C2(n19689), .A(n19679), .B(n19678), .ZN(
        P3_U2898) );
  AOI22_X1 U21875 ( .A1(n19997), .A2(n19685), .B1(n19979), .B2(n19684), .ZN(
        n19681) );
  AOI22_X1 U21876 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19981), .B1(
        n19906), .B2(n19686), .ZN(n19680) );
  OAI211_X1 U21877 ( .C1(n19972), .C2(n19689), .A(n19681), .B(n19680), .ZN(
        P3_U2890) );
  AOI22_X1 U21878 ( .A1(n19906), .A2(n19685), .B1(n19984), .B2(n19684), .ZN(
        n19683) );
  AOI22_X1 U21879 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19987), .B1(
        n19995), .B2(n19686), .ZN(n19682) );
  OAI211_X1 U21880 ( .C1(n19881), .C2(n19689), .A(n19683), .B(n19682), .ZN(
        P3_U2882) );
  AOI22_X1 U21881 ( .A1(n19995), .A2(n19685), .B1(n19993), .B2(n19684), .ZN(
        n19688) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19998), .B1(
        n19916), .B2(n19686), .ZN(n19687) );
  OAI211_X1 U21883 ( .C1(n19978), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P3_U2874) );
  OAI22_X1 U21884 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19897), .ZN(n19690) );
  INV_X1 U21885 ( .A(n19690), .ZN(U256) );
  NAND2_X1 U21886 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19901), .ZN(n19720) );
  NAND2_X1 U21887 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19901), .ZN(n19730) );
  INV_X1 U21888 ( .A(n19730), .ZN(n19717) );
  INV_X1 U21889 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21470) );
  NOR2_X2 U21890 ( .A1(n21470), .A2(n19902), .ZN(n19725) );
  AOI22_X1 U21891 ( .A1(n19921), .A2(n19717), .B1(n19903), .B2(n19725), .ZN(
        n19694) );
  INV_X1 U21892 ( .A(n19691), .ZN(n19904) );
  NOR2_X2 U21893 ( .A1(n19692), .A2(n19904), .ZN(n19727) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19907), .B1(
        n19906), .B2(n19727), .ZN(n19693) );
  OAI211_X1 U21895 ( .C1(n20002), .C2(n19720), .A(n19694), .B(n19693), .ZN(
        P3_U2993) );
  INV_X1 U21896 ( .A(n19720), .ZN(n19726) );
  AOI22_X1 U21897 ( .A1(n19921), .A2(n19726), .B1(n19910), .B2(n19725), .ZN(
        n19696) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19911), .B1(
        n19995), .B2(n19727), .ZN(n19695) );
  OAI211_X1 U21899 ( .C1(n19914), .C2(n19730), .A(n19696), .B(n19695), .ZN(
        P3_U2985) );
  AOI22_X1 U21900 ( .A1(n19933), .A2(n19717), .B1(n19915), .B2(n19725), .ZN(
        n19698) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19727), .ZN(n19697) );
  OAI211_X1 U21902 ( .C1(n19914), .C2(n19720), .A(n19698), .B(n19697), .ZN(
        P3_U2977) );
  AOI22_X1 U21903 ( .A1(n19933), .A2(n19726), .B1(n19920), .B2(n19725), .ZN(
        n19700) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19727), .ZN(n19699) );
  OAI211_X1 U21905 ( .C1(n19931), .C2(n19730), .A(n19700), .B(n19699), .ZN(
        P3_U2969) );
  AOI22_X1 U21906 ( .A1(n19939), .A2(n19726), .B1(n19926), .B2(n19725), .ZN(
        n19702) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19928), .B1(
        n19927), .B2(n19727), .ZN(n19701) );
  OAI211_X1 U21908 ( .C1(n19937), .C2(n19730), .A(n19702), .B(n19701), .ZN(
        P3_U2961) );
  AOI22_X1 U21909 ( .A1(n19945), .A2(n19726), .B1(n19932), .B2(n19725), .ZN(
        n19704) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19934), .B1(
        n19933), .B2(n19727), .ZN(n19703) );
  OAI211_X1 U21911 ( .C1(n19943), .C2(n19730), .A(n19704), .B(n19703), .ZN(
        P3_U2953) );
  AOI22_X1 U21912 ( .A1(n19957), .A2(n19717), .B1(n19938), .B2(n19725), .ZN(
        n19706) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19727), .ZN(n19705) );
  OAI211_X1 U21914 ( .C1(n19943), .C2(n19720), .A(n19706), .B(n19705), .ZN(
        P3_U2945) );
  AOI22_X1 U21915 ( .A1(n19957), .A2(n19726), .B1(n19944), .B2(n19725), .ZN(
        n19708) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n19727), .ZN(n19707) );
  OAI211_X1 U21917 ( .C1(n19874), .C2(n19730), .A(n19708), .B(n19707), .ZN(
        P3_U2937) );
  AOI22_X1 U21918 ( .A1(n19963), .A2(n19726), .B1(n19950), .B2(n19725), .ZN(
        n19710) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n19727), .ZN(n19709) );
  OAI211_X1 U21920 ( .C1(n19955), .C2(n19730), .A(n19710), .B(n19709), .ZN(
        P3_U2929) );
  AOI22_X1 U21921 ( .A1(n19968), .A2(n19726), .B1(n19956), .B2(n19725), .ZN(
        n19712) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19958), .B1(
        n19957), .B2(n19727), .ZN(n19711) );
  OAI211_X1 U21923 ( .C1(n19961), .C2(n19730), .A(n19712), .B(n19711), .ZN(
        P3_U2921) );
  AOI22_X1 U21924 ( .A1(n19974), .A2(n19726), .B1(n19962), .B2(n19725), .ZN(
        n19714) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19964), .B1(
        n19963), .B2(n19727), .ZN(n19713) );
  OAI211_X1 U21926 ( .C1(n19972), .C2(n19730), .A(n19714), .B(n19713), .ZN(
        P3_U2913) );
  AOI22_X1 U21927 ( .A1(n19980), .A2(n19726), .B1(n19967), .B2(n19725), .ZN(
        n19716) );
  AOI22_X1 U21928 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19969), .B1(
        n19968), .B2(n19727), .ZN(n19715) );
  OAI211_X1 U21929 ( .C1(n19881), .C2(n19730), .A(n19716), .B(n19715), .ZN(
        P3_U2905) );
  AOI22_X1 U21930 ( .A1(n19997), .A2(n19717), .B1(n19973), .B2(n19725), .ZN(
        n19719) );
  AOI22_X1 U21931 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n19727), .ZN(n19718) );
  OAI211_X1 U21932 ( .C1(n19881), .C2(n19720), .A(n19719), .B(n19718), .ZN(
        P3_U2897) );
  AOI22_X1 U21933 ( .A1(n19997), .A2(n19726), .B1(n19979), .B2(n19725), .ZN(
        n19722) );
  AOI22_X1 U21934 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19981), .B1(
        n19980), .B2(n19727), .ZN(n19721) );
  OAI211_X1 U21935 ( .C1(n19991), .C2(n19730), .A(n19722), .B(n19721), .ZN(
        P3_U2889) );
  AOI22_X1 U21936 ( .A1(n19906), .A2(n19726), .B1(n19984), .B2(n19725), .ZN(
        n19724) );
  AOI22_X1 U21937 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19987), .B1(
        n19986), .B2(n19727), .ZN(n19723) );
  OAI211_X1 U21938 ( .C1(n19896), .C2(n19730), .A(n19724), .B(n19723), .ZN(
        P3_U2881) );
  AOI22_X1 U21939 ( .A1(n19995), .A2(n19726), .B1(n19993), .B2(n19725), .ZN(
        n19729) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19998), .B1(
        n19997), .B2(n19727), .ZN(n19728) );
  OAI211_X1 U21941 ( .C1(n20002), .C2(n19730), .A(n19729), .B(n19728), .ZN(
        P3_U2873) );
  OAI22_X1 U21942 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19897), .ZN(n19731) );
  INV_X1 U21943 ( .A(n19731), .ZN(U255) );
  INV_X1 U21944 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19732) );
  NOR2_X1 U21945 ( .A1(n19732), .A2(n19653), .ZN(n19762) );
  INV_X1 U21946 ( .A(n19762), .ZN(n19771) );
  NAND2_X1 U21947 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19901), .ZN(n19765) );
  INV_X1 U21948 ( .A(n19765), .ZN(n19767) );
  AND2_X1 U21949 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n19854), .ZN(n19766) );
  AOI22_X1 U21950 ( .A1(n19921), .A2(n19767), .B1(n19903), .B2(n19766), .ZN(
        n19735) );
  NOR2_X2 U21951 ( .A1(n19733), .A2(n19904), .ZN(n19768) );
  AOI22_X1 U21952 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19907), .B1(
        n19906), .B2(n19768), .ZN(n19734) );
  OAI211_X1 U21953 ( .C1(n20002), .C2(n19771), .A(n19735), .B(n19734), .ZN(
        P3_U2992) );
  AOI22_X1 U21954 ( .A1(n19921), .A2(n19762), .B1(n19910), .B2(n19766), .ZN(
        n19737) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19911), .B1(
        n19995), .B2(n19768), .ZN(n19736) );
  OAI211_X1 U21956 ( .C1(n19914), .C2(n19765), .A(n19737), .B(n19736), .ZN(
        P3_U2984) );
  AOI22_X1 U21957 ( .A1(n19927), .A2(n19762), .B1(n19915), .B2(n19766), .ZN(
        n19739) );
  AOI22_X1 U21958 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19768), .ZN(n19738) );
  OAI211_X1 U21959 ( .C1(n19925), .C2(n19765), .A(n19739), .B(n19738), .ZN(
        P3_U2976) );
  AOI22_X1 U21960 ( .A1(n19939), .A2(n19767), .B1(n19920), .B2(n19766), .ZN(
        n19741) );
  AOI22_X1 U21961 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19768), .ZN(n19740) );
  OAI211_X1 U21962 ( .C1(n19925), .C2(n19771), .A(n19741), .B(n19740), .ZN(
        P3_U2968) );
  AOI22_X1 U21963 ( .A1(n19945), .A2(n19767), .B1(n19926), .B2(n19766), .ZN(
        n19743) );
  AOI22_X1 U21964 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19928), .B1(
        n19927), .B2(n19768), .ZN(n19742) );
  OAI211_X1 U21965 ( .C1(n19931), .C2(n19771), .A(n19743), .B(n19742), .ZN(
        P3_U2960) );
  AOI22_X1 U21966 ( .A1(n19951), .A2(n19767), .B1(n19932), .B2(n19766), .ZN(
        n19745) );
  AOI22_X1 U21967 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19934), .B1(
        n19933), .B2(n19768), .ZN(n19744) );
  OAI211_X1 U21968 ( .C1(n19937), .C2(n19771), .A(n19745), .B(n19744), .ZN(
        P3_U2952) );
  AOI22_X1 U21969 ( .A1(n19957), .A2(n19767), .B1(n19938), .B2(n19766), .ZN(
        n19747) );
  AOI22_X1 U21970 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19768), .ZN(n19746) );
  OAI211_X1 U21971 ( .C1(n19943), .C2(n19771), .A(n19747), .B(n19746), .ZN(
        P3_U2944) );
  AOI22_X1 U21972 ( .A1(n19957), .A2(n19762), .B1(n19944), .B2(n19766), .ZN(
        n19749) );
  AOI22_X1 U21973 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n19768), .ZN(n19748) );
  OAI211_X1 U21974 ( .C1(n19874), .C2(n19765), .A(n19749), .B(n19748), .ZN(
        P3_U2936) );
  AOI22_X1 U21975 ( .A1(n19950), .A2(n19766), .B1(n19968), .B2(n19767), .ZN(
        n19751) );
  AOI22_X1 U21976 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n19768), .ZN(n19750) );
  OAI211_X1 U21977 ( .C1(n19874), .C2(n19771), .A(n19751), .B(n19750), .ZN(
        P3_U2928) );
  AOI22_X1 U21978 ( .A1(n19974), .A2(n19767), .B1(n19956), .B2(n19766), .ZN(
        n19753) );
  AOI22_X1 U21979 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19958), .B1(
        n19957), .B2(n19768), .ZN(n19752) );
  OAI211_X1 U21980 ( .C1(n19955), .C2(n19771), .A(n19753), .B(n19752), .ZN(
        P3_U2920) );
  AOI22_X1 U21981 ( .A1(n19980), .A2(n19767), .B1(n19962), .B2(n19766), .ZN(
        n19755) );
  AOI22_X1 U21982 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19964), .B1(
        n19963), .B2(n19768), .ZN(n19754) );
  OAI211_X1 U21983 ( .C1(n19961), .C2(n19771), .A(n19755), .B(n19754), .ZN(
        P3_U2912) );
  AOI22_X1 U21984 ( .A1(n19980), .A2(n19762), .B1(n19967), .B2(n19766), .ZN(
        n19757) );
  AOI22_X1 U21985 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19969), .B1(
        n19968), .B2(n19768), .ZN(n19756) );
  OAI211_X1 U21986 ( .C1(n19881), .C2(n19765), .A(n19757), .B(n19756), .ZN(
        P3_U2904) );
  AOI22_X1 U21987 ( .A1(n19986), .A2(n19762), .B1(n19973), .B2(n19766), .ZN(
        n19759) );
  AOI22_X1 U21988 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n19768), .ZN(n19758) );
  OAI211_X1 U21989 ( .C1(n19978), .C2(n19765), .A(n19759), .B(n19758), .ZN(
        P3_U2896) );
  AOI22_X1 U21990 ( .A1(n19997), .A2(n19762), .B1(n19979), .B2(n19766), .ZN(
        n19761) );
  AOI22_X1 U21991 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19981), .B1(
        n19980), .B2(n19768), .ZN(n19760) );
  OAI211_X1 U21992 ( .C1(n19991), .C2(n19765), .A(n19761), .B(n19760), .ZN(
        P3_U2888) );
  AOI22_X1 U21993 ( .A1(n19906), .A2(n19762), .B1(n19984), .B2(n19766), .ZN(
        n19764) );
  AOI22_X1 U21994 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19987), .B1(
        n19986), .B2(n19768), .ZN(n19763) );
  OAI211_X1 U21995 ( .C1(n19896), .C2(n19765), .A(n19764), .B(n19763), .ZN(
        P3_U2880) );
  AOI22_X1 U21996 ( .A1(n19916), .A2(n19767), .B1(n19993), .B2(n19766), .ZN(
        n19770) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19998), .B1(
        n19997), .B2(n19768), .ZN(n19769) );
  OAI211_X1 U21998 ( .C1(n19896), .C2(n19771), .A(n19770), .B(n19769), .ZN(
        P3_U2872) );
  OAI22_X1 U21999 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19897), .ZN(n19772) );
  INV_X1 U22000 ( .A(n19772), .ZN(U254) );
  NAND2_X1 U22001 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19901), .ZN(n19805) );
  NAND2_X1 U22002 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19901), .ZN(n19811) );
  INV_X1 U22003 ( .A(n19811), .ZN(n19802) );
  INV_X1 U22004 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21480) );
  NOR2_X2 U22005 ( .A1(n21480), .A2(n19902), .ZN(n19806) );
  AOI22_X1 U22006 ( .A1(n19916), .A2(n19802), .B1(n19903), .B2(n19806), .ZN(
        n19775) );
  NOR2_X2 U22007 ( .A1(n19773), .A2(n19904), .ZN(n19808) );
  AOI22_X1 U22008 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19907), .B1(
        n19906), .B2(n19808), .ZN(n19774) );
  OAI211_X1 U22009 ( .C1(n19818), .C2(n19805), .A(n19775), .B(n19774), .ZN(
        P3_U2991) );
  INV_X1 U22010 ( .A(n19805), .ZN(n19807) );
  AOI22_X1 U22011 ( .A1(n19927), .A2(n19807), .B1(n19910), .B2(n19806), .ZN(
        n19777) );
  AOI22_X1 U22012 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19911), .B1(
        n19995), .B2(n19808), .ZN(n19776) );
  OAI211_X1 U22013 ( .C1(n19818), .C2(n19811), .A(n19777), .B(n19776), .ZN(
        P3_U2983) );
  AOI22_X1 U22014 ( .A1(n19933), .A2(n19807), .B1(n19915), .B2(n19806), .ZN(
        n19779) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19808), .ZN(n19778) );
  OAI211_X1 U22016 ( .C1(n19914), .C2(n19811), .A(n19779), .B(n19778), .ZN(
        P3_U2975) );
  AOI22_X1 U22017 ( .A1(n19933), .A2(n19802), .B1(n19920), .B2(n19806), .ZN(
        n19781) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19808), .ZN(n19780) );
  OAI211_X1 U22019 ( .C1(n19931), .C2(n19805), .A(n19781), .B(n19780), .ZN(
        P3_U2967) );
  AOI22_X1 U22020 ( .A1(n19945), .A2(n19807), .B1(n19926), .B2(n19806), .ZN(
        n19783) );
  AOI22_X1 U22021 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19928), .B1(
        n19927), .B2(n19808), .ZN(n19782) );
  OAI211_X1 U22022 ( .C1(n19931), .C2(n19811), .A(n19783), .B(n19782), .ZN(
        P3_U2959) );
  AOI22_X1 U22023 ( .A1(n19951), .A2(n19807), .B1(n19932), .B2(n19806), .ZN(
        n19785) );
  AOI22_X1 U22024 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19934), .B1(
        n19933), .B2(n19808), .ZN(n19784) );
  OAI211_X1 U22025 ( .C1(n19937), .C2(n19811), .A(n19785), .B(n19784), .ZN(
        P3_U2951) );
  AOI22_X1 U22026 ( .A1(n19957), .A2(n19807), .B1(n19938), .B2(n19806), .ZN(
        n19787) );
  AOI22_X1 U22027 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19808), .ZN(n19786) );
  OAI211_X1 U22028 ( .C1(n19943), .C2(n19811), .A(n19787), .B(n19786), .ZN(
        P3_U2943) );
  AOI22_X1 U22029 ( .A1(n19963), .A2(n19807), .B1(n19944), .B2(n19806), .ZN(
        n19789) );
  AOI22_X1 U22030 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n19808), .ZN(n19788) );
  OAI211_X1 U22031 ( .C1(n19949), .C2(n19811), .A(n19789), .B(n19788), .ZN(
        P3_U2935) );
  AOI22_X1 U22032 ( .A1(n19950), .A2(n19806), .B1(n19968), .B2(n19807), .ZN(
        n19791) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n19808), .ZN(n19790) );
  OAI211_X1 U22034 ( .C1(n19874), .C2(n19811), .A(n19791), .B(n19790), .ZN(
        P3_U2927) );
  AOI22_X1 U22035 ( .A1(n19974), .A2(n19807), .B1(n19956), .B2(n19806), .ZN(
        n19793) );
  AOI22_X1 U22036 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19958), .B1(
        n19957), .B2(n19808), .ZN(n19792) );
  OAI211_X1 U22037 ( .C1(n19955), .C2(n19811), .A(n19793), .B(n19792), .ZN(
        P3_U2919) );
  AOI22_X1 U22038 ( .A1(n19974), .A2(n19802), .B1(n19962), .B2(n19806), .ZN(
        n19795) );
  AOI22_X1 U22039 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19964), .B1(
        n19963), .B2(n19808), .ZN(n19794) );
  OAI211_X1 U22040 ( .C1(n19972), .C2(n19805), .A(n19795), .B(n19794), .ZN(
        P3_U2911) );
  AOI22_X1 U22041 ( .A1(n19980), .A2(n19802), .B1(n19967), .B2(n19806), .ZN(
        n19797) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19969), .B1(
        n19968), .B2(n19808), .ZN(n19796) );
  OAI211_X1 U22043 ( .C1(n19881), .C2(n19805), .A(n19797), .B(n19796), .ZN(
        P3_U2903) );
  AOI22_X1 U22044 ( .A1(n19997), .A2(n19807), .B1(n19973), .B2(n19806), .ZN(
        n19799) );
  AOI22_X1 U22045 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n19808), .ZN(n19798) );
  OAI211_X1 U22046 ( .C1(n19881), .C2(n19811), .A(n19799), .B(n19798), .ZN(
        P3_U2895) );
  AOI22_X1 U22047 ( .A1(n19997), .A2(n19802), .B1(n19979), .B2(n19806), .ZN(
        n19801) );
  AOI22_X1 U22048 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19981), .B1(
        n19980), .B2(n19808), .ZN(n19800) );
  OAI211_X1 U22049 ( .C1(n19991), .C2(n19805), .A(n19801), .B(n19800), .ZN(
        P3_U2887) );
  AOI22_X1 U22050 ( .A1(n19906), .A2(n19802), .B1(n19984), .B2(n19806), .ZN(
        n19804) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19987), .B1(
        n19986), .B2(n19808), .ZN(n19803) );
  OAI211_X1 U22052 ( .C1(n19896), .C2(n19805), .A(n19804), .B(n19803), .ZN(
        P3_U2879) );
  AOI22_X1 U22053 ( .A1(n19916), .A2(n19807), .B1(n19993), .B2(n19806), .ZN(
        n19810) );
  AOI22_X1 U22054 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19998), .B1(
        n19997), .B2(n19808), .ZN(n19809) );
  OAI211_X1 U22055 ( .C1(n19896), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P3_U2871) );
  OAI22_X1 U22056 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19897), .ZN(n19812) );
  INV_X1 U22057 ( .A(n19812), .ZN(U253) );
  NAND2_X1 U22058 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n19901), .ZN(n19852) );
  NAND2_X1 U22059 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19901), .ZN(n19844) );
  INV_X1 U22060 ( .A(n19844), .ZN(n19848) );
  INV_X1 U22061 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21485) );
  NOR2_X2 U22062 ( .A1(n21485), .A2(n19902), .ZN(n19847) );
  AOI22_X1 U22063 ( .A1(n19921), .A2(n19848), .B1(n19903), .B2(n19847), .ZN(
        n19815) );
  NOR2_X2 U22064 ( .A1(n19813), .A2(n19904), .ZN(n19849) );
  AOI22_X1 U22065 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19907), .B1(
        n19906), .B2(n19849), .ZN(n19814) );
  OAI211_X1 U22066 ( .C1(n20002), .C2(n19852), .A(n19815), .B(n19814), .ZN(
        P3_U2990) );
  AOI22_X1 U22067 ( .A1(n19927), .A2(n19848), .B1(n19910), .B2(n19847), .ZN(
        n19817) );
  AOI22_X1 U22068 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19911), .B1(
        n19995), .B2(n19849), .ZN(n19816) );
  OAI211_X1 U22069 ( .C1(n19818), .C2(n19852), .A(n19817), .B(n19816), .ZN(
        P3_U2982) );
  INV_X1 U22070 ( .A(n19852), .ZN(n19841) );
  AOI22_X1 U22071 ( .A1(n19927), .A2(n19841), .B1(n19915), .B2(n19847), .ZN(
        n19820) );
  AOI22_X1 U22072 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19849), .ZN(n19819) );
  OAI211_X1 U22073 ( .C1(n19925), .C2(n19844), .A(n19820), .B(n19819), .ZN(
        P3_U2974) );
  AOI22_X1 U22074 ( .A1(n19939), .A2(n19848), .B1(n19920), .B2(n19847), .ZN(
        n19822) );
  AOI22_X1 U22075 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19849), .ZN(n19821) );
  OAI211_X1 U22076 ( .C1(n19925), .C2(n19852), .A(n19822), .B(n19821), .ZN(
        P3_U2966) );
  AOI22_X1 U22077 ( .A1(n19945), .A2(n19848), .B1(n19926), .B2(n19847), .ZN(
        n19824) );
  AOI22_X1 U22078 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19928), .B1(
        n19927), .B2(n19849), .ZN(n19823) );
  OAI211_X1 U22079 ( .C1(n19931), .C2(n19852), .A(n19824), .B(n19823), .ZN(
        P3_U2958) );
  AOI22_X1 U22080 ( .A1(n19945), .A2(n19841), .B1(n19932), .B2(n19847), .ZN(
        n19826) );
  AOI22_X1 U22081 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19934), .B1(
        n19933), .B2(n19849), .ZN(n19825) );
  OAI211_X1 U22082 ( .C1(n19943), .C2(n19844), .A(n19826), .B(n19825), .ZN(
        P3_U2950) );
  AOI22_X1 U22083 ( .A1(n19957), .A2(n19848), .B1(n19938), .B2(n19847), .ZN(
        n19828) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19849), .ZN(n19827) );
  OAI211_X1 U22085 ( .C1(n19943), .C2(n19852), .A(n19828), .B(n19827), .ZN(
        P3_U2942) );
  AOI22_X1 U22086 ( .A1(n19957), .A2(n19841), .B1(n19944), .B2(n19847), .ZN(
        n19830) );
  AOI22_X1 U22087 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n19849), .ZN(n19829) );
  OAI211_X1 U22088 ( .C1(n19874), .C2(n19844), .A(n19830), .B(n19829), .ZN(
        P3_U2934) );
  AOI22_X1 U22089 ( .A1(n19963), .A2(n19841), .B1(n19950), .B2(n19847), .ZN(
        n19832) );
  AOI22_X1 U22090 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n19849), .ZN(n19831) );
  OAI211_X1 U22091 ( .C1(n19955), .C2(n19844), .A(n19832), .B(n19831), .ZN(
        P3_U2926) );
  AOI22_X1 U22092 ( .A1(n19968), .A2(n19841), .B1(n19956), .B2(n19847), .ZN(
        n19834) );
  AOI22_X1 U22093 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19958), .B1(
        n19957), .B2(n19849), .ZN(n19833) );
  OAI211_X1 U22094 ( .C1(n19961), .C2(n19844), .A(n19834), .B(n19833), .ZN(
        P3_U2918) );
  AOI22_X1 U22095 ( .A1(n19980), .A2(n19848), .B1(n19962), .B2(n19847), .ZN(
        n19836) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19964), .B1(
        n19963), .B2(n19849), .ZN(n19835) );
  OAI211_X1 U22097 ( .C1(n19961), .C2(n19852), .A(n19836), .B(n19835), .ZN(
        P3_U2910) );
  AOI22_X1 U22098 ( .A1(n19980), .A2(n19841), .B1(n19967), .B2(n19847), .ZN(
        n19838) );
  AOI22_X1 U22099 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19969), .B1(
        n19968), .B2(n19849), .ZN(n19837) );
  OAI211_X1 U22100 ( .C1(n19881), .C2(n19844), .A(n19838), .B(n19837), .ZN(
        P3_U2902) );
  AOI22_X1 U22101 ( .A1(n19997), .A2(n19848), .B1(n19973), .B2(n19847), .ZN(
        n19840) );
  AOI22_X1 U22102 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n19849), .ZN(n19839) );
  OAI211_X1 U22103 ( .C1(n19881), .C2(n19852), .A(n19840), .B(n19839), .ZN(
        P3_U2894) );
  AOI22_X1 U22104 ( .A1(n19997), .A2(n19841), .B1(n19979), .B2(n19847), .ZN(
        n19843) );
  AOI22_X1 U22105 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19981), .B1(
        n19980), .B2(n19849), .ZN(n19842) );
  OAI211_X1 U22106 ( .C1(n19991), .C2(n19844), .A(n19843), .B(n19842), .ZN(
        P3_U2886) );
  AOI22_X1 U22107 ( .A1(n19995), .A2(n19848), .B1(n19984), .B2(n19847), .ZN(
        n19846) );
  AOI22_X1 U22108 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19987), .B1(
        n19986), .B2(n19849), .ZN(n19845) );
  OAI211_X1 U22109 ( .C1(n19991), .C2(n19852), .A(n19846), .B(n19845), .ZN(
        P3_U2878) );
  AOI22_X1 U22110 ( .A1(n19916), .A2(n19848), .B1(n19993), .B2(n19847), .ZN(
        n19851) );
  AOI22_X1 U22111 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19998), .B1(
        n19997), .B2(n19849), .ZN(n19850) );
  OAI211_X1 U22112 ( .C1(n19896), .C2(n19852), .A(n19851), .B(n19850), .ZN(
        P3_U2870) );
  OAI22_X1 U22113 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19897), .ZN(n19853) );
  INV_X1 U22114 ( .A(n19853), .ZN(U252) );
  NAND2_X1 U22115 ( .A1(n19901), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U22116 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19901), .ZN(n19885) );
  INV_X1 U22117 ( .A(n19885), .ZN(n19891) );
  AND2_X1 U22118 ( .A1(n19854), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U22119 ( .A1(n19921), .A2(n19891), .B1(n19903), .B2(n19890), .ZN(
        n19857) );
  NOR2_X2 U22120 ( .A1(n19855), .A2(n19904), .ZN(n19892) );
  AOI22_X1 U22121 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19907), .B1(
        n19906), .B2(n19892), .ZN(n19856) );
  OAI211_X1 U22122 ( .C1(n20002), .C2(n19895), .A(n19857), .B(n19856), .ZN(
        P3_U2989) );
  INV_X1 U22123 ( .A(n19895), .ZN(n19882) );
  AOI22_X1 U22124 ( .A1(n19921), .A2(n19882), .B1(n19910), .B2(n19890), .ZN(
        n19859) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19911), .B1(
        n19995), .B2(n19892), .ZN(n19858) );
  OAI211_X1 U22126 ( .C1(n19914), .C2(n19885), .A(n19859), .B(n19858), .ZN(
        P3_U2981) );
  AOI22_X1 U22127 ( .A1(n19933), .A2(n19891), .B1(n19915), .B2(n19890), .ZN(
        n19861) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19892), .ZN(n19860) );
  OAI211_X1 U22129 ( .C1(n19914), .C2(n19895), .A(n19861), .B(n19860), .ZN(
        P3_U2973) );
  AOI22_X1 U22130 ( .A1(n19933), .A2(n19882), .B1(n19920), .B2(n19890), .ZN(
        n19863) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19892), .ZN(n19862) );
  OAI211_X1 U22132 ( .C1(n19931), .C2(n19885), .A(n19863), .B(n19862), .ZN(
        P3_U2965) );
  AOI22_X1 U22133 ( .A1(n19939), .A2(n19882), .B1(n19926), .B2(n19890), .ZN(
        n19865) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19928), .B1(
        n19927), .B2(n19892), .ZN(n19864) );
  OAI211_X1 U22135 ( .C1(n19937), .C2(n19885), .A(n19865), .B(n19864), .ZN(
        P3_U2957) );
  AOI22_X1 U22136 ( .A1(n19945), .A2(n19882), .B1(n19932), .B2(n19890), .ZN(
        n19867) );
  AOI22_X1 U22137 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19934), .B1(
        n19933), .B2(n19892), .ZN(n19866) );
  OAI211_X1 U22138 ( .C1(n19943), .C2(n19885), .A(n19867), .B(n19866), .ZN(
        P3_U2949) );
  AOI22_X1 U22139 ( .A1(n19951), .A2(n19882), .B1(n19938), .B2(n19890), .ZN(
        n19869) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19892), .ZN(n19868) );
  OAI211_X1 U22141 ( .C1(n19949), .C2(n19885), .A(n19869), .B(n19868), .ZN(
        P3_U2941) );
  AOI22_X1 U22142 ( .A1(n19963), .A2(n19891), .B1(n19944), .B2(n19890), .ZN(
        n19871) );
  AOI22_X1 U22143 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n19892), .ZN(n19870) );
  OAI211_X1 U22144 ( .C1(n19949), .C2(n19895), .A(n19871), .B(n19870), .ZN(
        P3_U2933) );
  AOI22_X1 U22145 ( .A1(n19950), .A2(n19890), .B1(n19968), .B2(n19891), .ZN(
        n19873) );
  AOI22_X1 U22146 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n19892), .ZN(n19872) );
  OAI211_X1 U22147 ( .C1(n19874), .C2(n19895), .A(n19873), .B(n19872), .ZN(
        P3_U2925) );
  AOI22_X1 U22148 ( .A1(n19968), .A2(n19882), .B1(n19956), .B2(n19890), .ZN(
        n19876) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19958), .B1(
        n19957), .B2(n19892), .ZN(n19875) );
  OAI211_X1 U22150 ( .C1(n19961), .C2(n19885), .A(n19876), .B(n19875), .ZN(
        P3_U2917) );
  AOI22_X1 U22151 ( .A1(n19980), .A2(n19891), .B1(n19962), .B2(n19890), .ZN(
        n19878) );
  AOI22_X1 U22152 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19964), .B1(
        n19963), .B2(n19892), .ZN(n19877) );
  OAI211_X1 U22153 ( .C1(n19961), .C2(n19895), .A(n19878), .B(n19877), .ZN(
        P3_U2909) );
  AOI22_X1 U22154 ( .A1(n19980), .A2(n19882), .B1(n19967), .B2(n19890), .ZN(
        n19880) );
  AOI22_X1 U22155 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19969), .B1(
        n19968), .B2(n19892), .ZN(n19879) );
  OAI211_X1 U22156 ( .C1(n19881), .C2(n19885), .A(n19880), .B(n19879), .ZN(
        P3_U2901) );
  AOI22_X1 U22157 ( .A1(n19986), .A2(n19882), .B1(n19973), .B2(n19890), .ZN(
        n19884) );
  AOI22_X1 U22158 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n19892), .ZN(n19883) );
  OAI211_X1 U22159 ( .C1(n19978), .C2(n19885), .A(n19884), .B(n19883), .ZN(
        P3_U2893) );
  AOI22_X1 U22160 ( .A1(n19906), .A2(n19891), .B1(n19979), .B2(n19890), .ZN(
        n19887) );
  AOI22_X1 U22161 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19981), .B1(
        n19980), .B2(n19892), .ZN(n19886) );
  OAI211_X1 U22162 ( .C1(n19978), .C2(n19895), .A(n19887), .B(n19886), .ZN(
        P3_U2885) );
  AOI22_X1 U22163 ( .A1(n19995), .A2(n19891), .B1(n19984), .B2(n19890), .ZN(
        n19889) );
  AOI22_X1 U22164 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19987), .B1(
        n19986), .B2(n19892), .ZN(n19888) );
  OAI211_X1 U22165 ( .C1(n19991), .C2(n19895), .A(n19889), .B(n19888), .ZN(
        P3_U2877) );
  AOI22_X1 U22166 ( .A1(n19916), .A2(n19891), .B1(n19993), .B2(n19890), .ZN(
        n19894) );
  AOI22_X1 U22167 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19998), .B1(
        n19997), .B2(n19892), .ZN(n19893) );
  OAI211_X1 U22168 ( .C1(n19896), .C2(n19895), .A(n19894), .B(n19893), .ZN(
        P3_U2869) );
  OAI22_X1 U22169 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19897), .ZN(n19899) );
  INV_X1 U22170 ( .A(n19899), .ZN(U251) );
  INV_X1 U22171 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19900) );
  NOR2_X1 U22172 ( .A1(n19653), .A2(n19900), .ZN(n19994) );
  INV_X1 U22173 ( .A(n19994), .ZN(n19990) );
  NAND2_X1 U22174 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19901), .ZN(n20001) );
  INV_X1 U22175 ( .A(n20001), .ZN(n19985) );
  INV_X1 U22176 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n21600) );
  NOR2_X2 U22177 ( .A1(n19902), .A2(n21600), .ZN(n19992) );
  AOI22_X1 U22178 ( .A1(n19921), .A2(n19985), .B1(n19903), .B2(n19992), .ZN(
        n19909) );
  NOR2_X2 U22179 ( .A1(n19905), .A2(n19904), .ZN(n19996) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19907), .B1(
        n19906), .B2(n19996), .ZN(n19908) );
  OAI211_X1 U22181 ( .C1(n20002), .C2(n19990), .A(n19909), .B(n19908), .ZN(
        P3_U2988) );
  AOI22_X1 U22182 ( .A1(n19921), .A2(n19994), .B1(n19910), .B2(n19992), .ZN(
        n19913) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19911), .B1(
        n19995), .B2(n19996), .ZN(n19912) );
  OAI211_X1 U22184 ( .C1(n19914), .C2(n20001), .A(n19913), .B(n19912), .ZN(
        P3_U2980) );
  AOI22_X1 U22185 ( .A1(n19927), .A2(n19994), .B1(n19915), .B2(n19992), .ZN(
        n19919) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19917), .B1(
        n19916), .B2(n19996), .ZN(n19918) );
  OAI211_X1 U22187 ( .C1(n19925), .C2(n20001), .A(n19919), .B(n19918), .ZN(
        P3_U2972) );
  AOI22_X1 U22188 ( .A1(n19939), .A2(n19985), .B1(n19920), .B2(n19992), .ZN(
        n19924) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n19996), .ZN(n19923) );
  OAI211_X1 U22190 ( .C1(n19925), .C2(n19990), .A(n19924), .B(n19923), .ZN(
        P3_U2964) );
  AOI22_X1 U22191 ( .A1(n19945), .A2(n19985), .B1(n19926), .B2(n19992), .ZN(
        n19930) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19928), .B1(
        n19927), .B2(n19996), .ZN(n19929) );
  OAI211_X1 U22193 ( .C1(n19931), .C2(n19990), .A(n19930), .B(n19929), .ZN(
        P3_U2956) );
  AOI22_X1 U22194 ( .A1(n19951), .A2(n19985), .B1(n19932), .B2(n19992), .ZN(
        n19936) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19934), .B1(
        n19933), .B2(n19996), .ZN(n19935) );
  OAI211_X1 U22196 ( .C1(n19937), .C2(n19990), .A(n19936), .B(n19935), .ZN(
        P3_U2948) );
  AOI22_X1 U22197 ( .A1(n19957), .A2(n19985), .B1(n19938), .B2(n19992), .ZN(
        n19942) );
  AOI22_X1 U22198 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19940), .B1(
        n19939), .B2(n19996), .ZN(n19941) );
  OAI211_X1 U22199 ( .C1(n19943), .C2(n19990), .A(n19942), .B(n19941), .ZN(
        P3_U2940) );
  AOI22_X1 U22200 ( .A1(n19963), .A2(n19985), .B1(n19944), .B2(n19992), .ZN(
        n19948) );
  AOI22_X1 U22201 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19946), .B1(
        n19945), .B2(n19996), .ZN(n19947) );
  OAI211_X1 U22202 ( .C1(n19949), .C2(n19990), .A(n19948), .B(n19947), .ZN(
        P3_U2932) );
  AOI22_X1 U22203 ( .A1(n19963), .A2(n19994), .B1(n19950), .B2(n19992), .ZN(
        n19954) );
  AOI22_X1 U22204 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19952), .B1(
        n19951), .B2(n19996), .ZN(n19953) );
  OAI211_X1 U22205 ( .C1(n19955), .C2(n20001), .A(n19954), .B(n19953), .ZN(
        P3_U2924) );
  AOI22_X1 U22206 ( .A1(n19968), .A2(n19994), .B1(n19956), .B2(n19992), .ZN(
        n19960) );
  AOI22_X1 U22207 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19958), .B1(
        n19957), .B2(n19996), .ZN(n19959) );
  OAI211_X1 U22208 ( .C1(n19961), .C2(n20001), .A(n19960), .B(n19959), .ZN(
        P3_U2916) );
  AOI22_X1 U22209 ( .A1(n19974), .A2(n19994), .B1(n19962), .B2(n19992), .ZN(
        n19966) );
  AOI22_X1 U22210 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19964), .B1(
        n19963), .B2(n19996), .ZN(n19965) );
  OAI211_X1 U22211 ( .C1(n19972), .C2(n20001), .A(n19966), .B(n19965), .ZN(
        P3_U2908) );
  AOI22_X1 U22212 ( .A1(n19986), .A2(n19985), .B1(n19967), .B2(n19992), .ZN(
        n19971) );
  AOI22_X1 U22213 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19969), .B1(
        n19968), .B2(n19996), .ZN(n19970) );
  OAI211_X1 U22214 ( .C1(n19972), .C2(n19990), .A(n19971), .B(n19970), .ZN(
        P3_U2900) );
  AOI22_X1 U22215 ( .A1(n19986), .A2(n19994), .B1(n19973), .B2(n19992), .ZN(
        n19977) );
  AOI22_X1 U22216 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n19996), .ZN(n19976) );
  OAI211_X1 U22217 ( .C1(n19978), .C2(n20001), .A(n19977), .B(n19976), .ZN(
        P3_U2892) );
  AOI22_X1 U22218 ( .A1(n19997), .A2(n19994), .B1(n19979), .B2(n19992), .ZN(
        n19983) );
  AOI22_X1 U22219 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19981), .B1(
        n19980), .B2(n19996), .ZN(n19982) );
  OAI211_X1 U22220 ( .C1(n19991), .C2(n20001), .A(n19983), .B(n19982), .ZN(
        P3_U2884) );
  AOI22_X1 U22221 ( .A1(n19995), .A2(n19985), .B1(n19984), .B2(n19992), .ZN(
        n19989) );
  AOI22_X1 U22222 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19987), .B1(
        n19986), .B2(n19996), .ZN(n19988) );
  OAI211_X1 U22223 ( .C1(n19991), .C2(n19990), .A(n19989), .B(n19988), .ZN(
        P3_U2876) );
  AOI22_X1 U22224 ( .A1(n19995), .A2(n19994), .B1(n19993), .B2(n19992), .ZN(
        n20000) );
  AOI22_X1 U22225 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19998), .B1(
        n19997), .B2(n19996), .ZN(n19999) );
  OAI211_X1 U22226 ( .C1(n20002), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P3_U2868) );
  AOI22_X1 U22227 ( .A1(n20004), .A2(n20459), .B1(BUF2_REG_31__SCAN_IN), .B2(
        n20003), .ZN(n20007) );
  AOI22_X1 U22228 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n20457), .B1(n20005), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n20006) );
  NAND2_X1 U22229 ( .A1(n20007), .A2(n20006), .ZN(P2_U2888) );
  INV_X1 U22230 ( .A(n20008), .ZN(n20010) );
  OAI222_X1 U22231 ( .A1(n20013), .A2(n20209), .B1(n20012), .B2(n20513), .C1(
        n20011), .C2(n20465), .ZN(P2_U2904) );
  OAI222_X1 U22232 ( .A1(n20016), .A2(n20209), .B1(n20015), .B2(n20513), .C1(
        n20465), .C2(n20014), .ZN(P2_U2905) );
  INV_X1 U22233 ( .A(n20209), .ZN(n20253) );
  AOI22_X1 U22234 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n20457), .B1(n20017), 
        .B2(n20253), .ZN(n20018) );
  OAI21_X1 U22235 ( .B1(n20019), .B2(n20465), .A(n20018), .ZN(P2_U2906) );
  OAI222_X1 U22236 ( .A1(n20022), .A2(n20209), .B1(n20021), .B2(n20513), .C1(
        n20465), .C2(n20020), .ZN(P2_U2907) );
  INV_X1 U22237 ( .A(n20465), .ZN(n20522) );
  AOI22_X1 U22238 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n20457), .B1(n20023), 
        .B2(n20522), .ZN(n20024) );
  OAI21_X1 U22239 ( .B1(n20209), .B2(n20025), .A(n20024), .ZN(P2_U2908) );
  OAI222_X1 U22240 ( .A1(n20028), .A2(n20209), .B1(n20027), .B2(n20513), .C1(
        n20465), .C2(n20026), .ZN(P2_U2909) );
  AOI22_X1 U22241 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n20457), .B1(n20029), .B2(
        n20253), .ZN(n20030) );
  OAI21_X1 U22242 ( .B1(n20031), .B2(n20465), .A(n20030), .ZN(P2_U2910) );
  OAI222_X1 U22243 ( .A1(n20034), .A2(n20209), .B1(n20033), .B2(n20513), .C1(
        n20465), .C2(n20032), .ZN(P2_U2911) );
  AOI22_X1 U22244 ( .A1(P2_EAX_REG_7__SCAN_IN), .A2(n20457), .B1(n20035), .B2(
        n20253), .ZN(n20036) );
  OAI21_X1 U22245 ( .B1(n20037), .B2(n20465), .A(n20036), .ZN(P2_U2912) );
  NOR2_X1 U22246 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20038), .ZN(
        n20537) );
  AOI22_X1 U22247 ( .A1(n20191), .A2(n20471), .B1(n20190), .B2(n20537), .ZN(
        n20049) );
  AOI21_X1 U22248 ( .B1(n20549), .B2(n20543), .A(n22411), .ZN(n20039) );
  NOR2_X1 U22249 ( .A1(n20039), .A2(n20192), .ZN(n20044) );
  INV_X1 U22250 ( .A(n20040), .ZN(n20045) );
  AOI21_X1 U22251 ( .B1(n20045), .B2(n20196), .A(n20195), .ZN(n20041) );
  AOI21_X1 U22252 ( .B1(n20044), .B2(n20042), .A(n20041), .ZN(n20043) );
  OAI21_X1 U22253 ( .B1(n20537), .B2(n20544), .A(n20044), .ZN(n20047) );
  OAI21_X1 U22254 ( .B1(n20045), .B2(n20537), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20046) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20540), .B1(
        n15512), .B2(n20539), .ZN(n20048) );
  OAI211_X1 U22256 ( .C1(n20207), .C2(n20549), .A(n20049), .B(n20048), .ZN(
        P2_U3167) );
  NAND2_X1 U22257 ( .A1(n20126), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20057) );
  INV_X1 U22258 ( .A(n20050), .ZN(n20054) );
  INV_X1 U22259 ( .A(n20060), .ZN(n20052) );
  NOR2_X1 U22260 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20051), .ZN(
        n20550) );
  OAI21_X1 U22261 ( .B1(n20052), .B2(n20550), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20053) );
  OAI21_X1 U22262 ( .B1(n20057), .B2(n20054), .A(n20053), .ZN(n20551) );
  AOI22_X1 U22263 ( .A1(n20551), .A2(n15512), .B1(n20550), .B2(n20190), .ZN(
        n20064) );
  OAI21_X1 U22264 ( .B1(n20055), .B2(n20552), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20056) );
  OAI21_X1 U22265 ( .B1(n20058), .B2(n20057), .A(n20056), .ZN(n20062) );
  AOI21_X1 U22266 ( .B1(n20550), .B2(n20199), .A(n20195), .ZN(n20059) );
  OAI21_X1 U22267 ( .B1(n20060), .B2(n20180), .A(n20059), .ZN(n20061) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20191), .ZN(n20063) );
  OAI211_X1 U22269 ( .C1(n20207), .C2(n20561), .A(n20064), .B(n20063), .ZN(
        P2_U3151) );
  INV_X1 U22270 ( .A(n20065), .ZN(n20066) );
  NAND3_X1 U22271 ( .A1(n20146), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20077) );
  INV_X1 U22272 ( .A(n20077), .ZN(n20071) );
  NAND2_X1 U22273 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20071), .ZN(
        n20067) );
  INV_X1 U22274 ( .A(n20067), .ZN(n20556) );
  NOR2_X1 U22275 ( .A1(n20066), .A2(n20556), .ZN(n20068) );
  OAI22_X1 U22276 ( .A1(n20068), .A2(n20103), .B1(n20077), .B2(n20192), .ZN(
        n20557) );
  AOI22_X1 U22277 ( .A1(n20557), .A2(n15512), .B1(n20190), .B2(n20556), .ZN(
        n20073) );
  NOR2_X1 U22278 ( .A1(n20262), .A2(n20148), .ZN(n20070) );
  OAI22_X1 U22279 ( .A1(n20068), .A2(n20180), .B1(n20525), .B2(n20067), .ZN(
        n20069) );
  OAI22_X1 U22280 ( .A1(n20071), .A2(n20070), .B1(n20195), .B2(n20069), .ZN(
        n20558) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20185), .ZN(n20072) );
  OAI211_X1 U22282 ( .C1(n20188), .C2(n20561), .A(n20073), .B(n20072), .ZN(
        P2_U3143) );
  INV_X1 U22283 ( .A(n20569), .ZN(n20075) );
  INV_X1 U22284 ( .A(n20563), .ZN(n20074) );
  AOI21_X1 U22285 ( .B1(n20075), .B2(n20074), .A(n22411), .ZN(n20076) );
  NOR3_X1 U22286 ( .A1(n20145), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20101) );
  NAND2_X1 U22287 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20101), .ZN(
        n20093) );
  NOR2_X1 U22288 ( .A1(n20077), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20562) );
  INV_X1 U22289 ( .A(n20562), .ZN(n20081) );
  NAND2_X1 U22290 ( .A1(n20093), .A2(n20081), .ZN(n20084) );
  AOI21_X1 U22291 ( .B1(n11915), .B2(n20081), .A(n20103), .ZN(n20078) );
  INV_X1 U22292 ( .A(n15512), .ZN(n20099) );
  AOI22_X1 U22293 ( .A1(n20185), .A2(n20569), .B1(n20190), .B2(n20562), .ZN(
        n20087) );
  INV_X1 U22294 ( .A(n20079), .ZN(n20085) );
  INV_X1 U22295 ( .A(n11915), .ZN(n20080) );
  NAND2_X1 U22296 ( .A1(n20080), .A2(n20165), .ZN(n20082) );
  AOI21_X1 U22297 ( .B1(n20082), .B2(n20081), .A(n20525), .ZN(n20083) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20191), .ZN(n20086) );
  OAI211_X1 U22299 ( .C1(n20567), .C2(n20099), .A(n20087), .B(n20086), .ZN(
        P2_U3135) );
  OAI21_X1 U22300 ( .B1(n20092), .B2(n20178), .A(n20167), .ZN(n20096) );
  INV_X1 U22301 ( .A(n20101), .ZN(n20088) );
  OR2_X1 U22302 ( .A1(n20096), .A2(n20088), .ZN(n20091) );
  NAND2_X1 U22303 ( .A1(n11236), .A2(n20093), .ZN(n20089) );
  NAND2_X1 U22304 ( .A1(n20089), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20090) );
  INV_X1 U22305 ( .A(n20093), .ZN(n20568) );
  AOI22_X1 U22306 ( .A1(n20185), .A2(n20576), .B1(n20190), .B2(n20568), .ZN(
        n20098) );
  AOI21_X1 U22307 ( .B1(n20093), .B2(n20192), .A(n20525), .ZN(n20095) );
  NOR2_X1 U22308 ( .A1(n11236), .A2(n20180), .ZN(n20094) );
  OAI22_X1 U22309 ( .A1(n20096), .A2(n20101), .B1(n20095), .B2(n20094), .ZN(
        n20570) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20570), .B1(
        n20569), .B2(n20191), .ZN(n20097) );
  OAI211_X1 U22311 ( .C1(n20574), .C2(n20099), .A(n20098), .B(n20097), .ZN(
        P2_U3127) );
  AND2_X1 U22312 ( .A1(n20122), .A2(n20101), .ZN(n20575) );
  AOI22_X1 U22313 ( .A1(n20191), .A2(n20576), .B1(n20190), .B2(n20575), .ZN(
        n20111) );
  AOI21_X1 U22314 ( .B1(n20487), .B2(n20581), .A(n22411), .ZN(n20102) );
  NOR2_X1 U22315 ( .A1(n20102), .A2(n20192), .ZN(n20106) );
  NOR2_X1 U22316 ( .A1(n20147), .A2(n20132), .ZN(n20582) );
  INV_X1 U22317 ( .A(n20582), .ZN(n20116) );
  INV_X1 U22318 ( .A(n11927), .ZN(n20107) );
  OAI21_X1 U22319 ( .B1(n20107), .B2(n20103), .A(n20165), .ZN(n20104) );
  AOI21_X1 U22320 ( .B1(n20106), .B2(n20116), .A(n20104), .ZN(n20105) );
  OAI21_X1 U22321 ( .B1(n20582), .B2(n20575), .A(n20106), .ZN(n20109) );
  OAI21_X1 U22322 ( .B1(n20107), .B2(n20575), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20108) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n15512), .ZN(n20110) );
  OAI211_X1 U22324 ( .C1(n20207), .C2(n20581), .A(n20111), .B(n20110), .ZN(
        P2_U3119) );
  INV_X1 U22325 ( .A(n20132), .ZN(n20134) );
  NAND2_X1 U22326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20134), .ZN(
        n20114) );
  INV_X1 U22327 ( .A(n20117), .ZN(n20112) );
  OAI21_X1 U22328 ( .B1(n20112), .B2(n20582), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20113) );
  OAI21_X1 U22329 ( .B1(n20114), .B2(n20192), .A(n20113), .ZN(n20583) );
  AOI22_X1 U22330 ( .A1(n20583), .A2(n15512), .B1(n20190), .B2(n20582), .ZN(
        n20121) );
  OAI22_X1 U22331 ( .A1(n20115), .A2(n22411), .B1(n20132), .B2(n20150), .ZN(
        n20119) );
  OAI211_X1 U22332 ( .C1(n20117), .C2(n20180), .A(n20192), .B(n20116), .ZN(
        n20118) );
  NAND3_X1 U22333 ( .A1(n20119), .A2(n20199), .A3(n20118), .ZN(n20585) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20585), .B1(
        n20584), .B2(n20191), .ZN(n20120) );
  OAI211_X1 U22335 ( .C1(n20207), .C2(n20594), .A(n20121), .B(n20120), .ZN(
        P2_U3111) );
  INV_X1 U22336 ( .A(n11919), .ZN(n20123) );
  NAND2_X1 U22337 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20122), .ZN(
        n20160) );
  NOR2_X1 U22338 ( .A1(n20160), .A2(n20132), .ZN(n20588) );
  OAI21_X1 U22339 ( .B1(n20123), .B2(n20588), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20124) );
  OAI21_X1 U22340 ( .B1(n20132), .B2(n20162), .A(n20124), .ZN(n20589) );
  AOI22_X1 U22341 ( .A1(n20589), .A2(n15512), .B1(n20190), .B2(n20588), .ZN(
        n20131) );
  OAI21_X1 U22342 ( .B1(n20488), .B2(n20590), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20125) );
  OAI21_X1 U22343 ( .B1(n20126), .B2(n20132), .A(n20125), .ZN(n20129) );
  AOI21_X1 U22344 ( .B1(n20588), .B2(n20199), .A(n20195), .ZN(n20127) );
  OAI21_X1 U22345 ( .B1(n11919), .B2(n20180), .A(n20127), .ZN(n20128) );
  NAND2_X1 U22346 ( .A1(n20129), .A2(n20128), .ZN(n20591) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20591), .B1(
        n20488), .B2(n20191), .ZN(n20130) );
  OAI211_X1 U22348 ( .C1(n20207), .C2(n20600), .A(n20131), .B(n20130), .ZN(
        P2_U3103) );
  NAND2_X1 U22349 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20150), .ZN(
        n20175) );
  NOR2_X1 U22350 ( .A1(n20175), .A2(n20132), .ZN(n20595) );
  AOI22_X1 U22351 ( .A1(n20185), .A2(n20602), .B1(n20190), .B2(n20595), .ZN(
        n20143) );
  OAI21_X1 U22352 ( .B1(n20133), .B2(n20178), .A(n20167), .ZN(n20141) );
  NAND2_X1 U22353 ( .A1(n20150), .A2(n20134), .ZN(n20140) );
  INV_X1 U22354 ( .A(n20140), .ZN(n20137) );
  OAI21_X1 U22355 ( .B1(n20167), .B2(n20595), .A(n20199), .ZN(n20135) );
  OAI21_X1 U22356 ( .B1(n11912), .B2(n20180), .A(n20135), .ZN(n20136) );
  OAI21_X1 U22357 ( .B1(n20141), .B2(n20137), .A(n20136), .ZN(n20597) );
  INV_X1 U22358 ( .A(n11912), .ZN(n20138) );
  OAI21_X1 U22359 ( .B1(n20138), .B2(n20595), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20139) );
  OAI21_X1 U22360 ( .B1(n20141), .B2(n20140), .A(n20139), .ZN(n20596) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20597), .B1(
        n15512), .B2(n20596), .ZN(n20142) );
  OAI211_X1 U22362 ( .C1(n20188), .C2(n20600), .A(n20143), .B(n20142), .ZN(
        P2_U3095) );
  NAND2_X1 U22363 ( .A1(n20146), .A2(n20145), .ZN(n20174) );
  NOR2_X1 U22364 ( .A1(n20147), .A2(n20174), .ZN(n20609) );
  AOI22_X1 U22365 ( .A1(n20191), .A2(n20603), .B1(n20190), .B2(n20609), .ZN(
        n20159) );
  OAI21_X1 U22366 ( .B1(n20149), .B2(n20148), .A(n20167), .ZN(n20157) );
  NOR2_X1 U22367 ( .A1(n20150), .A2(n20174), .ZN(n20153) );
  OAI21_X1 U22368 ( .B1(n20167), .B2(n20609), .A(n20199), .ZN(n20151) );
  OAI21_X1 U22369 ( .B1(n11918), .B2(n20180), .A(n20151), .ZN(n20152) );
  OAI21_X1 U22370 ( .B1(n20157), .B2(n20153), .A(n20152), .ZN(n20612) );
  INV_X1 U22371 ( .A(n20153), .ZN(n20156) );
  INV_X1 U22372 ( .A(n11918), .ZN(n20154) );
  OAI21_X1 U22373 ( .B1(n20154), .B2(n20609), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20155) );
  OAI21_X1 U22374 ( .B1(n20157), .B2(n20156), .A(n20155), .ZN(n20611) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20612), .B1(
        n15512), .B2(n20611), .ZN(n20158) );
  OAI211_X1 U22376 ( .C1(n20207), .C2(n20622), .A(n20159), .B(n20158), .ZN(
        P2_U3079) );
  INV_X1 U22377 ( .A(n11931), .ZN(n20166) );
  NOR2_X1 U22378 ( .A1(n20160), .A2(n20174), .ZN(n20616) );
  OAI21_X1 U22379 ( .B1(n20166), .B2(n20616), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20161) );
  AOI22_X1 U22380 ( .A1(n20617), .A2(n15512), .B1(n20190), .B2(n20616), .ZN(
        n20173) );
  NOR2_X1 U22381 ( .A1(n20162), .A2(n20174), .ZN(n20171) );
  NOR2_X2 U22382 ( .A1(n20184), .A2(n20163), .ZN(n20626) );
  INV_X1 U22383 ( .A(n20626), .ZN(n20400) );
  AOI21_X1 U22384 ( .B1(n20622), .B2(n20400), .A(n20164), .ZN(n20170) );
  AOI21_X1 U22385 ( .B1(n20166), .B2(n20165), .A(n20616), .ZN(n20168) );
  NOR3_X1 U22386 ( .A1(n20168), .A2(n20167), .A3(n20525), .ZN(n20169) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20185), .ZN(n20172) );
  OAI211_X1 U22388 ( .C1(n20188), .C2(n20622), .A(n20173), .B(n20172), .ZN(
        P2_U3071) );
  OR2_X1 U22389 ( .A1(n20174), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20189) );
  INV_X1 U22390 ( .A(n11924), .ZN(n20176) );
  NOR2_X1 U22391 ( .A1(n20175), .A2(n20174), .ZN(n20624) );
  OAI21_X1 U22392 ( .B1(n20176), .B2(n20624), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20177) );
  OAI21_X1 U22393 ( .B1(n20189), .B2(n20192), .A(n20177), .ZN(n20625) );
  AOI22_X1 U22394 ( .A1(n20625), .A2(n15512), .B1(n20190), .B2(n20624), .ZN(
        n20187) );
  OAI21_X1 U22395 ( .B1(n20184), .B2(n20178), .A(n20189), .ZN(n20182) );
  AOI21_X1 U22396 ( .B1(n20624), .B2(n20199), .A(n20195), .ZN(n20179) );
  OAI21_X1 U22397 ( .B1(n11924), .B2(n20180), .A(n20179), .ZN(n20181) );
  NAND2_X1 U22398 ( .A1(n20182), .A2(n20181), .ZN(n20627) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20627), .B1(
        n20633), .B2(n20185), .ZN(n20186) );
  OAI211_X1 U22400 ( .C1(n20188), .C2(n20400), .A(n20187), .B(n20186), .ZN(
        P2_U3063) );
  NOR2_X1 U22401 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20189), .ZN(
        n20631) );
  AOI22_X1 U22402 ( .A1(n20191), .A2(n20633), .B1(n20190), .B2(n20631), .ZN(
        n20206) );
  AOI21_X1 U22403 ( .B1(n20640), .B2(n20630), .A(n22411), .ZN(n20193) );
  NOR2_X1 U22404 ( .A1(n20193), .A2(n20192), .ZN(n20201) );
  INV_X1 U22405 ( .A(n20194), .ZN(n20202) );
  AOI21_X1 U22406 ( .B1(n20202), .B2(n20196), .A(n20195), .ZN(n20197) );
  AOI21_X1 U22407 ( .B1(n20201), .B2(n20198), .A(n20197), .ZN(n20200) );
  OAI21_X1 U22408 ( .B1(n20529), .B2(n20631), .A(n20201), .ZN(n20204) );
  OAI21_X1 U22409 ( .B1(n20202), .B2(n20631), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20203) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20637), .B1(
        n15512), .B2(n20636), .ZN(n20205) );
  OAI211_X1 U22411 ( .C1(n20207), .C2(n20640), .A(n20206), .B(n20205), .ZN(
        P2_U3055) );
  OAI222_X1 U22412 ( .A1(n20210), .A2(n20209), .B1(n20208), .B2(n20513), .C1(
        n20465), .C2(n20213), .ZN(P2_U2913) );
  OAI22_X2 U22413 ( .A1(n20913), .A2(n20212), .B1(n21496), .B2(n20211), .ZN(
        n20249) );
  INV_X1 U22414 ( .A(n20249), .ZN(n20245) );
  NOR2_X2 U22415 ( .A1(n11732), .A2(n20527), .ZN(n20248) );
  AOI22_X1 U22416 ( .A1(n20530), .A2(n20214), .B1(n20529), .B2(n20248), .ZN(
        n20216) );
  AOI22_X1 U22417 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20531), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20532), .ZN(n20252) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20534), .B1(
        n20471), .B2(n20242), .ZN(n20215) );
  OAI211_X1 U22419 ( .C1(n20245), .C2(n20640), .A(n20216), .B(n20215), .ZN(
        P2_U3174) );
  AOI22_X1 U22420 ( .A1(n20249), .A2(n20471), .B1(n20248), .B2(n20537), .ZN(
        n20218) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20540), .B1(
        n20214), .B2(n20539), .ZN(n20217) );
  OAI211_X1 U22422 ( .C1(n20252), .C2(n20549), .A(n20218), .B(n20217), .ZN(
        P2_U3166) );
  AOI22_X1 U22423 ( .A1(n20545), .A2(n20214), .B1(n20544), .B2(n20248), .ZN(
        n20220) );
  AOI22_X1 U22424 ( .A1(n20552), .A2(n20242), .B1(n20538), .B2(n20249), .ZN(
        n20219) );
  OAI211_X1 U22425 ( .C1(n20422), .C2(n11935), .A(n20220), .B(n20219), .ZN(
        P2_U3158) );
  AOI22_X1 U22426 ( .A1(n20551), .A2(n20214), .B1(n20550), .B2(n20248), .ZN(
        n20222) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20249), .ZN(n20221) );
  OAI211_X1 U22428 ( .C1(n20252), .C2(n20561), .A(n20222), .B(n20221), .ZN(
        P2_U3150) );
  AOI22_X1 U22429 ( .A1(n20557), .A2(n20214), .B1(n20248), .B2(n20556), .ZN(
        n20224) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20242), .ZN(n20223) );
  OAI211_X1 U22431 ( .C1(n20245), .C2(n20561), .A(n20224), .B(n20223), .ZN(
        P2_U3142) );
  INV_X1 U22432 ( .A(n20214), .ZN(n20229) );
  AOI22_X1 U22433 ( .A1(n20249), .A2(n20563), .B1(n20248), .B2(n20562), .ZN(
        n20226) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20564), .B1(
        n20569), .B2(n20242), .ZN(n20225) );
  OAI211_X1 U22435 ( .C1(n20567), .C2(n20229), .A(n20226), .B(n20225), .ZN(
        P2_U3134) );
  AOI22_X1 U22436 ( .A1(n20249), .A2(n20569), .B1(n20248), .B2(n20568), .ZN(
        n20228) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20570), .B1(
        n20576), .B2(n20242), .ZN(n20227) );
  OAI211_X1 U22438 ( .C1(n20574), .C2(n20229), .A(n20228), .B(n20227), .ZN(
        P2_U3126) );
  AOI22_X1 U22439 ( .A1(n20242), .A2(n20584), .B1(n20248), .B2(n20575), .ZN(
        n20231) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20214), .ZN(n20230) );
  OAI211_X1 U22441 ( .C1(n20245), .C2(n20487), .A(n20231), .B(n20230), .ZN(
        P2_U3118) );
  AOI22_X1 U22442 ( .A1(n20583), .A2(n20214), .B1(n20582), .B2(n20248), .ZN(
        n20233) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20585), .B1(
        n20488), .B2(n20242), .ZN(n20232) );
  OAI211_X1 U22444 ( .C1(n20245), .C2(n20581), .A(n20233), .B(n20232), .ZN(
        P2_U3110) );
  AOI22_X1 U22445 ( .A1(n20589), .A2(n20214), .B1(n20588), .B2(n20248), .ZN(
        n20235) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20591), .B1(
        n20488), .B2(n20249), .ZN(n20234) );
  OAI211_X1 U22447 ( .C1(n20252), .C2(n20600), .A(n20235), .B(n20234), .ZN(
        P2_U3102) );
  AOI22_X1 U22448 ( .A1(n20242), .A2(n20602), .B1(n20595), .B2(n20248), .ZN(
        n20237) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20597), .B1(
        n20214), .B2(n20596), .ZN(n20236) );
  OAI211_X1 U22450 ( .C1(n20245), .C2(n20600), .A(n20237), .B(n20236), .ZN(
        P2_U3094) );
  AOI22_X1 U22451 ( .A1(n20249), .A2(n20602), .B1(n20601), .B2(n20248), .ZN(
        n20239) );
  AOI22_X1 U22452 ( .A1(n20214), .A2(n20604), .B1(n20603), .B2(n20242), .ZN(
        n20238) );
  OAI211_X1 U22453 ( .C1(n20608), .C2(n11928), .A(n20239), .B(n20238), .ZN(
        P2_U3086) );
  AOI22_X1 U22454 ( .A1(n20249), .A2(n20603), .B1(n20609), .B2(n20248), .ZN(
        n20241) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20612), .B1(
        n20214), .B2(n20611), .ZN(n20240) );
  OAI211_X1 U22456 ( .C1(n20252), .C2(n20622), .A(n20241), .B(n20240), .ZN(
        P2_U3078) );
  AOI22_X1 U22457 ( .A1(n20617), .A2(n20214), .B1(n20248), .B2(n20616), .ZN(
        n20244) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20242), .ZN(n20243) );
  OAI211_X1 U22459 ( .C1(n20245), .C2(n20622), .A(n20244), .B(n20243), .ZN(
        P2_U3070) );
  AOI22_X1 U22460 ( .A1(n20625), .A2(n20214), .B1(n20248), .B2(n20624), .ZN(
        n20247) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20627), .B1(
        n20626), .B2(n20249), .ZN(n20246) );
  OAI211_X1 U22462 ( .C1(n20252), .C2(n20630), .A(n20247), .B(n20246), .ZN(
        P2_U3062) );
  AOI22_X1 U22463 ( .A1(n20249), .A2(n20633), .B1(n20248), .B2(n20631), .ZN(
        n20251) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20214), .ZN(n20250) );
  OAI211_X1 U22465 ( .C1(n20252), .C2(n20640), .A(n20251), .B(n20250), .ZN(
        P2_U3054) );
  AOI22_X1 U22466 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n20457), .B1(n20254), .B2(
        n20253), .ZN(n20267) );
  NOR2_X1 U22467 ( .A1(n20255), .A2(n20458), .ZN(n20258) );
  AOI21_X1 U22468 ( .B1(n20255), .B2(n20458), .A(n20258), .ZN(n20460) );
  INV_X1 U22469 ( .A(n20460), .ZN(n20256) );
  NOR2_X1 U22470 ( .A1(n20519), .A2(n20518), .ZN(n20516) );
  NOR2_X1 U22471 ( .A1(n20256), .A2(n20516), .ZN(n20257) );
  NOR2_X1 U22472 ( .A1(n20258), .A2(n20257), .ZN(n20259) );
  XOR2_X1 U22473 ( .A(n20408), .B(n20259), .Z(n20410) );
  INV_X1 U22474 ( .A(n20410), .ZN(n20261) );
  NAND2_X1 U22475 ( .A1(n20259), .A2(n20408), .ZN(n20260) );
  OAI21_X1 U22476 ( .B1(n20261), .B2(n20409), .A(n20260), .ZN(n20360) );
  XNOR2_X1 U22477 ( .A(n20262), .B(n20263), .ZN(n20361) );
  NOR2_X1 U22478 ( .A1(n20360), .A2(n20361), .ZN(n20359) );
  AOI21_X1 U22479 ( .B1(n20263), .B2(n20262), .A(n20359), .ZN(n20265) );
  INV_X1 U22480 ( .A(n20310), .ZN(n20264) );
  NOR2_X1 U22481 ( .A1(n20265), .A2(n20264), .ZN(n20312) );
  OR3_X1 U22482 ( .A1(n20312), .A2(n20313), .A3(n20517), .ZN(n20266) );
  OAI211_X1 U22483 ( .C1(n20268), .C2(n20465), .A(n20267), .B(n20266), .ZN(
        P2_U2914) );
  AOI22_X1 U22484 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20531), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20532), .ZN(n20300) );
  NOR2_X2 U22485 ( .A1(n20268), .A2(n20525), .ZN(n20306) );
  AOI22_X1 U22486 ( .A1(n20530), .A2(n20306), .B1(n20529), .B2(n20270), .ZN(
        n20272) );
  AOI22_X1 U22487 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20531), .ZN(n20309) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20534), .B1(
        n20533), .B2(n20297), .ZN(n20271) );
  OAI211_X1 U22489 ( .C1(n20300), .C2(n20543), .A(n20272), .B(n20271), .ZN(
        P2_U3173) );
  AOI22_X1 U22490 ( .A1(n20297), .A2(n20471), .B1(n20270), .B2(n20537), .ZN(
        n20274) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20540), .B1(
        n20306), .B2(n20539), .ZN(n20273) );
  OAI211_X1 U22492 ( .C1(n20300), .C2(n20549), .A(n20274), .B(n20273), .ZN(
        P2_U3165) );
  INV_X1 U22493 ( .A(n20552), .ZN(n20373) );
  AOI22_X1 U22494 ( .A1(n20545), .A2(n20306), .B1(n20544), .B2(n20270), .ZN(
        n20276) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20546), .B1(
        n20538), .B2(n20297), .ZN(n20275) );
  OAI211_X1 U22496 ( .C1(n20300), .C2(n20373), .A(n20276), .B(n20275), .ZN(
        P2_U3157) );
  AOI22_X1 U22497 ( .A1(n20551), .A2(n20306), .B1(n20550), .B2(n20270), .ZN(
        n20278) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20297), .ZN(n20277) );
  OAI211_X1 U22499 ( .C1(n20300), .C2(n20561), .A(n20278), .B(n20277), .ZN(
        P2_U3149) );
  AOI22_X1 U22500 ( .A1(n20557), .A2(n20306), .B1(n20270), .B2(n20556), .ZN(
        n20280) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20305), .ZN(n20279) );
  OAI211_X1 U22502 ( .C1(n20309), .C2(n20561), .A(n20280), .B(n20279), .ZN(
        P2_U3141) );
  INV_X1 U22503 ( .A(n20306), .ZN(n20285) );
  AOI22_X1 U22504 ( .A1(n20305), .A2(n20569), .B1(n20270), .B2(n20562), .ZN(
        n20282) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20297), .ZN(n20281) );
  OAI211_X1 U22506 ( .C1(n20567), .C2(n20285), .A(n20282), .B(n20281), .ZN(
        P2_U3133) );
  AOI22_X1 U22507 ( .A1(n20297), .A2(n20569), .B1(n20270), .B2(n20568), .ZN(
        n20284) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20570), .B1(
        n20576), .B2(n20305), .ZN(n20283) );
  OAI211_X1 U22509 ( .C1(n20574), .C2(n20285), .A(n20284), .B(n20283), .ZN(
        P2_U3125) );
  AOI22_X1 U22510 ( .A1(n20305), .A2(n20584), .B1(n20270), .B2(n20575), .ZN(
        n20287) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20306), .ZN(n20286) );
  OAI211_X1 U22512 ( .C1(n20309), .C2(n20487), .A(n20287), .B(n20286), .ZN(
        P2_U3117) );
  AOI22_X1 U22513 ( .A1(n20583), .A2(n20306), .B1(n20582), .B2(n20270), .ZN(
        n20289) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20585), .B1(
        n20584), .B2(n20297), .ZN(n20288) );
  OAI211_X1 U22515 ( .C1(n20300), .C2(n20594), .A(n20289), .B(n20288), .ZN(
        P2_U3109) );
  AOI22_X1 U22516 ( .A1(n20589), .A2(n20306), .B1(n20588), .B2(n20270), .ZN(
        n20291) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20591), .B1(
        n20488), .B2(n20297), .ZN(n20290) );
  OAI211_X1 U22518 ( .C1(n20300), .C2(n20600), .A(n20291), .B(n20290), .ZN(
        P2_U3101) );
  AOI22_X1 U22519 ( .A1(n20305), .A2(n20602), .B1(n20595), .B2(n20270), .ZN(
        n20293) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20597), .B1(
        n20306), .B2(n20596), .ZN(n20292) );
  OAI211_X1 U22521 ( .C1(n20309), .C2(n20600), .A(n20293), .B(n20292), .ZN(
        P2_U3093) );
  INV_X1 U22522 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n20296) );
  AOI22_X1 U22523 ( .A1(n20297), .A2(n20602), .B1(n20601), .B2(n20270), .ZN(
        n20295) );
  AOI22_X1 U22524 ( .A1(n20306), .A2(n20604), .B1(n20603), .B2(n20305), .ZN(
        n20294) );
  OAI211_X1 U22525 ( .C1(n20608), .C2(n20296), .A(n20295), .B(n20294), .ZN(
        P2_U3085) );
  AOI22_X1 U22526 ( .A1(n20297), .A2(n20603), .B1(n20609), .B2(n20270), .ZN(
        n20299) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20612), .B1(
        n20306), .B2(n20611), .ZN(n20298) );
  OAI211_X1 U22528 ( .C1(n20300), .C2(n20622), .A(n20299), .B(n20298), .ZN(
        P2_U3077) );
  AOI22_X1 U22529 ( .A1(n20617), .A2(n20306), .B1(n20270), .B2(n20616), .ZN(
        n20302) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20305), .ZN(n20301) );
  OAI211_X1 U22531 ( .C1(n20309), .C2(n20622), .A(n20302), .B(n20301), .ZN(
        P2_U3069) );
  AOI22_X1 U22532 ( .A1(n20625), .A2(n20306), .B1(n20270), .B2(n20624), .ZN(
        n20304) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20627), .B1(
        n20633), .B2(n20305), .ZN(n20303) );
  OAI211_X1 U22534 ( .C1(n20309), .C2(n20400), .A(n20304), .B(n20303), .ZN(
        P2_U3061) );
  AOI22_X1 U22535 ( .A1(n20305), .A2(n20533), .B1(n20270), .B2(n20631), .ZN(
        n20308) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20306), .ZN(n20307) );
  OAI211_X1 U22537 ( .C1(n20309), .C2(n20630), .A(n20308), .B(n20307), .ZN(
        P2_U3053) );
  OAI22_X1 U22538 ( .A1(n20310), .A2(n20515), .B1(n20513), .B2(n18247), .ZN(
        n20311) );
  INV_X1 U22539 ( .A(n20311), .ZN(n20316) );
  XOR2_X1 U22540 ( .A(n20313), .B(n20312), .Z(n20314) );
  NAND2_X1 U22541 ( .A1(n20314), .A2(n20461), .ZN(n20315) );
  OAI211_X1 U22542 ( .C1(n20317), .C2(n20465), .A(n20316), .B(n20315), .ZN(
        P2_U2915) );
  AOI22_X1 U22543 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20531), .ZN(n20351) );
  NOR2_X2 U22544 ( .A1(n20317), .A2(n20525), .ZN(n20354) );
  NOR2_X2 U22545 ( .A1(n11725), .A2(n20527), .ZN(n20352) );
  AOI22_X1 U22546 ( .A1(n20530), .A2(n20354), .B1(n20529), .B2(n20352), .ZN(
        n20319) );
  AOI22_X1 U22547 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20531), .ZN(n20357) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20534), .B1(
        n20533), .B2(n20348), .ZN(n20318) );
  OAI211_X1 U22549 ( .C1(n20351), .C2(n20543), .A(n20319), .B(n20318), .ZN(
        P2_U3172) );
  AOI22_X1 U22550 ( .A1(n20348), .A2(n20471), .B1(n20352), .B2(n20537), .ZN(
        n20321) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20540), .B1(
        n20354), .B2(n20539), .ZN(n20320) );
  OAI211_X1 U22552 ( .C1(n20351), .C2(n20549), .A(n20321), .B(n20320), .ZN(
        P2_U3164) );
  AOI22_X1 U22553 ( .A1(n20545), .A2(n20354), .B1(n20544), .B2(n20352), .ZN(
        n20323) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20546), .B1(
        n20538), .B2(n20348), .ZN(n20322) );
  OAI211_X1 U22555 ( .C1(n20351), .C2(n20373), .A(n20323), .B(n20322), .ZN(
        P2_U3156) );
  AOI22_X1 U22556 ( .A1(n20551), .A2(n20354), .B1(n20550), .B2(n20352), .ZN(
        n20325) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20348), .ZN(n20324) );
  OAI211_X1 U22558 ( .C1(n20351), .C2(n20561), .A(n20325), .B(n20324), .ZN(
        P2_U3148) );
  AOI22_X1 U22559 ( .A1(n20557), .A2(n20354), .B1(n20352), .B2(n20556), .ZN(
        n20327) );
  INV_X1 U22560 ( .A(n20351), .ZN(n20353) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20353), .ZN(n20326) );
  OAI211_X1 U22562 ( .C1(n20357), .C2(n20561), .A(n20327), .B(n20326), .ZN(
        P2_U3140) );
  INV_X1 U22563 ( .A(n20354), .ZN(n20332) );
  AOI22_X1 U22564 ( .A1(n20348), .A2(n20563), .B1(n20352), .B2(n20562), .ZN(
        n20329) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20564), .B1(
        n20569), .B2(n20353), .ZN(n20328) );
  OAI211_X1 U22566 ( .C1(n20567), .C2(n20332), .A(n20329), .B(n20328), .ZN(
        P2_U3132) );
  AOI22_X1 U22567 ( .A1(n20348), .A2(n20569), .B1(n20352), .B2(n20568), .ZN(
        n20331) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20570), .B1(
        n20576), .B2(n20353), .ZN(n20330) );
  OAI211_X1 U22569 ( .C1(n20574), .C2(n20332), .A(n20331), .B(n20330), .ZN(
        P2_U3124) );
  AOI22_X1 U22570 ( .A1(n20348), .A2(n20576), .B1(n20352), .B2(n20575), .ZN(
        n20334) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20354), .ZN(n20333) );
  OAI211_X1 U22572 ( .C1(n20351), .C2(n20581), .A(n20334), .B(n20333), .ZN(
        P2_U3116) );
  AOI22_X1 U22573 ( .A1(n20583), .A2(n20354), .B1(n20582), .B2(n20352), .ZN(
        n20336) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20585), .B1(
        n20488), .B2(n20353), .ZN(n20335) );
  OAI211_X1 U22575 ( .C1(n20357), .C2(n20581), .A(n20336), .B(n20335), .ZN(
        P2_U3108) );
  AOI22_X1 U22576 ( .A1(n20589), .A2(n20354), .B1(n20588), .B2(n20352), .ZN(
        n20338) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20591), .B1(
        n20488), .B2(n20348), .ZN(n20337) );
  OAI211_X1 U22578 ( .C1(n20351), .C2(n20600), .A(n20338), .B(n20337), .ZN(
        P2_U3100) );
  AOI22_X1 U22579 ( .A1(n20348), .A2(n20590), .B1(n20352), .B2(n20595), .ZN(
        n20340) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20597), .B1(
        n20354), .B2(n20596), .ZN(n20339) );
  OAI211_X1 U22581 ( .C1(n20351), .C2(n20495), .A(n20340), .B(n20339), .ZN(
        P2_U3092) );
  INV_X1 U22582 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n20343) );
  AOI22_X1 U22583 ( .A1(n20348), .A2(n20602), .B1(n20601), .B2(n20352), .ZN(
        n20342) );
  AOI22_X1 U22584 ( .A1(n20354), .A2(n20604), .B1(n20603), .B2(n20353), .ZN(
        n20341) );
  OAI211_X1 U22585 ( .C1(n20608), .C2(n20343), .A(n20342), .B(n20341), .ZN(
        P2_U3084) );
  AOI22_X1 U22586 ( .A1(n20348), .A2(n20603), .B1(n20609), .B2(n20352), .ZN(
        n20345) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20612), .B1(
        n20354), .B2(n20611), .ZN(n20344) );
  OAI211_X1 U22588 ( .C1(n20351), .C2(n20622), .A(n20345), .B(n20344), .ZN(
        P2_U3076) );
  AOI22_X1 U22589 ( .A1(n20617), .A2(n20354), .B1(n20352), .B2(n20616), .ZN(
        n20347) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20353), .ZN(n20346) );
  OAI211_X1 U22591 ( .C1(n20357), .C2(n20622), .A(n20347), .B(n20346), .ZN(
        P2_U3068) );
  AOI22_X1 U22592 ( .A1(n20625), .A2(n20354), .B1(n20352), .B2(n20624), .ZN(
        n20350) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20627), .B1(
        n20626), .B2(n20348), .ZN(n20349) );
  OAI211_X1 U22594 ( .C1(n20351), .C2(n20630), .A(n20350), .B(n20349), .ZN(
        P2_U3060) );
  AOI22_X1 U22595 ( .A1(n20353), .A2(n20533), .B1(n20352), .B2(n20631), .ZN(
        n20356) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20354), .ZN(n20355) );
  OAI211_X1 U22597 ( .C1(n20357), .C2(n20630), .A(n20356), .B(n20355), .ZN(
        P2_U3052) );
  AOI22_X1 U22598 ( .A1(n20459), .A2(n20358), .B1(n20457), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n20364) );
  AOI21_X1 U22599 ( .B1(n20361), .B2(n20360), .A(n20359), .ZN(n20362) );
  OR2_X1 U22600 ( .A1(n20362), .A2(n20517), .ZN(n20363) );
  OAI211_X1 U22601 ( .C1(n20365), .C2(n20465), .A(n20364), .B(n20363), .ZN(
        P2_U2916) );
  INV_X1 U22602 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20368) );
  NOR2_X2 U22603 ( .A1(n20365), .A2(n20525), .ZN(n20404) );
  NOR2_X2 U22604 ( .A1(n11728), .A2(n20527), .ZN(n20402) );
  AOI22_X1 U22605 ( .A1(n20530), .A2(n20404), .B1(n20529), .B2(n20402), .ZN(
        n20367) );
  AOI22_X1 U22606 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20531), .ZN(n20401) );
  AOI22_X1 U22607 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20531), .ZN(n20407) );
  INV_X1 U22608 ( .A(n20407), .ZN(n20397) );
  AOI22_X1 U22609 ( .A1(n20533), .A2(n20403), .B1(n20471), .B2(n20397), .ZN(
        n20366) );
  OAI211_X1 U22610 ( .C1(n20470), .C2(n20368), .A(n20367), .B(n20366), .ZN(
        P2_U3171) );
  AOI22_X1 U22611 ( .A1(n20403), .A2(n20471), .B1(n20402), .B2(n20537), .ZN(
        n20370) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20540), .B1(
        n20404), .B2(n20539), .ZN(n20369) );
  OAI211_X1 U22613 ( .C1(n20407), .C2(n20549), .A(n20370), .B(n20369), .ZN(
        P2_U3163) );
  AOI22_X1 U22614 ( .A1(n20545), .A2(n20404), .B1(n20544), .B2(n20402), .ZN(
        n20372) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20546), .B1(
        n20538), .B2(n20403), .ZN(n20371) );
  OAI211_X1 U22616 ( .C1(n20407), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P2_U3155) );
  AOI22_X1 U22617 ( .A1(n20551), .A2(n20404), .B1(n20550), .B2(n20402), .ZN(
        n20375) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20403), .ZN(n20374) );
  OAI211_X1 U22619 ( .C1(n20407), .C2(n20561), .A(n20375), .B(n20374), .ZN(
        P2_U3147) );
  AOI22_X1 U22620 ( .A1(n20557), .A2(n20404), .B1(n20402), .B2(n20556), .ZN(
        n20377) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20397), .ZN(n20376) );
  OAI211_X1 U22622 ( .C1(n20401), .C2(n20561), .A(n20377), .B(n20376), .ZN(
        P2_U3139) );
  INV_X1 U22623 ( .A(n20404), .ZN(n20382) );
  AOI22_X1 U22624 ( .A1(n20403), .A2(n20563), .B1(n20402), .B2(n20562), .ZN(
        n20379) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20564), .B1(
        n20569), .B2(n20397), .ZN(n20378) );
  OAI211_X1 U22626 ( .C1(n20567), .C2(n20382), .A(n20379), .B(n20378), .ZN(
        P2_U3131) );
  AOI22_X1 U22627 ( .A1(n20397), .A2(n20576), .B1(n20402), .B2(n20568), .ZN(
        n20381) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20570), .B1(
        n20569), .B2(n20403), .ZN(n20380) );
  OAI211_X1 U22629 ( .C1(n20574), .C2(n20382), .A(n20381), .B(n20380), .ZN(
        P2_U3123) );
  AOI22_X1 U22630 ( .A1(n20403), .A2(n20576), .B1(n20402), .B2(n20575), .ZN(
        n20384) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20404), .ZN(n20383) );
  OAI211_X1 U22632 ( .C1(n20407), .C2(n20581), .A(n20384), .B(n20383), .ZN(
        P2_U3115) );
  AOI22_X1 U22633 ( .A1(n20583), .A2(n20404), .B1(n20582), .B2(n20402), .ZN(
        n20386) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20585), .B1(
        n20584), .B2(n20403), .ZN(n20385) );
  OAI211_X1 U22635 ( .C1(n20407), .C2(n20594), .A(n20386), .B(n20385), .ZN(
        P2_U3107) );
  AOI22_X1 U22636 ( .A1(n20589), .A2(n20404), .B1(n20588), .B2(n20402), .ZN(
        n20388) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20591), .B1(
        n20488), .B2(n20403), .ZN(n20387) );
  OAI211_X1 U22638 ( .C1(n20407), .C2(n20600), .A(n20388), .B(n20387), .ZN(
        P2_U3099) );
  AOI22_X1 U22639 ( .A1(n20397), .A2(n20602), .B1(n20595), .B2(n20402), .ZN(
        n20390) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20597), .B1(
        n20404), .B2(n20596), .ZN(n20389) );
  OAI211_X1 U22641 ( .C1(n20401), .C2(n20600), .A(n20390), .B(n20389), .ZN(
        P2_U3091) );
  AOI22_X1 U22642 ( .A1(n20403), .A2(n20602), .B1(n20601), .B2(n20402), .ZN(
        n20392) );
  AOI22_X1 U22643 ( .A1(n20404), .A2(n20604), .B1(n20603), .B2(n20397), .ZN(
        n20391) );
  OAI211_X1 U22644 ( .C1(n20608), .C2(n11902), .A(n20392), .B(n20391), .ZN(
        P2_U3083) );
  AOI22_X1 U22645 ( .A1(n20403), .A2(n20603), .B1(n20609), .B2(n20402), .ZN(
        n20394) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20612), .B1(
        n20404), .B2(n20611), .ZN(n20393) );
  OAI211_X1 U22647 ( .C1(n20407), .C2(n20622), .A(n20394), .B(n20393), .ZN(
        P2_U3075) );
  AOI22_X1 U22648 ( .A1(n20617), .A2(n20404), .B1(n20402), .B2(n20616), .ZN(
        n20396) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20397), .ZN(n20395) );
  OAI211_X1 U22650 ( .C1(n20401), .C2(n20622), .A(n20396), .B(n20395), .ZN(
        P2_U3067) );
  AOI22_X1 U22651 ( .A1(n20625), .A2(n20404), .B1(n20402), .B2(n20624), .ZN(
        n20399) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20627), .B1(
        n20633), .B2(n20397), .ZN(n20398) );
  OAI211_X1 U22653 ( .C1(n20401), .C2(n20400), .A(n20399), .B(n20398), .ZN(
        P2_U3059) );
  AOI22_X1 U22654 ( .A1(n20403), .A2(n20633), .B1(n20402), .B2(n20631), .ZN(
        n20406) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20404), .ZN(n20405) );
  OAI211_X1 U22656 ( .C1(n20407), .C2(n20640), .A(n20406), .B(n20405), .ZN(
        P2_U3051) );
  AOI22_X1 U22657 ( .A1(n20408), .A2(n20459), .B1(n20457), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n20413) );
  XNOR2_X1 U22658 ( .A(n20410), .B(n20409), .ZN(n20411) );
  NAND2_X1 U22659 ( .A1(n20411), .A2(n20461), .ZN(n20412) );
  OAI211_X1 U22660 ( .C1(n20414), .C2(n20465), .A(n20413), .B(n20412), .ZN(
        P2_U2917) );
  AOI22_X1 U22661 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20531), .ZN(n20450) );
  NOR2_X2 U22662 ( .A1(n20414), .A2(n20525), .ZN(n20453) );
  NOR2_X2 U22663 ( .A1(n11727), .A2(n20527), .ZN(n20451) );
  AOI22_X1 U22664 ( .A1(n20530), .A2(n20453), .B1(n20529), .B2(n20451), .ZN(
        n20416) );
  AOI22_X1 U22665 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20531), .ZN(n20456) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20534), .B1(
        n20533), .B2(n20447), .ZN(n20415) );
  OAI211_X1 U22667 ( .C1(n20450), .C2(n20543), .A(n20416), .B(n20415), .ZN(
        P2_U3170) );
  AOI22_X1 U22668 ( .A1(n20447), .A2(n20471), .B1(n20451), .B2(n20537), .ZN(
        n20418) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20540), .B1(
        n20453), .B2(n20539), .ZN(n20417) );
  OAI211_X1 U22670 ( .C1(n20450), .C2(n20549), .A(n20418), .B(n20417), .ZN(
        P2_U3162) );
  INV_X1 U22671 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U22672 ( .A1(n20545), .A2(n20453), .B1(n20544), .B2(n20451), .ZN(
        n20420) );
  AOI22_X1 U22673 ( .A1(n20552), .A2(n20452), .B1(n20538), .B2(n20447), .ZN(
        n20419) );
  OAI211_X1 U22674 ( .C1(n20422), .C2(n20421), .A(n20420), .B(n20419), .ZN(
        P2_U3154) );
  AOI22_X1 U22675 ( .A1(n20551), .A2(n20453), .B1(n20550), .B2(n20451), .ZN(
        n20424) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20447), .ZN(n20423) );
  OAI211_X1 U22677 ( .C1(n20450), .C2(n20561), .A(n20424), .B(n20423), .ZN(
        P2_U3146) );
  AOI22_X1 U22678 ( .A1(n20557), .A2(n20453), .B1(n20451), .B2(n20556), .ZN(
        n20426) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20452), .ZN(n20425) );
  OAI211_X1 U22680 ( .C1(n20456), .C2(n20561), .A(n20426), .B(n20425), .ZN(
        P2_U3138) );
  INV_X1 U22681 ( .A(n20453), .ZN(n20431) );
  AOI22_X1 U22682 ( .A1(n20452), .A2(n20569), .B1(n20451), .B2(n20562), .ZN(
        n20428) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20447), .ZN(n20427) );
  OAI211_X1 U22684 ( .C1(n20567), .C2(n20431), .A(n20428), .B(n20427), .ZN(
        P2_U3130) );
  AOI22_X1 U22685 ( .A1(n20447), .A2(n20569), .B1(n20451), .B2(n20568), .ZN(
        n20430) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20570), .B1(
        n20576), .B2(n20452), .ZN(n20429) );
  OAI211_X1 U22687 ( .C1(n20574), .C2(n20431), .A(n20430), .B(n20429), .ZN(
        P2_U3122) );
  AOI22_X1 U22688 ( .A1(n20452), .A2(n20584), .B1(n20451), .B2(n20575), .ZN(
        n20433) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20453), .ZN(n20432) );
  OAI211_X1 U22690 ( .C1(n20456), .C2(n20487), .A(n20433), .B(n20432), .ZN(
        P2_U3114) );
  AOI22_X1 U22691 ( .A1(n20583), .A2(n20453), .B1(n20582), .B2(n20451), .ZN(
        n20435) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20585), .B1(
        n20584), .B2(n20447), .ZN(n20434) );
  OAI211_X1 U22693 ( .C1(n20450), .C2(n20594), .A(n20435), .B(n20434), .ZN(
        P2_U3106) );
  AOI22_X1 U22694 ( .A1(n20589), .A2(n20453), .B1(n20588), .B2(n20451), .ZN(
        n20437) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20591), .B1(
        n20488), .B2(n20447), .ZN(n20436) );
  OAI211_X1 U22696 ( .C1(n20450), .C2(n20600), .A(n20437), .B(n20436), .ZN(
        P2_U3098) );
  AOI22_X1 U22697 ( .A1(n20447), .A2(n20590), .B1(n20595), .B2(n20451), .ZN(
        n20439) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20597), .B1(
        n20453), .B2(n20596), .ZN(n20438) );
  OAI211_X1 U22699 ( .C1(n20450), .C2(n20495), .A(n20439), .B(n20438), .ZN(
        P2_U3090) );
  INV_X1 U22700 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U22701 ( .A1(n20447), .A2(n20602), .B1(n20601), .B2(n20451), .ZN(
        n20441) );
  AOI22_X1 U22702 ( .A1(n20453), .A2(n20604), .B1(n20603), .B2(n20452), .ZN(
        n20440) );
  OAI211_X1 U22703 ( .C1(n20608), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P2_U3082) );
  AOI22_X1 U22704 ( .A1(n20452), .A2(n20610), .B1(n20609), .B2(n20451), .ZN(
        n20444) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20612), .B1(
        n20453), .B2(n20611), .ZN(n20443) );
  OAI211_X1 U22706 ( .C1(n20456), .C2(n20615), .A(n20444), .B(n20443), .ZN(
        P2_U3074) );
  AOI22_X1 U22707 ( .A1(n20617), .A2(n20453), .B1(n20451), .B2(n20616), .ZN(
        n20446) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20452), .ZN(n20445) );
  OAI211_X1 U22709 ( .C1(n20456), .C2(n20622), .A(n20446), .B(n20445), .ZN(
        P2_U3066) );
  AOI22_X1 U22710 ( .A1(n20625), .A2(n20453), .B1(n20451), .B2(n20624), .ZN(
        n20449) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20627), .B1(
        n20626), .B2(n20447), .ZN(n20448) );
  OAI211_X1 U22712 ( .C1(n20450), .C2(n20630), .A(n20449), .B(n20448), .ZN(
        P2_U3058) );
  AOI22_X1 U22713 ( .A1(n20452), .A2(n20533), .B1(n20451), .B2(n20631), .ZN(
        n20455) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20453), .ZN(n20454) );
  OAI211_X1 U22715 ( .C1(n20456), .C2(n20630), .A(n20455), .B(n20454), .ZN(
        P2_U3050) );
  AOI22_X1 U22716 ( .A1(n20459), .A2(n20458), .B1(n20457), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n20464) );
  XOR2_X1 U22717 ( .A(n20516), .B(n20460), .Z(n20462) );
  NAND2_X1 U22718 ( .A1(n20462), .A2(n20461), .ZN(n20463) );
  OAI211_X1 U22719 ( .C1(n20466), .C2(n20465), .A(n20464), .B(n20463), .ZN(
        P2_U2918) );
  INV_X1 U22720 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20469) );
  NOR2_X2 U22721 ( .A1(n20466), .A2(n20525), .ZN(n20509) );
  NOR2_X2 U22722 ( .A1(n12819), .A2(n20527), .ZN(n20507) );
  AOI22_X1 U22723 ( .A1(n20530), .A2(n20509), .B1(n20529), .B2(n20507), .ZN(
        n20468) );
  AOI22_X1 U22724 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20531), .ZN(n20512) );
  AOI22_X1 U22725 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20531), .ZN(n20506) );
  AOI22_X1 U22726 ( .A1(n20533), .A2(n20503), .B1(n20471), .B2(n20508), .ZN(
        n20467) );
  OAI211_X1 U22727 ( .C1(n20470), .C2(n20469), .A(n20468), .B(n20467), .ZN(
        P2_U3169) );
  AOI22_X1 U22728 ( .A1(n20503), .A2(n20471), .B1(n20507), .B2(n20537), .ZN(
        n20473) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20540), .B1(
        n20509), .B2(n20539), .ZN(n20472) );
  OAI211_X1 U22730 ( .C1(n20506), .C2(n20549), .A(n20473), .B(n20472), .ZN(
        P2_U3161) );
  AOI22_X1 U22731 ( .A1(n20545), .A2(n20509), .B1(n20544), .B2(n20507), .ZN(
        n20475) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20546), .B1(
        n20552), .B2(n20508), .ZN(n20474) );
  OAI211_X1 U22733 ( .C1(n20512), .C2(n20549), .A(n20475), .B(n20474), .ZN(
        P2_U3153) );
  AOI22_X1 U22734 ( .A1(n20551), .A2(n20509), .B1(n20550), .B2(n20507), .ZN(
        n20477) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20503), .ZN(n20476) );
  OAI211_X1 U22736 ( .C1(n20506), .C2(n20561), .A(n20477), .B(n20476), .ZN(
        P2_U3145) );
  AOI22_X1 U22737 ( .A1(n20557), .A2(n20509), .B1(n20507), .B2(n20556), .ZN(
        n20479) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20508), .ZN(n20478) );
  OAI211_X1 U22739 ( .C1(n20512), .C2(n20561), .A(n20479), .B(n20478), .ZN(
        P2_U3137) );
  INV_X1 U22740 ( .A(n20509), .ZN(n20484) );
  AOI22_X1 U22741 ( .A1(n20508), .A2(n20569), .B1(n20507), .B2(n20562), .ZN(
        n20481) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20503), .ZN(n20480) );
  OAI211_X1 U22743 ( .C1(n20567), .C2(n20484), .A(n20481), .B(n20480), .ZN(
        P2_U3129) );
  AOI22_X1 U22744 ( .A1(n20503), .A2(n20569), .B1(n20507), .B2(n20568), .ZN(
        n20483) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20570), .B1(
        n20576), .B2(n20508), .ZN(n20482) );
  OAI211_X1 U22746 ( .C1(n20574), .C2(n20484), .A(n20483), .B(n20482), .ZN(
        P2_U3121) );
  AOI22_X1 U22747 ( .A1(n20508), .A2(n20584), .B1(n20507), .B2(n20575), .ZN(
        n20486) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20509), .ZN(n20485) );
  OAI211_X1 U22749 ( .C1(n20512), .C2(n20487), .A(n20486), .B(n20485), .ZN(
        P2_U3113) );
  AOI22_X1 U22750 ( .A1(n20583), .A2(n20509), .B1(n20582), .B2(n20507), .ZN(
        n20490) );
  AOI22_X1 U22751 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20585), .B1(
        n20488), .B2(n20508), .ZN(n20489) );
  OAI211_X1 U22752 ( .C1(n20512), .C2(n20581), .A(n20490), .B(n20489), .ZN(
        P2_U3105) );
  AOI22_X1 U22753 ( .A1(n20589), .A2(n20509), .B1(n20588), .B2(n20507), .ZN(
        n20492) );
  AOI22_X1 U22754 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20591), .B1(
        n20590), .B2(n20508), .ZN(n20491) );
  OAI211_X1 U22755 ( .C1(n20512), .C2(n20594), .A(n20492), .B(n20491), .ZN(
        P2_U3097) );
  AOI22_X1 U22756 ( .A1(n20503), .A2(n20590), .B1(n20595), .B2(n20507), .ZN(
        n20494) );
  AOI22_X1 U22757 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20597), .B1(
        n20509), .B2(n20596), .ZN(n20493) );
  OAI211_X1 U22758 ( .C1(n20506), .C2(n20495), .A(n20494), .B(n20493), .ZN(
        P2_U3089) );
  AOI22_X1 U22759 ( .A1(n20503), .A2(n20602), .B1(n20601), .B2(n20507), .ZN(
        n20497) );
  AOI22_X1 U22760 ( .A1(n20509), .A2(n20604), .B1(n20603), .B2(n20508), .ZN(
        n20496) );
  OAI211_X1 U22761 ( .C1(n20608), .C2(n20498), .A(n20497), .B(n20496), .ZN(
        P2_U3081) );
  AOI22_X1 U22762 ( .A1(n20503), .A2(n20603), .B1(n20609), .B2(n20507), .ZN(
        n20500) );
  AOI22_X1 U22763 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20612), .B1(
        n20509), .B2(n20611), .ZN(n20499) );
  OAI211_X1 U22764 ( .C1(n20506), .C2(n20622), .A(n20500), .B(n20499), .ZN(
        P2_U3073) );
  AOI22_X1 U22765 ( .A1(n20617), .A2(n20509), .B1(n20507), .B2(n20616), .ZN(
        n20502) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20508), .ZN(n20501) );
  OAI211_X1 U22767 ( .C1(n20512), .C2(n20622), .A(n20502), .B(n20501), .ZN(
        P2_U3065) );
  AOI22_X1 U22768 ( .A1(n20625), .A2(n20509), .B1(n20507), .B2(n20624), .ZN(
        n20505) );
  AOI22_X1 U22769 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20627), .B1(
        n20626), .B2(n20503), .ZN(n20504) );
  OAI211_X1 U22770 ( .C1(n20506), .C2(n20630), .A(n20505), .B(n20504), .ZN(
        P2_U3057) );
  AOI22_X1 U22771 ( .A1(n20508), .A2(n20533), .B1(n20507), .B2(n20631), .ZN(
        n20511) );
  AOI22_X1 U22772 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20509), .ZN(n20510) );
  OAI211_X1 U22773 ( .C1(n20512), .C2(n20630), .A(n20511), .B(n20510), .ZN(
        P2_U3049) );
  INV_X1 U22774 ( .A(n20526), .ZN(n20523) );
  OAI22_X1 U22775 ( .A1(n20515), .A2(n20518), .B1(n20514), .B2(n20513), .ZN(
        n20521) );
  AOI211_X1 U22776 ( .C1(n20519), .C2(n20518), .A(n20517), .B(n20516), .ZN(
        n20520) );
  AOI211_X1 U22777 ( .C1(n20523), .C2(n20522), .A(n20521), .B(n20520), .ZN(
        n20524) );
  INV_X1 U22778 ( .A(n20524), .ZN(P2_U2919) );
  AOI22_X1 U22779 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20531), .ZN(n20641) );
  NOR2_X2 U22780 ( .A1(n20526), .A2(n20525), .ZN(n20635) );
  AOI22_X1 U22781 ( .A1(n20530), .A2(n20635), .B1(n20529), .B2(n11154), .ZN(
        n20536) );
  AOI22_X1 U22782 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20532), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20531), .ZN(n20623) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20534), .B1(
        n20533), .B2(n20634), .ZN(n20535) );
  OAI211_X1 U22784 ( .C1(n20641), .C2(n20543), .A(n20536), .B(n20535), .ZN(
        P2_U3168) );
  AOI22_X1 U22785 ( .A1(n20618), .A2(n20538), .B1(n11154), .B2(n20537), .ZN(
        n20542) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20540), .B1(
        n20635), .B2(n20539), .ZN(n20541) );
  OAI211_X1 U22787 ( .C1(n20623), .C2(n20543), .A(n20542), .B(n20541), .ZN(
        P2_U3160) );
  AOI22_X1 U22788 ( .A1(n20545), .A2(n20635), .B1(n20544), .B2(n11154), .ZN(
        n20548) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20546), .B1(
        n20552), .B2(n20618), .ZN(n20547) );
  OAI211_X1 U22790 ( .C1(n20623), .C2(n20549), .A(n20548), .B(n20547), .ZN(
        P2_U3152) );
  AOI22_X1 U22791 ( .A1(n20551), .A2(n20635), .B1(n20550), .B2(n11154), .ZN(
        n20555) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20553), .B1(
        n20552), .B2(n20634), .ZN(n20554) );
  OAI211_X1 U22793 ( .C1(n20641), .C2(n20561), .A(n20555), .B(n20554), .ZN(
        P2_U3144) );
  AOI22_X1 U22794 ( .A1(n20557), .A2(n20635), .B1(n11154), .B2(n20556), .ZN(
        n20560) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20558), .B1(
        n20563), .B2(n20618), .ZN(n20559) );
  OAI211_X1 U22796 ( .C1(n20623), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P2_U3136) );
  INV_X1 U22797 ( .A(n20635), .ZN(n20573) );
  AOI22_X1 U22798 ( .A1(n20618), .A2(n20569), .B1(n11154), .B2(n20562), .ZN(
        n20566) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20564), .B1(
        n20563), .B2(n20634), .ZN(n20565) );
  OAI211_X1 U22800 ( .C1(n20567), .C2(n20573), .A(n20566), .B(n20565), .ZN(
        P2_U3128) );
  AOI22_X1 U22801 ( .A1(n20618), .A2(n20576), .B1(n11154), .B2(n20568), .ZN(
        n20572) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20570), .B1(
        n20569), .B2(n20634), .ZN(n20571) );
  OAI211_X1 U22803 ( .C1(n20574), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P2_U3120) );
  AOI22_X1 U22804 ( .A1(n20634), .A2(n20576), .B1(n11154), .B2(n20575), .ZN(
        n20580) );
  AOI22_X1 U22805 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20635), .ZN(n20579) );
  OAI211_X1 U22806 ( .C1(n20641), .C2(n20581), .A(n20580), .B(n20579), .ZN(
        P2_U3112) );
  AOI22_X1 U22807 ( .A1(n20583), .A2(n20635), .B1(n20582), .B2(n11154), .ZN(
        n20587) );
  AOI22_X1 U22808 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20585), .B1(
        n20584), .B2(n20634), .ZN(n20586) );
  OAI211_X1 U22809 ( .C1(n20641), .C2(n20594), .A(n20587), .B(n20586), .ZN(
        P2_U3104) );
  AOI22_X1 U22810 ( .A1(n20589), .A2(n20635), .B1(n20588), .B2(n11154), .ZN(
        n20593) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20591), .B1(
        n20590), .B2(n20618), .ZN(n20592) );
  OAI211_X1 U22812 ( .C1(n20623), .C2(n20594), .A(n20593), .B(n20592), .ZN(
        P2_U3096) );
  AOI22_X1 U22813 ( .A1(n20618), .A2(n20602), .B1(n20595), .B2(n11154), .ZN(
        n20599) );
  AOI22_X1 U22814 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20597), .B1(
        n20635), .B2(n20596), .ZN(n20598) );
  OAI211_X1 U22815 ( .C1(n20623), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        P2_U3088) );
  INV_X1 U22816 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n20607) );
  AOI22_X1 U22817 ( .A1(n20634), .A2(n20602), .B1(n20601), .B2(n11154), .ZN(
        n20606) );
  AOI22_X1 U22818 ( .A1(n20635), .A2(n20604), .B1(n20603), .B2(n20618), .ZN(
        n20605) );
  OAI211_X1 U22819 ( .C1(n20608), .C2(n20607), .A(n20606), .B(n20605), .ZN(
        P2_U3080) );
  AOI22_X1 U22820 ( .A1(n20618), .A2(n20610), .B1(n20609), .B2(n11154), .ZN(
        n20614) );
  AOI22_X1 U22821 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20612), .B1(
        n20635), .B2(n20611), .ZN(n20613) );
  OAI211_X1 U22822 ( .C1(n20623), .C2(n20615), .A(n20614), .B(n20613), .ZN(
        P2_U3072) );
  AOI22_X1 U22823 ( .A1(n20617), .A2(n20635), .B1(n11154), .B2(n20616), .ZN(
        n20621) );
  AOI22_X1 U22824 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20619), .B1(
        n20626), .B2(n20618), .ZN(n20620) );
  OAI211_X1 U22825 ( .C1(n20623), .C2(n20622), .A(n20621), .B(n20620), .ZN(
        P2_U3064) );
  AOI22_X1 U22826 ( .A1(n20625), .A2(n20635), .B1(n11154), .B2(n20624), .ZN(
        n20629) );
  AOI22_X1 U22827 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20627), .B1(
        n20626), .B2(n20634), .ZN(n20628) );
  OAI211_X1 U22828 ( .C1(n20641), .C2(n20630), .A(n20629), .B(n20628), .ZN(
        P2_U3056) );
  AOI22_X1 U22829 ( .A1(n20634), .A2(n20633), .B1(n11154), .B2(n20631), .ZN(
        n20639) );
  AOI22_X1 U22830 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20637), .B1(
        n20636), .B2(n20635), .ZN(n20638) );
  OAI211_X1 U22831 ( .C1(n20641), .C2(n20640), .A(n20639), .B(n20638), .ZN(
        P2_U3048) );
  INV_X1 U22832 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20931) );
  INV_X1 U22833 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20642) );
  AOI222_X1 U22834 ( .A1(n20931), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20934), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20642), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20643) );
  OAI22_X1 U22835 ( .A1(n20693), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n20696), .ZN(n20644) );
  INV_X1 U22836 ( .A(n20644), .ZN(U376) );
  OAI22_X1 U22837 ( .A1(n20693), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20696), .ZN(n20645) );
  INV_X1 U22838 ( .A(n20645), .ZN(U365) );
  OAI22_X1 U22839 ( .A1(n20693), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20643), .ZN(n20646) );
  INV_X1 U22840 ( .A(n20646), .ZN(U354) );
  OAI22_X1 U22841 ( .A1(n20693), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20643), .ZN(n20647) );
  INV_X1 U22842 ( .A(n20647), .ZN(U353) );
  OAI22_X1 U22843 ( .A1(n20693), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20643), .ZN(n20648) );
  INV_X1 U22844 ( .A(n20648), .ZN(U352) );
  OAI22_X1 U22845 ( .A1(n20693), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n20643), .ZN(n20649) );
  INV_X1 U22846 ( .A(n20649), .ZN(U351) );
  INV_X2 U22847 ( .A(n20693), .ZN(n20696) );
  OAI22_X1 U22848 ( .A1(n20693), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20696), .ZN(n20650) );
  INV_X1 U22849 ( .A(n20650), .ZN(U350) );
  AOI22_X1 U22850 ( .A1(n20696), .A2(n20652), .B1(n20651), .B2(n20693), .ZN(
        U349) );
  AOI22_X1 U22851 ( .A1(n20696), .A2(n20654), .B1(n20653), .B2(n20693), .ZN(
        U348) );
  OAI22_X1 U22852 ( .A1(n20693), .A2(P3_ADDRESS_REG_9__SCAN_IN), .B1(
        P2_ADDRESS_REG_9__SCAN_IN), .B2(n20696), .ZN(n20655) );
  INV_X1 U22853 ( .A(n20655), .ZN(U347) );
  OAI22_X1 U22854 ( .A1(n20693), .A2(P3_ADDRESS_REG_10__SCAN_IN), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(n20696), .ZN(n20656) );
  INV_X1 U22855 ( .A(n20656), .ZN(U375) );
  AOI22_X1 U22856 ( .A1(n20696), .A2(n20658), .B1(n20657), .B2(n20693), .ZN(
        U374) );
  AOI22_X1 U22857 ( .A1(n20696), .A2(n20660), .B1(n20659), .B2(n20693), .ZN(
        U373) );
  AOI22_X1 U22858 ( .A1(n20696), .A2(n20662), .B1(n20661), .B2(n20693), .ZN(
        U372) );
  AOI22_X1 U22859 ( .A1(n20696), .A2(n20664), .B1(n20663), .B2(n20693), .ZN(
        U371) );
  AOI22_X1 U22860 ( .A1(n20696), .A2(n20666), .B1(n20665), .B2(n20693), .ZN(
        U370) );
  AOI22_X1 U22861 ( .A1(n20696), .A2(n20668), .B1(n20667), .B2(n20693), .ZN(
        U369) );
  AOI22_X1 U22862 ( .A1(n20696), .A2(n20670), .B1(n20669), .B2(n20693), .ZN(
        U368) );
  AOI22_X1 U22863 ( .A1(n20696), .A2(n20672), .B1(n20671), .B2(n20693), .ZN(
        U367) );
  AOI22_X1 U22864 ( .A1(n20696), .A2(n20674), .B1(n20673), .B2(n20693), .ZN(
        U366) );
  AOI22_X1 U22865 ( .A1(n20696), .A2(n20676), .B1(n20675), .B2(n20693), .ZN(
        U364) );
  AOI22_X1 U22866 ( .A1(n20696), .A2(n20678), .B1(n20677), .B2(n20693), .ZN(
        U363) );
  AOI22_X1 U22867 ( .A1(n20696), .A2(n20680), .B1(n20679), .B2(n20693), .ZN(
        U362) );
  AOI22_X1 U22868 ( .A1(n20696), .A2(n20682), .B1(n20681), .B2(n20693), .ZN(
        U361) );
  AOI22_X1 U22869 ( .A1(n20696), .A2(n20684), .B1(n20683), .B2(n20693), .ZN(
        U360) );
  AOI22_X1 U22870 ( .A1(n20696), .A2(n20686), .B1(n20685), .B2(n20693), .ZN(
        U359) );
  AOI22_X1 U22871 ( .A1(n20696), .A2(n20688), .B1(n20687), .B2(n20693), .ZN(
        U358) );
  AOI22_X1 U22872 ( .A1(n20696), .A2(n20690), .B1(n20689), .B2(n20693), .ZN(
        U357) );
  AOI22_X1 U22873 ( .A1(n20696), .A2(n20692), .B1(n20691), .B2(n20693), .ZN(
        U356) );
  AOI22_X1 U22874 ( .A1(n20696), .A2(n20695), .B1(n20694), .B2(n20693), .ZN(
        U355) );
  AOI22_X1 U22875 ( .A1(n22130), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20698) );
  OAI21_X1 U22876 ( .B1(n20699), .B2(n20718), .A(n20698), .ZN(P1_U2936) );
  AOI22_X1 U22877 ( .A1(n20708), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20700) );
  OAI21_X1 U22878 ( .B1(n13512), .B2(n20718), .A(n20700), .ZN(P1_U2935) );
  AOI22_X1 U22879 ( .A1(n20708), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20701) );
  OAI21_X1 U22880 ( .B1(n13505), .B2(n20718), .A(n20701), .ZN(P1_U2934) );
  AOI22_X1 U22881 ( .A1(n20708), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20702) );
  OAI21_X1 U22882 ( .B1(n13534), .B2(n20718), .A(n20702), .ZN(P1_U2933) );
  AOI22_X1 U22883 ( .A1(n20708), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20703) );
  OAI21_X1 U22884 ( .B1(n20704), .B2(n20718), .A(n20703), .ZN(P1_U2932) );
  AOI22_X1 U22885 ( .A1(n20708), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20705) );
  OAI21_X1 U22886 ( .B1(n15656), .B2(n20718), .A(n20705), .ZN(P1_U2931) );
  AOI22_X1 U22887 ( .A1(n20708), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20706) );
  OAI21_X1 U22888 ( .B1(n13562), .B2(n20718), .A(n20706), .ZN(P1_U2930) );
  AOI22_X1 U22889 ( .A1(n22130), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20707) );
  OAI21_X1 U22890 ( .B1(n15676), .B2(n20718), .A(n20707), .ZN(P1_U2929) );
  AOI22_X1 U22891 ( .A1(n20708), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20709) );
  OAI21_X1 U22892 ( .B1(n16297), .B2(n20718), .A(n20709), .ZN(P1_U2928) );
  AOI22_X1 U22893 ( .A1(n22130), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20710) );
  OAI21_X1 U22894 ( .B1(n16339), .B2(n20718), .A(n20710), .ZN(P1_U2927) );
  AOI22_X1 U22895 ( .A1(n22130), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20712) );
  OAI21_X1 U22896 ( .B1(n16361), .B2(n20718), .A(n20712), .ZN(P1_U2926) );
  AOI22_X1 U22897 ( .A1(n22130), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20713) );
  OAI21_X1 U22898 ( .B1(n16792), .B2(n20718), .A(n20713), .ZN(P1_U2925) );
  AOI22_X1 U22899 ( .A1(n22130), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20714) );
  OAI21_X1 U22900 ( .B1(n16788), .B2(n20718), .A(n20714), .ZN(P1_U2924) );
  AOI22_X1 U22901 ( .A1(n22130), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20715) );
  OAI21_X1 U22902 ( .B1(n16784), .B2(n20718), .A(n20715), .ZN(P1_U2923) );
  AOI22_X1 U22903 ( .A1(n22130), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20716) );
  OAI21_X1 U22904 ( .B1(n16780), .B2(n20718), .A(n20716), .ZN(P1_U2922) );
  AOI22_X1 U22905 ( .A1(n22130), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20711), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20717) );
  OAI21_X1 U22906 ( .B1(n20719), .B2(n20718), .A(n20717), .ZN(P1_U2921) );
  OAI222_X1 U22907 ( .A1(n20772), .A2(n20722), .B1(n20721), .B2(n22787), .C1(
        n20724), .C2(n20776), .ZN(P1_U3197) );
  INV_X1 U22908 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20723) );
  OAI222_X1 U22909 ( .A1(n20772), .A2(n20724), .B1(n20723), .B2(n22787), .C1(
        n20726), .C2(n20776), .ZN(P1_U3198) );
  INV_X1 U22910 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20725) );
  INV_X1 U22911 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n22247) );
  OAI222_X1 U22912 ( .A1(n20772), .A2(n20726), .B1(n20725), .B2(n22787), .C1(
        n22247), .C2(n20776), .ZN(P1_U3199) );
  INV_X1 U22913 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20727) );
  OAI222_X1 U22914 ( .A1(n20772), .A2(n22247), .B1(n20727), .B2(n22787), .C1(
        n22273), .C2(n20776), .ZN(P1_U3200) );
  INV_X1 U22915 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20728) );
  INV_X1 U22916 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n22282) );
  OAI222_X1 U22917 ( .A1(n20772), .A2(n22273), .B1(n20728), .B2(n22787), .C1(
        n22282), .C2(n20776), .ZN(P1_U3201) );
  INV_X1 U22918 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20729) );
  OAI222_X1 U22919 ( .A1(n20776), .A2(n22295), .B1(n20729), .B2(n22787), .C1(
        n22282), .C2(n20772), .ZN(P1_U3202) );
  INV_X1 U22920 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20730) );
  OAI222_X1 U22921 ( .A1(n20776), .A2(n20731), .B1(n20730), .B2(n22787), .C1(
        n22295), .C2(n20772), .ZN(P1_U3203) );
  INV_X1 U22922 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20732) );
  OAI222_X1 U22923 ( .A1(n20776), .A2(n20734), .B1(n20732), .B2(n22787), .C1(
        n20731), .C2(n20772), .ZN(P1_U3204) );
  INV_X1 U22924 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20733) );
  OAI222_X1 U22925 ( .A1(n20772), .A2(n20734), .B1(n20733), .B2(n22787), .C1(
        n20735), .C2(n20776), .ZN(P1_U3205) );
  INV_X1 U22926 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20736) );
  OAI222_X1 U22927 ( .A1(n20776), .A2(n22317), .B1(n20736), .B2(n22787), .C1(
        n20735), .C2(n20772), .ZN(P1_U3206) );
  INV_X1 U22928 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20737) );
  OAI222_X1 U22929 ( .A1(n20776), .A2(n16950), .B1(n20737), .B2(n22787), .C1(
        n22317), .C2(n20772), .ZN(P1_U3207) );
  INV_X1 U22930 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20738) );
  OAI222_X1 U22931 ( .A1(n20772), .A2(n16950), .B1(n20738), .B2(n22787), .C1(
        n20740), .C2(n20776), .ZN(P1_U3208) );
  INV_X1 U22932 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20739) );
  OAI222_X1 U22933 ( .A1(n20772), .A2(n20740), .B1(n20739), .B2(n22787), .C1(
        n20742), .C2(n20776), .ZN(P1_U3209) );
  INV_X1 U22934 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U22935 ( .A1(n20772), .A2(n20742), .B1(n20741), .B2(n22787), .C1(
        n20744), .C2(n20776), .ZN(P1_U3210) );
  INV_X1 U22936 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20743) );
  OAI222_X1 U22937 ( .A1(n20772), .A2(n20744), .B1(n20743), .B2(n22787), .C1(
        n20746), .C2(n20776), .ZN(P1_U3211) );
  INV_X1 U22938 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20745) );
  OAI222_X1 U22939 ( .A1(n20772), .A2(n20746), .B1(n20745), .B2(n22787), .C1(
        n20747), .C2(n20776), .ZN(P1_U3212) );
  INV_X1 U22940 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20748) );
  OAI222_X1 U22941 ( .A1(n20776), .A2(n20750), .B1(n20748), .B2(n22787), .C1(
        n20747), .C2(n20772), .ZN(P1_U3213) );
  INV_X1 U22942 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20749) );
  OAI222_X1 U22943 ( .A1(n20772), .A2(n20750), .B1(n20749), .B2(n22787), .C1(
        n20751), .C2(n20776), .ZN(P1_U3214) );
  INV_X1 U22944 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20752) );
  OAI222_X1 U22945 ( .A1(n20776), .A2(n20754), .B1(n20752), .B2(n22787), .C1(
        n20751), .C2(n20772), .ZN(P1_U3215) );
  INV_X1 U22946 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20753) );
  OAI222_X1 U22947 ( .A1(n20772), .A2(n20754), .B1(n20753), .B2(n22787), .C1(
        n22369), .C2(n20776), .ZN(P1_U3216) );
  INV_X1 U22948 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20755) );
  OAI222_X1 U22949 ( .A1(n20776), .A2(n20756), .B1(n20755), .B2(n22787), .C1(
        n22369), .C2(n20772), .ZN(P1_U3217) );
  INV_X1 U22950 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20757) );
  OAI222_X1 U22951 ( .A1(n20776), .A2(n20759), .B1(n20757), .B2(n22787), .C1(
        n20756), .C2(n20772), .ZN(P1_U3218) );
  INV_X1 U22952 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20758) );
  OAI222_X1 U22953 ( .A1(n20772), .A2(n20759), .B1(n20758), .B2(n22787), .C1(
        n20761), .C2(n20776), .ZN(P1_U3219) );
  INV_X1 U22954 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20760) );
  OAI222_X1 U22955 ( .A1(n20772), .A2(n20761), .B1(n20760), .B2(n22787), .C1(
        n20762), .C2(n20776), .ZN(P1_U3220) );
  INV_X1 U22956 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20763) );
  OAI222_X1 U22957 ( .A1(n20776), .A2(n20765), .B1(n20763), .B2(n22787), .C1(
        n20762), .C2(n20772), .ZN(P1_U3221) );
  INV_X1 U22958 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20764) );
  OAI222_X1 U22959 ( .A1(n20772), .A2(n20765), .B1(n20764), .B2(n22787), .C1(
        n20767), .C2(n20776), .ZN(P1_U3222) );
  INV_X1 U22960 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20766) );
  INV_X1 U22961 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20768) );
  OAI222_X1 U22962 ( .A1(n20772), .A2(n20767), .B1(n20766), .B2(n22787), .C1(
        n20768), .C2(n20776), .ZN(P1_U3223) );
  INV_X1 U22963 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20769) );
  OAI222_X1 U22964 ( .A1(n20776), .A2(n20771), .B1(n20769), .B2(n22787), .C1(
        n20768), .C2(n20772), .ZN(P1_U3224) );
  INV_X1 U22965 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20770) );
  INV_X1 U22966 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20773) );
  OAI222_X1 U22967 ( .A1(n20772), .A2(n20771), .B1(n20770), .B2(n22787), .C1(
        n20773), .C2(n20776), .ZN(P1_U3225) );
  INV_X1 U22968 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20774) );
  OAI222_X1 U22969 ( .A1(n20776), .A2(n20775), .B1(n20774), .B2(n22787), .C1(
        n20773), .C2(n20772), .ZN(P1_U3226) );
  OAI22_X1 U22970 ( .A1(n22784), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22787), .ZN(n20777) );
  INV_X1 U22971 ( .A(n20777), .ZN(P1_U3458) );
  NOR4_X1 U22972 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20781) );
  NOR4_X1 U22973 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20780) );
  NOR4_X1 U22974 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20779) );
  NOR4_X1 U22975 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20778) );
  NAND4_X1 U22976 ( .A1(n20781), .A2(n20780), .A3(n20779), .A4(n20778), .ZN(
        n20787) );
  NOR4_X1 U22977 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20785) );
  AOI211_X1 U22978 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20784) );
  NOR4_X1 U22979 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20783) );
  NOR4_X1 U22980 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20782) );
  NAND4_X1 U22981 ( .A1(n20785), .A2(n20784), .A3(n20783), .A4(n20782), .ZN(
        n20786) );
  NOR2_X1 U22982 ( .A1(n20787), .A2(n20786), .ZN(n20804) );
  NOR3_X1 U22983 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20797) );
  NOR2_X1 U22984 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20793) );
  OAI21_X1 U22985 ( .B1(n20797), .B2(n20793), .A(n20804), .ZN(n20788) );
  OAI21_X1 U22986 ( .B1(n20804), .B2(n20789), .A(n20788), .ZN(P1_U2808) );
  OAI22_X1 U22987 ( .A1(n22784), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22787), .ZN(n20790) );
  INV_X1 U22988 ( .A(n20790), .ZN(P1_U3459) );
  NOR3_X1 U22989 ( .A1(n20792), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20791) );
  AOI221_X1 U22990 ( .B1(n20793), .B2(n20792), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20791), .ZN(n20795) );
  INV_X1 U22991 ( .A(n20804), .ZN(n20801) );
  AOI22_X1 U22992 ( .A1(n20804), .A2(n20795), .B1(n20794), .B2(n20801), .ZN(
        P1_U3481) );
  OAI22_X1 U22993 ( .A1(n22784), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22787), .ZN(n20796) );
  INV_X1 U22994 ( .A(n20796), .ZN(P1_U3460) );
  OAI21_X1 U22995 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20797), .A(n20804), .ZN(
        n20798) );
  OAI21_X1 U22996 ( .B1(n20804), .B2(n20799), .A(n20798), .ZN(P1_U2807) );
  OAI22_X1 U22997 ( .A1(n22784), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22787), .ZN(n20800) );
  INV_X1 U22998 ( .A(n20800), .ZN(P1_U3461) );
  NOR2_X1 U22999 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20803) );
  AOI22_X1 U23000 ( .A1(n20804), .A2(n20803), .B1(n20802), .B2(n20801), .ZN(
        P1_U3482) );
  INV_X1 U23001 ( .A(n20805), .ZN(n20827) );
  AOI22_X1 U23002 ( .A1(n20861), .A2(n20827), .B1(n20806), .B2(n20826), .ZN(
        n20807) );
  OAI21_X1 U23003 ( .B1(n20830), .B2(n20808), .A(n20807), .ZN(P1_U2855) );
  INV_X1 U23004 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n22341) );
  INV_X1 U23005 ( .A(n20809), .ZN(n22346) );
  AOI22_X1 U23006 ( .A1(n22346), .A2(n20827), .B1(n20826), .B2(n22345), .ZN(
        n20810) );
  OAI21_X1 U23007 ( .B1(n20830), .B2(n22341), .A(n20810), .ZN(P1_U2857) );
  INV_X1 U23008 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n20813) );
  OAI22_X1 U23009 ( .A1(n22380), .A2(n20805), .B1(n22378), .B2(n20820), .ZN(
        n20811) );
  INV_X1 U23010 ( .A(n20811), .ZN(n20812) );
  OAI21_X1 U23011 ( .B1(n20830), .B2(n20813), .A(n20812), .ZN(P1_U2851) );
  INV_X1 U23012 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U23013 ( .A1(n22361), .A2(n20827), .B1(n22358), .B2(n20826), .ZN(
        n20814) );
  OAI21_X1 U23014 ( .B1(n20830), .B2(n20815), .A(n20814), .ZN(P1_U2853) );
  INV_X1 U23015 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n22289) );
  AND2_X1 U23016 ( .A1(n20817), .A2(n20816), .ZN(n20818) );
  OR2_X1 U23017 ( .A1(n20819), .A2(n20818), .ZN(n22198) );
  NOR2_X1 U23018 ( .A1(n22198), .A2(n20820), .ZN(n20821) );
  AOI21_X1 U23019 ( .B1(n22298), .B2(n20827), .A(n20821), .ZN(n20822) );
  OAI21_X1 U23020 ( .B1(n20830), .B2(n22289), .A(n20822), .ZN(P1_U2865) );
  NAND2_X1 U23021 ( .A1(n15256), .A2(n20823), .ZN(n20824) );
  AND2_X1 U23022 ( .A1(n20825), .A2(n20824), .ZN(n22261) );
  AOI22_X1 U23023 ( .A1(n22271), .A2(n20827), .B1(n20826), .B2(n22261), .ZN(
        n20828) );
  OAI21_X1 U23024 ( .B1(n20830), .B2(n20829), .A(n20828), .ZN(P1_U2867) );
  AOI22_X1 U23025 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22241), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20857), .ZN(n20836) );
  OAI21_X1 U23026 ( .B1(n20833), .B2(n20832), .A(n20831), .ZN(n20834) );
  INV_X1 U23027 ( .A(n20834), .ZN(n22170) );
  AOI22_X1 U23028 ( .A1(n22170), .A2(n20853), .B1(n20860), .B2(n22257), .ZN(
        n20835) );
  OAI211_X1 U23029 ( .C1(n20856), .C2(n22260), .A(n20836), .B(n20835), .ZN(
        P1_U2995) );
  AOI22_X1 U23030 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22241), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20857), .ZN(n20842) );
  OAI21_X1 U23031 ( .B1(n20839), .B2(n20838), .A(n20837), .ZN(n20840) );
  INV_X1 U23032 ( .A(n20840), .ZN(n22193) );
  AOI22_X1 U23033 ( .A1(n22193), .A2(n20853), .B1(n20860), .B2(n22271), .ZN(
        n20841) );
  OAI211_X1 U23034 ( .C1(n20856), .C2(n22264), .A(n20842), .B(n20841), .ZN(
        P1_U2994) );
  AOI22_X1 U23035 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22241), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20857), .ZN(n20848) );
  OAI21_X1 U23036 ( .B1(n20845), .B2(n20844), .A(n20843), .ZN(n20846) );
  INV_X1 U23037 ( .A(n20846), .ZN(n22189) );
  AOI22_X1 U23038 ( .A1(n22189), .A2(n20853), .B1(n20860), .B2(n22284), .ZN(
        n20847) );
  OAI211_X1 U23039 ( .C1(n20856), .C2(n22287), .A(n20848), .B(n20847), .ZN(
        P1_U2993) );
  AOI22_X1 U23040 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22241), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20857), .ZN(n20855) );
  OAI21_X1 U23041 ( .B1(n20851), .B2(n20850), .A(n20849), .ZN(n20852) );
  INV_X1 U23042 ( .A(n20852), .ZN(n22202) );
  AOI22_X1 U23043 ( .A1(n22202), .A2(n20853), .B1(n20860), .B2(n22298), .ZN(
        n20854) );
  OAI211_X1 U23044 ( .C1(n20856), .C2(n22300), .A(n20855), .B(n20854), .ZN(
        P1_U2992) );
  AOI22_X1 U23045 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22241), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20857), .ZN(n20863) );
  AOI22_X1 U23046 ( .A1(n20861), .A2(n20860), .B1(n20859), .B2(n20858), .ZN(
        n20862) );
  OAI211_X1 U23047 ( .C1(n20864), .C2(n22386), .A(n20863), .B(n20862), .ZN(
        P1_U2982) );
  NAND2_X1 U23048 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20865), .ZN(n20868) );
  OAI21_X1 U23049 ( .B1(n20866), .B2(n22406), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20867) );
  OAI21_X1 U23050 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20868), .A(n20867), 
        .ZN(P1_U2803) );
  INV_X1 U23051 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U23052 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n11164), .ZN(n20870) );
  OAI21_X1 U23053 ( .B1(n20871), .B2(n20933), .A(n20870), .ZN(U247) );
  INV_X1 U23054 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U23055 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n11164), .ZN(n20872) );
  OAI21_X1 U23056 ( .B1(n20873), .B2(n20933), .A(n20872), .ZN(U246) );
  INV_X1 U23057 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20875) );
  AOI22_X1 U23058 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n11164), .ZN(n20874) );
  OAI21_X1 U23059 ( .B1(n20875), .B2(n20933), .A(n20874), .ZN(U245) );
  INV_X1 U23060 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20877) );
  AOI22_X1 U23061 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n11164), .ZN(n20876) );
  OAI21_X1 U23062 ( .B1(n20877), .B2(n20933), .A(n20876), .ZN(U244) );
  INV_X1 U23063 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U23064 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n11164), .ZN(n20878) );
  OAI21_X1 U23065 ( .B1(n20879), .B2(n20933), .A(n20878), .ZN(U243) );
  INV_X1 U23066 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U23067 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n11164), .ZN(n20880) );
  OAI21_X1 U23068 ( .B1(n20881), .B2(n20933), .A(n20880), .ZN(U242) );
  AOI22_X1 U23069 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n11164), .ZN(n20882) );
  OAI21_X1 U23070 ( .B1(n20883), .B2(n20933), .A(n20882), .ZN(U241) );
  INV_X1 U23071 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20885) );
  AOI22_X1 U23072 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n11164), .ZN(n20884) );
  OAI21_X1 U23073 ( .B1(n20885), .B2(n20933), .A(n20884), .ZN(U240) );
  INV_X1 U23074 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20887) );
  AOI22_X1 U23075 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n11164), .ZN(n20886) );
  OAI21_X1 U23076 ( .B1(n20887), .B2(n20933), .A(n20886), .ZN(U239) );
  INV_X1 U23077 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U23078 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n11164), .ZN(n20888) );
  OAI21_X1 U23079 ( .B1(n20889), .B2(n20933), .A(n20888), .ZN(U238) );
  AOI22_X1 U23080 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n11164), .ZN(n20890) );
  OAI21_X1 U23081 ( .B1(n14596), .B2(n20933), .A(n20890), .ZN(U237) );
  INV_X1 U23082 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U23083 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n11164), .ZN(n20891) );
  OAI21_X1 U23084 ( .B1(n20892), .B2(n20933), .A(n20891), .ZN(U236) );
  AOI22_X1 U23085 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11164), .ZN(n20893) );
  OAI21_X1 U23086 ( .B1(n20894), .B2(n20933), .A(n20893), .ZN(U235) );
  AOI22_X1 U23087 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n11164), .ZN(n20895) );
  OAI21_X1 U23088 ( .B1(n14614), .B2(n20933), .A(n20895), .ZN(U234) );
  INV_X1 U23089 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20897) );
  AOI22_X1 U23090 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11164), .ZN(n20896) );
  OAI21_X1 U23091 ( .B1(n20897), .B2(n20933), .A(n20896), .ZN(U233) );
  INV_X1 U23092 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20899) );
  AOI22_X1 U23093 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n11164), .ZN(n20898) );
  OAI21_X1 U23094 ( .B1(n20899), .B2(n20933), .A(n20898), .ZN(U232) );
  AOI22_X1 U23095 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11164), .ZN(n20900) );
  OAI21_X1 U23096 ( .B1(n20901), .B2(n20933), .A(n20900), .ZN(U231) );
  AOI22_X1 U23097 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11164), .ZN(n20902) );
  OAI21_X1 U23098 ( .B1(n20903), .B2(n20933), .A(n20902), .ZN(U230) );
  AOI22_X1 U23099 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n11164), .ZN(n20904) );
  OAI21_X1 U23100 ( .B1(n20905), .B2(n20933), .A(n20904), .ZN(U229) );
  AOI22_X1 U23101 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n11164), .ZN(n20906) );
  OAI21_X1 U23102 ( .B1(n20907), .B2(n20933), .A(n20906), .ZN(U228) );
  AOI22_X1 U23103 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n11164), .ZN(n20908) );
  OAI21_X1 U23104 ( .B1(n20909), .B2(n20933), .A(n20908), .ZN(U227) );
  AOI22_X1 U23105 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n11164), .ZN(n20910) );
  OAI21_X1 U23106 ( .B1(n20911), .B2(n20933), .A(n20910), .ZN(U226) );
  AOI22_X1 U23107 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n11164), .ZN(n20912) );
  OAI21_X1 U23108 ( .B1(n20913), .B2(n20933), .A(n20912), .ZN(U225) );
  AOI22_X1 U23109 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n11164), .ZN(n20914) );
  OAI21_X1 U23110 ( .B1(n20915), .B2(n20933), .A(n20914), .ZN(U224) );
  AOI22_X1 U23111 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n11164), .ZN(n20916) );
  OAI21_X1 U23112 ( .B1(n20917), .B2(n20933), .A(n20916), .ZN(U223) );
  AOI22_X1 U23113 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n11164), .ZN(n20918) );
  OAI21_X1 U23114 ( .B1(n20919), .B2(n20933), .A(n20918), .ZN(U222) );
  AOI22_X1 U23115 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n11164), .ZN(n20921) );
  OAI21_X1 U23116 ( .B1(n20922), .B2(n20933), .A(n20921), .ZN(U221) );
  AOI22_X1 U23117 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n11164), .ZN(n20923) );
  OAI21_X1 U23118 ( .B1(n20924), .B2(n20933), .A(n20923), .ZN(U220) );
  AOI22_X1 U23119 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n11164), .ZN(n20925) );
  OAI21_X1 U23120 ( .B1(n20926), .B2(n20933), .A(n20925), .ZN(U219) );
  AOI22_X1 U23121 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n11164), .ZN(n20927) );
  OAI21_X1 U23122 ( .B1(n20928), .B2(n20933), .A(n20927), .ZN(U218) );
  AOI22_X1 U23123 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20920), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n11164), .ZN(n20929) );
  OAI21_X1 U23124 ( .B1(n20930), .B2(n20933), .A(n20929), .ZN(U217) );
  OAI222_X1 U23125 ( .A1(U212), .A2(n20934), .B1(n20933), .B2(n20932), .C1(
        U214), .C2(n20931), .ZN(U216) );
  AOI22_X1 U23126 ( .A1(n22787), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20935), 
        .B2(n22784), .ZN(P1_U3483) );
  OAI21_X1 U23127 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20937), .A(n20936), 
        .ZN(n20938) );
  INV_X1 U23128 ( .A(n20941), .ZN(n22453) );
  AOI211_X1 U23129 ( .C1(n20939), .C2(n20938), .A(n22453), .B(n22091), .ZN(
        n20940) );
  OAI21_X1 U23130 ( .B1(n20940), .B2(n22113), .A(n22102), .ZN(n20946) );
  AND2_X1 U23131 ( .A1(n20941), .A2(n22057), .ZN(n20943) );
  AOI211_X1 U23132 ( .C1(n20944), .C2(n22088), .A(n20943), .B(n20942), .ZN(
        n20945) );
  MUX2_X1 U23133 ( .A(n20946), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20945), 
        .Z(P3_U3296) );
  INV_X1 U23134 ( .A(n20948), .ZN(n20950) );
  AOI22_X1 U23135 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20998), .ZN(n20952) );
  OAI21_X1 U23136 ( .B1(n20953), .B2(n21004), .A(n20952), .ZN(P3_U2768) );
  AOI22_X1 U23137 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20998), .ZN(n20954) );
  OAI21_X1 U23138 ( .B1(n20955), .B2(n21004), .A(n20954), .ZN(P3_U2769) );
  AOI22_X1 U23139 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20998), .ZN(n20956) );
  OAI21_X1 U23140 ( .B1(n20957), .B2(n21004), .A(n20956), .ZN(P3_U2770) );
  AOI22_X1 U23141 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20998), .ZN(n20958) );
  OAI21_X1 U23142 ( .B1(n21503), .B2(n21004), .A(n20958), .ZN(P3_U2771) );
  AOI22_X1 U23143 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20998), .ZN(n20959) );
  OAI21_X1 U23144 ( .B1(n20960), .B2(n21004), .A(n20959), .ZN(P3_U2772) );
  AOI22_X1 U23145 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20998), .ZN(n20961) );
  OAI21_X1 U23146 ( .B1(n21519), .B2(n21004), .A(n20961), .ZN(P3_U2773) );
  AOI22_X1 U23147 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20998), .ZN(n20962) );
  OAI21_X1 U23148 ( .B1(n21520), .B2(n21004), .A(n20962), .ZN(P3_U2774) );
  AOI22_X1 U23149 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20998), .ZN(n20963) );
  OAI21_X1 U23150 ( .B1(n20964), .B2(n21004), .A(n20963), .ZN(P3_U2775) );
  AOI22_X1 U23151 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20998), .ZN(n20965) );
  OAI21_X1 U23152 ( .B1(n20966), .B2(n21004), .A(n20965), .ZN(P3_U2776) );
  AOI22_X1 U23153 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20998), .ZN(n20967) );
  OAI21_X1 U23154 ( .B1(n20968), .B2(n21004), .A(n20967), .ZN(P3_U2777) );
  AOI22_X1 U23155 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20998), .ZN(n20969) );
  OAI21_X1 U23156 ( .B1(n21527), .B2(n21004), .A(n20969), .ZN(P3_U2778) );
  AOI22_X1 U23157 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20998), .ZN(n20970) );
  OAI21_X1 U23158 ( .B1(n20971), .B2(n21004), .A(n20970), .ZN(P3_U2779) );
  AOI22_X1 U23159 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20998), .ZN(n20972) );
  OAI21_X1 U23160 ( .B1(n21548), .B2(n21004), .A(n20972), .ZN(P3_U2780) );
  AOI22_X1 U23161 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20998), .ZN(n20973) );
  OAI21_X1 U23162 ( .B1(n20974), .B2(n21004), .A(n20973), .ZN(P3_U2781) );
  AOI22_X1 U23163 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20990), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20998), .ZN(n20975) );
  OAI21_X1 U23164 ( .B1(n21540), .B2(n21004), .A(n20975), .ZN(P3_U2782) );
  AOI22_X1 U23165 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20998), .ZN(n20976) );
  OAI21_X1 U23166 ( .B1(n21605), .B2(n21004), .A(n20976), .ZN(P3_U2783) );
  AOI22_X1 U23167 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20998), .ZN(n20977) );
  OAI21_X1 U23168 ( .B1(n20978), .B2(n21004), .A(n20977), .ZN(P3_U2784) );
  AOI22_X1 U23169 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20998), .ZN(n20979) );
  OAI21_X1 U23170 ( .B1(n21476), .B2(n21004), .A(n20979), .ZN(P3_U2785) );
  AOI22_X1 U23171 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20998), .ZN(n20980) );
  OAI21_X1 U23172 ( .B1(n20981), .B2(n21004), .A(n20980), .ZN(P3_U2786) );
  AOI22_X1 U23173 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n21001), .ZN(n20982) );
  OAI21_X1 U23174 ( .B1(n21431), .B2(n21004), .A(n20982), .ZN(P3_U2787) );
  AOI22_X1 U23175 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n21001), .ZN(n20983) );
  OAI21_X1 U23176 ( .B1(n21430), .B2(n21004), .A(n20983), .ZN(P3_U2788) );
  AOI22_X1 U23177 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n21001), .ZN(n20984) );
  OAI21_X1 U23178 ( .B1(n21458), .B2(n21004), .A(n20984), .ZN(P3_U2789) );
  AOI22_X1 U23179 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21002), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n21001), .ZN(n20985) );
  OAI21_X1 U23180 ( .B1(n20986), .B2(n21004), .A(n20985), .ZN(P3_U2790) );
  AOI22_X1 U23181 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n21001), .ZN(n20987) );
  OAI21_X1 U23182 ( .B1(n21585), .B2(n21004), .A(n20987), .ZN(P3_U2791) );
  AOI22_X1 U23183 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n21001), .ZN(n20988) );
  OAI21_X1 U23184 ( .B1(n20989), .B2(n21004), .A(n20988), .ZN(P3_U2792) );
  AOI22_X1 U23185 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20990), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n21001), .ZN(n20991) );
  OAI21_X1 U23186 ( .B1(n20992), .B2(n21004), .A(n20991), .ZN(P3_U2793) );
  AOI22_X1 U23187 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21002), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n21001), .ZN(n20993) );
  OAI21_X1 U23188 ( .B1(n21438), .B2(n21004), .A(n20993), .ZN(P3_U2794) );
  AOI22_X1 U23189 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21002), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n21001), .ZN(n20994) );
  OAI21_X1 U23190 ( .B1(n20995), .B2(n21004), .A(n20994), .ZN(P3_U2795) );
  AOI22_X1 U23191 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21002), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n21001), .ZN(n20996) );
  OAI21_X1 U23192 ( .B1(n20997), .B2(n21004), .A(n20996), .ZN(P3_U2796) );
  AOI22_X1 U23193 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21002), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20998), .ZN(n20999) );
  OAI21_X1 U23194 ( .B1(n21000), .B2(n21004), .A(n20999), .ZN(P3_U2797) );
  AOI22_X1 U23195 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n21002), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n21001), .ZN(n21003) );
  OAI21_X1 U23196 ( .B1(n21580), .B2(n21004), .A(n21003), .ZN(P3_U2798) );
  NAND2_X1 U23197 ( .A1(n21005), .A2(n21638), .ZN(n21611) );
  OAI22_X1 U23198 ( .A1(n21385), .A2(n21006), .B1(n21016), .B2(n21306), .ZN(
        n21007) );
  INV_X1 U23199 ( .A(n21007), .ZN(n21014) );
  AOI21_X1 U23200 ( .B1(n21199), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n22096), .ZN(n21169) );
  NAND2_X1 U23201 ( .A1(n21199), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21008) );
  OAI21_X1 U23202 ( .B1(n22096), .B2(n21008), .A(n21375), .ZN(n21011) );
  OAI22_X1 U23203 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n21349), .B1(n21377), 
        .B2(n21009), .ZN(n21010) );
  AOI221_X1 U23204 ( .B1(n21169), .B2(n21012), .C1(n21011), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n21010), .ZN(n21013) );
  OAI211_X1 U23205 ( .C1(n21611), .C2(n21423), .A(n21014), .B(n21013), .ZN(
        P3_U2670) );
  NAND2_X1 U23206 ( .A1(n21391), .A2(n21214), .ZN(n21136) );
  NAND2_X1 U23207 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21638), .ZN(
        n21631) );
  NAND2_X1 U23208 ( .A1(n21015), .A2(n21631), .ZN(n21626) );
  NOR2_X1 U23209 ( .A1(n21017), .A2(n21016), .ZN(n21031) );
  AOI211_X1 U23210 ( .C1(n21017), .C2(n21016), .A(n21031), .B(n21349), .ZN(
        n21020) );
  OAI22_X1 U23211 ( .A1(n21018), .A2(n21375), .B1(n21017), .B2(n21306), .ZN(
        n21019) );
  AOI211_X1 U23212 ( .C1(n21021), .C2(n21626), .A(n21020), .B(n21019), .ZN(
        n21029) );
  INV_X1 U23213 ( .A(n21030), .ZN(n21023) );
  OAI21_X1 U23214 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21022), .A(
        n21199), .ZN(n21039) );
  AOI211_X1 U23215 ( .C1(n21023), .C2(n21200), .A(n22096), .B(n21039), .ZN(
        n21027) );
  AOI211_X1 U23216 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n21025), .A(n21024), .B(
        n21385), .ZN(n21026) );
  AOI211_X1 U23217 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n21420), .A(n21027), .B(
        n21026), .ZN(n21028) );
  OAI211_X1 U23218 ( .C1(n21030), .C2(n21136), .A(n21029), .B(n21028), .ZN(
        P3_U2669) );
  AOI21_X1 U23219 ( .B1(n21339), .B2(n21031), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n21043) );
  AOI21_X1 U23220 ( .B1(n21339), .B2(n21052), .A(n21416), .ZN(n21061) );
  AOI211_X1 U23221 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n21032), .A(n21046), .B(
        n21385), .ZN(n21037) );
  NOR2_X1 U23222 ( .A1(n21033), .A2(n21622), .ZN(n21625) );
  AOI21_X1 U23223 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21625), .A(
        n21656), .ZN(n21644) );
  NOR2_X1 U23224 ( .A1(n21034), .A2(n21644), .ZN(n21635) );
  OAI22_X1 U23225 ( .A1(n21635), .A2(n21423), .B1(n21377), .B2(n21035), .ZN(
        n21036) );
  AOI211_X1 U23226 ( .C1(n21399), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n21037), .B(n21036), .ZN(n21042) );
  AOI21_X1 U23227 ( .B1(n21040), .B2(n21039), .A(n22096), .ZN(n21038) );
  OAI21_X1 U23228 ( .B1(n21040), .B2(n21039), .A(n21038), .ZN(n21041) );
  OAI211_X1 U23229 ( .C1(n21043), .C2(n21061), .A(n21042), .B(n21041), .ZN(
        P3_U2668) );
  AOI21_X1 U23230 ( .B1(n11234), .B2(n21044), .A(n21423), .ZN(n21055) );
  OAI22_X1 U23231 ( .A1(n21377), .A2(n21045), .B1(n21057), .B2(n21375), .ZN(
        n21054) );
  NAND2_X1 U23232 ( .A1(n21339), .A2(n21060), .ZN(n21051) );
  OAI211_X1 U23233 ( .C1(n21046), .C2(n21045), .A(n21419), .B(n21062), .ZN(
        n21050) );
  AOI21_X1 U23234 ( .B1(n21047), .B2(n21415), .A(n21214), .ZN(n21067) );
  NAND3_X1 U23235 ( .A1(n21391), .A2(n21067), .A3(n21048), .ZN(n21049) );
  OAI211_X1 U23236 ( .C1(n21052), .C2(n21051), .A(n21050), .B(n21049), .ZN(
        n21053) );
  NOR4_X1 U23237 ( .A1(n22043), .A2(n21055), .A3(n21054), .A4(n21053), .ZN(
        n21059) );
  OAI211_X1 U23238 ( .C1(n21057), .C2(n21214), .A(n21056), .B(n21169), .ZN(
        n21058) );
  OAI211_X1 U23239 ( .C1(n21061), .C2(n21060), .A(n21059), .B(n21058), .ZN(
        P3_U2667) );
  AOI211_X1 U23240 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n21062), .A(n21081), .B(
        n21385), .ZN(n21063) );
  AOI21_X1 U23241 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n21420), .A(n21063), .ZN(
        n21072) );
  INV_X1 U23242 ( .A(n21064), .ZN(n21073) );
  NOR2_X1 U23243 ( .A1(n21073), .A2(n21349), .ZN(n21068) );
  AOI22_X1 U23244 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n21399), .B1(
        n21065), .B2(n21068), .ZN(n21071) );
  XNOR2_X1 U23245 ( .A(n21067), .B(n21066), .ZN(n21069) );
  OR2_X1 U23246 ( .A1(n21416), .A2(n21068), .ZN(n21090) );
  AOI22_X1 U23247 ( .A1(n21391), .A2(n21069), .B1(P3_REIP_REG_5__SCAN_IN), 
        .B2(n21090), .ZN(n21070) );
  NAND4_X1 U23248 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n18767), .ZN(
        P3_U2666) );
  NOR2_X1 U23249 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n21349), .ZN(n21091) );
  AOI21_X1 U23250 ( .B1(n21073), .B2(n21091), .A(n22043), .ZN(n21085) );
  NOR2_X1 U23251 ( .A1(n21074), .A2(n21200), .ZN(n21092) );
  NAND2_X1 U23252 ( .A1(n21391), .A2(n21199), .ZN(n21116) );
  NOR3_X1 U23253 ( .A1(n21078), .A2(n21092), .A3(n21116), .ZN(n21077) );
  OAI22_X1 U23254 ( .A1(n21377), .A2(n21080), .B1(n21075), .B2(n21375), .ZN(
        n21076) );
  AOI211_X1 U23255 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n21090), .A(n21077), .B(
        n21076), .ZN(n21084) );
  OAI211_X1 U23256 ( .C1(n21079), .C2(n21214), .A(n21078), .B(n21169), .ZN(
        n21083) );
  OAI211_X1 U23257 ( .C1(n21081), .C2(n21080), .A(n21419), .B(n21086), .ZN(
        n21082) );
  NAND4_X1 U23258 ( .A1(n21085), .A2(n21084), .A3(n21083), .A4(n21082), .ZN(
        P3_U2665) );
  AOI22_X1 U23259 ( .A1(n21420), .A2(P3_EBX_REG_7__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n21399), .ZN(n21099) );
  NOR2_X1 U23260 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21349), .ZN(n21088) );
  AOI211_X1 U23261 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n21086), .A(n21111), .B(
        n21385), .ZN(n21087) );
  AOI211_X1 U23262 ( .C1(n21089), .C2(n21088), .A(n22043), .B(n21087), .ZN(
        n21098) );
  OAI21_X1 U23263 ( .B1(n21091), .B2(n21090), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n21097) );
  INV_X1 U23264 ( .A(n21092), .ZN(n21103) );
  NAND2_X1 U23265 ( .A1(n14024), .A2(n21103), .ZN(n21094) );
  AOI21_X1 U23266 ( .B1(n21095), .B2(n21094), .A(n22096), .ZN(n21093) );
  OAI21_X1 U23267 ( .B1(n21095), .B2(n21094), .A(n21093), .ZN(n21096) );
  NAND4_X1 U23268 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        P3_U2664) );
  NOR2_X1 U23269 ( .A1(n21349), .A2(n21125), .ZN(n21100) );
  NOR2_X1 U23270 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n21100), .ZN(n21108) );
  OAI21_X1 U23271 ( .B1(n21349), .B2(n21101), .A(n21306), .ZN(n21102) );
  INV_X1 U23272 ( .A(n21102), .ZN(n21131) );
  OAI21_X1 U23273 ( .B1(n21104), .B2(n21103), .A(n21199), .ZN(n21105) );
  XOR2_X1 U23274 ( .A(n21106), .B(n21105), .Z(n21107) );
  OAI22_X1 U23275 ( .A1(n21108), .A2(n21131), .B1(n22096), .B2(n21107), .ZN(
        n21109) );
  AOI211_X1 U23276 ( .C1(n21420), .C2(P3_EBX_REG_8__SCAN_IN), .A(n22043), .B(
        n21109), .ZN(n21113) );
  OAI211_X1 U23277 ( .C1(n21111), .C2(n21110), .A(n21419), .B(n21117), .ZN(
        n21112) );
  OAI211_X1 U23278 ( .C1(n21375), .C2(n21114), .A(n21113), .B(n21112), .ZN(
        P3_U2663) );
  NOR2_X1 U23279 ( .A1(n21115), .A2(n21200), .ZN(n21134) );
  INV_X1 U23280 ( .A(n21116), .ZN(n21408) );
  NAND2_X1 U23281 ( .A1(n21408), .A2(n21121), .ZN(n21129) );
  AOI211_X1 U23282 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n21117), .A(n21141), .B(
        n21385), .ZN(n21124) );
  AOI22_X1 U23283 ( .A1(n21420), .A2(P3_EBX_REG_9__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n21399), .ZN(n21118) );
  INV_X1 U23284 ( .A(n21118), .ZN(n21123) );
  OAI21_X1 U23285 ( .B1(n21119), .B2(n21214), .A(n21169), .ZN(n21120) );
  OAI22_X1 U23286 ( .A1(n21130), .A2(n21131), .B1(n21121), .B2(n21120), .ZN(
        n21122) );
  NOR4_X1 U23287 ( .A1(n22043), .A2(n21124), .A3(n21123), .A4(n21122), .ZN(
        n21128) );
  NAND2_X1 U23288 ( .A1(n21157), .A2(n21130), .ZN(n21127) );
  OAI211_X1 U23289 ( .C1(n21134), .C2(n21129), .A(n21128), .B(n21127), .ZN(
        P3_U2662) );
  AOI22_X1 U23290 ( .A1(n21420), .A2(P3_EBX_REG_10__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n21399), .ZN(n21144) );
  INV_X1 U23291 ( .A(n21157), .ZN(n21132) );
  NOR2_X1 U23292 ( .A1(n21130), .A2(n21132), .ZN(n21145) );
  OAI21_X1 U23293 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n21132), .A(n21131), .ZN(
        n21139) );
  OAI21_X1 U23294 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21133), .A(
        n21199), .ZN(n21148) );
  OAI21_X1 U23295 ( .B1(n21134), .B2(n21137), .A(n21391), .ZN(n21135) );
  AOI22_X1 U23296 ( .A1(n21137), .A2(n21148), .B1(n21136), .B2(n21135), .ZN(
        n21138) );
  AOI221_X1 U23297 ( .B1(n21145), .B2(n22041), .C1(n21139), .C2(
        P3_REIP_REG_10__SCAN_IN), .A(n21138), .ZN(n21143) );
  OAI211_X1 U23298 ( .C1(n21141), .C2(n21140), .A(n21419), .B(n21146), .ZN(
        n21142) );
  NAND4_X1 U23299 ( .A1(n21144), .A2(n21143), .A3(n18767), .A4(n21142), .ZN(
        P3_U2661) );
  AOI21_X1 U23300 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n21145), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n21156) );
  AOI21_X1 U23301 ( .B1(n21339), .B2(n21185), .A(n21416), .ZN(n21172) );
  AOI211_X1 U23302 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n21146), .A(n21163), .B(
        n21385), .ZN(n21154) );
  OAI21_X1 U23303 ( .B1(n21147), .B2(n21200), .A(n21199), .ZN(n21158) );
  INV_X1 U23304 ( .A(n21158), .ZN(n21160) );
  OAI221_X1 U23305 ( .B1(n21150), .B2(n21160), .C1(n21149), .C2(n21148), .A(
        n21391), .ZN(n21151) );
  OAI211_X1 U23306 ( .C1(n21377), .C2(n21152), .A(n18767), .B(n21151), .ZN(
        n21153) );
  AOI211_X1 U23307 ( .C1(n21399), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21154), .B(n21153), .ZN(n21155) );
  OAI21_X1 U23308 ( .B1(n21156), .B2(n21172), .A(n21155), .ZN(P3_U2660) );
  NAND4_X1 U23309 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_11__SCAN_IN), .A4(n21157), .ZN(n21197) );
  INV_X1 U23310 ( .A(n21161), .ZN(n21159) );
  AOI221_X1 U23311 ( .B1(n21161), .B2(n21160), .C1(n21159), .C2(n21158), .A(
        n22096), .ZN(n21167) );
  OAI211_X1 U23312 ( .C1(n21163), .C2(n21162), .A(n21419), .B(n21173), .ZN(
        n21164) );
  OAI211_X1 U23313 ( .C1(n21165), .C2(n21375), .A(n18767), .B(n21164), .ZN(
        n21166) );
  AOI211_X1 U23314 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n21420), .A(n21167), .B(
        n21166), .ZN(n21168) );
  OAI221_X1 U23315 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n21197), .C1(n21171), 
        .C2(n21172), .A(n21168), .ZN(P3_U2659) );
  OAI21_X1 U23316 ( .B1(n21170), .B2(n21214), .A(n21169), .ZN(n21182) );
  NOR2_X1 U23317 ( .A1(n21171), .A2(n21197), .ZN(n21184) );
  OAI21_X1 U23318 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n21197), .A(n21172), 
        .ZN(n21179) );
  AOI211_X1 U23319 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n21173), .A(n21193), .B(
        n21385), .ZN(n21174) );
  AOI211_X1 U23320 ( .C1(n21420), .C2(P3_EBX_REG_13__SCAN_IN), .A(n22043), .B(
        n21174), .ZN(n21176) );
  OAI211_X1 U23321 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n21186), .A(
        n21408), .B(n21183), .ZN(n21175) );
  OAI211_X1 U23322 ( .C1(n21375), .C2(n21177), .A(n21176), .B(n21175), .ZN(
        n21178) );
  AOI221_X1 U23323 ( .B1(n21184), .B2(n21180), .C1(n21179), .C2(
        P3_REIP_REG_13__SCAN_IN), .A(n21178), .ZN(n21181) );
  OAI21_X1 U23324 ( .B1(n21183), .B2(n21182), .A(n21181), .ZN(P3_U2658) );
  AOI21_X1 U23325 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n21184), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n21190) );
  AOI221_X1 U23326 ( .B1(n21198), .B2(n21339), .C1(n21185), .C2(n21339), .A(
        n21416), .ZN(n21228) );
  OAI21_X1 U23327 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21186), .A(
        n21199), .ZN(n21187) );
  XOR2_X1 U23328 ( .A(n21188), .B(n21187), .Z(n21189) );
  OAI22_X1 U23329 ( .A1(n21190), .A2(n21228), .B1(n22096), .B2(n21189), .ZN(
        n21191) );
  AOI211_X1 U23330 ( .C1(n21420), .C2(P3_EBX_REG_14__SCAN_IN), .A(n22043), .B(
        n21191), .ZN(n21195) );
  OAI211_X1 U23331 ( .C1(n21193), .C2(n21192), .A(n21419), .B(n21205), .ZN(
        n21194) );
  OAI211_X1 U23332 ( .C1(n21375), .C2(n21196), .A(n21195), .B(n21194), .ZN(
        P3_U2657) );
  NOR2_X1 U23333 ( .A1(n21198), .A2(n21197), .ZN(n21224) );
  INV_X1 U23334 ( .A(n21224), .ZN(n21230) );
  INV_X1 U23335 ( .A(n21202), .ZN(n21204) );
  OAI21_X1 U23336 ( .B1(n21201), .B2(n21200), .A(n21199), .ZN(n21213) );
  INV_X1 U23337 ( .A(n21213), .ZN(n21203) );
  AOI221_X1 U23338 ( .B1(n21204), .B2(n21203), .C1(n21202), .C2(n21213), .A(
        n22096), .ZN(n21210) );
  AOI211_X1 U23339 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n21205), .A(n21219), .B(
        n21385), .ZN(n21209) );
  OAI22_X1 U23340 ( .A1(n21377), .A2(n21207), .B1(n21206), .B2(n21375), .ZN(
        n21208) );
  NOR4_X1 U23341 ( .A1(n22043), .A2(n21210), .A3(n21209), .A4(n21208), .ZN(
        n21211) );
  OAI221_X1 U23342 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n21230), .C1(n21212), 
        .C2(n21228), .A(n21211), .ZN(P3_U2656) );
  OAI21_X1 U23343 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n21214), .A(
        n21213), .ZN(n21216) );
  OAI21_X1 U23344 ( .B1(n21217), .B2(n21216), .A(n21391), .ZN(n21215) );
  AOI21_X1 U23345 ( .B1(n21217), .B2(n21216), .A(n21215), .ZN(n21223) );
  OAI211_X1 U23346 ( .C1(n21219), .C2(n21218), .A(n21419), .B(n21232), .ZN(
        n21220) );
  OAI211_X1 U23347 ( .C1(n21221), .C2(n21375), .A(n18767), .B(n21220), .ZN(
        n21222) );
  AOI211_X1 U23348 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n21420), .A(n21223), .B(
        n21222), .ZN(n21226) );
  OAI211_X1 U23349 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n21224), .B(n21231), .ZN(n21225) );
  OAI211_X1 U23350 ( .C1(n21228), .C2(n21227), .A(n21226), .B(n21225), .ZN(
        P3_U2655) );
  NAND2_X1 U23351 ( .A1(n21267), .A2(n21306), .ZN(n21229) );
  NAND2_X1 U23352 ( .A1(n21418), .A2(n21229), .ZN(n21262) );
  AOI211_X1 U23353 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n21232), .A(n21247), .B(
        n21385), .ZN(n21239) );
  OAI211_X1 U23354 ( .C1(n21235), .C2(n21234), .A(n21391), .B(n21233), .ZN(
        n21236) );
  OAI211_X1 U23355 ( .C1(n21377), .C2(n21237), .A(n18767), .B(n21236), .ZN(
        n21238) );
  AOI211_X1 U23356 ( .C1(n21399), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n21239), .B(n21238), .ZN(n21240) );
  OAI221_X1 U23357 ( .B1(n21262), .B2(n21242), .C1(n21262), .C2(n21241), .A(
        n21240), .ZN(P3_U2654) );
  INV_X1 U23358 ( .A(n21279), .ZN(n21253) );
  AOI22_X1 U23359 ( .A1(n21420), .A2(P3_EBX_REG_18__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21399), .ZN(n21250) );
  OAI211_X1 U23360 ( .C1(n21245), .C2(n21244), .A(n21391), .B(n21243), .ZN(
        n21249) );
  OAI211_X1 U23361 ( .C1(n21247), .C2(n21246), .A(n21419), .B(n21254), .ZN(
        n21248) );
  AND4_X1 U23362 ( .A1(n21250), .A2(n18767), .A3(n21249), .A4(n21248), .ZN(
        n21251) );
  OAI221_X1 U23363 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n21253), .C1(n21252), 
        .C2(n21262), .A(n21251), .ZN(P3_U2653) );
  AOI211_X1 U23364 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n21254), .A(n21274), .B(
        n21385), .ZN(n21266) );
  OAI22_X1 U23365 ( .A1(n21377), .A2(n21256), .B1(n21255), .B2(n21375), .ZN(
        n21265) );
  OAI211_X1 U23366 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(P3_REIP_REG_19__SCAN_IN), .A(n21279), .B(n21268), .ZN(n21261) );
  OAI211_X1 U23367 ( .C1(n21259), .C2(n21258), .A(n21391), .B(n21257), .ZN(
        n21260) );
  OAI211_X1 U23368 ( .C1(n21263), .C2(n21262), .A(n21261), .B(n21260), .ZN(
        n21264) );
  OR4_X1 U23369 ( .A1(n22043), .A2(n21266), .A3(n21265), .A4(n21264), .ZN(
        P3_U2652) );
  AOI22_X1 U23370 ( .A1(n21420), .A2(P3_EBX_REG_20__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21399), .ZN(n21278) );
  OAI221_X1 U23371 ( .B1(n21349), .B2(n21280), .C1(n21349), .C2(n21267), .A(
        n21306), .ZN(n21293) );
  NOR2_X1 U23372 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n21268), .ZN(n21269) );
  AOI22_X1 U23373 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n21293), .B1(n21279), 
        .B2(n21269), .ZN(n21277) );
  OAI211_X1 U23374 ( .C1(n21272), .C2(n21271), .A(n21391), .B(n21270), .ZN(
        n21276) );
  OAI211_X1 U23375 ( .C1(n21274), .C2(n21273), .A(n21419), .B(n21281), .ZN(
        n21275) );
  NAND4_X1 U23376 ( .A1(n21278), .A2(n21277), .A3(n21276), .A4(n21275), .ZN(
        P3_U2651) );
  NAND2_X1 U23377 ( .A1(n21280), .A2(n21279), .ZN(n21317) );
  AOI211_X1 U23378 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n21281), .A(n21298), .B(
        n21385), .ZN(n21285) );
  OAI22_X1 U23379 ( .A1(n21377), .A2(n21283), .B1(n21282), .B2(n21375), .ZN(
        n21284) );
  AOI211_X1 U23380 ( .C1(n21293), .C2(P3_REIP_REG_21__SCAN_IN), .A(n21285), 
        .B(n21284), .ZN(n21290) );
  OAI211_X1 U23381 ( .C1(n21288), .C2(n21287), .A(n21391), .B(n21286), .ZN(
        n21289) );
  OAI211_X1 U23382 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n21317), .A(n21290), 
        .B(n21289), .ZN(P3_U2650) );
  AOI22_X1 U23383 ( .A1(n21420), .A2(P3_EBX_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21399), .ZN(n21302) );
  AOI211_X1 U23384 ( .C1(n21291), .C2(n21680), .A(n21304), .B(n21317), .ZN(
        n21292) );
  AOI21_X1 U23385 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n21293), .A(n21292), 
        .ZN(n21301) );
  OAI211_X1 U23386 ( .C1(n21296), .C2(n21295), .A(n21391), .B(n21294), .ZN(
        n21300) );
  OAI211_X1 U23387 ( .C1(n21298), .C2(n21297), .A(n21419), .B(n21307), .ZN(
        n21299) );
  NAND4_X1 U23388 ( .A1(n21302), .A2(n21301), .A3(n21300), .A4(n21299), .ZN(
        P3_U2649) );
  NAND2_X1 U23389 ( .A1(n21304), .A2(n21303), .ZN(n21318) );
  INV_X1 U23390 ( .A(n21305), .ZN(n21320) );
  OAI21_X1 U23391 ( .B1(n21320), .B2(n21349), .A(n21306), .ZN(n21333) );
  AOI211_X1 U23392 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n21307), .A(n21319), .B(
        n21385), .ZN(n21311) );
  OAI22_X1 U23393 ( .A1(n21377), .A2(n21309), .B1(n21308), .B2(n21375), .ZN(
        n21310) );
  AOI211_X1 U23394 ( .C1(n21333), .C2(P3_REIP_REG_23__SCAN_IN), .A(n21311), 
        .B(n21310), .ZN(n21316) );
  OAI211_X1 U23395 ( .C1(n21314), .C2(n21313), .A(n21391), .B(n21312), .ZN(
        n21315) );
  OAI211_X1 U23396 ( .C1(n21318), .C2(n21317), .A(n21316), .B(n21315), .ZN(
        P3_U2648) );
  OAI21_X1 U23397 ( .B1(n21319), .B2(n21326), .A(n21330), .ZN(n21329) );
  NOR2_X1 U23398 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21349), .ZN(n21332) );
  AOI22_X1 U23399 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n21399), .B1(
        n21320), .B2(n21332), .ZN(n21325) );
  OAI211_X1 U23400 ( .C1(n21323), .C2(n21322), .A(n21391), .B(n21321), .ZN(
        n21324) );
  OAI211_X1 U23401 ( .C1(n21326), .C2(n21377), .A(n21325), .B(n21324), .ZN(
        n21327) );
  AOI21_X1 U23402 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21333), .A(n21327), 
        .ZN(n21328) );
  OAI21_X1 U23403 ( .B1(n21385), .B2(n21329), .A(n21328), .ZN(P3_U2647) );
  AOI22_X1 U23404 ( .A1(n21420), .A2(P3_EBX_REG_25__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21399), .ZN(n21343) );
  AOI211_X1 U23405 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n21330), .A(n21345), .B(
        n21385), .ZN(n21331) );
  AOI221_X1 U23406 ( .B1(n21333), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n21332), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n21331), .ZN(n21342) );
  OAI211_X1 U23407 ( .C1(n21336), .C2(n21335), .A(n21391), .B(n21334), .ZN(
        n21341) );
  NAND3_X1 U23408 ( .A1(n21339), .A2(n21338), .A3(n21337), .ZN(n21340) );
  NAND4_X1 U23409 ( .A1(n21343), .A2(n21342), .A3(n21341), .A4(n21340), .ZN(
        P3_U2646) );
  NAND2_X1 U23410 ( .A1(n21418), .A2(n21344), .ZN(n21370) );
  OAI21_X1 U23411 ( .B1(n21346), .B2(n21345), .A(n21419), .ZN(n21347) );
  INV_X1 U23412 ( .A(n21347), .ZN(n21353) );
  NOR3_X1 U23413 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n21349), .A3(n21348), 
        .ZN(n21352) );
  AOI22_X1 U23414 ( .A1(n21420), .A2(P3_EBX_REG_26__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21399), .ZN(n21350) );
  INV_X1 U23415 ( .A(n21350), .ZN(n21351) );
  AOI211_X1 U23416 ( .C1(n21353), .C2(n21360), .A(n21352), .B(n21351), .ZN(
        n21358) );
  OAI211_X1 U23417 ( .C1(n21356), .C2(n21355), .A(n21391), .B(n21354), .ZN(
        n21357) );
  OAI211_X1 U23418 ( .C1(n21370), .C2(n21359), .A(n21358), .B(n21357), .ZN(
        P3_U2645) );
  AOI211_X1 U23419 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n21360), .A(n21371), .B(
        n21385), .ZN(n21363) );
  AOI22_X1 U23420 ( .A1(n21420), .A2(P3_EBX_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21399), .ZN(n21361) );
  INV_X1 U23421 ( .A(n21361), .ZN(n21362) );
  AOI211_X1 U23422 ( .C1(n21364), .C2(n21862), .A(n21363), .B(n21362), .ZN(
        n21369) );
  OAI211_X1 U23423 ( .C1(n21367), .C2(n21366), .A(n21391), .B(n21365), .ZN(
        n21368) );
  OAI211_X1 U23424 ( .C1(n21370), .C2(n21862), .A(n21369), .B(n21368), .ZN(
        P3_U2644) );
  OAI21_X1 U23425 ( .B1(n21371), .B2(n21376), .A(n21387), .ZN(n21386) );
  NOR2_X1 U23426 ( .A1(n21373), .A2(n21372), .ZN(n21379) );
  INV_X1 U23427 ( .A(n21374), .ZN(n21394) );
  OAI22_X1 U23428 ( .A1(n21377), .A2(n21376), .B1(n11349), .B2(n21375), .ZN(
        n21378) );
  AOI221_X1 U23429 ( .B1(n21379), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n21394), 
        .C2(n21940), .A(n21378), .ZN(n21384) );
  OAI211_X1 U23430 ( .C1(n21382), .C2(n21381), .A(n21391), .B(n21380), .ZN(
        n21383) );
  OAI211_X1 U23431 ( .C1(n21386), .C2(n21385), .A(n21384), .B(n21383), .ZN(
        P3_U2643) );
  AOI22_X1 U23432 ( .A1(n21420), .A2(P3_EBX_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21399), .ZN(n21398) );
  NAND2_X1 U23433 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n21387), .ZN(n21388) );
  AOI22_X1 U23434 ( .A1(n21389), .A2(n21388), .B1(P3_REIP_REG_29__SCAN_IN), 
        .B2(n21400), .ZN(n21397) );
  OAI211_X1 U23435 ( .C1(n21393), .C2(n21392), .A(n21391), .B(n21390), .ZN(
        n21396) );
  NAND3_X1 U23436 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n21394), .A3(n21898), 
        .ZN(n21395) );
  NAND4_X1 U23437 ( .A1(n21398), .A2(n21397), .A3(n21396), .A4(n21395), .ZN(
        P3_U2642) );
  AOI22_X1 U23438 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21420), .B1(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21399), .ZN(n21414) );
  INV_X1 U23439 ( .A(n21400), .ZN(n21401) );
  NAND2_X1 U23440 ( .A1(n21402), .A2(n21401), .ZN(n21405) );
  AOI22_X1 U23441 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21405), .B1(n21404), 
        .B2(n21403), .ZN(n21413) );
  NAND3_X1 U23442 ( .A1(n21408), .A2(n21407), .A3(n21406), .ZN(n21412) );
  NAND3_X1 U23443 ( .A1(n21410), .A2(P3_REIP_REG_30__SCAN_IN), .A3(n21409), 
        .ZN(n21411) );
  NAND4_X1 U23444 ( .A1(n21414), .A2(n21413), .A3(n21412), .A4(n21411), .ZN(
        P3_U2640) );
  NOR3_X1 U23445 ( .A1(n21416), .A2(n21652), .A3(n21415), .ZN(n21417) );
  AOI21_X1 U23446 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n21418), .A(n21417), .ZN(
        n21422) );
  OAI21_X1 U23447 ( .B1(n21420), .B2(n21419), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n21421) );
  OAI211_X1 U23448 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n21423), .A(
        n21422), .B(n21421), .ZN(P3_U2671) );
  OAI22_X1 U23449 ( .A1(n21427), .A2(n21426), .B1(n21425), .B2(n21424), .ZN(
        n21428) );
  NAND2_X1 U23450 ( .A1(n22115), .A2(n21428), .ZN(n21592) );
  NAND2_X1 U23451 ( .A1(n21429), .A2(n21604), .ZN(n21601) );
  INV_X1 U23452 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n21436) );
  NAND4_X1 U23453 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n21456) );
  NOR2_X1 U23454 ( .A1(n21431), .A2(n21430), .ZN(n21457) );
  NAND3_X1 U23455 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n21433) );
  NAND3_X1 U23456 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .ZN(n21432) );
  NOR2_X1 U23457 ( .A1(n21521), .A2(n21587), .ZN(n21586) );
  NAND3_X1 U23458 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n21586), .ZN(n21437) );
  NOR2_X1 U23459 ( .A1(n21433), .A2(n21437), .ZN(n21441) );
  AOI21_X1 U23460 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n21588), .A(n21441), .ZN(
        n21435) );
  NAND2_X2 U23461 ( .A1(n21607), .A2(n21604), .ZN(n21544) );
  OAI222_X1 U23462 ( .A1(n21601), .A2(n21436), .B1(n21575), .B2(n21435), .C1(
        n21544), .C2(n21434), .ZN(P3_U2722) );
  INV_X1 U23463 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21442) );
  INV_X1 U23464 ( .A(n21437), .ZN(n21454) );
  NAND2_X1 U23465 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21454), .ZN(n21448) );
  NOR2_X1 U23466 ( .A1(n21438), .A2(n21448), .ZN(n21446) );
  AOI21_X1 U23467 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n21588), .A(n21446), .ZN(
        n21440) );
  OAI222_X1 U23468 ( .A1(n21601), .A2(n21442), .B1(n21441), .B2(n21440), .C1(
        n21544), .C2(n21439), .ZN(P3_U2723) );
  INV_X1 U23469 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21447) );
  INV_X1 U23470 ( .A(n21448), .ZN(n21443) );
  AOI21_X1 U23471 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n21588), .A(n21443), .ZN(
        n21445) );
  OAI222_X1 U23472 ( .A1(n21601), .A2(n21447), .B1(n21446), .B2(n21445), .C1(
        n21544), .C2(n21444), .ZN(P3_U2724) );
  NAND2_X1 U23473 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21593), .ZN(n21450) );
  OAI211_X1 U23474 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n21454), .A(n21588), .B(
        n21448), .ZN(n21449) );
  OAI211_X1 U23475 ( .C1(n21451), .C2(n21544), .A(n21450), .B(n21449), .ZN(
        P3_U2725) );
  INV_X1 U23476 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21455) );
  AOI22_X1 U23477 ( .A1(n21586), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n21588), .ZN(n21453) );
  OAI222_X1 U23478 ( .A1(n21601), .A2(n21455), .B1(n21454), .B2(n21453), .C1(
        n21544), .C2(n21452), .ZN(P3_U2726) );
  NOR2_X1 U23479 ( .A1(n21521), .A2(n21592), .ZN(n21595) );
  NOR2_X1 U23480 ( .A1(n21456), .A2(n21606), .ZN(n21479) );
  NAND2_X1 U23481 ( .A1(n21457), .A2(n21479), .ZN(n21462) );
  NOR2_X1 U23482 ( .A1(n21458), .A2(n21462), .ZN(n21465) );
  AOI21_X1 U23483 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21588), .A(n21465), .ZN(
        n21460) );
  OAI222_X1 U23484 ( .A1(n21601), .A2(n21461), .B1(n21586), .B2(n21460), .C1(
        n21544), .C2(n21459), .ZN(P3_U2728) );
  INV_X1 U23485 ( .A(n21462), .ZN(n21469) );
  AOI21_X1 U23486 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21588), .A(n21469), .ZN(
        n21464) );
  OAI222_X1 U23487 ( .A1(n21466), .A2(n21601), .B1(n21465), .B2(n21464), .C1(
        n21544), .C2(n21463), .ZN(P3_U2729) );
  AOI22_X1 U23488 ( .A1(n21479), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n21588), .ZN(n21468) );
  OAI222_X1 U23489 ( .A1(n21470), .A2(n21601), .B1(n21469), .B2(n21468), .C1(
        n21544), .C2(n21467), .ZN(P3_U2730) );
  NAND2_X1 U23490 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21593), .ZN(n21474) );
  NAND2_X1 U23491 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n21479), .ZN(n21471) );
  OAI211_X1 U23492 ( .C1(n21472), .C2(P3_EAX_REG_4__SCAN_IN), .A(n21588), .B(
        n21471), .ZN(n21473) );
  OAI211_X1 U23493 ( .C1(n21475), .C2(n21544), .A(n21474), .B(n21473), .ZN(
        P3_U2731) );
  NAND2_X1 U23494 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n21594) );
  NOR3_X1 U23495 ( .A1(n21594), .A2(n21476), .A3(n21606), .ZN(n21484) );
  AOI21_X1 U23496 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21588), .A(n21484), .ZN(
        n21478) );
  OAI222_X1 U23497 ( .A1(n21480), .A2(n21601), .B1(n21479), .B2(n21478), .C1(
        n21544), .C2(n21477), .ZN(P3_U2732) );
  NOR2_X1 U23498 ( .A1(n21594), .A2(n21606), .ZN(n21481) );
  AOI21_X1 U23499 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n21588), .A(n21481), .ZN(
        n21483) );
  OAI222_X1 U23500 ( .A1(n21485), .A2(n21601), .B1(n21484), .B2(n21483), .C1(
        n21544), .C2(n21482), .ZN(P3_U2733) );
  NOR2_X2 U23501 ( .A1(n21486), .A2(n21588), .ZN(n21570) );
  NOR2_X2 U23502 ( .A1(n21487), .A2(n21588), .ZN(n21569) );
  AOI22_X1 U23503 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n21569), .ZN(n21490) );
  NAND2_X1 U23504 ( .A1(n21575), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n21581) );
  NOR2_X2 U23505 ( .A1(n21581), .A2(n21580), .ZN(n21579) );
  NOR2_X1 U23506 ( .A1(n21521), .A2(n21571), .ZN(n21514) );
  NAND2_X1 U23507 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21514), .ZN(n21513) );
  NAND2_X1 U23508 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21502), .ZN(n21492) );
  NAND2_X1 U23509 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n21488), .ZN(n21501) );
  OAI211_X1 U23510 ( .C1(n21488), .C2(P3_EAX_REG_21__SCAN_IN), .A(n21588), .B(
        n21501), .ZN(n21489) );
  OAI211_X1 U23511 ( .C1(n21491), .C2(n21544), .A(n21490), .B(n21489), .ZN(
        P3_U2714) );
  AOI22_X1 U23512 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n21569), .ZN(n21494) );
  OAI211_X1 U23513 ( .C1(n21502), .C2(P3_EAX_REG_20__SCAN_IN), .A(n21588), .B(
        n21492), .ZN(n21493) );
  OAI211_X1 U23514 ( .C1(n21495), .C2(n21544), .A(n21494), .B(n21493), .ZN(
        P3_U2715) );
  NAND3_X1 U23515 ( .A1(n21588), .A2(P3_EAX_REG_22__SCAN_IN), .A3(n21501), 
        .ZN(n21500) );
  INV_X1 U23516 ( .A(n21569), .ZN(n21535) );
  OAI22_X1 U23517 ( .A1(n21497), .A2(n21544), .B1(n21496), .B2(n21535), .ZN(
        n21498) );
  AOI21_X1 U23518 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n21570), .A(n21498), .ZN(
        n21499) );
  OAI211_X1 U23519 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n21501), .A(n21500), .B(
        n21499), .ZN(P3_U2713) );
  AOI22_X1 U23520 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21569), .ZN(n21506) );
  AOI211_X1 U23521 ( .C1(n21503), .C2(n21508), .A(n21502), .B(n21546), .ZN(
        n21504) );
  INV_X1 U23522 ( .A(n21504), .ZN(n21505) );
  OAI211_X1 U23523 ( .C1(n21507), .C2(n21544), .A(n21506), .B(n21505), .ZN(
        P3_U2716) );
  AOI22_X1 U23524 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21569), .ZN(n21511) );
  OAI211_X1 U23525 ( .C1(n21509), .C2(P3_EAX_REG_18__SCAN_IN), .A(n21588), .B(
        n21508), .ZN(n21510) );
  OAI211_X1 U23526 ( .C1(n21512), .C2(n21544), .A(n21511), .B(n21510), .ZN(
        P3_U2717) );
  AOI22_X1 U23527 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21569), .ZN(n21516) );
  OAI211_X1 U23528 ( .C1(n21514), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21588), .B(
        n21513), .ZN(n21515) );
  OAI211_X1 U23529 ( .C1(n21517), .C2(n21544), .A(n21516), .B(n21515), .ZN(
        P3_U2718) );
  AOI22_X1 U23530 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21569), .ZN(n21524) );
  NAND4_X1 U23531 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n21518)
         );
  NAND2_X1 U23532 ( .A1(n21565), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21564) );
  NAND2_X1 U23533 ( .A1(n21558), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21559) );
  OAI211_X1 U23534 ( .C1(n21522), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21588), .B(
        n21526), .ZN(n21523) );
  OAI211_X1 U23535 ( .C1(n21525), .C2(n21544), .A(n21524), .B(n21523), .ZN(
        P3_U2710) );
  AOI22_X1 U23536 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n21569), .ZN(n21530) );
  NOR2_X4 U23537 ( .A1(n21526), .A2(n21527), .ZN(n21554) );
  AOI211_X1 U23538 ( .C1(n21527), .C2(n21526), .A(n21554), .B(n21546), .ZN(
        n21528) );
  INV_X1 U23539 ( .A(n21528), .ZN(n21529) );
  OAI211_X1 U23540 ( .C1(n21531), .C2(n21544), .A(n21530), .B(n21529), .ZN(
        P3_U2709) );
  NAND2_X1 U23541 ( .A1(n21547), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n21541) );
  OR2_X1 U23542 ( .A1(n21541), .A2(n21540), .ZN(n21534) );
  NAND2_X1 U23543 ( .A1(n21588), .A2(n21541), .ZN(n21539) );
  OAI21_X1 U23544 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n21606), .A(n21539), .ZN(
        n21532) );
  AOI22_X1 U23545 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21569), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n21532), .ZN(n21533) );
  OAI21_X1 U23546 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n21534), .A(n21533), .ZN(
        P3_U2704) );
  OAI22_X1 U23547 ( .A1(n21536), .A2(n21544), .B1(n12999), .B2(n21535), .ZN(
        n21537) );
  AOI21_X1 U23548 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n21570), .A(n21537), .ZN(
        n21538) );
  OAI221_X1 U23549 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n21541), .C1(n21540), 
        .C2(n21539), .A(n21538), .ZN(P3_U2705) );
  AOI22_X1 U23550 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n21569), .ZN(n21543) );
  OAI211_X1 U23551 ( .C1(n21547), .C2(P3_EAX_REG_29__SCAN_IN), .A(n21588), .B(
        n21541), .ZN(n21542) );
  OAI211_X1 U23552 ( .C1(n21545), .C2(n21544), .A(n21543), .B(n21542), .ZN(
        P3_U2706) );
  AOI22_X1 U23553 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n21569), .ZN(n21551) );
  AOI211_X1 U23554 ( .C1(n21548), .C2(n21553), .A(n21547), .B(n21546), .ZN(
        n21549) );
  INV_X1 U23555 ( .A(n21549), .ZN(n21550) );
  OAI211_X1 U23556 ( .C1(n21552), .C2(n21544), .A(n21551), .B(n21550), .ZN(
        P3_U2707) );
  AOI22_X1 U23557 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n21569), .ZN(n21556) );
  OAI211_X1 U23558 ( .C1(n21554), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21588), .B(
        n21553), .ZN(n21555) );
  OAI211_X1 U23559 ( .C1(n21557), .C2(n21544), .A(n21556), .B(n21555), .ZN(
        P3_U2708) );
  AOI22_X1 U23560 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n21569), .ZN(n21562) );
  CLKBUF_X1 U23561 ( .A(n21558), .Z(n21560) );
  OAI211_X1 U23562 ( .C1(n21560), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21588), .B(
        n21559), .ZN(n21561) );
  OAI211_X1 U23563 ( .C1(n21563), .C2(n21544), .A(n21562), .B(n21561), .ZN(
        P3_U2711) );
  AOI22_X1 U23564 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21569), .ZN(n21567) );
  OAI211_X1 U23565 ( .C1(n21565), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21588), .B(
        n21564), .ZN(n21566) );
  OAI211_X1 U23566 ( .C1(n21568), .C2(n21544), .A(n21567), .B(n21566), .ZN(
        P3_U2712) );
  AOI22_X1 U23567 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21570), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21569), .ZN(n21573) );
  OAI211_X1 U23568 ( .C1(n21579), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21588), .B(
        n21571), .ZN(n21572) );
  OAI211_X1 U23569 ( .C1(n21574), .C2(n21544), .A(n21573), .B(n21572), .ZN(
        P3_U2719) );
  NAND2_X1 U23570 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21593), .ZN(n21577) );
  OAI211_X1 U23571 ( .C1(n21575), .C2(P3_EAX_REG_14__SCAN_IN), .A(n21588), .B(
        n21581), .ZN(n21576) );
  OAI211_X1 U23572 ( .C1(n21578), .C2(n21544), .A(n21577), .B(n21576), .ZN(
        P3_U2721) );
  AOI21_X1 U23573 ( .B1(n21581), .B2(n21580), .A(n21579), .ZN(n21582) );
  AOI22_X1 U23574 ( .A1(n21593), .A2(BUF2_REG_15__SCAN_IN), .B1(n21582), .B2(
        n21588), .ZN(n21583) );
  OAI21_X1 U23575 ( .B1(n21584), .B2(n21544), .A(n21583), .ZN(P3_U2720) );
  AOI22_X1 U23576 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21593), .B1(n21586), .B2(
        n21585), .ZN(n21590) );
  NAND3_X1 U23577 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21588), .A3(n21587), .ZN(
        n21589) );
  OAI211_X1 U23578 ( .C1(n21591), .C2(n21544), .A(n21590), .B(n21589), .ZN(
        P3_U2727) );
  AOI22_X1 U23579 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21593), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n21592), .ZN(n21597) );
  OAI211_X1 U23580 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(P3_EAX_REG_1__SCAN_IN), 
        .A(n21595), .B(n21594), .ZN(n21596) );
  OAI211_X1 U23581 ( .C1(n21598), .C2(n21544), .A(n21597), .B(n21596), .ZN(
        P3_U2734) );
  OAI22_X1 U23582 ( .A1(n21601), .A2(n21600), .B1(n21544), .B2(n21599), .ZN(
        n21602) );
  INV_X1 U23583 ( .A(n21602), .ZN(n21603) );
  OAI221_X1 U23584 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21606), .C1(n21605), 
        .C2(n21604), .A(n21603), .ZN(P3_U2735) );
  INV_X1 U23585 ( .A(n21654), .ZN(n21657) );
  NOR2_X1 U23586 ( .A1(n21607), .A2(n21791), .ZN(n21610) );
  AOI22_X1 U23587 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21884), .B1(
        n21610), .B2(n21609), .ZN(n22071) );
  AOI222_X1 U23588 ( .A1(n21767), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n22071), 
        .B2(n21652), .C1(n21609), .C2(n22105), .ZN(n21608) );
  AOI22_X1 U23589 ( .A1(n21657), .A2(n21609), .B1(n21608), .B2(n21654), .ZN(
        P3_U3290) );
  AOI21_X1 U23590 ( .B1(n21791), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n22022), .ZN(n21615) );
  OAI22_X1 U23591 ( .A1(n21610), .A2(n21611), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21615), .ZN(n22070) );
  INV_X1 U23592 ( .A(n21611), .ZN(n21613) );
  OAI22_X1 U23593 ( .A1(n21694), .A2(n21913), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21627) );
  NOR2_X1 U23594 ( .A1(n21612), .A2(n21767), .ZN(n21629) );
  AOI222_X1 U23595 ( .A1(n22070), .A2(n21652), .B1(n21613), .B2(n22105), .C1(
        n21627), .C2(n21629), .ZN(n21614) );
  AOI22_X1 U23596 ( .A1(n21657), .A2(n21622), .B1(n21614), .B2(n21654), .ZN(
        P3_U3289) );
  NOR2_X1 U23597 ( .A1(n21622), .A2(n21615), .ZN(n21636) );
  AOI21_X1 U23598 ( .B1(n21616), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n21636), .ZN(n21624) );
  OAI22_X1 U23599 ( .A1(n21620), .A2(n21619), .B1(n21618), .B2(n21617), .ZN(
        n21645) );
  AOI211_X1 U23600 ( .C1(n21622), .C2(n21621), .A(n21642), .B(n21645), .ZN(
        n21623) );
  OAI222_X1 U23601 ( .A1(n21626), .A2(n16106), .B1(n21625), .B2(n21624), .C1(
        n21631), .C2(n21623), .ZN(n22067) );
  INV_X1 U23602 ( .A(n21627), .ZN(n21630) );
  AOI222_X1 U23603 ( .A1(n22067), .A2(n21652), .B1(n21630), .B2(n21629), .C1(
        n21628), .C2(n22105), .ZN(n21634) );
  INV_X1 U23604 ( .A(n21631), .ZN(n21632) );
  AOI22_X1 U23605 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21657), .B1(
        n22105), .B2(n21632), .ZN(n21633) );
  OAI21_X1 U23606 ( .B1(n21657), .B2(n21634), .A(n21633), .ZN(P3_U3288) );
  INV_X1 U23607 ( .A(n21635), .ZN(n21653) );
  INV_X1 U23608 ( .A(n21636), .ZN(n21650) );
  NOR2_X1 U23609 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21656), .ZN(
        n21643) );
  AOI211_X1 U23610 ( .C1(n21639), .C2(n21638), .A(n21637), .B(n16106), .ZN(
        n21641) );
  AOI22_X1 U23611 ( .A1(n21643), .A2(n21642), .B1(n21641), .B2(n21640), .ZN(
        n21649) );
  AOI21_X1 U23612 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n21656), .ZN(n21647) );
  AOI22_X1 U23613 ( .A1(n21647), .A2(n21646), .B1(n21645), .B2(n21644), .ZN(
        n21648) );
  OAI211_X1 U23614 ( .C1(n21651), .C2(n21650), .A(n21649), .B(n21648), .ZN(
        n22065) );
  AOI22_X1 U23615 ( .A1(n22105), .A2(n21653), .B1(n21652), .B2(n22065), .ZN(
        n21655) );
  AOI22_X1 U23616 ( .A1(n21657), .A2(n21656), .B1(n21655), .B2(n21654), .ZN(
        P3_U3285) );
  AOI22_X1 U23617 ( .A1(n22117), .A2(n21659), .B1(n21967), .B2(n21658), .ZN(
        n21672) );
  INV_X1 U23618 ( .A(n21660), .ZN(n21762) );
  NAND3_X1 U23619 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21739), .A3(
        n21762), .ZN(n21793) );
  NOR2_X1 U23620 ( .A1(n21661), .A2(n21793), .ZN(n21987) );
  NAND2_X1 U23621 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21987), .ZN(
        n21809) );
  NOR2_X1 U23622 ( .A1(n21662), .A2(n21809), .ZN(n21886) );
  AOI21_X1 U23623 ( .B1(n21987), .B2(n21663), .A(n21884), .ZN(n21664) );
  INV_X1 U23624 ( .A(n21664), .ZN(n21667) );
  NAND3_X1 U23625 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21738), .A3(
        n21762), .ZN(n21768) );
  NAND2_X1 U23626 ( .A1(n21985), .A2(n21665), .ZN(n21988) );
  NOR2_X1 U23627 ( .A1(n21768), .A2(n21988), .ZN(n21993) );
  NAND2_X1 U23628 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21993), .ZN(
        n21867) );
  NAND2_X1 U23629 ( .A1(n21893), .A2(n21867), .ZN(n21666) );
  OAI211_X1 U23630 ( .C1(n21888), .C2(n21886), .A(n21667), .B(n21666), .ZN(
        n21971) );
  AOI21_X1 U23631 ( .B1(n21888), .B2(n16106), .A(n21668), .ZN(n21669) );
  AOI211_X1 U23632 ( .C1(n22022), .C2(n21670), .A(n21971), .B(n21669), .ZN(
        n21671) );
  NAND2_X1 U23633 ( .A1(n21672), .A2(n21671), .ZN(n21826) );
  OAI21_X1 U23634 ( .B1(n22044), .B2(n21826), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21681) );
  NAND2_X1 U23635 ( .A1(n22119), .A2(n21673), .ZN(n21922) );
  NAND2_X1 U23636 ( .A1(n21985), .A2(n21675), .ZN(n21676) );
  AOI22_X1 U23637 ( .A1(n21674), .A2(n22117), .B1(n21967), .B2(n21769), .ZN(
        n21763) );
  INV_X1 U23638 ( .A(n21867), .ZN(n21837) );
  AND2_X1 U23639 ( .A1(n21675), .A2(n21987), .ZN(n21866) );
  AOI22_X1 U23640 ( .A1(n21893), .A2(n21837), .B1(n21699), .B2(n21866), .ZN(
        n21879) );
  OAI21_X1 U23641 ( .B1(n21676), .B2(n21763), .A(n21879), .ZN(n21949) );
  INV_X1 U23642 ( .A(n21949), .ZN(n21825) );
  NOR2_X1 U23643 ( .A1(n21825), .A2(n22044), .ZN(n21980) );
  AOI22_X1 U23644 ( .A1(n22039), .A2(n21678), .B1(n21677), .B2(n21980), .ZN(
        n21679) );
  OAI221_X1 U23645 ( .B1(n22043), .B2(n21681), .C1(n18767), .C2(n21680), .A(
        n21679), .ZN(P3_U2841) );
  NAND2_X1 U23646 ( .A1(n21888), .A2(n16106), .ZN(n21975) );
  AOI221_X1 U23647 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n22022), .C1(
        n21767), .C2(n21975), .A(n21682), .ZN(n21684) );
  AOI22_X1 U23648 ( .A1(n22043), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21941), .ZN(n21683) );
  OAI21_X1 U23649 ( .B1(n21684), .B2(n22044), .A(n21683), .ZN(P3_U2862) );
  NAND2_X1 U23650 ( .A1(n22043), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n21693) );
  INV_X1 U23651 ( .A(n21911), .ZN(n22015) );
  NOR2_X1 U23652 ( .A1(n21685), .A2(n22015), .ZN(n21687) );
  AND2_X1 U23653 ( .A1(n21767), .A2(n21975), .ZN(n21686) );
  MUX2_X1 U23654 ( .A(n21687), .B(n21686), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21691) );
  OAI22_X1 U23655 ( .A1(n21689), .A2(n21930), .B1(n21745), .B2(n21688), .ZN(
        n21690) );
  OAI21_X1 U23656 ( .B1(n21691), .B2(n21690), .A(n22027), .ZN(n21692) );
  OAI211_X1 U23657 ( .C1(n21950), .C2(n21694), .A(n21693), .B(n21692), .ZN(
        P3_U2861) );
  NAND2_X1 U23658 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21696) );
  INV_X1 U23659 ( .A(n21998), .ZN(n21996) );
  OAI21_X1 U23660 ( .B1(n21871), .B2(n21694), .A(n21996), .ZN(n21695) );
  OAI21_X1 U23661 ( .B1(n21696), .B2(n16106), .A(n21695), .ZN(n21697) );
  AOI22_X1 U23662 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21697), .B1(
        n21893), .B2(n21708), .ZN(n21701) );
  NAND3_X1 U23663 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21699), .A3(
        n21698), .ZN(n21700) );
  OAI211_X1 U23664 ( .C1(n21702), .C2(n21745), .A(n21701), .B(n21700), .ZN(
        n21703) );
  AOI22_X1 U23665 ( .A1(n22027), .A2(n21703), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21941), .ZN(n21705) );
  OAI211_X1 U23666 ( .C1(n21706), .C2(n21805), .A(n21705), .B(n21704), .ZN(
        P3_U2860) );
  AOI22_X1 U23667 ( .A1(n21708), .A2(n21893), .B1(n21707), .B2(n21996), .ZN(
        n21709) );
  NAND3_X1 U23668 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21709), .A3(
        n21986), .ZN(n21718) );
  OAI21_X1 U23669 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21710), .A(
        n21718), .ZN(n21711) );
  OAI21_X1 U23670 ( .B1(n21712), .B2(n21745), .A(n21711), .ZN(n21713) );
  AOI22_X1 U23671 ( .A1(n22027), .A2(n21713), .B1(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21941), .ZN(n21715) );
  OAI211_X1 U23672 ( .C1(n21716), .C2(n21805), .A(n21715), .B(n21714), .ZN(
        P3_U2859) );
  NAND2_X1 U23673 ( .A1(n22043), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n21724) );
  INV_X1 U23674 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21717) );
  NOR2_X1 U23675 ( .A1(n21727), .A2(n21717), .ZN(n21720) );
  AND2_X1 U23676 ( .A1(n21911), .A2(n21718), .ZN(n21719) );
  MUX2_X1 U23677 ( .A(n21720), .B(n21719), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n21721) );
  OAI21_X1 U23678 ( .B1(n21722), .B2(n21721), .A(n22027), .ZN(n21723) );
  OAI211_X1 U23679 ( .C1(n21950), .C2(n21725), .A(n21724), .B(n21723), .ZN(
        P3_U2858) );
  INV_X1 U23680 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21736) );
  NAND2_X1 U23681 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21726) );
  NOR2_X1 U23682 ( .A1(n21727), .A2(n21726), .ZN(n21729) );
  MUX2_X1 U23683 ( .A(n21729), .B(n21728), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n21733) );
  OAI22_X1 U23684 ( .A1(n21745), .A2(n21731), .B1(n21930), .B2(n21730), .ZN(
        n21732) );
  OAI21_X1 U23685 ( .B1(n21733), .B2(n21732), .A(n22027), .ZN(n21734) );
  OAI211_X1 U23686 ( .C1(n21950), .C2(n21736), .A(n21735), .B(n21734), .ZN(
        P3_U2857) );
  INV_X1 U23687 ( .A(n21737), .ZN(n21746) );
  NAND2_X1 U23688 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21738), .ZN(
        n21742) );
  NAND2_X1 U23689 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21739), .ZN(
        n21741) );
  OAI22_X1 U23690 ( .A1(n16106), .A2(n21742), .B1(n21740), .B2(n21741), .ZN(
        n21761) );
  AOI22_X1 U23691 ( .A1(n21893), .A2(n21742), .B1(n21996), .B2(n21741), .ZN(
        n21743) );
  NAND3_X1 U23692 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21743), .A3(
        n21986), .ZN(n21751) );
  OAI21_X1 U23693 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21761), .A(
        n21751), .ZN(n21744) );
  OAI21_X1 U23694 ( .B1(n21746), .B2(n21745), .A(n21744), .ZN(n21747) );
  AOI22_X1 U23695 ( .A1(n22027), .A2(n21747), .B1(n21941), .B2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21749) );
  NAND2_X1 U23696 ( .A1(n22043), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n21748) );
  OAI211_X1 U23697 ( .C1(n21750), .C2(n21805), .A(n21749), .B(n21748), .ZN(
        P3_U2855) );
  AOI22_X1 U23698 ( .A1(n22043), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n21941), 
        .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21759) );
  NAND3_X1 U23699 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21911), .A3(
        n21751), .ZN(n21754) );
  NAND3_X1 U23700 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21752), .A3(
        n21761), .ZN(n21753) );
  OAI211_X1 U23701 ( .C1(n21755), .C2(n21928), .A(n21754), .B(n21753), .ZN(
        n21757) );
  AOI22_X1 U23702 ( .A1(n22027), .A2(n21757), .B1(n21853), .B2(n21756), .ZN(
        n21758) );
  OAI211_X1 U23703 ( .C1(n21760), .C2(n22055), .A(n21759), .B(n21758), .ZN(
        P3_U2854) );
  NAND2_X1 U23704 ( .A1(n21762), .A2(n21761), .ZN(n21817) );
  AOI22_X1 U23705 ( .A1(n22043), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n22050), 
        .B2(n21764), .ZN(n21775) );
  NAND2_X1 U23706 ( .A1(n21893), .A2(n21765), .ZN(n21794) );
  NOR2_X1 U23707 ( .A1(n21893), .A2(n21793), .ZN(n21766) );
  AOI22_X1 U23708 ( .A1(n21884), .A2(n21794), .B1(n21771), .B2(n21766), .ZN(
        n21779) );
  NOR2_X1 U23709 ( .A1(n21767), .A2(n21793), .ZN(n21777) );
  INV_X1 U23710 ( .A(n21777), .ZN(n22046) );
  NOR2_X1 U23711 ( .A1(n22117), .A2(n21967), .ZN(n21992) );
  NAND2_X1 U23712 ( .A1(n21893), .A2(n21768), .ZN(n21806) );
  OAI21_X1 U23713 ( .B1(n21769), .B2(n21928), .A(n21806), .ZN(n21770) );
  AOI21_X1 U23714 ( .B1(n22117), .B2(n21990), .A(n21770), .ZN(n22048) );
  OAI211_X1 U23715 ( .C1(n21771), .C2(n21992), .A(n22048), .B(n21950), .ZN(
        n21772) );
  AOI221_X1 U23716 ( .B1(n22049), .B2(n21791), .C1(n22046), .C2(n21791), .A(
        n21772), .ZN(n22034) );
  OAI21_X1 U23717 ( .B1(n21888), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n22034), .ZN(n21773) );
  OAI211_X1 U23718 ( .C1(n21779), .C2(n21773), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18767), .ZN(n21774) );
  OAI211_X1 U23719 ( .C1(n21776), .C2(n22055), .A(n21775), .B(n21774), .ZN(
        P3_U2851) );
  NAND2_X1 U23720 ( .A1(n21778), .A2(n21777), .ZN(n21790) );
  OAI211_X1 U23721 ( .C1(n21884), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n21888), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21783) );
  AOI21_X1 U23722 ( .B1(n22117), .B2(n21780), .A(n21779), .ZN(n21781) );
  OAI211_X1 U23723 ( .C1(n21782), .C2(n21928), .A(n21781), .B(n21806), .ZN(
        n22029) );
  AOI21_X1 U23724 ( .B1(n21790), .B2(n21783), .A(n22029), .ZN(n21789) );
  AOI22_X1 U23725 ( .A1(n22027), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n22050), .B2(n21784), .ZN(n21788) );
  AOI22_X1 U23726 ( .A1(n21941), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n22039), .B2(n21785), .ZN(n21787) );
  OAI211_X1 U23727 ( .C1(n21789), .C2(n21788), .A(n21787), .B(n21786), .ZN(
        P3_U2850) );
  AOI22_X1 U23728 ( .A1(n22043), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n21941), 
        .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21803) );
  AOI22_X1 U23729 ( .A1(n21893), .A2(n22023), .B1(n21791), .B2(n21790), .ZN(
        n22026) );
  AOI22_X1 U23730 ( .A1(n22022), .A2(n21819), .B1(n21792), .B2(n21975), .ZN(
        n21795) );
  NAND2_X1 U23731 ( .A1(n22022), .A2(n21793), .ZN(n22033) );
  AND4_X1 U23732 ( .A1(n21795), .A2(n21806), .A3(n21794), .A4(n22033), .ZN(
        n21799) );
  NOR2_X1 U23733 ( .A1(n21819), .A2(n21817), .ZN(n21796) );
  AOI22_X1 U23734 ( .A1(n21797), .A2(n21967), .B1(n21796), .B2(n21818), .ZN(
        n21798) );
  OAI221_X1 U23735 ( .B1(n21818), .B2(n22026), .C1(n21818), .C2(n21799), .A(
        n21798), .ZN(n21801) );
  AOI22_X1 U23736 ( .A1(n22027), .A2(n21801), .B1(n22039), .B2(n21800), .ZN(
        n21802) );
  OAI211_X1 U23737 ( .C1(n21805), .C2(n21804), .A(n21803), .B(n21802), .ZN(
        P3_U2848) );
  NAND2_X1 U23738 ( .A1(n21888), .A2(n22033), .ZN(n22045) );
  AOI21_X1 U23739 ( .B1(n21807), .B2(n21806), .A(n22035), .ZN(n21808) );
  AOI211_X1 U23740 ( .C1(n21809), .C2(n22045), .A(n21813), .B(n21808), .ZN(
        n22013) );
  NOR2_X1 U23741 ( .A1(n21810), .A2(n21928), .ZN(n21989) );
  OAI21_X1 U23742 ( .B1(n21811), .B2(n21930), .A(n22027), .ZN(n21812) );
  NOR2_X1 U23743 ( .A1(n21989), .A2(n21812), .ZN(n22014) );
  AOI211_X1 U23744 ( .C1(n22013), .C2(n22014), .A(n22043), .B(n21813), .ZN(
        n21814) );
  AOI211_X1 U23745 ( .C1(n21853), .C2(n21816), .A(n21815), .B(n21814), .ZN(
        n21823) );
  NOR4_X1 U23746 ( .A1(n22013), .A2(n21819), .A3(n21818), .A4(n21817), .ZN(
        n21821) );
  OAI221_X1 U23747 ( .B1(n21821), .B2(n21989), .C1(n21821), .C2(n21820), .A(
        n22027), .ZN(n21822) );
  OAI211_X1 U23748 ( .C1(n21824), .C2(n22055), .A(n21823), .B(n21822), .ZN(
        P3_U2847) );
  NOR2_X1 U23749 ( .A1(n21825), .A2(n21835), .ZN(n21855) );
  OAI21_X1 U23750 ( .B1(n22015), .B2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21827) );
  OAI22_X1 U23751 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21855), .B1(
        n21827), .B2(n21826), .ZN(n21832) );
  OAI22_X1 U23752 ( .A1(n21950), .A2(n21836), .B1(n22055), .B2(n21828), .ZN(
        n21829) );
  INV_X1 U23753 ( .A(n21829), .ZN(n21831) );
  OAI211_X1 U23754 ( .C1(n22044), .C2(n21832), .A(n21831), .B(n21830), .ZN(
        P3_U2840) );
  AOI22_X1 U23755 ( .A1(n21853), .A2(n21834), .B1(n22039), .B2(n21833), .ZN(
        n21846) );
  NOR2_X1 U23756 ( .A1(n21836), .A2(n21835), .ZN(n21951) );
  NAND3_X1 U23757 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n21951), .ZN(n21864) );
  NOR3_X1 U23758 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21879), .A3(
        n21864), .ZN(n21842) );
  NAND2_X1 U23759 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21838) );
  OAI221_X1 U23760 ( .B1(n21998), .B2(n21866), .C1(n21998), .C2(n21951), .A(
        n21986), .ZN(n21945) );
  AOI21_X1 U23761 ( .B1(n21837), .B2(n21951), .A(n16106), .ZN(n21948) );
  AOI211_X1 U23762 ( .C1(n21911), .C2(n21838), .A(n21945), .B(n21948), .ZN(
        n21849) );
  OAI22_X1 U23763 ( .A1(n21849), .A2(n21840), .B1(n21928), .B2(n21839), .ZN(
        n21841) );
  OAI21_X1 U23764 ( .B1(n21842), .B2(n21841), .A(n22027), .ZN(n21844) );
  NAND2_X1 U23765 ( .A1(n21941), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21843) );
  NAND4_X1 U23766 ( .A1(n21846), .A2(n21845), .A3(n21844), .A4(n21843), .ZN(
        P3_U2837) );
  INV_X1 U23767 ( .A(n21847), .ZN(n21861) );
  NAND2_X1 U23768 ( .A1(n21967), .A2(n21848), .ZN(n21868) );
  OAI211_X1 U23769 ( .C1(n22015), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n21849), .B(n21868), .ZN(n21851) );
  NOR2_X1 U23770 ( .A1(n21851), .A2(n21850), .ZN(n21854) );
  NAND2_X1 U23771 ( .A1(n21853), .A2(n21852), .ZN(n21872) );
  OAI21_X1 U23772 ( .B1(n21854), .B2(n22044), .A(n21872), .ZN(n21858) );
  NAND2_X1 U23773 ( .A1(n21856), .A2(n21855), .ZN(n21957) );
  NOR2_X1 U23774 ( .A1(n21957), .A2(n21857), .ZN(n21863) );
  AOI222_X1 U23775 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21858), 
        .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21941), .C1(n21858), 
        .C2(n21863), .ZN(n21860) );
  NAND2_X1 U23776 ( .A1(n22043), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21859) );
  OAI211_X1 U23777 ( .C1(n21861), .C2(n22055), .A(n21860), .B(n21859), .ZN(
        P3_U2836) );
  NOR2_X1 U23778 ( .A1(n18767), .A2(n21862), .ZN(n21875) );
  INV_X1 U23779 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21935) );
  NAND2_X1 U23780 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21863), .ZN(
        n21936) );
  OR2_X1 U23781 ( .A1(n21865), .A2(n21864), .ZN(n21880) );
  NOR2_X1 U23782 ( .A1(n21935), .A2(n21880), .ZN(n21887) );
  AND2_X1 U23783 ( .A1(n21866), .A2(n21887), .ZN(n21883) );
  NOR2_X1 U23784 ( .A1(n21996), .A2(n21935), .ZN(n21869) );
  OAI21_X1 U23785 ( .B1(n21867), .B2(n21880), .A(n21893), .ZN(n21885) );
  OAI211_X1 U23786 ( .C1(n21883), .C2(n21869), .A(n21868), .B(n21885), .ZN(
        n21870) );
  OAI21_X1 U23787 ( .B1(n21871), .B2(n21870), .A(n22027), .ZN(n21873) );
  AOI22_X1 U23788 ( .A1(n21935), .A2(n21936), .B1(n21873), .B2(n21872), .ZN(
        n21874) );
  AOI211_X1 U23789 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n21941), .A(
        n21875), .B(n21874), .ZN(n21876) );
  OAI21_X1 U23790 ( .B1(n21877), .B2(n22055), .A(n21876), .ZN(P3_U2835) );
  AOI22_X1 U23791 ( .A1(n21941), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n22039), .B2(n21878), .ZN(n21897) );
  AOI22_X1 U23792 ( .A1(n22117), .A2(n21931), .B1(n21967), .B2(n21929), .ZN(
        n21882) );
  OR3_X1 U23793 ( .A1(n21881), .A2(n21880), .A3(n21879), .ZN(n21907) );
  NAND2_X1 U23794 ( .A1(n21882), .A2(n21907), .ZN(n21903) );
  NOR2_X1 U23795 ( .A1(n21884), .A2(n21883), .ZN(n21890) );
  OAI221_X1 U23796 ( .B1(n21888), .B2(n21887), .C1(n21888), .C2(n21886), .A(
        n21885), .ZN(n21889) );
  NOR2_X1 U23797 ( .A1(n21890), .A2(n21889), .ZN(n21927) );
  OAI22_X1 U23798 ( .A1(n21892), .A2(n21930), .B1(n21891), .B2(n21928), .ZN(
        n21900) );
  AOI21_X1 U23799 ( .B1(n21911), .B2(n21925), .A(n21900), .ZN(n21894) );
  NAND2_X1 U23800 ( .A1(n21893), .A2(n21935), .ZN(n21926) );
  NAND4_X1 U23801 ( .A1(n21927), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n21894), .A4(n21926), .ZN(n21895) );
  OAI211_X1 U23802 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n21903), .A(
        n22027), .B(n21895), .ZN(n21896) );
  OAI211_X1 U23803 ( .C1(n21898), .C2(n18767), .A(n21897), .B(n21896), .ZN(
        P3_U2833) );
  OAI21_X1 U23804 ( .B1(n22015), .B2(n21899), .A(n21927), .ZN(n21909) );
  NOR2_X1 U23805 ( .A1(n21909), .A2(n21900), .ZN(n21901) );
  AOI21_X1 U23806 ( .B1(n21901), .B2(n22027), .A(n21910), .ZN(n21902) );
  AOI22_X1 U23807 ( .A1(n22043), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21902), 
        .B2(n18767), .ZN(n21905) );
  NAND4_X1 U23808 ( .A1(n22027), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n21910), .A4(n21903), .ZN(n21904) );
  OAI211_X1 U23809 ( .C1(n21906), .C2(n22055), .A(n21905), .B(n21904), .ZN(
        P3_U2832) );
  NOR4_X1 U23810 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21910), .A3(
        n21908), .A4(n21907), .ZN(n21916) );
  AOI21_X1 U23811 ( .B1(n21911), .B2(n21910), .A(n21909), .ZN(n21914) );
  OAI22_X1 U23812 ( .A1(n21914), .A2(n21913), .B1(n21930), .B2(n21912), .ZN(
        n21915) );
  AOI211_X1 U23813 ( .C1(n21917), .C2(n21967), .A(n21916), .B(n21915), .ZN(
        n21921) );
  AOI22_X1 U23814 ( .A1(n21941), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n22039), .B2(n21918), .ZN(n21920) );
  OAI211_X1 U23815 ( .C1(n21921), .C2(n22044), .A(n21920), .B(n21919), .ZN(
        P3_U2831) );
  OAI22_X1 U23816 ( .A1(n21931), .A2(n21930), .B1(n21929), .B2(n21928), .ZN(
        n21937) );
  AOI21_X1 U23817 ( .B1(n21942), .B2(n22117), .A(n21941), .ZN(n21943) );
  INV_X1 U23818 ( .A(n21943), .ZN(n21944) );
  AOI211_X1 U23819 ( .C1(n21967), .C2(n21946), .A(n21945), .B(n21944), .ZN(
        n21960) );
  NAND2_X1 U23820 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21960), .ZN(
        n21947) );
  OAI21_X1 U23821 ( .B1(n21948), .B2(n21947), .A(n18767), .ZN(n21958) );
  NAND3_X1 U23822 ( .A1(n21951), .A2(n21950), .A3(n21949), .ZN(n21955) );
  AOI21_X1 U23823 ( .B1(n21953), .B2(n22039), .A(n21952), .ZN(n21954) );
  OAI221_X1 U23824 ( .B1(n21958), .B2(n21956), .C1(n21958), .C2(n21955), .A(
        n21954), .ZN(P3_U2839) );
  NOR3_X1 U23825 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n22044), .A3(
        n21957), .ZN(n21962) );
  AOI211_X1 U23826 ( .C1(n22015), .C2(n21960), .A(n21959), .B(n21958), .ZN(
        n21961) );
  AOI211_X1 U23827 ( .C1(n22039), .C2(n21963), .A(n21962), .B(n21961), .ZN(
        n21964) );
  OAI21_X1 U23828 ( .B1(n18767), .B2(n21965), .A(n21964), .ZN(P3_U2838) );
  AOI22_X1 U23829 ( .A1(n22117), .A2(n21968), .B1(n21967), .B2(n21966), .ZN(
        n21969) );
  NAND2_X1 U23830 ( .A1(n22027), .A2(n21969), .ZN(n21970) );
  OAI21_X1 U23831 ( .B1(n21971), .B2(n21970), .A(n18767), .ZN(n21977) );
  AOI22_X1 U23832 ( .A1(n22039), .A2(n21972), .B1(n21980), .B2(n21976), .ZN(
        n21974) );
  OAI211_X1 U23833 ( .C1(n21976), .C2(n21977), .A(n21974), .B(n21973), .ZN(
        P3_U2843) );
  NAND3_X1 U23834 ( .A1(n21976), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n21975), 
        .ZN(n21978) );
  NAND2_X1 U23835 ( .A1(n21978), .A2(n21977), .ZN(n21981) );
  AOI22_X1 U23836 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21981), .B1(
        n21980), .B2(n21979), .ZN(n21983) );
  OAI211_X1 U23837 ( .C1(n21984), .C2(n22055), .A(n21983), .B(n21982), .ZN(
        P3_U2842) );
  NAND2_X1 U23838 ( .A1(n21985), .A2(n22050), .ZN(n22020) );
  NAND3_X1 U23839 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21987), .A3(
        n21986), .ZN(n21995) );
  NOR3_X1 U23840 ( .A1(n21990), .A2(n21989), .A3(n21988), .ZN(n21991) );
  OAI22_X1 U23841 ( .A1(n21993), .A2(n16106), .B1(n21992), .B2(n21991), .ZN(
        n21994) );
  AOI211_X1 U23842 ( .C1(n21996), .C2(n21995), .A(n22044), .B(n21994), .ZN(
        n22005) );
  AOI221_X1 U23843 ( .B1(n21998), .B2(n22005), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n22005), .A(n21997), .ZN(
        n21999) );
  AOI22_X1 U23844 ( .A1(n22000), .A2(n22039), .B1(n21999), .B2(n18767), .ZN(
        n22002) );
  NAND2_X1 U23845 ( .A1(n22043), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n22001) );
  OAI211_X1 U23846 ( .C1(n22003), .C2(n22020), .A(n22002), .B(n22001), .ZN(
        P3_U2844) );
  INV_X1 U23847 ( .A(n22020), .ZN(n22008) );
  NOR3_X1 U23848 ( .A1(n22043), .A2(n22005), .A3(n22004), .ZN(n22006) );
  AOI211_X1 U23849 ( .C1(n22009), .C2(n22008), .A(n22007), .B(n22006), .ZN(
        n22010) );
  OAI21_X1 U23850 ( .B1(n22011), .B2(n22055), .A(n22010), .ZN(P3_U2845) );
  AOI221_X1 U23851 ( .B1(n22015), .B2(n22014), .C1(n22013), .C2(n22014), .A(
        n22012), .ZN(n22016) );
  AOI22_X1 U23852 ( .A1(n22017), .A2(n22039), .B1(n22016), .B2(n18767), .ZN(
        n22019) );
  OAI211_X1 U23853 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n22020), .A(
        n22019), .B(n22018), .ZN(P3_U2846) );
  AOI22_X1 U23854 ( .A1(n22043), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n22050), 
        .B2(n22021), .ZN(n22031) );
  OAI21_X1 U23855 ( .B1(n22024), .B2(n22023), .A(n22022), .ZN(n22025) );
  NAND3_X1 U23856 ( .A1(n22027), .A2(n22026), .A3(n22025), .ZN(n22028) );
  OAI211_X1 U23857 ( .C1(n22029), .C2(n22028), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18767), .ZN(n22030) );
  OAI211_X1 U23858 ( .C1(n22032), .C2(n22055), .A(n22031), .B(n22030), .ZN(
        P3_U2849) );
  OAI211_X1 U23859 ( .C1(n22035), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n22034), .B(n22033), .ZN(n22036) );
  NAND2_X1 U23860 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n22036), .ZN(
        n22042) );
  NOR2_X1 U23861 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n22049), .ZN(
        n22037) );
  AOI22_X1 U23862 ( .A1(n22039), .A2(n22038), .B1(n22050), .B2(n22037), .ZN(
        n22040) );
  OAI221_X1 U23863 ( .B1(n22043), .B2(n22042), .C1(n18767), .C2(n22041), .A(
        n22040), .ZN(P3_U2852) );
  AOI21_X1 U23864 ( .B1(n22046), .B2(n22045), .A(n22044), .ZN(n22047) );
  AOI21_X1 U23865 ( .B1(n22048), .B2(n22047), .A(n22043), .ZN(n22051) );
  AOI22_X1 U23866 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n22051), .B1(
        n22050), .B2(n22049), .ZN(n22054) );
  INV_X1 U23867 ( .A(n22052), .ZN(n22053) );
  OAI211_X1 U23868 ( .C1(n22056), .C2(n22055), .A(n22054), .B(n22053), .ZN(
        P3_U2853) );
  NAND2_X1 U23869 ( .A1(n22453), .A2(n22057), .ZN(n22103) );
  INV_X1 U23870 ( .A(n22058), .ZN(n22095) );
  NOR2_X1 U23871 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .ZN(
        n22087) );
  NAND3_X1 U23872 ( .A1(n22063), .A2(n22060), .A3(n22059), .ZN(n22114) );
  OAI22_X1 U23873 ( .A1(n22063), .A2(n22062), .B1(n22061), .B2(n16106), .ZN(
        n22120) );
  AOI211_X1 U23874 ( .C1(n22074), .C2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n22064), .B(n22120), .ZN(n22086) );
  INV_X1 U23875 ( .A(n22074), .ZN(n22066) );
  AOI22_X1 U23876 ( .A1(n22074), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n22065), .B2(n22066), .ZN(n22083) );
  MUX2_X1 U23877 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n22067), .S(
        n22066), .Z(n22078) );
  AOI222_X1 U23878 ( .A1(n22071), .A2(n22070), .B1(n22071), .B2(n22069), .C1(
        n22070), .C2(n22068), .ZN(n22073) );
  OAI21_X1 U23879 ( .B1(n22074), .B2(n22073), .A(n22072), .ZN(n22077) );
  AND2_X1 U23880 ( .A1(n22078), .A2(n22077), .ZN(n22075) );
  OAI221_X1 U23881 ( .B1(n22078), .B2(n22077), .C1(n22076), .C2(n22075), .A(
        n22080), .ZN(n22082) );
  AOI21_X1 U23882 ( .B1(n22080), .B2(n22079), .A(n22078), .ZN(n22081) );
  AOI222_X1 U23883 ( .A1(n22083), .A2(n22082), .B1(n22083), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n22082), .C2(n22081), .ZN(
        n22084) );
  NOR3_X1 U23884 ( .A1(n22119), .A2(n22117), .A3(n22084), .ZN(n22085) );
  OAI211_X1 U23885 ( .C1(n22087), .C2(n22114), .A(n22086), .B(n22085), .ZN(
        n22109) );
  AOI211_X1 U23886 ( .C1(n22090), .C2(n22089), .A(n22088), .B(n22109), .ZN(
        n22097) );
  AOI21_X1 U23887 ( .B1(n22453), .B2(n22091), .A(n22097), .ZN(n22112) );
  NAND3_X1 U23888 ( .A1(n22093), .A2(n22112), .A3(n22092), .ZN(n22094) );
  NAND4_X1 U23889 ( .A1(n22096), .A2(n22103), .A3(n22095), .A4(n22094), .ZN(
        P3_U2997) );
  NOR2_X1 U23890 ( .A1(n22097), .A2(n22113), .ZN(n22101) );
  INV_X1 U23891 ( .A(n22098), .ZN(n22099) );
  OAI21_X1 U23892 ( .B1(n22101), .B2(n22100), .A(n22099), .ZN(P3_U3282) );
  INV_X1 U23893 ( .A(n22102), .ZN(n22106) );
  INV_X1 U23894 ( .A(n22103), .ZN(n22104) );
  AOI211_X1 U23895 ( .C1(n22106), .C2(n22105), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n22104), .ZN(n22107) );
  AOI211_X1 U23896 ( .C1(n22115), .C2(n22109), .A(n22108), .B(n22107), .ZN(
        n22110) );
  OAI221_X1 U23897 ( .B1(n22113), .B2(n22112), .C1(n22113), .C2(n22111), .A(
        n22110), .ZN(P3_U2996) );
  INV_X1 U23898 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n22123) );
  NAND2_X1 U23899 ( .A1(n22115), .A2(n22114), .ZN(n22125) );
  AOI22_X1 U23900 ( .A1(n22119), .A2(n22118), .B1(n22117), .B2(n22116), .ZN(
        n22122) );
  NOR2_X1 U23901 ( .A1(n22125), .A2(n22120), .ZN(n22121) );
  AOI22_X1 U23902 ( .A1(n22123), .A2(n22125), .B1(n22122), .B2(n22121), .ZN(
        P3_U3295) );
  AOI21_X1 U23903 ( .B1(n22125), .B2(P3_FLUSH_REG_SCAN_IN), .A(n22124), .ZN(
        n22126) );
  INV_X1 U23904 ( .A(n22126), .ZN(P3_U2637) );
  AOI211_X1 U23905 ( .C1(n22130), .C2(n22129), .A(n22128), .B(n22127), .ZN(
        n22136) );
  OAI211_X1 U23906 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n22132), .A(n22131), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n22133) );
  AOI21_X1 U23907 ( .B1(n22133), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n22401), 
        .ZN(n22135) );
  NAND2_X1 U23908 ( .A1(n22136), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n22134) );
  OAI21_X1 U23909 ( .B1(n22136), .B2(n22135), .A(n22134), .ZN(P1_U3485) );
  NOR4_X1 U23910 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n22139), .A3(
        n22138), .A4(n22137), .ZN(n22140) );
  AOI21_X1 U23911 ( .B1(n22241), .B2(P1_REIP_REG_14__SCAN_IN), .A(n22140), 
        .ZN(n22145) );
  INV_X1 U23912 ( .A(n22141), .ZN(n22142) );
  AOI22_X1 U23913 ( .A1(n22143), .A2(n22239), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n22142), .ZN(n22144) );
  OAI211_X1 U23914 ( .C1(n22245), .C2(n22146), .A(n22145), .B(n22144), .ZN(
        P1_U3017) );
  NAND2_X1 U23915 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n22160), .ZN(
        n22159) );
  NOR3_X1 U23916 ( .A1(n14389), .A2(n22148), .A3(n22151), .ZN(n22147) );
  AOI211_X1 U23917 ( .C1(n22148), .C2(n22166), .A(n22147), .B(n22163), .ZN(
        n22157) );
  AND3_X1 U23918 ( .A1(n22150), .A2(n22149), .A3(n22239), .ZN(n22155) );
  NOR2_X1 U23919 ( .A1(n22151), .A2(n22162), .ZN(n22164) );
  NOR2_X1 U23920 ( .A1(n22245), .A2(n22152), .ZN(n22153) );
  NOR4_X1 U23921 ( .A1(n22155), .A2(n22164), .A3(n22154), .A4(n22153), .ZN(
        n22156) );
  OAI221_X1 U23922 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n22159), .C1(
        n22158), .C2(n22157), .A(n22156), .ZN(P1_U3029) );
  AOI22_X1 U23923 ( .A1(n22225), .A2(n22162), .B1(n22161), .B2(n22160), .ZN(
        n22206) );
  NOR3_X1 U23924 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n22206), .A3(
        n22179), .ZN(n22169) );
  AOI211_X1 U23925 ( .C1(n22166), .C2(n22165), .A(n22164), .B(n22163), .ZN(
        n22180) );
  OR2_X1 U23926 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n22206), .ZN(
        n22177) );
  AOI21_X1 U23927 ( .B1(n22180), .B2(n22177), .A(n22167), .ZN(n22168) );
  AOI211_X1 U23928 ( .C1(n22170), .C2(n22239), .A(n22169), .B(n22168), .ZN(
        n22172) );
  NAND2_X1 U23929 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22241), .ZN(n22171) );
  OAI211_X1 U23930 ( .C1(n22245), .C2(n22246), .A(n22172), .B(n22171), .ZN(
        P1_U3027) );
  NOR2_X1 U23931 ( .A1(n22173), .A2(n22226), .ZN(n22174) );
  AOI211_X1 U23932 ( .C1(n22231), .C2(n22176), .A(n22175), .B(n22174), .ZN(
        n22178) );
  OAI211_X1 U23933 ( .C1(n22180), .C2(n22179), .A(n22178), .B(n22177), .ZN(
        P1_U3028) );
  NAND2_X1 U23934 ( .A1(n22181), .A2(n22204), .ZN(n22187) );
  OAI21_X1 U23935 ( .B1(n22221), .B2(n22183), .A(n22182), .ZN(n22222) );
  INV_X1 U23936 ( .A(n22222), .ZN(n22201) );
  OAI21_X1 U23937 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n22184), .A(
        n22201), .ZN(n22185) );
  AOI21_X1 U23938 ( .B1(n22225), .B2(n22186), .A(n22185), .ZN(n22197) );
  OAI22_X1 U23939 ( .A1(n22206), .A2(n22187), .B1(n22197), .B2(n22204), .ZN(
        n22188) );
  AOI21_X1 U23940 ( .B1(n22189), .B2(n22239), .A(n22188), .ZN(n22191) );
  NAND2_X1 U23941 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22241), .ZN(n22190) );
  OAI211_X1 U23942 ( .C1(n22245), .C2(n22276), .A(n22191), .B(n22190), .ZN(
        P1_U3025) );
  OAI21_X1 U23943 ( .B1(n22203), .B2(n22206), .A(n22205), .ZN(n22192) );
  INV_X1 U23944 ( .A(n22192), .ZN(n22196) );
  AOI22_X1 U23945 ( .A1(n22193), .A2(n22239), .B1(n22231), .B2(n22261), .ZN(
        n22195) );
  NAND2_X1 U23946 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22241), .ZN(n22194) );
  OAI211_X1 U23947 ( .C1(n22197), .C2(n22196), .A(n22195), .B(n22194), .ZN(
        P1_U3026) );
  INV_X1 U23948 ( .A(n22198), .ZN(n22293) );
  AOI22_X1 U23949 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22241), .B1(n22231), 
        .B2(n22293), .ZN(n22209) );
  AOI21_X1 U23950 ( .B1(n22201), .B2(n22200), .A(n22199), .ZN(n22210) );
  AOI22_X1 U23951 ( .A1(n22202), .A2(n22239), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n22210), .ZN(n22208) );
  NOR4_X1 U23952 ( .A1(n22206), .A2(n22205), .A3(n22204), .A4(n22203), .ZN(
        n22218) );
  NAND2_X1 U23953 ( .A1(n22218), .A2(n22211), .ZN(n22207) );
  NAND3_X1 U23954 ( .A1(n22209), .A2(n22208), .A3(n22207), .ZN(P1_U3024) );
  NAND2_X1 U23955 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n22218), .ZN(
        n22217) );
  AOI21_X1 U23956 ( .B1(n22218), .B2(n22211), .A(n22210), .ZN(n22215) );
  INV_X1 U23957 ( .A(n22212), .ZN(n22213) );
  AOI222_X1 U23958 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22241), .B1(n22231), 
        .B2(n22302), .C1(n22239), .C2(n22213), .ZN(n22214) );
  OAI221_X1 U23959 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n22217), .C1(
        n22216), .C2(n22215), .A(n22214), .ZN(P1_U3023) );
  NAND2_X1 U23960 ( .A1(n22219), .A2(n22218), .ZN(n22237) );
  INV_X1 U23961 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n22233) );
  NOR2_X1 U23962 ( .A1(n22221), .A2(n22220), .ZN(n22223) );
  AOI211_X1 U23963 ( .C1(n22225), .C2(n22224), .A(n22223), .B(n22222), .ZN(
        n22234) );
  NOR2_X1 U23964 ( .A1(n22227), .A2(n22226), .ZN(n22228) );
  AOI211_X1 U23965 ( .C1(n22231), .C2(n22230), .A(n22229), .B(n22228), .ZN(
        n22232) );
  OAI221_X1 U23966 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n22237), .C1(
        n22233), .C2(n22234), .A(n22232), .ZN(P1_U3022) );
  XOR2_X1 U23967 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n22233), .Z(
        n22236) );
  OAI22_X1 U23968 ( .A1(n22237), .A2(n22236), .B1(n22235), .B2(n22234), .ZN(
        n22238) );
  AOI21_X1 U23969 ( .B1(n22240), .B2(n22239), .A(n22238), .ZN(n22243) );
  NAND2_X1 U23970 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n22241), .ZN(n22242) );
  OAI211_X1 U23971 ( .C1(n22245), .C2(n22244), .A(n22243), .B(n22242), .ZN(
        P1_U3021) );
  AND2_X1 U23972 ( .A1(n22262), .A2(n22333), .ZN(n22249) );
  OAI21_X1 U23973 ( .B1(n22279), .B2(n22262), .A(n22339), .ZN(n22274) );
  OAI22_X1 U23974 ( .A1(n22274), .A2(n22247), .B1(n22377), .B2(n22246), .ZN(
        n22248) );
  AOI21_X1 U23975 ( .B1(n22250), .B2(n22249), .A(n22248), .ZN(n22259) );
  INV_X1 U23976 ( .A(n22251), .ZN(n22255) );
  AOI21_X1 U23977 ( .B1(n22355), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22353), .ZN(n22253) );
  NAND2_X1 U23978 ( .A1(n22376), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n22252) );
  OAI211_X1 U23979 ( .C1(n22255), .C2(n22254), .A(n22253), .B(n22252), .ZN(
        n22256) );
  AOI21_X1 U23980 ( .B1(n22257), .B2(n22270), .A(n22256), .ZN(n22258) );
  OAI211_X1 U23981 ( .C1(n22260), .C2(n22384), .A(n22259), .B(n22258), .ZN(
        P1_U2836) );
  INV_X1 U23982 ( .A(n22261), .ZN(n22268) );
  NOR3_X1 U23983 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22373), .A3(n22262), .ZN(
        n22263) );
  AOI211_X1 U23984 ( .C1(n22355), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n22353), .B(n22263), .ZN(n22267) );
  INV_X1 U23985 ( .A(n22264), .ZN(n22265) );
  AOI22_X1 U23986 ( .A1(n22265), .A2(n22357), .B1(n22376), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n22266) );
  OAI211_X1 U23987 ( .C1(n22377), .C2(n22268), .A(n22267), .B(n22266), .ZN(
        n22269) );
  AOI21_X1 U23988 ( .B1(n22271), .B2(n22270), .A(n22269), .ZN(n22272) );
  OAI21_X1 U23989 ( .B1(n22274), .B2(n22273), .A(n22272), .ZN(P1_U2835) );
  OAI22_X1 U23990 ( .A1(n22377), .A2(n22276), .B1(n22342), .B2(n22275), .ZN(
        n22277) );
  AOI211_X1 U23991 ( .C1(n22355), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n22353), .B(n22277), .ZN(n22286) );
  NAND2_X1 U23992 ( .A1(n22333), .A2(n22278), .ZN(n22281) );
  AOI21_X1 U23993 ( .B1(n22333), .B2(n22280), .A(n22279), .ZN(n22296) );
  AOI21_X1 U23994 ( .B1(n22282), .B2(n22281), .A(n22296), .ZN(n22283) );
  AOI21_X1 U23995 ( .B1(n22284), .B2(n22360), .A(n22283), .ZN(n22285) );
  OAI211_X1 U23996 ( .C1(n22287), .C2(n22384), .A(n22286), .B(n22285), .ZN(
        P1_U2834) );
  AOI21_X1 U23997 ( .B1(n22355), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22353), .ZN(n22288) );
  OAI21_X1 U23998 ( .B1(n22342), .B2(n22289), .A(n22288), .ZN(n22292) );
  NOR2_X1 U23999 ( .A1(n22290), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n22291) );
  AOI211_X1 U24000 ( .C1(n22293), .C2(n22359), .A(n22292), .B(n22291), .ZN(
        n22294) );
  OAI21_X1 U24001 ( .B1(n22296), .B2(n22295), .A(n22294), .ZN(n22297) );
  AOI21_X1 U24002 ( .B1(n22298), .B2(n22360), .A(n22297), .ZN(n22299) );
  OAI21_X1 U24003 ( .B1(n22300), .B2(n22384), .A(n22299), .ZN(P1_U2833) );
  NOR2_X1 U24004 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22301), .ZN(n22312) );
  INV_X1 U24005 ( .A(n22302), .ZN(n22304) );
  OAI22_X1 U24006 ( .A1(n22304), .A2(n22377), .B1(n22342), .B2(n22303), .ZN(
        n22305) );
  AOI211_X1 U24007 ( .C1(n22355), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n22353), .B(n22305), .ZN(n22310) );
  OAI22_X1 U24008 ( .A1(n22307), .A2(n22379), .B1(n22306), .B2(n22384), .ZN(
        n22308) );
  INV_X1 U24009 ( .A(n22308), .ZN(n22309) );
  OAI211_X1 U24010 ( .C1(n22312), .C2(n22311), .A(n22310), .B(n22309), .ZN(
        P1_U2832) );
  NOR2_X1 U24011 ( .A1(n22373), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n22331) );
  AOI22_X1 U24012 ( .A1(n22331), .A2(n22313), .B1(n22376), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n22322) );
  INV_X1 U24013 ( .A(n22314), .ZN(n22318) );
  INV_X1 U24014 ( .A(n22330), .ZN(n22316) );
  OAI222_X1 U24015 ( .A1(n22377), .A2(n22318), .B1(n22317), .B2(n22316), .C1(
        n22315), .C2(n22370), .ZN(n22319) );
  AOI211_X1 U24016 ( .C1(n22320), .C2(n22360), .A(n22353), .B(n22319), .ZN(
        n22321) );
  OAI211_X1 U24017 ( .C1(n22323), .C2(n22384), .A(n22322), .B(n22321), .ZN(
        P1_U2829) );
  INV_X1 U24018 ( .A(n22324), .ZN(n22326) );
  OAI22_X1 U24019 ( .A1(n22326), .A2(n22377), .B1(n22342), .B2(n22325), .ZN(
        n22327) );
  AOI211_X1 U24020 ( .C1(n22355), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n22353), .B(n22327), .ZN(n22337) );
  AOI22_X1 U24021 ( .A1(n22329), .A2(n22357), .B1(n22360), .B2(n22328), .ZN(
        n22336) );
  OAI21_X1 U24022 ( .B1(n22331), .B2(n22330), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n22335) );
  NAND3_X1 U24023 ( .A1(n22333), .A2(n22332), .A3(n16950), .ZN(n22334) );
  NAND4_X1 U24024 ( .A1(n22337), .A2(n22336), .A3(n22335), .A4(n22334), .ZN(
        P1_U2828) );
  AOI21_X1 U24025 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n22339), .A(n22338), 
        .ZN(n22349) );
  OAI22_X1 U24026 ( .A1(n22342), .A2(n22341), .B1(n22340), .B2(n22370), .ZN(
        n22343) );
  AOI211_X1 U24027 ( .C1(n22357), .C2(n22344), .A(n22353), .B(n22343), .ZN(
        n22348) );
  AOI22_X1 U24028 ( .A1(n22346), .A2(n22360), .B1(n22359), .B2(n22345), .ZN(
        n22347) );
  OAI211_X1 U24029 ( .C1(n22350), .C2(n22349), .A(n22348), .B(n22347), .ZN(
        P1_U2825) );
  NOR3_X1 U24030 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n22352), .A3(n22351), 
        .ZN(n22354) );
  AOI211_X1 U24031 ( .C1(n22355), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n22354), .B(n22353), .ZN(n22367) );
  AOI22_X1 U24032 ( .A1(n22357), .A2(n22356), .B1(n22376), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n22366) );
  AOI22_X1 U24033 ( .A1(n22361), .A2(n22360), .B1(n22359), .B2(n22358), .ZN(
        n22365) );
  OAI21_X1 U24034 ( .B1(n22363), .B2(n22362), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n22364) );
  NAND4_X1 U24035 ( .A1(n22367), .A2(n22366), .A3(n22365), .A4(n22364), .ZN(
        P1_U2821) );
  OAI22_X1 U24036 ( .A1(n22370), .A2(n13810), .B1(n22369), .B2(n22368), .ZN(
        n22375) );
  INV_X1 U24037 ( .A(n22371), .ZN(n22372) );
  NOR3_X1 U24038 ( .A1(n22373), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n22372), 
        .ZN(n22374) );
  AOI211_X1 U24039 ( .C1(n22376), .C2(P1_EBX_REG_21__SCAN_IN), .A(n22375), .B(
        n22374), .ZN(n22383) );
  OAI22_X1 U24040 ( .A1(n22380), .A2(n22379), .B1(n22378), .B2(n22377), .ZN(
        n22381) );
  INV_X1 U24041 ( .A(n22381), .ZN(n22382) );
  OAI211_X1 U24042 ( .C1(n22385), .C2(n22384), .A(n22383), .B(n22382), .ZN(
        P1_U2819) );
  OAI21_X1 U24043 ( .B1(n22388), .B2(n22387), .A(n22386), .ZN(P1_U2806) );
  NOR2_X1 U24044 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22389), .ZN(n22392) );
  AOI21_X1 U24045 ( .B1(n22392), .B2(n22391), .A(n22390), .ZN(n22394) );
  OAI211_X1 U24046 ( .C1(n22397), .C2(n22489), .A(n22394), .B(n22393), .ZN(
        P1_U3163) );
  OAI22_X1 U24047 ( .A1(n22397), .A2(n15600), .B1(n22396), .B2(n22395), .ZN(
        P1_U3466) );
  INV_X1 U24048 ( .A(n22398), .ZN(n22407) );
  AOI21_X1 U24049 ( .B1(n22401), .B2(n22400), .A(n22399), .ZN(n22402) );
  OAI22_X1 U24050 ( .A1(n22404), .A2(n22403), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22402), .ZN(n22405) );
  OAI21_X1 U24051 ( .B1(n22407), .B2(n22406), .A(n22405), .ZN(P1_U3161) );
  INV_X1 U24052 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22409) );
  OAI21_X1 U24053 ( .B1(n22410), .B2(n22409), .A(n22408), .ZN(P1_U3465) );
  OAI21_X1 U24054 ( .B1(n22414), .B2(n22411), .A(n22412), .ZN(P2_U2818) );
  OAI21_X1 U24055 ( .B1(n22414), .B2(n22413), .A(n22412), .ZN(P2_U3592) );
  OAI21_X1 U24056 ( .B1(n22418), .B2(n22415), .A(n22416), .ZN(P3_U2636) );
  OAI21_X1 U24057 ( .B1(n22418), .B2(n22417), .A(n22416), .ZN(P3_U3281) );
  INV_X1 U24058 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22443) );
  NAND2_X1 U24059 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n22438) );
  INV_X1 U24060 ( .A(n22438), .ZN(n22441) );
  AOI211_X1 U24061 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n22443), .B(
        n22441), .ZN(n22420) );
  INV_X1 U24062 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22436) );
  AOI21_X1 U24063 ( .B1(n22453), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22436), 
        .ZN(n22458) );
  AOI21_X1 U24064 ( .B1(NA), .B2(n22419), .A(n22440), .ZN(n22450) );
  OAI22_X1 U24065 ( .A1(n22421), .A2(n22420), .B1(n22458), .B2(n22450), .ZN(
        P3_U3029) );
  INV_X1 U24066 ( .A(n22422), .ZN(n22428) );
  INV_X1 U24067 ( .A(n22423), .ZN(n22424) );
  AOI211_X1 U24068 ( .C1(NA), .C2(n22426), .A(n22425), .B(n22424), .ZN(n22427)
         );
  OAI22_X1 U24069 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22428), .B1(n22787), 
        .B2(n22427), .ZN(P1_U3194) );
  INV_X1 U24070 ( .A(n22429), .ZN(n22430) );
  AND3_X1 U24071 ( .A1(n18316), .A2(HOLD), .A3(n22430), .ZN(n22431) );
  AOI21_X1 U24072 ( .B1(n22433), .B2(n22432), .A(n22431), .ZN(n22434) );
  OAI21_X1 U24073 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n22435), .A(n22434), .ZN(P2_U3209) );
  NOR2_X1 U24074 ( .A1(n22436), .A2(n22443), .ZN(n22449) );
  AOI21_X1 U24075 ( .B1(n22449), .B2(n22438), .A(n22437), .ZN(n22448) );
  OAI21_X1 U24076 ( .B1(n22453), .B2(n22440), .A(n22439), .ZN(n22447) );
  AOI21_X1 U24077 ( .B1(n22443), .B2(n22442), .A(n22441), .ZN(n22445) );
  OAI211_X1 U24078 ( .C1(n22445), .C2(n22453), .A(P3_STATE_REG_1__SCAN_IN), 
        .B(n22444), .ZN(n22446) );
  OAI211_X1 U24079 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(n22448), .A(n22447), 
        .B(n22446), .ZN(P3_U3030) );
  AND2_X1 U24080 ( .A1(n22449), .A2(n22452), .ZN(n22451) );
  NOR2_X1 U24081 ( .A1(n22451), .A2(n22450), .ZN(n22457) );
  NAND2_X1 U24082 ( .A1(n22453), .A2(n22452), .ZN(n22454) );
  AOI21_X1 U24083 ( .B1(n22454), .B2(P3_STATE_REG_1__SCAN_IN), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22455) );
  OAI211_X1 U24084 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(n22455), .A(HOLD), .B(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22456) );
  OAI21_X1 U24085 ( .B1(n22458), .B2(n22457), .A(n22456), .ZN(P3_U3031) );
  NOR3_X1 U24086 ( .A1(n22715), .A2(n22778), .A3(n22534), .ZN(n22459) );
  NOR2_X1 U24087 ( .A1(n22534), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22536) );
  NOR2_X1 U24088 ( .A1(n22459), .A2(n22536), .ZN(n22467) );
  INV_X1 U24089 ( .A(n22467), .ZN(n22461) );
  NOR2_X1 U24090 ( .A1(n22485), .A2(n22518), .ZN(n22466) );
  INV_X1 U24091 ( .A(n22464), .ZN(n22460) );
  NOR2_X1 U24092 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22462), .ZN(
        n22714) );
  AOI22_X1 U24093 ( .A1(n22778), .A2(n22552), .B1(n22559), .B2(n22714), .ZN(
        n22469) );
  INV_X1 U24094 ( .A(n22714), .ZN(n22463) );
  AOI22_X1 U24095 ( .A1(n22464), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22463), .ZN(n22465) );
  OAI211_X1 U24096 ( .C1(n22467), .C2(n22466), .A(n22529), .B(n22465), .ZN(
        n22716) );
  AOI22_X1 U24097 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n22715), .B2(n22561), .ZN(n22468) );
  OAI211_X1 U24098 ( .C1(n22719), .C2(n22555), .A(n22469), .B(n22468), .ZN(
        P1_U3033) );
  NOR3_X1 U24099 ( .A1(n22722), .A2(n22729), .A3(n22534), .ZN(n22472) );
  NOR2_X1 U24100 ( .A1(n22472), .A2(n22536), .ZN(n22479) );
  INV_X1 U24101 ( .A(n22479), .ZN(n22474) );
  NOR2_X1 U24102 ( .A1(n22485), .A2(n11222), .ZN(n22478) );
  NOR2_X1 U24103 ( .A1(n22473), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22503) );
  NOR3_X1 U24104 ( .A1(n22475), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22493) );
  NAND2_X1 U24105 ( .A1(n22524), .A2(n22493), .ZN(n22720) );
  OAI22_X1 U24106 ( .A1(n22681), .A2(n22564), .B1(n22543), .B2(n22720), .ZN(
        n22476) );
  INV_X1 U24107 ( .A(n22476), .ZN(n22481) );
  NOR2_X1 U24108 ( .A1(n22503), .A2(n22489), .ZN(n22508) );
  AOI21_X1 U24109 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22720), .A(n22508), 
        .ZN(n22477) );
  AOI22_X1 U24110 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n22729), .B2(n22561), .ZN(n22480) );
  OAI211_X1 U24111 ( .C1(n22726), .C2(n22555), .A(n22481), .B(n22480), .ZN(
        P1_U3049) );
  INV_X1 U24112 ( .A(n22493), .ZN(n22488) );
  OAI21_X1 U24113 ( .B1(n22483), .B2(n22482), .A(n22494), .ZN(n22491) );
  OR2_X1 U24114 ( .A1(n22485), .A2(n22484), .ZN(n22487) );
  NOR2_X1 U24115 ( .A1(n22524), .A2(n22488), .ZN(n22727) );
  INV_X1 U24116 ( .A(n22727), .ZN(n22486) );
  AND2_X1 U24117 ( .A1(n22487), .A2(n22486), .ZN(n22496) );
  OAI22_X1 U24118 ( .A1(n22489), .A2(n22488), .B1(n22491), .B2(n22496), .ZN(
        n22490) );
  AOI22_X1 U24119 ( .A1(n22728), .A2(n22561), .B1(n22727), .B2(n22559), .ZN(
        n22500) );
  INV_X1 U24120 ( .A(n22491), .ZN(n22497) );
  OAI21_X1 U24121 ( .B1(n22494), .B2(n22493), .A(n22492), .ZN(n22495) );
  AOI21_X1 U24122 ( .B1(n22497), .B2(n22496), .A(n22495), .ZN(n22498) );
  AOI22_X1 U24123 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22552), .B2(n22729), .ZN(n22499) );
  OAI211_X1 U24124 ( .C1(n22733), .C2(n22555), .A(n22500), .B(n22499), .ZN(
        P1_U3057) );
  NOR2_X1 U24125 ( .A1(n22737), .A2(n22534), .ZN(n22501) );
  AOI21_X1 U24126 ( .B1(n22501), .B2(n22735), .A(n22536), .ZN(n22511) );
  INV_X1 U24127 ( .A(n22511), .ZN(n22504) );
  NOR2_X1 U24128 ( .A1(n22502), .A2(n11222), .ZN(n22510) );
  NOR3_X1 U24129 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n22505), .ZN(n22613) );
  INV_X1 U24130 ( .A(n22613), .ZN(n22734) );
  OAI22_X1 U24131 ( .A1(n22735), .A2(n22544), .B1(n22734), .B2(n22543), .ZN(
        n22506) );
  INV_X1 U24132 ( .A(n22506), .ZN(n22513) );
  AOI211_X1 U24133 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22734), .A(n22508), 
        .B(n22507), .ZN(n22509) );
  OAI21_X1 U24134 ( .B1(n22511), .B2(n22510), .A(n22509), .ZN(n22738) );
  AOI22_X1 U24135 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22552), .B2(n22737), .ZN(n22512) );
  OAI211_X1 U24136 ( .C1(n22741), .C2(n22555), .A(n22513), .B(n22512), .ZN(
        P1_U3081) );
  INV_X1 U24137 ( .A(n22514), .ZN(n22743) );
  AOI22_X1 U24138 ( .A1(n22743), .A2(n22560), .B1(n22559), .B2(n22742), .ZN(
        n22516) );
  AOI22_X1 U24139 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n22750), .B2(n22561), .ZN(n22515) );
  OAI211_X1 U24140 ( .C1(n22564), .C2(n22747), .A(n22516), .B(n22515), .ZN(
        P1_U3105) );
  NOR3_X1 U24141 ( .A1(n22750), .A2(n22749), .A3(n22534), .ZN(n22517) );
  NOR2_X1 U24142 ( .A1(n22517), .A2(n22536), .ZN(n22531) );
  INV_X1 U24143 ( .A(n22531), .ZN(n22522) );
  AND2_X1 U24144 ( .A1(n22519), .A2(n22518), .ZN(n22530) );
  NAND2_X1 U24145 ( .A1(n22524), .A2(n22523), .ZN(n22527) );
  INV_X1 U24146 ( .A(n22527), .ZN(n22748) );
  AOI22_X1 U24147 ( .A1(n22750), .A2(n22552), .B1(n22559), .B2(n22748), .ZN(
        n22533) );
  INV_X1 U24148 ( .A(n22525), .ZN(n22526) );
  AOI21_X1 U24149 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22527), .A(n22526), 
        .ZN(n22528) );
  OAI211_X1 U24150 ( .C1(n22531), .C2(n22530), .A(n22529), .B(n22528), .ZN(
        n22751) );
  AOI22_X1 U24151 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22749), .B2(n22561), .ZN(n22532) );
  OAI211_X1 U24152 ( .C1(n22754), .C2(n22555), .A(n22533), .B(n22532), .ZN(
        P1_U3113) );
  NOR2_X1 U24153 ( .A1(n22535), .A2(n22534), .ZN(n22537) );
  AOI21_X1 U24154 ( .B1(n22537), .B2(n22551), .A(n22536), .ZN(n22550) );
  INV_X1 U24155 ( .A(n22550), .ZN(n22541) );
  AND2_X1 U24156 ( .A1(n22538), .A2(n11222), .ZN(n22549) );
  OR2_X1 U24157 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22542), .ZN(
        n22756) );
  OAI22_X1 U24158 ( .A1(n22772), .A2(n22544), .B1(n22756), .B2(n22543), .ZN(
        n22545) );
  INV_X1 U24159 ( .A(n22545), .ZN(n22554) );
  AOI22_X1 U24160 ( .A1(n22546), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22756), .ZN(n22547) );
  OAI211_X1 U24161 ( .C1(n22550), .C2(n22549), .A(n22548), .B(n22547), .ZN(
        n22761) );
  AOI22_X1 U24162 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22552), .B2(n22759), .ZN(n22553) );
  OAI211_X1 U24163 ( .C1(n22765), .C2(n22555), .A(n22554), .B(n22553), .ZN(
        P1_U3129) );
  INV_X1 U24164 ( .A(n22556), .ZN(n22767) );
  AOI22_X1 U24165 ( .A1(n22767), .A2(n22560), .B1(n22559), .B2(n22766), .ZN(
        n22558) );
  AOI22_X1 U24166 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n22768), .B2(n22561), .ZN(n22557) );
  OAI211_X1 U24167 ( .C1(n22564), .C2(n22772), .A(n22558), .B(n22557), .ZN(
        P1_U3137) );
  AOI22_X1 U24168 ( .A1(n22776), .A2(n22560), .B1(n22774), .B2(n22559), .ZN(
        n22563) );
  AOI22_X1 U24169 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n22778), .B2(n22561), .ZN(n22562) );
  OAI211_X1 U24170 ( .C1(n22564), .C2(n22782), .A(n22563), .B(n22562), .ZN(
        P1_U3153) );
  AOI22_X1 U24171 ( .A1(n22778), .A2(n22582), .B1(n22575), .B2(n22714), .ZN(
        n22566) );
  AOI22_X1 U24172 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n22715), .B2(n22576), .ZN(n22565) );
  OAI211_X1 U24173 ( .C1(n22719), .C2(n22585), .A(n22566), .B(n22565), .ZN(
        P1_U3034) );
  NOR2_X1 U24174 ( .A1(n22579), .A2(n22720), .ZN(n22567) );
  AOI21_X1 U24175 ( .B1(n22729), .B2(n22576), .A(n22567), .ZN(n22569) );
  AOI22_X1 U24176 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22722), .B2(n22582), .ZN(n22568) );
  OAI211_X1 U24177 ( .C1(n22726), .C2(n22585), .A(n22569), .B(n22568), .ZN(
        P1_U3050) );
  AOI22_X1 U24178 ( .A1(n22728), .A2(n22576), .B1(n22727), .B2(n22575), .ZN(
        n22571) );
  AOI22_X1 U24179 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22729), .B2(n22582), .ZN(n22570) );
  OAI211_X1 U24180 ( .C1(n22733), .C2(n22585), .A(n22571), .B(n22570), .ZN(
        P1_U3058) );
  OAI22_X1 U24181 ( .A1(n22735), .A2(n22580), .B1(n22734), .B2(n22579), .ZN(
        n22572) );
  INV_X1 U24182 ( .A(n22572), .ZN(n22574) );
  AOI22_X1 U24183 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22737), .B2(n22582), .ZN(n22573) );
  OAI211_X1 U24184 ( .C1(n22741), .C2(n22585), .A(n22574), .B(n22573), .ZN(
        P1_U3082) );
  AOI22_X1 U24185 ( .A1(n22750), .A2(n22582), .B1(n22748), .B2(n22575), .ZN(
        n22578) );
  AOI22_X1 U24186 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n22749), .B2(n22576), .ZN(n22577) );
  OAI211_X1 U24187 ( .C1(n22754), .C2(n22585), .A(n22578), .B(n22577), .ZN(
        P1_U3114) );
  OAI22_X1 U24188 ( .A1(n22772), .A2(n22580), .B1(n22756), .B2(n22579), .ZN(
        n22581) );
  INV_X1 U24189 ( .A(n22581), .ZN(n22584) );
  AOI22_X1 U24190 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n22759), .B2(n22582), .ZN(n22583) );
  OAI211_X1 U24191 ( .C1(n22765), .C2(n22585), .A(n22584), .B(n22583), .ZN(
        P1_U3130) );
  AOI22_X1 U24192 ( .A1(n22778), .A2(n22602), .B1(n22595), .B2(n22714), .ZN(
        n22587) );
  AOI22_X1 U24193 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n22715), .B2(n22596), .ZN(n22586) );
  OAI211_X1 U24194 ( .C1(n22719), .C2(n22605), .A(n22587), .B(n22586), .ZN(
        P1_U3035) );
  NOR2_X1 U24195 ( .A1(n22599), .A2(n22720), .ZN(n22588) );
  AOI21_X1 U24196 ( .B1(n22729), .B2(n22596), .A(n22588), .ZN(n22590) );
  AOI22_X1 U24197 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22722), .B2(n22602), .ZN(n22589) );
  OAI211_X1 U24198 ( .C1(n22726), .C2(n22605), .A(n22590), .B(n22589), .ZN(
        P1_U3051) );
  AOI22_X1 U24199 ( .A1(n22728), .A2(n22596), .B1(n22727), .B2(n22595), .ZN(
        n22592) );
  AOI22_X1 U24200 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22729), .B2(n22602), .ZN(n22591) );
  OAI211_X1 U24201 ( .C1(n22733), .C2(n22605), .A(n22592), .B(n22591), .ZN(
        P1_U3059) );
  AOI22_X1 U24202 ( .A1(n22737), .A2(n22602), .B1(n22613), .B2(n22595), .ZN(
        n22594) );
  AOI22_X1 U24203 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22614), .B2(n22596), .ZN(n22593) );
  OAI211_X1 U24204 ( .C1(n22741), .C2(n22605), .A(n22594), .B(n22593), .ZN(
        P1_U3083) );
  AOI22_X1 U24205 ( .A1(n22750), .A2(n22602), .B1(n22748), .B2(n22595), .ZN(
        n22598) );
  AOI22_X1 U24206 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22749), .B2(n22596), .ZN(n22597) );
  OAI211_X1 U24207 ( .C1(n22754), .C2(n22605), .A(n22598), .B(n22597), .ZN(
        P1_U3115) );
  OAI22_X1 U24208 ( .A1(n22772), .A2(n22600), .B1(n22756), .B2(n22599), .ZN(
        n22601) );
  INV_X1 U24209 ( .A(n22601), .ZN(n22604) );
  AOI22_X1 U24210 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22759), .B2(n22602), .ZN(n22603) );
  OAI211_X1 U24211 ( .C1(n22765), .C2(n22605), .A(n22604), .B(n22603), .ZN(
        P1_U3131) );
  AOI22_X1 U24212 ( .A1(n22778), .A2(n22624), .B1(n22617), .B2(n22714), .ZN(
        n22607) );
  AOI22_X1 U24213 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n22715), .B2(n22618), .ZN(n22606) );
  OAI211_X1 U24214 ( .C1(n22719), .C2(n22627), .A(n22607), .B(n22606), .ZN(
        P1_U3036) );
  NOR2_X1 U24215 ( .A1(n22621), .A2(n22720), .ZN(n22608) );
  AOI21_X1 U24216 ( .B1(n22729), .B2(n22618), .A(n22608), .ZN(n22610) );
  AOI22_X1 U24217 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22722), .B2(n22624), .ZN(n22609) );
  OAI211_X1 U24218 ( .C1(n22726), .C2(n22627), .A(n22610), .B(n22609), .ZN(
        P1_U3052) );
  AOI22_X1 U24219 ( .A1(n22729), .A2(n22624), .B1(n22727), .B2(n22617), .ZN(
        n22612) );
  AOI22_X1 U24220 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22728), .B2(n22618), .ZN(n22611) );
  OAI211_X1 U24221 ( .C1(n22733), .C2(n22627), .A(n22612), .B(n22611), .ZN(
        P1_U3060) );
  AOI22_X1 U24222 ( .A1(n22737), .A2(n22624), .B1(n22613), .B2(n22617), .ZN(
        n22616) );
  AOI22_X1 U24223 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22614), .B2(n22618), .ZN(n22615) );
  OAI211_X1 U24224 ( .C1(n22741), .C2(n22627), .A(n22616), .B(n22615), .ZN(
        P1_U3084) );
  AOI22_X1 U24225 ( .A1(n22750), .A2(n22624), .B1(n22748), .B2(n22617), .ZN(
        n22620) );
  AOI22_X1 U24226 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22749), .B2(n22618), .ZN(n22619) );
  OAI211_X1 U24227 ( .C1(n22754), .C2(n22627), .A(n22620), .B(n22619), .ZN(
        P1_U3116) );
  OAI22_X1 U24228 ( .A1(n22772), .A2(n22622), .B1(n22756), .B2(n22621), .ZN(
        n22623) );
  INV_X1 U24229 ( .A(n22623), .ZN(n22626) );
  AOI22_X1 U24230 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22759), .B2(n22624), .ZN(n22625) );
  OAI211_X1 U24231 ( .C1(n22765), .C2(n22627), .A(n22626), .B(n22625), .ZN(
        P1_U3132) );
  AOI22_X1 U24232 ( .A1(n22778), .A2(n22646), .B1(n22639), .B2(n22714), .ZN(
        n22629) );
  AOI22_X1 U24233 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n22715), .B2(n22640), .ZN(n22628) );
  OAI211_X1 U24234 ( .C1(n22719), .C2(n22649), .A(n22629), .B(n22628), .ZN(
        P1_U3037) );
  OAI22_X1 U24235 ( .A1(n22681), .A2(n22630), .B1(n22720), .B2(n22643), .ZN(
        n22631) );
  INV_X1 U24236 ( .A(n22631), .ZN(n22633) );
  AOI22_X1 U24237 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n22729), .B2(n22640), .ZN(n22632) );
  OAI211_X1 U24238 ( .C1(n22726), .C2(n22649), .A(n22633), .B(n22632), .ZN(
        P1_U3053) );
  AOI22_X1 U24239 ( .A1(n22729), .A2(n22646), .B1(n22727), .B2(n22639), .ZN(
        n22635) );
  AOI22_X1 U24240 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22728), .B2(n22640), .ZN(n22634) );
  OAI211_X1 U24241 ( .C1(n22733), .C2(n22649), .A(n22635), .B(n22634), .ZN(
        P1_U3061) );
  OAI22_X1 U24242 ( .A1(n22735), .A2(n22644), .B1(n22734), .B2(n22643), .ZN(
        n22636) );
  INV_X1 U24243 ( .A(n22636), .ZN(n22638) );
  AOI22_X1 U24244 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22737), .B2(n22646), .ZN(n22637) );
  OAI211_X1 U24245 ( .C1(n22741), .C2(n22649), .A(n22638), .B(n22637), .ZN(
        P1_U3085) );
  AOI22_X1 U24246 ( .A1(n22750), .A2(n22646), .B1(n22748), .B2(n22639), .ZN(
        n22642) );
  AOI22_X1 U24247 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n22749), .B2(n22640), .ZN(n22641) );
  OAI211_X1 U24248 ( .C1(n22754), .C2(n22649), .A(n22642), .B(n22641), .ZN(
        P1_U3117) );
  OAI22_X1 U24249 ( .A1(n22772), .A2(n22644), .B1(n22756), .B2(n22643), .ZN(
        n22645) );
  INV_X1 U24250 ( .A(n22645), .ZN(n22648) );
  AOI22_X1 U24251 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22759), .B2(n22646), .ZN(n22647) );
  OAI211_X1 U24252 ( .C1(n22765), .C2(n22649), .A(n22648), .B(n22647), .ZN(
        P1_U3133) );
  AOI22_X1 U24253 ( .A1(n22778), .A2(n22668), .B1(n22661), .B2(n22714), .ZN(
        n22651) );
  AOI22_X1 U24254 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22715), .B2(n22662), .ZN(n22650) );
  OAI211_X1 U24255 ( .C1(n22719), .C2(n22671), .A(n22651), .B(n22650), .ZN(
        P1_U3038) );
  OAI22_X1 U24256 ( .A1(n22681), .A2(n22652), .B1(n22720), .B2(n22665), .ZN(
        n22653) );
  INV_X1 U24257 ( .A(n22653), .ZN(n22655) );
  AOI22_X1 U24258 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n22729), .B2(n22662), .ZN(n22654) );
  OAI211_X1 U24259 ( .C1(n22726), .C2(n22671), .A(n22655), .B(n22654), .ZN(
        P1_U3054) );
  AOI22_X1 U24260 ( .A1(n22728), .A2(n22662), .B1(n22727), .B2(n22661), .ZN(
        n22657) );
  AOI22_X1 U24261 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22729), .B2(n22668), .ZN(n22656) );
  OAI211_X1 U24262 ( .C1(n22733), .C2(n22671), .A(n22657), .B(n22656), .ZN(
        P1_U3062) );
  OAI22_X1 U24263 ( .A1(n22735), .A2(n22666), .B1(n22734), .B2(n22665), .ZN(
        n22658) );
  INV_X1 U24264 ( .A(n22658), .ZN(n22660) );
  AOI22_X1 U24265 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22737), .B2(n22668), .ZN(n22659) );
  OAI211_X1 U24266 ( .C1(n22741), .C2(n22671), .A(n22660), .B(n22659), .ZN(
        P1_U3086) );
  AOI22_X1 U24267 ( .A1(n22749), .A2(n22662), .B1(n22748), .B2(n22661), .ZN(
        n22664) );
  AOI22_X1 U24268 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22750), .B2(n22668), .ZN(n22663) );
  OAI211_X1 U24269 ( .C1(n22754), .C2(n22671), .A(n22664), .B(n22663), .ZN(
        P1_U3118) );
  OAI22_X1 U24270 ( .A1(n22772), .A2(n22666), .B1(n22756), .B2(n22665), .ZN(
        n22667) );
  INV_X1 U24271 ( .A(n22667), .ZN(n22670) );
  AOI22_X1 U24272 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22759), .B2(n22668), .ZN(n22669) );
  OAI211_X1 U24273 ( .C1(n22765), .C2(n22671), .A(n22670), .B(n22669), .ZN(
        P1_U3134) );
  AOI22_X1 U24274 ( .A1(n22778), .A2(n22709), .B1(n22697), .B2(n22714), .ZN(
        n22673) );
  AOI22_X1 U24275 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22716), .B1(
        n22715), .B2(n22698), .ZN(n22672) );
  OAI211_X1 U24276 ( .C1(n22719), .C2(n22706), .A(n22673), .B(n22672), .ZN(
        P1_U3039) );
  INV_X1 U24277 ( .A(n22674), .ZN(n22676) );
  AOI22_X1 U24278 ( .A1(n22676), .A2(n22691), .B1(n22697), .B2(n22675), .ZN(
        n22679) );
  AOI22_X1 U24279 ( .A1(n22677), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n22715), .B2(n22709), .ZN(n22678) );
  OAI211_X1 U24280 ( .C1(n22713), .C2(n22681), .A(n22679), .B(n22678), .ZN(
        P1_U3047) );
  OAI22_X1 U24281 ( .A1(n22681), .A2(n22680), .B1(n22720), .B2(n22705), .ZN(
        n22682) );
  INV_X1 U24282 ( .A(n22682), .ZN(n22684) );
  AOI22_X1 U24283 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n22698), .B2(n22729), .ZN(n22683) );
  OAI211_X1 U24284 ( .C1(n22726), .C2(n22706), .A(n22684), .B(n22683), .ZN(
        P1_U3055) );
  AOI22_X1 U24285 ( .A1(n22729), .A2(n22709), .B1(n22727), .B2(n22697), .ZN(
        n22686) );
  AOI22_X1 U24286 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22728), .B2(n22698), .ZN(n22685) );
  OAI211_X1 U24287 ( .C1(n22733), .C2(n22706), .A(n22686), .B(n22685), .ZN(
        P1_U3063) );
  OAI22_X1 U24288 ( .A1(n22735), .A2(n22713), .B1(n22705), .B2(n22734), .ZN(
        n22687) );
  INV_X1 U24289 ( .A(n22687), .ZN(n22689) );
  AOI22_X1 U24290 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22737), .B2(n22709), .ZN(n22688) );
  OAI211_X1 U24291 ( .C1(n22741), .C2(n22706), .A(n22689), .B(n22688), .ZN(
        P1_U3087) );
  AOI22_X1 U24292 ( .A1(n22692), .A2(n22691), .B1(n22697), .B2(n22690), .ZN(
        n22696) );
  AOI22_X1 U24293 ( .A1(n22694), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22693), .B2(n22709), .ZN(n22695) );
  OAI211_X1 U24294 ( .C1(n22713), .C2(n22747), .A(n22696), .B(n22695), .ZN(
        P1_U3103) );
  AOI22_X1 U24295 ( .A1(n22749), .A2(n22698), .B1(n22697), .B2(n22748), .ZN(
        n22700) );
  AOI22_X1 U24296 ( .A1(n22751), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n22750), .B2(n22709), .ZN(n22699) );
  OAI211_X1 U24297 ( .C1(n22754), .C2(n22706), .A(n22700), .B(n22699), .ZN(
        P1_U3119) );
  OAI22_X1 U24298 ( .A1(n22772), .A2(n22713), .B1(n22705), .B2(n22756), .ZN(
        n22701) );
  INV_X1 U24299 ( .A(n22701), .ZN(n22703) );
  AOI22_X1 U24300 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22759), .B2(n22709), .ZN(n22702) );
  OAI211_X1 U24301 ( .C1(n22765), .C2(n22706), .A(n22703), .B(n22702), .ZN(
        P1_U3135) );
  OAI22_X1 U24302 ( .A1(n22707), .A2(n22706), .B1(n22705), .B2(n22704), .ZN(
        n22708) );
  INV_X1 U24303 ( .A(n22708), .ZN(n22712) );
  AOI22_X1 U24304 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n22768), .B2(n22709), .ZN(n22711) );
  OAI211_X1 U24305 ( .C1(n22713), .C2(n22782), .A(n22712), .B(n22711), .ZN(
        P1_U3151) );
  AOI22_X1 U24306 ( .A1(n22778), .A2(n22760), .B1(n22773), .B2(n22714), .ZN(
        n22718) );
  AOI22_X1 U24307 ( .A1(n22716), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n22715), .B2(n22777), .ZN(n22717) );
  OAI211_X1 U24308 ( .C1(n22719), .C2(n22764), .A(n22718), .B(n22717), .ZN(
        P1_U3040) );
  NOR2_X1 U24309 ( .A1(n22755), .A2(n22720), .ZN(n22721) );
  AOI21_X1 U24310 ( .B1(n22729), .B2(n22777), .A(n22721), .ZN(n22725) );
  AOI22_X1 U24311 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22723), .B1(
        n22722), .B2(n22760), .ZN(n22724) );
  OAI211_X1 U24312 ( .C1(n22726), .C2(n22764), .A(n22725), .B(n22724), .ZN(
        P1_U3056) );
  AOI22_X1 U24313 ( .A1(n22728), .A2(n22777), .B1(n22727), .B2(n22773), .ZN(
        n22732) );
  AOI22_X1 U24314 ( .A1(n22730), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22760), .B2(n22729), .ZN(n22731) );
  OAI211_X1 U24315 ( .C1(n22733), .C2(n22764), .A(n22732), .B(n22731), .ZN(
        P1_U3064) );
  OAI22_X1 U24316 ( .A1(n22735), .A2(n22757), .B1(n22734), .B2(n22755), .ZN(
        n22736) );
  INV_X1 U24317 ( .A(n22736), .ZN(n22740) );
  AOI22_X1 U24318 ( .A1(n22738), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22760), .B2(n22737), .ZN(n22739) );
  OAI211_X1 U24319 ( .C1(n22741), .C2(n22764), .A(n22740), .B(n22739), .ZN(
        P1_U3088) );
  AOI22_X1 U24320 ( .A1(n22743), .A2(n22775), .B1(n22773), .B2(n22742), .ZN(
        n22746) );
  AOI22_X1 U24321 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n22750), .B2(n22777), .ZN(n22745) );
  OAI211_X1 U24322 ( .C1(n22783), .C2(n22747), .A(n22746), .B(n22745), .ZN(
        P1_U3112) );
  AOI22_X1 U24323 ( .A1(n22749), .A2(n22777), .B1(n22748), .B2(n22773), .ZN(
        n22753) );
  AOI22_X1 U24324 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22751), .B1(
        n22750), .B2(n22760), .ZN(n22752) );
  OAI211_X1 U24325 ( .C1(n22754), .C2(n22764), .A(n22753), .B(n22752), .ZN(
        P1_U3120) );
  OAI22_X1 U24326 ( .A1(n22772), .A2(n22757), .B1(n22756), .B2(n22755), .ZN(
        n22758) );
  INV_X1 U24327 ( .A(n22758), .ZN(n22763) );
  AOI22_X1 U24328 ( .A1(n22761), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n22760), .B2(n22759), .ZN(n22762) );
  OAI211_X1 U24329 ( .C1(n22765), .C2(n22764), .A(n22763), .B(n22762), .ZN(
        P1_U3136) );
  AOI22_X1 U24330 ( .A1(n22767), .A2(n22775), .B1(n22773), .B2(n22766), .ZN(
        n22771) );
  AOI22_X1 U24331 ( .A1(n22769), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n22768), .B2(n22777), .ZN(n22770) );
  OAI211_X1 U24332 ( .C1(n22783), .C2(n22772), .A(n22771), .B(n22770), .ZN(
        P1_U3144) );
  AOI22_X1 U24333 ( .A1(n22776), .A2(n22775), .B1(n22774), .B2(n22773), .ZN(
        n22781) );
  AOI22_X1 U24334 ( .A1(n22779), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22778), .B2(n22777), .ZN(n22780) );
  OAI211_X1 U24335 ( .C1(n22783), .C2(n22782), .A(n22781), .B(n22780), .ZN(
        P1_U3160) );
  INV_X1 U24336 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22786) );
  AOI22_X1 U24337 ( .A1(n22787), .A2(n22786), .B1(n22785), .B2(n22784), .ZN(
        P1_U3486) );
  CLKBUF_X1 U11270 ( .A(n13191), .Z(n11160) );
  CLKBUF_X1 U11273 ( .A(n11161), .Z(n13968) );
  CLKBUF_X1 U11294 ( .A(n13092), .Z(n14409) );
  INV_X1 U11297 ( .A(n20528), .ZN(n11304) );
  CLKBUF_X2 U11344 ( .A(n12402), .Z(n12560) );
  CLKBUF_X3 U11372 ( .A(n18408), .Z(n11159) );
  CLKBUF_X3 U11373 ( .A(n14092), .Z(n18621) );
  NOR2_X2 U11403 ( .A1(n16592), .A2(n16595), .ZN(n16593) );
  NAND2_X1 U11411 ( .A1(n16343), .A2(n16342), .ZN(n16341) );
  CLKBUF_X1 U11416 ( .A(n13516), .Z(n11212) );
  CLKBUF_X1 U11742 ( .A(n18251), .Z(n18265) );
  CLKBUF_X1 U11772 ( .A(n21001), .Z(n20998) );
  CLKBUF_X1 U12363 ( .A(n14705), .Z(n11222) );
  OR2_X1 U12460 ( .A1(n20528), .A2(n20527), .ZN(n22789) );
endmodule

