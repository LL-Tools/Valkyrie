

module b15_C_SARLock_k_64_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778;

  OR2_X2 U3429 ( .A1(n6610), .A2(n4145), .ZN(n5042) );
  BUF_X2 U3430 ( .A(n4156), .Z(n4157) );
  CLKBUF_X2 U3431 ( .A(n3310), .Z(n3953) );
  CLKBUF_X2 U3432 ( .A(n3255), .Z(n3944) );
  CLKBUF_X1 U3433 ( .A(n3440), .Z(n3390) );
  CLKBUF_X2 U3434 ( .A(n3355), .Z(n3871) );
  CLKBUF_X2 U3435 ( .A(n3254), .Z(n3945) );
  NAND2_X1 U3436 ( .A1(n3417), .A2(n3263), .ZN(n3272) );
  AND4_X1 U3437 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3153)
         );
  AND2_X2 U3438 ( .A1(n4377), .A2(n3129), .ZN(n3347) );
  INV_X2 U3439 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3450) );
  AND2_X1 U3440 ( .A1(n4448), .A2(n4377), .ZN(n3254) );
  NAND2_X1 U3441 ( .A1(n4491), .A2(n3288), .ZN(n5057) );
  INV_X1 U3442 ( .A(n3263), .ZN(n3155) );
  NAND2_X1 U3443 ( .A1(n3267), .A2(n5258), .ZN(n3294) );
  INV_X1 U3444 ( .A(n4157), .ZN(n5477) );
  AND2_X1 U34450 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U34460 ( .A1(n3425), .A2(n4427), .ZN(n3089) );
  AND2_X2 U34470 ( .A1(n3344), .A2(n3369), .ZN(n3418) );
  AND2_X1 U34480 ( .A1(n3271), .A2(n3288), .ZN(n4423) );
  NOR3_X1 U3449 ( .A1(n5315), .A2(REIP_REG_29__SCAN_IN), .A3(n6570), .ZN(n5302) );
  INV_X1 U3450 ( .A(n3271), .ZN(n4491) );
  NOR2_X1 U34510 ( .A1(n4865), .A2(n4864), .ZN(n4942) );
  INV_X1 U34520 ( .A(n5907), .ZN(n6258) );
  INV_X1 U34530 ( .A(n6027), .ZN(n6061) );
  INV_X1 U3454 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U34550 ( .A1(n4463), .A2(n4378), .ZN(n3315) );
  NOR2_X4 U34560 ( .A1(n6021), .A2(n6535), .ZN(n6017) );
  INV_X2 U3457 ( .A(n5360), .ZN(n3686) );
  NAND2_X2 U3458 ( .A1(n5401), .A2(n3091), .ZN(n5360) );
  NAND2_X4 U34590 ( .A1(n3154), .A2(n3153), .ZN(n3267) );
  NAND2_X2 U34600 ( .A1(n5306), .A2(n3939), .ZN(n5296) );
  INV_X2 U34610 ( .A(n5295), .ZN(n5306) );
  NAND2_X2 U34620 ( .A1(n3988), .A2(n3987), .ZN(n6197) );
  OAI21_X1 U34630 ( .B1(n5892), .B2(n3072), .A(n3070), .ZN(n5638) );
  NOR2_X2 U34640 ( .A1(n5563), .A2(n4068), .ZN(n2986) );
  NOR2_X2 U34650 ( .A1(n2989), .A2(n5596), .ZN(n5590) );
  NAND2_X1 U3466 ( .A1(n5603), .A2(n5572), .ZN(n5597) );
  NOR2_X1 U3467 ( .A1(n4865), .A2(n4864), .ZN(n2995) );
  NAND2_X1 U34680 ( .A1(n3448), .A2(n3447), .ZN(n4559) );
  NAND2_X1 U34690 ( .A1(n6074), .A2(n4436), .ZN(n5871) );
  NAND3_X1 U34700 ( .A1(n3293), .A2(n3155), .A3(n4123), .ZN(n4299) );
  NOR2_X1 U34710 ( .A1(n3294), .A2(n3295), .ZN(n4124) );
  AND2_X1 U34720 ( .A1(n3278), .A2(n4529), .ZN(n4338) );
  NAND3_X2 U34730 ( .A1(n3038), .A2(n3230), .A3(n3229), .ZN(n3271) );
  NOR2_X1 U34740 ( .A1(n3040), .A2(n3039), .ZN(n3038) );
  CLKBUF_X2 U3475 ( .A(n3144), .Z(n2997) );
  BUF_X2 U3476 ( .A(n3356), .Z(n3916) );
  CLKBUF_X2 U3477 ( .A(n3248), .Z(n3952) );
  CLKBUF_X2 U3478 ( .A(n3349), .Z(n3942) );
  CLKBUF_X2 U3479 ( .A(n3354), .Z(n3876) );
  INV_X1 U3480 ( .A(n3315), .ZN(n3144) );
  AND2_X2 U3481 ( .A1(n3129), .A2(n3128), .ZN(n3248) );
  AND2_X1 U3482 ( .A1(n4076), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3135)
         );
  INV_X2 U3483 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4395) );
  INV_X2 U3484 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n3407) );
  OR2_X1 U3485 ( .A1(n5582), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5574)
         );
  OR2_X1 U3486 ( .A1(n4070), .A2(n4069), .ZN(n3109) );
  OR2_X1 U3487 ( .A1(n5563), .A2(n4068), .ZN(n5559) );
  OR2_X1 U3488 ( .A1(n5439), .A2(n5255), .ZN(n5826) );
  NAND2_X1 U3489 ( .A1(n5605), .A2(n5604), .ZN(n5603) );
  NAND2_X1 U3490 ( .A1(n5571), .A2(n5570), .ZN(n5605) );
  OAI21_X1 U3491 ( .B1(n5568), .B2(n4065), .A(n3004), .ZN(n4067) );
  OR2_X1 U3492 ( .A1(n5569), .A2(n4064), .ZN(n5570) );
  CLKBUF_X1 U3493 ( .A(n5617), .Z(n2990) );
  INV_X1 U3494 ( .A(n5415), .ZN(n5416) );
  NAND2_X1 U3495 ( .A1(n4950), .A2(n4044), .ZN(n5075) );
  NAND2_X1 U3496 ( .A1(n3086), .A2(n3603), .ZN(n3618) );
  NAND2_X1 U3497 ( .A1(n4952), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U3498 ( .A1(n3605), .A2(n3604), .ZN(n3087) );
  NAND2_X1 U3499 ( .A1(n4668), .A2(n4034), .ZN(n4952) );
  NAND2_X1 U3500 ( .A1(n2995), .A2(n2996), .ZN(n3605) );
  NAND2_X1 U3501 ( .A1(n4670), .A2(n4669), .ZN(n4668) );
  AND2_X1 U3502 ( .A1(n4942), .A2(n3099), .ZN(n5165) );
  AND2_X1 U3503 ( .A1(n2991), .A2(n2992), .ZN(n4670) );
  NAND2_X2 U3504 ( .A1(n3510), .A2(n3509), .ZN(n4865) );
  NOR2_X1 U3505 ( .A1(n4713), .A2(n4773), .ZN(n6386) );
  AND3_X1 U3506 ( .A1(n6169), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n2988) );
  XNOR2_X1 U3507 ( .A(n3475), .B(n3476), .ZN(n4008) );
  INV_X1 U3508 ( .A(n3427), .ZN(n4418) );
  AND2_X1 U3509 ( .A1(n4419), .A2(n4420), .ZN(n3427) );
  OAI21_X1 U3510 ( .B1(n4476), .B2(n3564), .A(n3409), .ZN(n4419) );
  NAND2_X1 U3511 ( .A1(n3406), .A2(n3367), .ZN(n3429) );
  NAND3_X1 U3512 ( .A1(n3026), .A2(n3367), .A3(n3030), .ZN(n3406) );
  NAND2_X1 U3513 ( .A1(n3412), .A2(n3411), .ZN(n3416) );
  NAND2_X1 U3514 ( .A1(n3339), .A2(n3338), .ZN(n3367) );
  NAND2_X1 U3515 ( .A1(n3418), .A2(n6493), .ZN(n3410) );
  NAND2_X1 U3516 ( .A1(n4288), .A2(n4289), .ZN(n6610) );
  OR2_X1 U3517 ( .A1(n4487), .A2(n4299), .ZN(n4288) );
  NAND2_X1 U3518 ( .A1(n4382), .A2(n4416), .ZN(n4487) );
  NAND2_X2 U3519 ( .A1(n3046), .A2(n4121), .ZN(n4382) );
  AND2_X1 U3520 ( .A1(n3243), .A2(n4374), .ZN(n3292) );
  NOR2_X1 U3521 ( .A1(n5053), .A2(n4073), .ZN(n4106) );
  NOR2_X2 U3522 ( .A1(n3288), .A2(n3271), .ZN(n5053) );
  OR2_X1 U3523 ( .A1(n3333), .A2(n3332), .ZN(n4048) );
  AND2_X1 U3524 ( .A1(n3271), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4074) );
  INV_X1 U3525 ( .A(n3288), .ZN(n3298) );
  OR2_X1 U3526 ( .A1(n3362), .A2(n3361), .ZN(n3983) );
  INV_X1 U3527 ( .A(n3278), .ZN(n4533) );
  OR2_X2 U3528 ( .A1(n3240), .A2(n3239), .ZN(n4529) );
  AND2_X1 U3529 ( .A1(n3208), .A2(n3207), .ZN(n3214) );
  AND4_X1 U3530 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3154)
         );
  AND2_X2 U3531 ( .A1(n3112), .A2(n3260), .ZN(n3278) );
  AND4_X1 U3532 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3229)
         );
  AND4_X1 U3533 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n3230)
         );
  AND4_X1 U3534 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  AND4_X1 U3535 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3207)
         );
  AND4_X1 U3536 ( .A1(n3202), .A2(n3201), .A3(n3114), .A4(n3200), .ZN(n3208)
         );
  AND4_X1 U3537 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3215)
         );
  AND4_X1 U3538 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3140)
         );
  AND4_X1 U3539 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3141)
         );
  AND4_X1 U3540 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3142)
         );
  AND4_X1 U3541 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3143)
         );
  AND4_X1 U3542 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3260)
         );
  AND4_X1 U3543 ( .A1(n3111), .A2(n3190), .A3(n3189), .A4(n3188), .ZN(n3191)
         );
  AND4_X1 U3544 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3192)
         );
  AND4_X1 U3545 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3193)
         );
  AND4_X1 U3546 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3194)
         );
  AND4_X1 U3547 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3173)
         );
  AND4_X1 U3548 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n3175)
         );
  BUF_X2 U3549 ( .A(n3253), .Z(n3950) );
  CLKBUF_X2 U3550 ( .A(n3385), .Z(n3951) );
  AND2_X2 U3551 ( .A1(n3129), .A2(n4378), .ZN(n3247) );
  AND2_X2 U3552 ( .A1(n3135), .A2(n4448), .ZN(n3253) );
  AND2_X2 U3553 ( .A1(n3128), .A2(n4463), .ZN(n3348) );
  AND2_X2 U3554 ( .A1(n4448), .A2(n4378), .ZN(n3310) );
  AND2_X2 U3555 ( .A1(n3135), .A2(n3129), .ZN(n3355) );
  INV_X2 U3556 ( .A(n6620), .ZN(n6609) );
  AND2_X2 U3557 ( .A1(n4395), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3134)
         );
  AND2_X2 U3558 ( .A1(n4395), .A2(n3043), .ZN(n4448) );
  AND2_X2 U3559 ( .A1(n3450), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3129)
         );
  AND2_X2 U3560 ( .A1(n5266), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3128)
         );
  AND2_X2 U3561 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U3562 ( .A1(n4428), .A2(n4418), .ZN(n3088) );
  NAND2_X1 U3563 ( .A1(n4950), .A2(n2983), .ZN(n2980) );
  AND2_X1 U3564 ( .A1(n2980), .A2(n2981), .ZN(n5113) );
  OR2_X1 U3565 ( .A1(n2982), .A2(n5074), .ZN(n2981) );
  INV_X1 U3566 ( .A(n4053), .ZN(n2982) );
  AND2_X1 U3567 ( .A1(n4044), .A2(n4053), .ZN(n2983) );
  NAND2_X1 U3568 ( .A1(n5617), .A2(n3084), .ZN(n2984) );
  NAND2_X1 U3569 ( .A1(n5617), .A2(n3084), .ZN(n2985) );
  NAND2_X1 U3570 ( .A1(n5617), .A2(n3084), .ZN(n5569) );
  NAND2_X2 U3571 ( .A1(n4060), .A2(n3016), .ZN(n5617) );
  NOR2_X2 U3572 ( .A1(n5372), .A2(n6667), .ZN(n5966) );
  NAND2_X1 U3573 ( .A1(n5075), .A2(n5074), .ZN(n5073) );
  OAI21_X1 U3574 ( .B1(n3006), .B2(n5683), .A(n5532), .ZN(n5524) );
  NAND2_X1 U3576 ( .A1(n3274), .A2(n3273), .ZN(n3373) );
  NAND2_X1 U3577 ( .A1(n5590), .A2(n2988), .ZN(n5573) );
  AND2_X1 U3578 ( .A1(n6169), .A2(n5756), .ZN(n2989) );
  XNOR2_X1 U3579 ( .A(n4006), .B(n6279), .ZN(n4737) );
  NAND2_X1 U3580 ( .A1(n6185), .A2(n2994), .ZN(n2991) );
  OR2_X1 U3581 ( .A1(n2993), .A2(n4870), .ZN(n2992) );
  INV_X1 U3582 ( .A(n4025), .ZN(n2993) );
  AND2_X1 U3583 ( .A1(n4015), .A2(n4025), .ZN(n2994) );
  AND2_X1 U3584 ( .A1(n5217), .A2(n3099), .ZN(n2996) );
  AND2_X1 U3585 ( .A1(n3134), .A2(n4377), .ZN(n3255) );
  AOI21_X2 U3586 ( .B1(n4515), .B2(n4085), .A(n3992), .ZN(n6196) );
  NAND2_X2 U3587 ( .A1(n3686), .A2(n3033), .ZN(n5474) );
  AOI21_X1 U3588 ( .B1(n2987), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3378), 
        .ZN(n3380) );
  INV_X1 U3589 ( .A(n3428), .ZN(n3401) );
  NAND2_X1 U3590 ( .A1(n3400), .A2(n3399), .ZN(n3428) );
  AND2_X1 U3591 ( .A1(n3044), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U3592 ( .A1(n4005), .A2(n4004), .ZN(n4006) );
  NAND2_X2 U3593 ( .A1(n5415), .A2(n3618), .ZN(n5401) );
  AND4_X2 U3594 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3003)
         );
  AND2_X4 U3595 ( .A1(n3383), .A2(n4468), .ZN(n4385) );
  AND2_X1 U3596 ( .A1(n4074), .A2(n3244), .ZN(n4113) );
  AOI21_X1 U3597 ( .B1(n3244), .B2(n3271), .A(n6493), .ZN(n4118) );
  OAI21_X1 U3598 ( .B1(n3272), .B2(n3244), .A(n3246), .ZN(n4334) );
  BUF_X2 U3599 ( .A(n3989), .Z(n4515) );
  XNOR2_X2 U3600 ( .A(n3429), .B(n3401), .ZN(n3989) );
  OAI21_X2 U3601 ( .B1(n4517), .B2(n4104), .A(n3978), .ZN(n4311) );
  NAND2_X4 U3602 ( .A1(n3416), .A2(n3415), .ZN(n4517) );
  OAI21_X2 U3603 ( .B1(n5235), .B2(n5233), .A(n5231), .ZN(n5892) );
  NOR2_X2 U3604 ( .A1(n5458), .A2(n3095), .ZN(n5320) );
  NOR2_X2 U3605 ( .A1(n4438), .A2(n4552), .ZN(n4507) );
  NAND3_X2 U3606 ( .A1(n3024), .A2(n3088), .A3(n3089), .ZN(n4438) );
  AOI21_X1 U3607 ( .B1(n5275), .B2(n5296), .A(n5274), .ZN(n5528) );
  XNOR2_X1 U3608 ( .A(n5274), .B(n3976), .ZN(n4285) );
  NAND2_X2 U3609 ( .A1(n4143), .A2(n3298), .ZN(n4274) );
  NAND2_X2 U3611 ( .A1(n5466), .A2(n3740), .ZN(n5458) );
  NOR2_X4 U3612 ( .A1(n5474), .A2(n5475), .ZN(n5466) );
  OAI21_X1 U3613 ( .B1(n4476), .B2(n4104), .A(n3986), .ZN(n4481) );
  NAND2_X2 U3614 ( .A1(n3406), .A2(n3405), .ZN(n4476) );
  AOI21_X1 U3615 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6391), .A(n4112), 
        .ZN(n4117) );
  INV_X1 U3616 ( .A(n4109), .ZN(n4111) );
  NAND2_X1 U3617 ( .A1(n5257), .A2(n3032), .ZN(n3031) );
  INV_X1 U3618 ( .A(n5437), .ZN(n3032) );
  OR2_X1 U3619 ( .A1(n5258), .A2(n3407), .ZN(n3967) );
  AND2_X1 U3620 ( .A1(n3263), .A2(n3288), .ZN(n4085) );
  NAND2_X1 U3621 ( .A1(n4113), .A2(n4085), .ZN(n4119) );
  OR2_X1 U3622 ( .A1(n6484), .A2(n4144), .ZN(n4145) );
  OR2_X1 U3623 ( .A1(n6258), .A2(n6504), .ZN(n4144) );
  NAND2_X1 U3624 ( .A1(n3036), .A2(n3035), .ZN(n3491) );
  AND2_X1 U3625 ( .A1(n4559), .A2(n3476), .ZN(n3035) );
  NOR2_X1 U3626 ( .A1(n5267), .A2(n6493), .ZN(n3927) );
  NAND2_X1 U3627 ( .A1(n3407), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3663) );
  NAND2_X1 U3628 ( .A1(n3036), .A2(n4559), .ZN(n3475) );
  INV_X1 U3629 ( .A(n3885), .ZN(n3964) );
  NOR2_X2 U3630 ( .A1(n3267), .A2(n3407), .ZN(n3646) );
  AND2_X1 U3631 ( .A1(n5557), .A2(n5674), .ZN(n3083) );
  INV_X1 U3632 ( .A(n3398), .ZN(n3399) );
  NAND2_X1 U3633 ( .A1(n4385), .A2(n6493), .ZN(n3400) );
  NOR2_X1 U3634 ( .A1(n3009), .A2(n3048), .ZN(n3047) );
  OAI21_X1 U3635 ( .B1(n4119), .B2(n4137), .A(n3049), .ZN(n3048) );
  NAND2_X1 U3636 ( .A1(n6493), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3049) );
  NAND2_X1 U3637 ( .A1(n3435), .A2(n3434), .ZN(n4467) );
  XNOR2_X1 U3638 ( .A(n4468), .B(n4467), .ZN(n4445) );
  INV_X1 U3639 ( .A(n4423), .ZN(n4294) );
  NAND2_X1 U3640 ( .A1(n4231), .A2(n4157), .ZN(n4340) );
  INV_X1 U3641 ( .A(n5444), .ZN(n3848) );
  NAND2_X1 U3642 ( .A1(n4353), .A2(n4423), .ZN(n3059) );
  OR3_X1 U3643 ( .A1(n4487), .A2(READY_N), .A3(n4358), .ZN(n6124) );
  INV_X1 U3644 ( .A(n3967), .ZN(n3975) );
  NOR2_X2 U3645 ( .A1(n5296), .A2(n5275), .ZN(n5274) );
  NAND2_X1 U3646 ( .A1(n5279), .A2(n4157), .ZN(n5281) );
  AND2_X1 U3647 ( .A1(n6169), .A2(n5732), .ZN(n4068) );
  OAI21_X1 U3649 ( .B1(n5678), .B2(n6014), .A(n3108), .ZN(n3034) );
  INV_X1 U3650 ( .A(n3247), .ZN(n3384) );
  AOI22_X1 U3651 ( .A1(n3433), .A2(n4880), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3432), .ZN(n3306) );
  NAND2_X1 U3652 ( .A1(n3094), .A2(n5402), .ZN(n3093) );
  INV_X1 U3653 ( .A(n5390), .ZN(n3094) );
  INV_X1 U3654 ( .A(n5120), .ZN(n3566) );
  NOR2_X1 U3655 ( .A1(n5110), .A2(n3101), .ZN(n3100) );
  INV_X1 U3656 ( .A(n4944), .ZN(n3101) );
  XNOR2_X1 U3657 ( .A(n4047), .B(n3516), .ZN(n4035) );
  NAND2_X1 U3658 ( .A1(n3493), .A2(n3492), .ZN(n3511) );
  INV_X1 U3659 ( .A(n5349), .ZN(n3053) );
  NAND2_X1 U3660 ( .A1(n2984), .A2(n3000), .ZN(n5568) );
  NAND2_X1 U3661 ( .A1(n4423), .A2(n4157), .ZN(n4258) );
  OR2_X1 U3662 ( .A1(n3321), .A2(n3320), .ZN(n3982) );
  INV_X1 U3663 ( .A(n4085), .ZN(n4104) );
  INV_X1 U3664 ( .A(n4113), .ZN(n4094) );
  NAND2_X1 U3665 ( .A1(n5848), .A2(n3023), .ZN(n5340) );
  INV_X1 U3666 ( .A(n5379), .ZN(n5370) );
  NOR2_X1 U3667 ( .A1(n5442), .A2(n5262), .ZN(n5311) );
  OR2_X1 U3668 ( .A1(n3868), .A2(n3867), .ZN(n5437) );
  AND2_X1 U3669 ( .A1(n3299), .A2(n3278), .ZN(n4413) );
  BUF_X1 U3670 ( .A(n3294), .Z(n4325) );
  INV_X1 U3671 ( .A(n6499), .ZN(n4416) );
  XNOR2_X1 U3672 ( .A(n4132), .B(n4131), .ZN(n5034) );
  INV_X1 U3673 ( .A(n3663), .ZN(n3974) );
  INV_X1 U3674 ( .A(n5298), .ZN(n3939) );
  AOI21_X1 U3675 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n5305) );
  AND2_X1 U3676 ( .A1(n5815), .A2(n3885), .ZN(n3886) );
  NAND2_X1 U3677 ( .A1(n3096), .A2(n5332), .ZN(n3095) );
  INV_X1 U3678 ( .A(n3097), .ZN(n3096) );
  AND2_X1 U3679 ( .A1(n3706), .A2(n3685), .ZN(n3033) );
  INV_X1 U3680 ( .A(n5484), .ZN(n3706) );
  INV_X1 U3681 ( .A(n5417), .ZN(n3617) );
  AND2_X1 U3682 ( .A1(n3505), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3529)
         );
  NAND2_X1 U3683 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3451) );
  OR3_X1 U3684 ( .A1(n5540), .A2(n6169), .A3(n5723), .ZN(n5549) );
  NAND2_X1 U3685 ( .A1(n3118), .A2(n3012), .ZN(n5348) );
  OR2_X1 U3686 ( .A1(n6169), .A2(n5920), .ZN(n5649) );
  INV_X1 U3687 ( .A(n4059), .ZN(n3069) );
  NAND2_X1 U3688 ( .A1(n3037), .A2(n3075), .ZN(n5235) );
  AND2_X1 U3689 ( .A1(n3076), .A2(n4057), .ZN(n3075) );
  NAND2_X1 U3690 ( .A1(n3073), .A2(n5113), .ZN(n3037) );
  NAND2_X1 U3691 ( .A1(n5113), .A2(n5114), .ZN(n3081) );
  OR2_X1 U3692 ( .A1(n6169), .A2(n4054), .ZN(n6167) );
  AND2_X1 U3693 ( .A1(n4946), .A2(n4945), .ZN(n5986) );
  NAND2_X1 U3694 ( .A1(n4164), .A2(n4163), .ZN(n3060) );
  AND2_X1 U3695 ( .A1(n4352), .A2(n4344), .ZN(n5794) );
  INV_X1 U3696 ( .A(n3341), .ZN(n3342) );
  INV_X1 U3697 ( .A(n3340), .ZN(n3343) );
  NAND2_X1 U3698 ( .A1(n4445), .A2(n6493), .ZN(n3448) );
  OAI21_X1 U3699 ( .B1(n4115), .B2(n4114), .A(n3047), .ZN(n3046) );
  INV_X1 U3700 ( .A(n4543), .ZN(n4881) );
  AOI221_X1 U3701 ( .B1(n6569), .B2(n5379), .C1(n5835), .C2(n5379), .A(n5832), 
        .ZN(n5831) );
  NAND2_X1 U3702 ( .A1(n4423), .A2(n4268), .ZN(n6014) );
  AND2_X1 U3703 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4267), .ZN(n4268) );
  XNOR2_X1 U3704 ( .A(n4266), .B(n4265), .ZN(n5678) );
  OAI21_X1 U3705 ( .B1(n5309), .B2(n4264), .A(n5281), .ZN(n4266) );
  INV_X1 U3706 ( .A(n5497), .ZN(n6625) );
  AND2_X1 U3707 ( .A1(n6074), .A2(n5259), .ZN(n6068) );
  INV_X1 U3708 ( .A(n6074), .ZN(n6067) );
  OR2_X1 U3709 ( .A1(n6194), .A2(n4407), .ZN(n6204) );
  XNOR2_X1 U3710 ( .A(n4072), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5682)
         );
  NAND2_X1 U3711 ( .A1(n6469), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4102) );
  NAND2_X1 U3712 ( .A1(n4118), .A2(n3288), .ZN(n3045) );
  OR2_X1 U3713 ( .A1(n3468), .A2(n3467), .ZN(n4017) );
  INV_X1 U3714 ( .A(n3458), .ZN(n3036) );
  NOR2_X1 U3715 ( .A1(n4058), .A2(n3080), .ZN(n3079) );
  INV_X1 U3716 ( .A(n5208), .ZN(n3080) );
  NAND2_X1 U3717 ( .A1(n3493), .A2(n3042), .ZN(n4047) );
  AND2_X1 U3718 ( .A1(n3492), .A2(n3513), .ZN(n3042) );
  AOI21_X1 U3719 ( .B1(n3007), .B2(n3267), .A(n3278), .ZN(n3268) );
  OAI21_X1 U3720 ( .B1(n3044), .B2(n3267), .A(n3278), .ZN(n3262) );
  AOI22_X1 U3721 ( .A1(n3355), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3249) );
  NOR2_X1 U3722 ( .A1(n6533), .A2(n5063), .ZN(n4152) );
  NAND2_X1 U3723 ( .A1(n3098), .A2(n3759), .ZN(n3097) );
  INV_X1 U3724 ( .A(n5345), .ZN(n3098) );
  NAND2_X1 U3725 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3702)
         );
  INV_X1 U3726 ( .A(n3267), .ZN(n3417) );
  NAND2_X1 U3727 ( .A1(n3288), .A2(n4529), .ZN(n4156) );
  AND2_X1 U3728 ( .A1(n3085), .A2(n4061), .ZN(n3084) );
  NOR2_X1 U3729 ( .A1(n3113), .A2(n3017), .ZN(n3085) );
  AND2_X1 U3730 ( .A1(n6169), .A2(n5921), .ZN(n3113) );
  INV_X1 U3731 ( .A(n5404), .ZN(n3058) );
  INV_X1 U3732 ( .A(n5420), .ZN(n4207) );
  NAND2_X1 U3733 ( .A1(n3004), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4056) );
  NOR2_X1 U3734 ( .A1(n3078), .A2(n3074), .ZN(n3073) );
  INV_X1 U3735 ( .A(n5114), .ZN(n3074) );
  INV_X1 U3736 ( .A(n3079), .ZN(n3078) );
  NAND2_X1 U3737 ( .A1(n3079), .A2(n3077), .ZN(n3076) );
  INV_X1 U3738 ( .A(n5115), .ZN(n3077) );
  NOR2_X1 U3739 ( .A1(n5990), .A2(n5125), .ZN(n3065) );
  OR2_X1 U3740 ( .A1(n4513), .A2(n4671), .ZN(n3062) );
  OR2_X1 U3741 ( .A1(n3396), .A2(n3395), .ZN(n3999) );
  NAND2_X1 U3742 ( .A1(n3276), .A2(n3275), .ZN(n3340) );
  NAND2_X1 U3743 ( .A1(n3371), .A2(n3309), .ZN(n3368) );
  OR2_X1 U3744 ( .A1(n3446), .A2(n3445), .ZN(n4009) );
  OAI22_X1 U3745 ( .A1(n4108), .A2(n4107), .B1(n4113), .B2(n4140), .ZN(n4115)
         );
  AOI221_X1 U3746 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n4117), .C1(
        n4470), .C2(n4117), .A(n4116), .ZN(n4142) );
  AOI22_X1 U3747 ( .A1(n3347), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U3748 ( .A1(n3248), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3145) );
  INV_X1 U3749 ( .A(n4515), .ZN(n4770) );
  AND2_X1 U3750 ( .A1(n3303), .A2(n3375), .ZN(n4880) );
  OAI21_X1 U3751 ( .B1(n6615), .B2(n5803), .A(n6595), .ZN(n4524) );
  INV_X1 U3752 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U3753 ( .A1(n4281), .A2(n4282), .ZN(n4371) );
  INV_X1 U3754 ( .A(n4281), .ZN(n3293) );
  INV_X1 U3755 ( .A(n4143), .ZN(n4347) );
  INV_X1 U3756 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U3757 ( .A1(n6017), .A2(n3022), .ZN(n5991) );
  NAND2_X1 U3758 ( .A1(n6044), .A2(n4152), .ZN(n6021) );
  INV_X1 U3759 ( .A(n5055), .ZN(n6044) );
  AND2_X1 U3760 ( .A1(n5986), .A2(n3063), .ZN(n5220) );
  NOR2_X1 U3761 ( .A1(n3064), .A2(n5205), .ZN(n3063) );
  INV_X1 U3762 ( .A(n3065), .ZN(n3064) );
  AND2_X1 U3763 ( .A1(n3650), .A2(n3649), .ZN(n5390) );
  AND2_X1 U3764 ( .A1(n4129), .A2(n3936), .ZN(n5534) );
  NOR2_X1 U3765 ( .A1(n3906), .A2(n5552), .ZN(n3907) );
  NAND2_X1 U3766 ( .A1(n3866), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3906)
         );
  AND2_X1 U3767 ( .A1(n3843), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3844)
         );
  AND2_X1 U3768 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n3844), .ZN(n3866)
         );
  NOR2_X1 U3769 ( .A1(n3821), .A2(n5336), .ZN(n3843) );
  AND2_X1 U3771 ( .A1(n5337), .A2(n3885), .ZN(n3804) );
  AND2_X1 U3772 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3776), .ZN(n3777)
         );
  NOR2_X1 U3773 ( .A1(n3723), .A2(n5863), .ZN(n3724) );
  NAND2_X1 U3774 ( .A1(n3724), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3775)
         );
  NOR2_X1 U3775 ( .A1(n3702), .A2(n5368), .ZN(n3703) );
  NOR2_X1 U3776 ( .A1(n3093), .A2(n3092), .ZN(n3091) );
  INV_X1 U3777 ( .A(n5377), .ZN(n3092) );
  INV_X1 U3778 ( .A(n5401), .ZN(n3090) );
  NAND2_X1 U3779 ( .A1(n2990), .A2(n4061), .ZN(n5627) );
  NAND2_X1 U3780 ( .A1(n3633), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3651)
         );
  NAND2_X1 U3781 ( .A1(n3598), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3599)
         );
  NOR2_X1 U3782 ( .A1(n3582), .A2(n3581), .ZN(n3598) );
  INV_X1 U3783 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3581) );
  AND2_X1 U3784 ( .A1(n3015), .A2(n5166), .ZN(n3099) );
  NOR2_X1 U3785 ( .A1(n3550), .A2(n5992), .ZN(n3567) );
  NAND2_X1 U3786 ( .A1(n3534), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3550)
         );
  NOR2_X1 U3787 ( .A1(n3504), .A2(n4872), .ZN(n3505) );
  AOI21_X1 U3788 ( .B1(n4026), .B2(n3646), .A(n3508), .ZN(n4810) );
  NAND2_X1 U3789 ( .A1(n3490), .A2(n3489), .ZN(n4510) );
  CLKBUF_X1 U3790 ( .A(n4508), .Z(n4509) );
  AOI21_X1 U3791 ( .B1(n4008), .B2(n3646), .A(n3474), .ZN(n4552) );
  NOR2_X1 U3792 ( .A1(n3451), .A2(n4734), .ZN(n3470) );
  INV_X1 U3793 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4734) );
  INV_X1 U3794 ( .A(n3457), .ZN(n3024) );
  AOI21_X1 U3795 ( .B1(n3449), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3424), 
        .ZN(n4427) );
  AND2_X1 U3796 ( .A1(n3083), .A2(n3117), .ZN(n3082) );
  NAND2_X1 U3797 ( .A1(n5276), .A2(n4263), .ZN(n5279) );
  NOR2_X1 U3798 ( .A1(n3116), .A2(n4262), .ZN(n4263) );
  INV_X1 U3799 ( .A(n5276), .ZN(n5309) );
  AND2_X1 U3800 ( .A1(n5311), .A2(n5310), .ZN(n5276) );
  NAND2_X1 U3801 ( .A1(n5559), .A2(n3115), .ZN(n5530) );
  NAND2_X1 U3802 ( .A1(n3067), .A2(n3066), .ZN(n5442) );
  INV_X1 U3803 ( .A(n5440), .ZN(n3066) );
  AND2_X1 U3804 ( .A1(n3118), .A2(n3019), .ZN(n5335) );
  INV_X1 U3805 ( .A(n5333), .ZN(n3052) );
  NAND2_X1 U3806 ( .A1(n3118), .A2(n3013), .ZN(n5351) );
  NAND2_X1 U3807 ( .A1(n2985), .A2(n4063), .ZN(n5610) );
  NAND2_X1 U3808 ( .A1(n5392), .A2(n5381), .ZN(n5383) );
  INV_X1 U3809 ( .A(n3071), .ZN(n3070) );
  OAI21_X1 U3810 ( .B1(n3072), .B2(n5893), .A(n5649), .ZN(n3071) );
  NAND2_X1 U3811 ( .A1(n3021), .A2(n4059), .ZN(n3072) );
  AND2_X1 U3812 ( .A1(n4207), .A2(n3056), .ZN(n5392) );
  AND2_X1 U3813 ( .A1(n3014), .A2(n3057), .ZN(n3056) );
  INV_X1 U3814 ( .A(n5393), .ZN(n3057) );
  NAND2_X1 U3815 ( .A1(n4207), .A2(n3014), .ZN(n5406) );
  NAND2_X1 U3816 ( .A1(n4207), .A2(n4206), .ZN(n5418) );
  NAND2_X1 U3817 ( .A1(n5986), .A2(n3065), .ZN(n5204) );
  NAND2_X1 U3818 ( .A1(n5986), .A2(n4193), .ZN(n5987) );
  NOR2_X1 U3819 ( .A1(n4557), .A2(n3061), .ZN(n4946) );
  OR2_X1 U3820 ( .A1(n3062), .A2(n4867), .ZN(n3061) );
  OR2_X1 U3821 ( .A1(n4557), .A2(n3062), .ZN(n4866) );
  NAND2_X1 U3822 ( .A1(n4172), .A2(n4171), .ZN(n4441) );
  INV_X1 U3823 ( .A(n4432), .ZN(n4171) );
  NOR2_X1 U3824 ( .A1(n4441), .A2(n4440), .ZN(n4555) );
  INV_X1 U3825 ( .A(n5663), .ZN(n5238) );
  AND2_X1 U3826 ( .A1(n4676), .A2(n4675), .ZN(n6219) );
  NAND2_X1 U3827 ( .A1(n4352), .A2(n4345), .ZN(n6288) );
  OR2_X1 U3828 ( .A1(n3413), .A2(n4045), .ZN(n3027) );
  AND2_X1 U3829 ( .A1(n3411), .A2(n3029), .ZN(n3028) );
  NAND2_X1 U3830 ( .A1(n3337), .A2(n3336), .ZN(n3030) );
  NAND2_X1 U3831 ( .A1(n3429), .A2(n3428), .ZN(n3458) );
  OR2_X1 U3832 ( .A1(n3272), .A2(n3652), .ZN(n5267) );
  INV_X1 U3833 ( .A(n3380), .ZN(n3381) );
  AND2_X1 U3834 ( .A1(n4776), .A2(n6396), .ZN(n4778) );
  AND2_X1 U3835 ( .A1(n5812), .A2(n5140), .ZN(n6301) );
  AND2_X1 U3836 ( .A1(n4515), .A2(n4600), .ZN(n5809) );
  AND2_X1 U3837 ( .A1(n6395), .A2(n4476), .ZN(n4712) );
  AND2_X1 U3838 ( .A1(n4515), .A2(n4516), .ZN(n4525) );
  AND2_X1 U3839 ( .A1(n6587), .A2(n4524), .ZN(n4548) );
  CLKBUF_X1 U3840 ( .A(n4445), .Z(n6344) );
  INV_X1 U3841 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U3842 ( .A1(n6493), .A2(n4524), .ZN(n4543) );
  INV_X1 U3843 ( .A(n4517), .ZN(n4773) );
  AOI21_X1 U3844 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6460), .A(n4543), .ZN(
        n6402) );
  NAND2_X1 U3845 ( .A1(n5836), .A2(n4151), .ZN(n5830) );
  NOR2_X1 U3846 ( .A1(n5340), .A2(n6565), .ZN(n5836) );
  AOI21_X1 U3847 ( .B1(REIP_REG_23__SCAN_IN), .B2(n4154), .A(n5370), .ZN(n5832) );
  NOR2_X1 U3848 ( .A1(n5854), .A2(n6560), .ZN(n5848) );
  INV_X1 U3849 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5368) );
  INV_X1 U3850 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5395) );
  NOR2_X1 U3851 ( .A1(n4149), .A2(n5429), .ZN(n5397) );
  NOR2_X1 U3852 ( .A1(n5991), .A2(n5126), .ZN(n5980) );
  INV_X1 U3853 ( .A(n6056), .ZN(n5846) );
  AND2_X1 U3854 ( .A1(n5042), .A2(n5035), .ZN(n6027) );
  INV_X1 U3855 ( .A(n6014), .ZN(n6045) );
  NAND2_X1 U3856 ( .A1(n4324), .A2(n4148), .ZN(n5055) );
  NOR2_X1 U3857 ( .A1(n3051), .A2(n3050), .ZN(n4148) );
  NAND2_X1 U3858 ( .A1(n3271), .A2(n5036), .ZN(n3050) );
  AND2_X1 U3859 ( .A1(n5042), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6024) );
  INV_X1 U3860 ( .A(n5042), .ZN(n6054) );
  INV_X1 U3861 ( .A(n6024), .ZN(n6051) );
  AND2_X1 U3862 ( .A1(n5977), .A2(n5054), .ZN(n6026) );
  AND2_X1 U3863 ( .A1(n4417), .A2(n4416), .ZN(n5497) );
  INV_X1 U3864 ( .A(n6622), .ZN(n5499) );
  INV_X1 U3865 ( .A(n5871), .ZN(n6072) );
  NOR2_X1 U3866 ( .A1(n6067), .A2(n4436), .ZN(n6071) );
  NAND2_X1 U3867 ( .A1(n4283), .A2(n6124), .ZN(n6074) );
  OAI21_X1 U3868 ( .B1(n4366), .B2(n4280), .A(n4416), .ZN(n4283) );
  INV_X1 U3869 ( .A(n6071), .ZN(n5521) );
  INV_X1 U3870 ( .A(n6096), .ZN(n4492) );
  AOI21_X1 U3871 ( .B1(n5298), .B2(n5295), .A(n5297), .ZN(n5538) );
  AOI21_X1 U3872 ( .B1(n5308), .B2(n5307), .A(n5306), .ZN(n5547) );
  NAND2_X1 U3873 ( .A1(n3107), .A2(n3106), .ZN(n3105) );
  INV_X1 U3874 ( .A(n5257), .ZN(n3106) );
  INV_X1 U3875 ( .A(n5255), .ZN(n3107) );
  NAND2_X1 U3876 ( .A1(n5207), .A2(n5208), .ZN(n6168) );
  INV_X1 U3877 ( .A(n6204), .ZN(n5657) );
  NAND2_X1 U3878 ( .A1(n2986), .A2(n5557), .ZN(n5550) );
  AND2_X1 U3879 ( .A1(n3118), .A2(n4228), .ZN(n5462) );
  AOI21_X1 U3880 ( .B1(n5892), .B2(n5893), .A(n3069), .ZN(n3068) );
  AND2_X1 U3881 ( .A1(n5663), .A2(n4679), .ZN(n6281) );
  NAND2_X1 U3882 ( .A1(n4424), .A2(n4423), .ZN(n4422) );
  XNOR2_X1 U3883 ( .A(n3060), .B(n4353), .ZN(n4424) );
  CLKBUF_X1 U3884 ( .A(n4370), .Z(n6049) );
  NOR2_X1 U3885 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6593) );
  OAI21_X1 U3886 ( .B1(n5081), .B2(n6591), .A(n5009), .ZN(n5095) );
  INV_X1 U3887 ( .A(n6337), .ZN(n4593) );
  AND2_X1 U3888 ( .A1(DATAI_1_), .A2(n4881), .ZN(n6413) );
  INV_X1 U3889 ( .A(n4972), .ZN(n6411) );
  AND2_X1 U3890 ( .A1(DATAI_6_), .A2(n4881), .ZN(n6444) );
  AND2_X1 U3891 ( .A1(DATAI_7_), .A2(n4881), .ZN(n6454) );
  INV_X1 U3892 ( .A(n4965), .ZN(n6450) );
  NAND2_X1 U3893 ( .A1(n4272), .A2(REIP_REG_31__SCAN_IN), .ZN(n3055) );
  AOI21_X1 U3894 ( .B1(n4285), .B2(n6018), .A(n3034), .ZN(n3054) );
  OAI21_X1 U3895 ( .B1(n5818), .B2(n5977), .A(n3102), .ZN(U2800) );
  AOI21_X1 U3896 ( .B1(n3104), .B2(n5820), .A(n3103), .ZN(n3102) );
  OAI21_X1 U3897 ( .B1(n5817), .B2(n6014), .A(n3002), .ZN(n3103) );
  OR2_X1 U3898 ( .A1(n5819), .A2(REIP_REG_27__SCAN_IN), .ZN(n3104) );
  OAI21_X1 U3899 ( .B1(n5682), .B2(n6178), .A(n3001), .ZN(U2955) );
  AND2_X1 U3900 ( .A1(n4491), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2998) );
  INV_X1 U3901 ( .A(n5258), .ZN(n4421) );
  NAND2_X1 U3902 ( .A1(n4942), .A2(n4944), .ZN(n4943) );
  NOR2_X1 U3903 ( .A1(n3090), .A2(n3093), .ZN(n5376) );
  OR2_X1 U3904 ( .A1(n5458), .A2(n5459), .ZN(n5344) );
  AND2_X1 U3905 ( .A1(n4063), .A2(n4064), .ZN(n3000) );
  AND2_X1 U3906 ( .A1(n4136), .A2(n4135), .ZN(n3001) );
  AND2_X1 U3907 ( .A1(n4942), .A2(n3015), .ZN(n5121) );
  AND2_X1 U3908 ( .A1(n5821), .A2(n3020), .ZN(n3002) );
  INV_X1 U3909 ( .A(n3067), .ZN(n5445) );
  NOR2_X1 U3910 ( .A1(n5323), .A2(n5446), .ZN(n3067) );
  AND2_X1 U3911 ( .A1(n4047), .A2(n4046), .ZN(n3004) );
  NOR2_X1 U3912 ( .A1(n5458), .A2(n3097), .ZN(n5331) );
  AND2_X2 U3913 ( .A1(n3128), .A2(n4448), .ZN(n3349) );
  OR2_X1 U3914 ( .A1(n5627), .A2(n3113), .ZN(n3005) );
  AND2_X1 U3915 ( .A1(n2986), .A2(n3083), .ZN(n3006) );
  OAI21_X1 U3916 ( .B1(n3296), .B2(n3268), .A(n5053), .ZN(n3277) );
  AND2_X1 U3917 ( .A1(n3245), .A2(n3044), .ZN(n3007) );
  OR3_X1 U3918 ( .A1(n5289), .A2(REIP_REG_31__SCAN_IN), .A3(n6580), .ZN(n3008)
         );
  AND2_X1 U3919 ( .A1(n4142), .A2(n4118), .ZN(n3009) );
  NOR2_X1 U3920 ( .A1(n5438), .A2(n5437), .ZN(n5255) );
  NAND2_X1 U3921 ( .A1(n3263), .A2(n3044), .ZN(n3295) );
  AND2_X2 U3922 ( .A1(n3135), .A2(n4463), .ZN(n3356) );
  NAND3_X1 U3923 ( .A1(n4448), .A2(n4377), .A3(INSTQUEUE_REG_0__0__SCAN_IN), 
        .ZN(n3010) );
  INV_X1 U3924 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4076) );
  NAND2_X1 U3925 ( .A1(n5256), .A2(n5305), .ZN(n5295) );
  NAND2_X1 U3926 ( .A1(n3105), .A2(n5307), .ZN(n5818) );
  NAND3_X1 U3927 ( .A1(n3134), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .A3(n4377), 
        .ZN(n3011) );
  NAND3_X1 U3928 ( .A1(n3304), .A2(n3305), .A3(n3306), .ZN(n3371) );
  INV_X1 U3929 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3930 ( .A1(n3007), .A2(n5258), .ZN(n4281) );
  AND2_X2 U3931 ( .A1(n4378), .A2(n3134), .ZN(n3385) );
  NAND2_X1 U3932 ( .A1(n3686), .A2(n3685), .ZN(n5361) );
  INV_X1 U3933 ( .A(n3051), .ZN(n5052) );
  NAND2_X1 U3934 ( .A1(n5042), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3051) );
  NOR2_X1 U3935 ( .A1(n5383), .A2(n5366), .ZN(n5364) );
  INV_X1 U3936 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6493) );
  AND2_X1 U3937 ( .A1(n4228), .A2(n5461), .ZN(n3012) );
  AND2_X1 U3938 ( .A1(n3012), .A2(n3053), .ZN(n3013) );
  AND2_X1 U3939 ( .A1(n4206), .A2(n3058), .ZN(n3014) );
  NAND2_X1 U3940 ( .A1(n3081), .A2(n5115), .ZN(n5207) );
  INV_X1 U3941 ( .A(n3068), .ZN(n5648) );
  AND2_X1 U3942 ( .A1(n4338), .A2(n3271), .ZN(n4123) );
  NOR2_X1 U3943 ( .A1(n3365), .A2(n6493), .ZN(n4045) );
  INV_X1 U3944 ( .A(n4045), .ZN(n3029) );
  AND2_X1 U3945 ( .A1(n3100), .A2(n3566), .ZN(n3015) );
  NAND2_X1 U3946 ( .A1(n3618), .A2(n3087), .ZN(n5414) );
  OR2_X1 U3947 ( .A1(n6169), .A2(n5928), .ZN(n3016) );
  AND2_X1 U3948 ( .A1(n6169), .A2(n5771), .ZN(n3017) );
  NAND2_X1 U3949 ( .A1(n4942), .A2(n3100), .ZN(n3018) );
  NAND2_X1 U3950 ( .A1(n5335), .A2(n5324), .ZN(n5323) );
  AND2_X1 U3951 ( .A1(n3013), .A2(n3052), .ZN(n3019) );
  NAND2_X1 U3952 ( .A1(n3089), .A2(n3088), .ZN(n4426) );
  AOI21_X1 U3953 ( .B1(n4035), .B2(n3646), .A(n3518), .ZN(n4864) );
  OR2_X1 U3954 ( .A1(n5846), .A2(n5822), .ZN(n3020) );
  AND2_X1 U3955 ( .A1(n4413), .A2(n5053), .ZN(n4279) );
  NAND2_X1 U3956 ( .A1(n6169), .A2(n5920), .ZN(n3021) );
  INV_X1 U3957 ( .A(n5459), .ZN(n3759) );
  INV_X2 U3958 ( .A(n6173), .ZN(n5894) );
  OR2_X1 U3959 ( .A1(n4557), .A2(n4513), .ZN(n4511) );
  AND3_X1 U3960 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n3022) );
  AND2_X1 U3961 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n3023) );
  NOR2_X2 U3962 ( .A1(n6173), .A2(n6691), .ZN(n6451) );
  OR2_X1 U3963 ( .A1(n6511), .A2(n6400), .ZN(n6173) );
  OAI21_X1 U3964 ( .B1(n4439), .B2(n3024), .A(n4438), .ZN(n5072) );
  NAND2_X1 U3965 ( .A1(n3410), .A2(n3028), .ZN(n3025) );
  NAND2_X1 U3966 ( .A1(n3025), .A2(n3027), .ZN(n3404) );
  NAND2_X1 U3967 ( .A1(n3030), .A2(n3367), .ZN(n3403) );
  INV_X1 U3968 ( .A(n3404), .ZN(n3026) );
  NOR2_X2 U3969 ( .A1(n5438), .A2(n3031), .ZN(n5256) );
  NAND2_X1 U3970 ( .A1(n3248), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3041) );
  NAND4_X1 U3971 ( .A1(n3041), .A2(n3221), .A3(n3222), .A4(n3010), .ZN(n3039)
         );
  NAND4_X1 U3972 ( .A1(n3220), .A2(n3228), .A3(n3227), .A4(n3011), .ZN(n3040)
         );
  NOR2_X2 U3973 ( .A1(n5540), .A2(n5564), .ZN(n5563) );
  NAND2_X1 U3974 ( .A1(n4067), .A2(n4066), .ZN(n5540) );
  INV_X2 U3975 ( .A(n3244), .ZN(n3044) );
  NAND2_X1 U3976 ( .A1(n3045), .A2(n3263), .ZN(n4088) );
  NAND4_X4 U3977 ( .A1(n3003), .A2(n3174), .A3(n3175), .A4(n3173), .ZN(n3244)
         );
  NAND3_X1 U3978 ( .A1(n3008), .A2(n3055), .A3(n3054), .ZN(U2796) );
  NAND2_X1 U3979 ( .A1(n3060), .A2(n3059), .ZN(n4431) );
  INV_X1 U3980 ( .A(n5638), .ZN(n4060) );
  NAND2_X1 U3981 ( .A1(n2986), .A2(n3082), .ZN(n4071) );
  NAND3_X1 U3982 ( .A1(n3087), .A2(n3617), .A3(n3618), .ZN(n5415) );
  INV_X1 U3983 ( .A(n3605), .ZN(n3086) );
  NAND2_X1 U3984 ( .A1(n5401), .A2(n5402), .ZN(n5389) );
  NAND2_X1 U3985 ( .A1(n5320), .A2(n5322), .ZN(n5321) );
  AOI22_X1 U3986 ( .A1(n3346), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U3987 ( .A1(n3849), .A2(n3848), .ZN(n5438) );
  INV_X1 U3988 ( .A(n5321), .ZN(n3849) );
  CLKBUF_X1 U3989 ( .A(n5638), .Z(n5640) );
  AND2_X1 U3990 ( .A1(n4770), .A2(n3998), .ZN(n6395) );
  NOR2_X2 U3991 ( .A1(n5597), .A2(n5598), .ZN(n5596) );
  NAND2_X1 U3992 ( .A1(n4285), .A2(n4284), .ZN(n4287) );
  AND2_X1 U3993 ( .A1(n4270), .A2(n4269), .ZN(n3108) );
  OR2_X1 U3994 ( .A1(n5055), .A2(REIP_REG_30__SCAN_IN), .ZN(n3110) );
  INV_X1 U3995 ( .A(n3295), .ZN(n3242) );
  OR2_X2 U3996 ( .A1(n4487), .A2(n6476), .ZN(n6178) );
  OR2_X1 U3997 ( .A1(n3315), .A2(n4703), .ZN(n3111) );
  AND4_X1 U3998 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3112)
         );
  OR2_X1 U3999 ( .A1(n3315), .A2(n3199), .ZN(n3114) );
  OAI21_X1 U4000 ( .B1(n4094), .B2(n4911), .A(n3487), .ZN(n3492) );
  AND2_X1 U4001 ( .A1(n5556), .A2(n5706), .ZN(n3115) );
  NOR2_X1 U4002 ( .A1(n4340), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3116)
         );
  AND2_X1 U4003 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3117) );
  AND2_X1 U4004 ( .A1(n5364), .A2(n4222), .ZN(n3118) );
  OR2_X1 U4005 ( .A1(n3307), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3119)
         );
  OR2_X1 U4006 ( .A1(n4079), .A2(n4080), .ZN(n4092) );
  NAND2_X1 U4007 ( .A1(n4103), .A2(n4102), .ZN(n4109) );
  NAND2_X1 U4008 ( .A1(n3248), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3125) );
  INV_X1 U4009 ( .A(n5363), .ZN(n3685) );
  OR2_X1 U4010 ( .A1(n3315), .A2(n3160), .ZN(n3161) );
  NOR2_X1 U4011 ( .A1(n4111), .A2(n4110), .ZN(n4112) );
  OAI21_X1 U4012 ( .B1(n4094), .B2(n4906), .A(n3469), .ZN(n3476) );
  OR2_X1 U4013 ( .A1(n3486), .A2(n3485), .ZN(n4028) );
  INV_X1 U4014 ( .A(n5481), .ZN(n4222) );
  OR2_X1 U4015 ( .A1(n3503), .A2(n3502), .ZN(n4037) );
  NAND2_X1 U4016 ( .A1(n3242), .A2(n3241), .ZN(n4374) );
  NOR2_X1 U4017 ( .A1(n4529), .A2(n3263), .ZN(n3299) );
  OR2_X1 U4018 ( .A1(n3935), .A2(n3934), .ZN(n4129) );
  INV_X1 U4019 ( .A(n3775), .ZN(n3776) );
  NAND2_X1 U4020 ( .A1(n3567), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3582)
         );
  INV_X1 U4021 ( .A(n4810), .ZN(n3509) );
  NOR2_X1 U4022 ( .A1(n4294), .A2(EBX_REG_29__SCAN_IN), .ZN(n4262) );
  INV_X1 U4023 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4064) );
  INV_X1 U4024 ( .A(n5421), .ZN(n4206) );
  INV_X1 U4025 ( .A(n3414), .ZN(n3411) );
  INV_X1 U4026 ( .A(n5868), .ZN(n4150) );
  NAND2_X1 U4027 ( .A1(n3777), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3821)
         );
  AND2_X1 U4028 ( .A1(n3529), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3534)
         );
  NAND2_X1 U4029 ( .A1(n5966), .A2(n4150), .ZN(n5854) );
  INV_X1 U4030 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5992) );
  OR2_X1 U4031 ( .A1(n4487), .A2(n5271), .ZN(n4488) );
  NOR2_X1 U4032 ( .A1(n3651), .A2(n5395), .ZN(n3668) );
  NOR2_X1 U4033 ( .A1(n3599), .A2(n5424), .ZN(n3633) );
  OR2_X1 U4034 ( .A1(n6169), .A2(n4062), .ZN(n4063) );
  AND2_X1 U4035 ( .A1(n6167), .A2(n4056), .ZN(n4057) );
  OR2_X1 U4036 ( .A1(n4487), .A2(n4328), .ZN(n4329) );
  INV_X1 U4037 ( .A(n6286), .ZN(n6274) );
  OR2_X1 U4038 ( .A1(n5788), .A2(n5794), .ZN(n5663) );
  AND2_X1 U4039 ( .A1(n4352), .A2(n4456), .ZN(n5788) );
  AND2_X1 U4040 ( .A1(n3431), .A2(n4690), .ZN(n4879) );
  INV_X1 U4041 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6460) );
  INV_X1 U4042 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6501) );
  OR2_X1 U4043 ( .A1(n4291), .A2(n6499), .ZN(n4289) );
  INV_X1 U4044 ( .A(n5977), .ZN(n6018) );
  NAND2_X1 U4045 ( .A1(n5042), .A2(n5055), .ZN(n5379) );
  AND2_X1 U4046 ( .A1(n5497), .A2(n4421), .ZN(n6622) );
  NAND2_X1 U4047 ( .A1(n6166), .A2(n4488), .ZN(n4490) );
  OAI21_X1 U4048 ( .B1(n3281), .B2(n6612), .A(n4307), .ZN(n6149) );
  INV_X1 U4049 ( .A(n6113), .ZN(n6162) );
  NAND2_X1 U4050 ( .A1(n3703), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3723)
         );
  INV_X1 U4051 ( .A(n5627), .ZN(n5630) );
  NAND2_X1 U4052 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3470), .ZN(n3504)
         );
  INV_X1 U4053 ( .A(n6178), .ZN(n6199) );
  NAND2_X1 U4054 ( .A1(n5530), .A2(n5683), .ZN(n5532) );
  AND2_X1 U4055 ( .A1(n5911), .A2(n5672), .ZN(n5783) );
  AND2_X1 U4056 ( .A1(n5488), .A2(n5487), .ZN(n5971) );
  AND2_X1 U4057 ( .A1(n6281), .A2(n5660), .ZN(n5241) );
  AND2_X1 U4058 ( .A1(n6593), .A2(n6502), .ZN(n6206) );
  NAND2_X1 U4059 ( .A1(n4330), .A2(n4329), .ZN(n4352) );
  INV_X1 U4060 ( .A(n6208), .ZN(n6292) );
  AND2_X1 U4061 ( .A1(n4352), .A2(n4351), .ZN(n6286) );
  NAND2_X1 U4062 ( .A1(n6591), .A2(n3407), .ZN(n6400) );
  NAND2_X1 U4063 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4382), .ZN(n6595) );
  INV_X1 U4064 ( .A(n5029), .ZN(n4916) );
  INV_X1 U4065 ( .A(n6325), .ZN(n6329) );
  NAND2_X1 U4066 ( .A1(n4771), .A2(n4770), .ZN(n6300) );
  INV_X1 U4067 ( .A(n6344), .ZN(n5812) );
  INV_X1 U4068 ( .A(n5003), .ZN(n5100) );
  AND2_X1 U4069 ( .A1(n5809), .A2(n4569), .ZN(n6337) );
  INV_X1 U4070 ( .A(n6368), .ZN(n6376) );
  INV_X1 U4071 ( .A(n6390), .ZN(n6364) );
  INV_X1 U4072 ( .A(n4964), .ZN(n4992) );
  NOR2_X1 U4073 ( .A1(n4476), .A2(n4773), .ZN(n5137) );
  INV_X1 U4074 ( .A(n5183), .ZN(n6393) );
  INV_X1 U4075 ( .A(n5177), .ZN(n6423) );
  AND2_X1 U4076 ( .A1(n4525), .A2(n4517), .ZN(n4859) );
  INV_X1 U4077 ( .A(n4602), .ZN(n4650) );
  INV_X1 U4078 ( .A(n4982), .ZN(n6441) );
  AND2_X1 U4079 ( .A1(n6501), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4122) );
  INV_X1 U4080 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6528) );
  INV_X1 U4081 ( .A(n5547), .ZN(n5508) );
  INV_X1 U4082 ( .A(n5252), .ZN(n5230) );
  OR2_X1 U4083 ( .A1(n6096), .A2(n4491), .ZN(n6075) );
  NAND2_X1 U4084 ( .A1(n4490), .A2(n4489), .ZN(n6096) );
  INV_X1 U4085 ( .A(n6149), .ZN(n6113) );
  OR2_X2 U4086 ( .A1(n4487), .A2(n6490), .ZN(n6166) );
  NOR2_X1 U4087 ( .A1(n5795), .A2(n5241), .ZN(n6205) );
  NAND2_X1 U4088 ( .A1(n4352), .A2(n4333), .ZN(n6208) );
  INV_X1 U4089 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4775) );
  AND2_X1 U4090 ( .A1(n4883), .A2(n4882), .ZN(n5019) );
  OR2_X1 U4091 ( .A1(n4781), .A2(n4773), .ZN(n5029) );
  OR2_X1 U4092 ( .A1(n4781), .A2(n4517), .ZN(n5203) );
  OR2_X1 U4093 ( .A1(n6300), .A2(n5138), .ZN(n6325) );
  OR2_X1 U4094 ( .A1(n6300), .A2(n5000), .ZN(n6334) );
  NAND2_X1 U4095 ( .A1(n4712), .A2(n4773), .ZN(n4964) );
  NAND2_X1 U4096 ( .A1(n6395), .A2(n5137), .ZN(n6447) );
  NAND2_X1 U4097 ( .A1(n4525), .A2(n4773), .ZN(n4602) );
  INV_X1 U4098 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6591) );
  INV_X1 U4099 ( .A(n6586), .ZN(n6582) );
  NAND2_X1 U4100 ( .A1(n3144), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3123)
         );
  AND2_X4 U4101 ( .A1(n3128), .A2(n3134), .ZN(n3346) );
  NAND2_X1 U4102 ( .A1(n3346), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3122)
         );
  NAND2_X1 U4103 ( .A1(n3253), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3121) );
  NAND2_X1 U4104 ( .A1(n3356), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3120)
         );
  NAND2_X1 U4105 ( .A1(n3348), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3127)
         );
  NOR2_X4 U4106 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U4107 ( .A1(n3347), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3126) );
  NAND2_X1 U4108 ( .A1(n3385), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3124)
         );
  NAND2_X1 U4109 ( .A1(n3355), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4110 ( .A1(n3349), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U4111 ( .A1(n3247), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4112 ( .A1(n3310), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4113 ( .A1(n3255), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3139) );
  AND2_X4 U4114 ( .A1(n3135), .A2(n3134), .ZN(n3354) );
  NAND2_X1 U4115 ( .A1(n3354), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4116 ( .A1(n3254), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U4118 ( .A1(n3440), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3136)
         );
  NAND4_X4 U4119 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n3263)
         );
  AOI22_X1 U4120 ( .A1(n3255), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3144), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4121 ( .A1(n3355), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4122 ( .A1(n3385), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4123 ( .A1(n3356), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4124 ( .A1(n3348), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4125 ( .A1(n3155), .A2(n3267), .ZN(n3245) );
  NAND2_X1 U4126 ( .A1(n3354), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U4127 ( .A1(n3355), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4128 ( .A1(n3247), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U4129 ( .A1(n3310), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3156) );
  NAND2_X1 U4130 ( .A1(n3255), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4131 ( .A1(n3253), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4132 ( .A1(n3356), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3162)
         );
  INV_X1 U4133 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3160) );
  AND4_X2 U4134 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3174)
         );
  NAND2_X1 U4135 ( .A1(n3248), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U4136 ( .A1(n3348), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3167)
         );
  NAND2_X1 U4137 ( .A1(n3385), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3166)
         );
  NAND2_X1 U4138 ( .A1(n3349), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4139 ( .A1(n3347), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4140 ( .A1(n3346), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3171)
         );
  NAND2_X1 U4141 ( .A1(n3254), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4142 ( .A1(n3440), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3169)
         );
  NAND2_X1 U4143 ( .A1(n3348), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3179)
         );
  NAND2_X1 U4144 ( .A1(n3355), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U4145 ( .A1(n3248), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U4146 ( .A1(n3385), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3176)
         );
  NAND2_X1 U4147 ( .A1(n3354), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4148 ( .A1(n3347), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4149 ( .A1(n3349), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U4150 ( .A1(n3247), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U4151 ( .A1(n3255), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3187) );
  NAND2_X1 U4152 ( .A1(n3346), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3186)
         );
  NAND2_X1 U4153 ( .A1(n3253), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U4154 ( .A1(n3254), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4155 ( .A1(n3440), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3190)
         );
  NAND2_X1 U4156 ( .A1(n3356), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3189)
         );
  NAND2_X1 U4157 ( .A1(n3310), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3188) );
  NAND4_X4 U4158 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n5258)
         );
  NAND2_X1 U4159 ( .A1(n3255), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4160 ( .A1(n3346), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4161 ( .A1(n3356), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4162 ( .A1(n3254), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4163 ( .A1(n3354), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4164 ( .A1(n3347), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3201) );
  INV_X1 U4165 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4166 ( .A1(n3440), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3200)
         );
  NAND2_X1 U4167 ( .A1(n3355), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4168 ( .A1(n3385), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4169 ( .A1(n3348), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3204)
         );
  NAND2_X1 U4170 ( .A1(n3310), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4171 ( .A1(n3247), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4172 ( .A1(n3253), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4173 ( .A1(n3248), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4174 ( .A1(n3349), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3209) );
  NAND3_X4 U4175 ( .A1(n3215), .A2(n3214), .A3(n3213), .ZN(n3288) );
  NAND2_X1 U4176 ( .A1(n3253), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4177 ( .A1(n3346), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3218)
         );
  NAND2_X1 U4178 ( .A1(n3347), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4179 ( .A1(n3440), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4180 ( .A1(n3247), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4181 ( .A1(n3385), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3221)
         );
  NAND2_X1 U4182 ( .A1(n3349), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4183 ( .A1(n3354), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4184 ( .A1(n3355), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4185 ( .A1(n3348), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3224)
         );
  NAND2_X1 U4186 ( .A1(n3310), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4187 ( .A1(n3144), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4188 ( .A1(n3356), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3227)
         );
  AND2_X4 U4189 ( .A1(n3298), .A2(n3271), .ZN(n3281) );
  NAND2_X1 U4190 ( .A1(n4281), .A2(n3281), .ZN(n3243) );
  AOI22_X1 U4191 ( .A1(n3346), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4192 ( .A1(n3248), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3385), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4193 ( .A1(n3356), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3144), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4194 ( .A1(n3247), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3231) );
  NAND4_X1 U4195 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3240)
         );
  AOI22_X1 U4196 ( .A1(n3255), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4197 ( .A1(n3348), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4198 ( .A1(n3354), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4199 ( .A1(n3253), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3235) );
  NAND4_X1 U4200 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3239)
         );
  INV_X1 U4201 ( .A(n4156), .ZN(n3241) );
  AND2_X1 U4202 ( .A1(n3245), .A2(n5258), .ZN(n3246) );
  XNOR2_X1 U4203 ( .A(n6528), .B(STATE_REG_1__SCAN_IN), .ZN(n4147) );
  NOR2_X1 U4204 ( .A1(n3288), .A2(n4147), .ZN(n3301) );
  AOI22_X1 U4205 ( .A1(n3385), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4206 ( .A1(n3248), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4207 ( .A1(n3354), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4208 ( .A1(n3346), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4209 ( .A1(n3356), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4210 ( .A1(n3347), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4211 ( .A1(n3144), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3256) );
  OAI211_X1 U4212 ( .C1(n3301), .C2(n3263), .A(n4338), .B(n5057), .ZN(n3261)
         );
  NOR2_X1 U4213 ( .A1(n4334), .A2(n3261), .ZN(n3269) );
  NAND2_X1 U4214 ( .A1(n3262), .A2(n5258), .ZN(n3265) );
  INV_X1 U4215 ( .A(n3294), .ZN(n3300) );
  NAND2_X1 U4216 ( .A1(n3300), .A2(n3155), .ZN(n3264) );
  NAND2_X1 U4217 ( .A1(n3265), .A2(n3264), .ZN(n3266) );
  NAND2_X1 U4218 ( .A1(n3272), .A2(n4529), .ZN(n3282) );
  NAND2_X1 U4219 ( .A1(n3266), .A2(n3282), .ZN(n3296) );
  NAND3_X1 U4220 ( .A1(n3277), .A2(n3269), .A3(n3292), .ZN(n3270) );
  NAND2_X1 U4221 ( .A1(n3270), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4222 ( .A1(n4113), .A2(n3272), .ZN(n3273) );
  NAND2_X1 U4223 ( .A1(n3373), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4224 ( .A1(n6593), .A2(n6493), .ZN(n4125) );
  MUX2_X1 U4225 ( .A(n4122), .B(n4125), .S(n6460), .Z(n3275) );
  NOR2_X1 U4226 ( .A1(n4533), .A2(n3267), .ZN(n3279) );
  INV_X1 U4227 ( .A(n4529), .ZN(n4159) );
  NAND4_X1 U4228 ( .A1(n3279), .A2(n4159), .A3(n3244), .A4(n5258), .ZN(n4450)
         );
  INV_X1 U4229 ( .A(n4450), .ZN(n3280) );
  NAND2_X1 U4230 ( .A1(n6593), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6500) );
  NOR2_X1 U4231 ( .A1(n3280), .A2(n6500), .ZN(n3286) );
  NAND2_X1 U4232 ( .A1(n3282), .A2(n3281), .ZN(n3285) );
  INV_X1 U4233 ( .A(n5057), .ZN(n3284) );
  NOR2_X1 U4234 ( .A1(n3278), .A2(n4491), .ZN(n3283) );
  AOI21_X1 U4235 ( .B1(n3284), .B2(n3295), .A(n3283), .ZN(n4335) );
  AND3_X1 U4236 ( .A1(n3286), .A2(n3285), .A3(n4335), .ZN(n3291) );
  NAND2_X1 U4237 ( .A1(n3272), .A2(n3244), .ZN(n3287) );
  NAND2_X1 U4238 ( .A1(n3287), .A2(n4529), .ZN(n3289) );
  OAI21_X1 U4239 ( .B1(n4334), .B2(n3289), .A(n3288), .ZN(n3290) );
  NAND4_X1 U4240 ( .A1(n3292), .A2(n3277), .A3(n3291), .A4(n3290), .ZN(n3341)
         );
  NAND2_X2 U4241 ( .A1(n3340), .A2(n3341), .ZN(n3369) );
  NAND2_X1 U4242 ( .A1(n3373), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4243 ( .A1(n4124), .A2(n4491), .ZN(n3297) );
  NOR2_X2 U4244 ( .A1(n3297), .A2(n3296), .ZN(n4143) );
  NAND2_X1 U4245 ( .A1(n4279), .A2(n3300), .ZN(n4350) );
  OAI211_X1 U4246 ( .C1(n3301), .C2(n4299), .A(n4274), .B(n4350), .ZN(n3302)
         );
  NAND2_X1 U4247 ( .A1(n3302), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3305) );
  INV_X1 U4248 ( .A(n4125), .ZN(n3433) );
  NAND2_X1 U4249 ( .A1(n6460), .A2(n4775), .ZN(n3303) );
  NAND2_X1 U4250 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3375) );
  INV_X1 U4251 ( .A(n4122), .ZN(n3432) );
  INV_X1 U4252 ( .A(n3305), .ZN(n3308) );
  INV_X1 U4253 ( .A(n3306), .ZN(n3307) );
  NAND2_X1 U4254 ( .A1(n3308), .A2(n3119), .ZN(n3309) );
  XNOR2_X1 U4255 ( .A(n3369), .B(n3368), .ZN(n4370) );
  AOI22_X1 U4256 ( .A1(n3871), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4257 ( .A1(n3952), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4258 ( .A1(n3385), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4259 ( .A1(n3876), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4260 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3321)
         );
  AOI22_X1 U4261 ( .A1(n3941), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3319) );
  INV_X1 U4262 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6700) );
  AOI22_X1 U4263 ( .A1(n3916), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4264 ( .A1(n3327), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4265 ( .A1(n3944), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3316) );
  NAND4_X1 U4266 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3320)
         );
  NAND2_X1 U4267 ( .A1(n2999), .A2(n3982), .ZN(n3322) );
  OAI21_X2 U4268 ( .B1(n4370), .B2(STATE2_REG_0__SCAN_IN), .A(n3322), .ZN(
        n3339) );
  INV_X1 U4269 ( .A(n3339), .ZN(n3337) );
  INV_X1 U4270 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4891) );
  AOI22_X1 U4272 ( .A1(n3871), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4273 ( .A1(n3248), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4274 ( .A1(n3385), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4275 ( .A1(n3354), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3323) );
  NAND4_X1 U4276 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3333)
         );
  AOI22_X1 U4277 ( .A1(n3346), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4278 ( .A1(n3916), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3330) );
  BUF_X1 U4279 ( .A(n3347), .Z(n3327) );
  AOI22_X1 U4280 ( .A1(n3327), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4281 ( .A1(n3255), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3328) );
  NAND4_X1 U4282 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3332)
         );
  INV_X1 U4283 ( .A(n4048), .ZN(n3334) );
  NAND2_X1 U4284 ( .A1(n2999), .A2(n3334), .ZN(n3345) );
  NAND2_X1 U4285 ( .A1(n2998), .A2(n3982), .ZN(n3335) );
  OAI211_X1 U4286 ( .C1(n4094), .C2(n4891), .A(n3345), .B(n3335), .ZN(n3338)
         );
  INV_X1 U4287 ( .A(n3338), .ZN(n3336) );
  NAND2_X1 U4288 ( .A1(n3343), .A2(n3342), .ZN(n3344) );
  INV_X1 U4289 ( .A(n3345), .ZN(n3364) );
  NAND2_X1 U4290 ( .A1(n3044), .A2(n4048), .ZN(n3365) );
  AOI22_X1 U4292 ( .A1(n3941), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4293 ( .A1(n3327), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4294 ( .A1(n3248), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4295 ( .A1(n3944), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3350) );
  NAND4_X1 U4296 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3362)
         );
  AOI22_X1 U4297 ( .A1(n3247), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3385), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4298 ( .A1(n3354), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4299 ( .A1(n3871), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4300 ( .A1(n3916), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3357) );
  NAND4_X1 U4301 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  INV_X1 U4302 ( .A(n3983), .ZN(n3363) );
  MUX2_X1 U4303 ( .A(n3364), .B(n4045), .S(n3363), .Z(n3414) );
  INV_X1 U4304 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4901) );
  AOI21_X1 U4305 ( .B1(n4491), .B2(n3983), .A(n6493), .ZN(n3366) );
  OAI211_X1 U4306 ( .C1(n4094), .C2(n4901), .A(n3366), .B(n3365), .ZN(n3413)
         );
  INV_X1 U4307 ( .A(n3368), .ZN(n3370) );
  NAND2_X1 U4308 ( .A1(n3370), .A2(n3369), .ZN(n3372) );
  NAND2_X1 U4309 ( .A1(n3372), .A2(n3371), .ZN(n3379) );
  INV_X1 U4310 ( .A(n3375), .ZN(n3374) );
  NAND2_X1 U4311 ( .A1(n3374), .A2(n6469), .ZN(n6392) );
  NAND2_X1 U4312 ( .A1(n3375), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4313 ( .A1(n6392), .A2(n3376), .ZN(n4606) );
  NAND2_X1 U4314 ( .A1(n3433), .A2(n4606), .ZN(n3377) );
  OAI21_X1 U4315 ( .B1(n4122), .B2(n6469), .A(n3377), .ZN(n3378) );
  NAND2_X1 U4316 ( .A1(n3379), .A2(n3380), .ZN(n3383) );
  INV_X1 U4317 ( .A(n3379), .ZN(n3382) );
  NAND2_X2 U4318 ( .A1(n3382), .A2(n3381), .ZN(n4468) );
  INV_X1 U4319 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4896) );
  AOI22_X1 U4320 ( .A1(n3871), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3389) );
  INV_X2 U4321 ( .A(n3384), .ZN(n3943) );
  AOI22_X1 U4322 ( .A1(n3952), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4323 ( .A1(n3385), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4324 ( .A1(n3876), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3386) );
  NAND4_X1 U4325 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3396)
         );
  AOI22_X1 U4326 ( .A1(n3941), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4327 ( .A1(n3916), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4328 ( .A1(n3327), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4329 ( .A1(n3944), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4330 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3395)
         );
  NAND2_X1 U4331 ( .A1(n4118), .A2(n3999), .ZN(n3397) );
  OAI21_X1 U4332 ( .B1(n4094), .B2(n4896), .A(n3397), .ZN(n3398) );
  NAND2_X1 U4333 ( .A1(n3989), .A2(n3646), .ZN(n3402) );
  NAND2_X1 U4334 ( .A1(n3402), .A2(n3663), .ZN(n3426) );
  NAND2_X1 U4335 ( .A1(n3403), .A2(n3404), .ZN(n3405) );
  INV_X1 U4336 ( .A(n3646), .ZN(n3564) );
  NOR2_X1 U4337 ( .A1(n4325), .A2(n3407), .ZN(n3449) );
  INV_X1 U4338 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4437) );
  OAI22_X1 U4339 ( .A1(n3967), .A2(n4437), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6050), .ZN(n3408) );
  AOI21_X1 U4340 ( .B1(n3449), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3408), 
        .ZN(n3409) );
  NOR2_X2 U4341 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3885) );
  NAND2_X1 U4342 ( .A1(n3410), .A2(n3413), .ZN(n3412) );
  NAND2_X1 U4343 ( .A1(n3414), .A2(n3413), .ZN(n3415) );
  AOI21_X1 U4344 ( .B1(n4517), .B2(n3417), .A(n3407), .ZN(n4404) );
  INV_X1 U4345 ( .A(n3418), .ZN(n6343) );
  INV_X1 U4346 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3419) );
  INV_X1 U4347 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5105) );
  OAI22_X1 U4348 ( .A1(n3967), .A2(n3419), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5105), .ZN(n3420) );
  AOI21_X1 U4349 ( .B1(n3449), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3420), 
        .ZN(n3421) );
  OAI21_X1 U4350 ( .B1(n6343), .B2(n3564), .A(n3421), .ZN(n4403) );
  NAND2_X1 U4351 ( .A1(n3426), .A2(n3427), .ZN(n3425) );
  INV_X1 U4352 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3423) );
  OAI21_X1 U4353 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3451), .ZN(n6203) );
  AOI22_X1 U4354 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3885), 
        .B2(n6203), .ZN(n3422) );
  OAI21_X1 U4355 ( .B1(n3967), .B2(n3423), .A(n3422), .ZN(n3424) );
  INV_X1 U4356 ( .A(n3426), .ZN(n4428) );
  NAND2_X1 U4357 ( .A1(n2987), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3435) );
  NAND3_X1 U4358 ( .A1(n6391), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6349) );
  INV_X1 U4359 ( .A(n6349), .ZN(n3430) );
  NAND2_X1 U4360 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3430), .ZN(n6341) );
  NAND2_X1 U4361 ( .A1(n6391), .A2(n6341), .ZN(n3431) );
  NAND3_X1 U4362 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4695) );
  INV_X1 U4363 ( .A(n4695), .ZN(n4692) );
  NAND2_X1 U4364 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4692), .ZN(n4690) );
  AOI22_X1 U4365 ( .A1(n3433), .A2(n4879), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3432), .ZN(n3434) );
  AOI22_X1 U4366 ( .A1(n3944), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4367 ( .A1(n3941), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4368 ( .A1(n3871), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4369 ( .A1(n3952), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3436) );
  NAND4_X1 U4370 ( .A1(n3439), .A2(n3438), .A3(n3437), .A4(n3436), .ZN(n3446)
         );
  AOI22_X1 U4371 ( .A1(n3943), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3385), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4372 ( .A1(n3876), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4373 ( .A1(n3940), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4374 ( .A1(n3945), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4375 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  AOI22_X1 U4376 ( .A1(n4113), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4118), 
        .B2(n4009), .ZN(n3447) );
  XNOR2_X2 U4377 ( .A(n3458), .B(n4559), .ZN(n3998) );
  INV_X1 U4378 ( .A(n3449), .ZN(n3472) );
  INV_X1 U4379 ( .A(n3451), .ZN(n3453) );
  INV_X1 U4380 ( .A(n3470), .ZN(n3452) );
  OAI21_X1 U4381 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3453), .A(n3452), 
        .ZN(n5068) );
  AOI22_X1 U4382 ( .A1(n3885), .A2(n5068), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4383 ( .A1(n3975), .A2(EAX_REG_3__SCAN_IN), .ZN(n3454) );
  OAI211_X1 U4384 ( .C1(n3472), .C2(n3450), .A(n3455), .B(n3454), .ZN(n3456)
         );
  AOI21_X1 U4385 ( .B1(n3998), .B2(n3646), .A(n3456), .ZN(n3457) );
  INV_X1 U4386 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4906) );
  AOI22_X1 U4387 ( .A1(n3871), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4388 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3952), .B1(n3943), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4389 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3942), .B1(n3385), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4390 ( .A1(n3876), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3459) );
  NAND4_X1 U4391 ( .A1(n3462), .A2(n3461), .A3(n3460), .A4(n3459), .ZN(n3468)
         );
  AOI22_X1 U4392 ( .A1(n3941), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4393 ( .A1(n3916), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4394 ( .A1(n3327), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4395 ( .A1(n3944), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4396 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3467)
         );
  NAND2_X1 U4397 ( .A1(n4118), .A2(n4017), .ZN(n3469) );
  OAI21_X1 U4398 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3470), .A(n3504), 
        .ZN(n6193) );
  INV_X1 U4399 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U4400 ( .A1(n3975), .A2(EAX_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3407), .ZN(n3471) );
  OAI21_X1 U4401 ( .B1(n3472), .B2(n4470), .A(n3471), .ZN(n3473) );
  MUX2_X1 U4402 ( .A(n6193), .B(n3473), .S(n3964), .Z(n3474) );
  INV_X1 U4403 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U4404 ( .A1(n3950), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4405 ( .A1(n3943), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4406 ( .A1(n3944), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4407 ( .A1(n3876), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4408 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3486)
         );
  AOI22_X1 U4409 ( .A1(n3871), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4410 ( .A1(n3385), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4411 ( .A1(n3941), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4412 ( .A1(n3327), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4413 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485)
         );
  NAND2_X1 U4414 ( .A1(n4118), .A2(n4028), .ZN(n3487) );
  XNOR2_X1 U4415 ( .A(n3491), .B(n3492), .ZN(n4016) );
  NAND2_X1 U4416 ( .A1(n4016), .A2(n3646), .ZN(n3490) );
  XNOR2_X1 U4417 ( .A(n3504), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6028) );
  INV_X1 U4418 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4872) );
  OAI22_X1 U4419 ( .A1(n6028), .A2(n3964), .B1(n3663), .B2(n4872), .ZN(n3488)
         );
  AOI21_X1 U4420 ( .B1(n3975), .B2(EAX_REG_5__SCAN_IN), .A(n3488), .ZN(n3489)
         );
  NAND2_X1 U4421 ( .A1(n4507), .A2(n4510), .ZN(n4508) );
  INV_X1 U4422 ( .A(n4508), .ZN(n3510) );
  INV_X1 U4423 ( .A(n3491), .ZN(n3493) );
  AOI22_X1 U4424 ( .A1(n3871), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4425 ( .A1(n3952), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4426 ( .A1(n3951), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4427 ( .A1(n3876), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3494) );
  NAND4_X1 U4428 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3503)
         );
  AOI22_X1 U4429 ( .A1(n3941), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4430 ( .A1(n3916), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4431 ( .A1(n3327), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4432 ( .A1(n3944), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3498) );
  NAND4_X1 U4433 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3502)
         );
  AOI22_X1 U4434 ( .A1(n4113), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4118), 
        .B2(n4037), .ZN(n3512) );
  NAND2_X1 U4435 ( .A1(n3511), .A2(n3512), .ZN(n4026) );
  INV_X1 U4436 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4811) );
  NOR2_X1 U4437 ( .A1(n3505), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3506)
         );
  OR2_X1 U4438 ( .A1(n3529), .A2(n3506), .ZN(n6184) );
  AOI22_X1 U4439 ( .A1(n6184), .A2(n3885), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3507) );
  OAI21_X1 U4440 ( .B1(n3967), .B2(n4811), .A(n3507), .ZN(n3508) );
  INV_X1 U4441 ( .A(n3512), .ZN(n3513) );
  INV_X1 U4442 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4443 ( .A1(n4118), .A2(n4048), .ZN(n3514) );
  OAI21_X1 U4444 ( .B1(n4094), .B2(n3515), .A(n3514), .ZN(n3516) );
  INV_X1 U4445 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4957) );
  XNOR2_X1 U4446 ( .A(n3529), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5048) );
  AOI22_X1 U4447 ( .A1(n5048), .A2(n3885), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3517) );
  OAI21_X1 U4448 ( .B1(n3967), .B2(n4957), .A(n3517), .ZN(n3518) );
  AOI22_X1 U4449 ( .A1(n3876), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4450 ( .A1(n3943), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4451 ( .A1(n3944), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4452 ( .A1(n3916), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4453 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3528)
         );
  AOI22_X1 U4454 ( .A1(n3941), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4455 ( .A1(n3871), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4456 ( .A1(n3952), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4457 ( .A1(n3390), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3523) );
  NAND4_X1 U4458 ( .A1(n3526), .A2(n3525), .A3(n3524), .A4(n3523), .ZN(n3527)
         );
  OAI21_X1 U4459 ( .B1(n3528), .B2(n3527), .A(n3646), .ZN(n3533) );
  XNOR2_X1 U4460 ( .A(n3534), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U4461 ( .A1(n6005), .A2(n3885), .ZN(n3532) );
  NAND2_X1 U4462 ( .A1(n3975), .A2(EAX_REG_8__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4463 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3530)
         );
  NAND4_X1 U4464 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n4944)
         );
  XNOR2_X1 U4465 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3550), .ZN(n5996) );
  INV_X1 U4466 ( .A(n5996), .ZN(n3549) );
  AOI22_X1 U4467 ( .A1(n3327), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4468 ( .A1(n3952), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4469 ( .A1(n3941), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4470 ( .A1(n3876), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4471 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AOI22_X1 U4472 ( .A1(n3871), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4473 ( .A1(n3951), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4474 ( .A1(n3944), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4475 ( .A1(n3916), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4476 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  NOR2_X1 U4477 ( .A1(n3544), .A2(n3543), .ZN(n3547) );
  NAND2_X1 U4478 ( .A1(n3975), .A2(EAX_REG_9__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4479 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3545)
         );
  OAI211_X1 U4480 ( .C1(n3564), .C2(n3547), .A(n3546), .B(n3545), .ZN(n3548)
         );
  AOI21_X1 U4481 ( .B1(n3549), .B2(n3885), .A(n3548), .ZN(n5110) );
  XNOR2_X1 U4482 ( .A(n3567), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5212)
         );
  AOI22_X1 U4483 ( .A1(n3327), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4484 ( .A1(n3876), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4485 ( .A1(n3952), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4486 ( .A1(n3944), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4487 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3560)
         );
  AOI22_X1 U4488 ( .A1(n3951), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4489 ( .A1(n3941), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4490 ( .A1(n3950), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4491 ( .A1(n3871), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3555) );
  NAND4_X1 U4492 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3559)
         );
  NOR2_X1 U4493 ( .A1(n3560), .A2(n3559), .ZN(n3563) );
  NAND2_X1 U4494 ( .A1(n3975), .A2(EAX_REG_10__SCAN_IN), .ZN(n3562) );
  NAND2_X1 U4495 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3561)
         );
  OAI211_X1 U4496 ( .C1(n3564), .C2(n3563), .A(n3562), .B(n3561), .ZN(n3565)
         );
  AOI21_X1 U4497 ( .B1(n5212), .B2(n3885), .A(n3565), .ZN(n5120) );
  XNOR2_X1 U4498 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3582), .ZN(n5976)
         );
  AOI22_X1 U4499 ( .A1(n3871), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4500 ( .A1(n3248), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4501 ( .A1(n3941), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4502 ( .A1(n3950), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3568) );
  NAND4_X1 U4503 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3577)
         );
  AOI22_X1 U4504 ( .A1(n3327), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4505 ( .A1(n3940), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4506 ( .A1(n3944), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4507 ( .A1(n3876), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3572) );
  NAND4_X1 U4508 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3576)
         );
  OR2_X1 U4509 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  AOI22_X1 U4510 ( .A1(n3646), .A2(n3578), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4511 ( .A1(n3975), .A2(EAX_REG_11__SCAN_IN), .ZN(n3579) );
  OAI211_X1 U4512 ( .C1(n5976), .C2(n3964), .A(n3580), .B(n3579), .ZN(n5166)
         );
  XNOR2_X1 U4513 ( .A(n3598), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5250)
         );
  INV_X1 U4514 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3583) );
  AOI21_X1 U4515 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3583), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3585) );
  INV_X1 U4516 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U4517 ( .A1(n3967), .A2(n5229), .ZN(n3584) );
  OAI22_X1 U4518 ( .A1(n5250), .A2(n3964), .B1(n3585), .B2(n3584), .ZN(n3597)
         );
  AOI22_X1 U4519 ( .A1(n3876), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4520 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3942), .B1(n3951), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4521 ( .A1(n3916), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4522 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3940), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4523 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3595)
         );
  AOI22_X1 U4524 ( .A1(n3941), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4525 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3248), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4526 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3944), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4527 ( .A1(n3871), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3590) );
  NAND4_X1 U4528 ( .A1(n3593), .A2(n3592), .A3(n3591), .A4(n3590), .ZN(n3594)
         );
  OAI21_X1 U4529 ( .B1(n3595), .B2(n3594), .A(n3646), .ZN(n3596) );
  NAND2_X1 U4530 ( .A1(n3597), .A2(n3596), .ZN(n5217) );
  INV_X1 U4531 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5522) );
  INV_X1 U4532 ( .A(n3599), .ZN(n3601) );
  INV_X1 U4533 ( .A(n3633), .ZN(n3600) );
  OAI21_X1 U4534 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3601), .A(n3600), 
        .ZN(n5898) );
  AOI22_X1 U4535 ( .A1(n3885), .A2(n5898), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3602) );
  OAI21_X1 U4536 ( .B1(n3967), .B2(n5522), .A(n3602), .ZN(n3603) );
  INV_X1 U4537 ( .A(n3603), .ZN(n3604) );
  AOI22_X1 U4538 ( .A1(n3876), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4539 ( .A1(n3871), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4540 ( .A1(n3952), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4541 ( .A1(n3941), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3606) );
  NAND4_X1 U4542 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3615)
         );
  AOI22_X1 U4543 ( .A1(n3950), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4544 ( .A1(n3940), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4545 ( .A1(n3944), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4546 ( .A1(n3390), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3610) );
  NAND4_X1 U4547 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3614)
         );
  OR2_X1 U4548 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  NAND2_X1 U4549 ( .A1(n3646), .A2(n3616), .ZN(n5417) );
  INV_X1 U4550 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5520) );
  AOI22_X1 U4551 ( .A1(n3871), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4552 ( .A1(n3248), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4553 ( .A1(n3951), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4554 ( .A1(n3941), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4555 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3628)
         );
  AOI22_X1 U4556 ( .A1(n3950), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4557 ( .A1(n3327), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4558 ( .A1(n3876), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4559 ( .A1(n3944), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4560 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  OR2_X1 U4561 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  NAND2_X1 U4562 ( .A1(n3646), .A2(n3629), .ZN(n3632) );
  XOR2_X1 U4563 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3633), .Z(n5656) );
  INV_X1 U4564 ( .A(n5656), .ZN(n3630) );
  AOI22_X1 U4565 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3885), 
        .B2(n3630), .ZN(n3631) );
  OAI211_X1 U4566 ( .C1(n5520), .C2(n3967), .A(n3632), .B(n3631), .ZN(n5402)
         );
  INV_X1 U4567 ( .A(EAX_REG_15__SCAN_IN), .ZN(n3636) );
  INV_X1 U4568 ( .A(n3651), .ZN(n3634) );
  XNOR2_X1 U4569 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3634), .ZN(n5643)
         );
  AOI22_X1 U4570 ( .A1(n3885), .A2(n5643), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3635) );
  OAI21_X1 U4571 ( .B1(n3967), .B2(n3636), .A(n3635), .ZN(n3637) );
  INV_X1 U4572 ( .A(n3637), .ZN(n3650) );
  AOI22_X1 U4573 ( .A1(n3941), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4574 ( .A1(n3871), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4575 ( .A1(n3952), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4576 ( .A1(n3327), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4577 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3648)
         );
  AOI22_X1 U4578 ( .A1(n3951), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4579 ( .A1(n3916), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4580 ( .A1(n3876), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4581 ( .A1(n3944), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4582 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3647)
         );
  OAI21_X1 U4583 ( .B1(n3648), .B2(n3647), .A(n3646), .ZN(n3649) );
  XOR2_X1 U4584 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3668), .Z(n5636) );
  NAND2_X1 U4585 ( .A1(n3244), .A2(n5258), .ZN(n3652) );
  AOI22_X1 U4586 ( .A1(n3950), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4587 ( .A1(n3871), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4588 ( .A1(n3944), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4589 ( .A1(n3876), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4590 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3662)
         );
  AOI22_X1 U4591 ( .A1(n3952), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4592 ( .A1(n3951), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4593 ( .A1(n3941), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4594 ( .A1(n3327), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3657) );
  NAND4_X1 U4595 ( .A1(n3660), .A2(n3659), .A3(n3658), .A4(n3657), .ZN(n3661)
         );
  OR2_X1 U4596 ( .A1(n3662), .A2(n3661), .ZN(n3666) );
  INV_X1 U4597 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3664) );
  INV_X1 U4598 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5632) );
  OAI22_X1 U4599 ( .A1(n3967), .A2(n3664), .B1(n3663), .B2(n5632), .ZN(n3665)
         );
  AOI21_X1 U4600 ( .B1(n3927), .B2(n3666), .A(n3665), .ZN(n3667) );
  OAI21_X1 U4601 ( .B1(n5636), .B2(n3964), .A(n3667), .ZN(n5377) );
  XNOR2_X1 U4602 ( .A(n3702), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5620)
         );
  NAND2_X1 U4603 ( .A1(n5620), .A2(n3885), .ZN(n3684) );
  AOI22_X1 U4604 ( .A1(n3346), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4605 ( .A1(n3950), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4606 ( .A1(n3943), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4607 ( .A1(n3952), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4608 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3680)
         );
  AOI22_X1 U4609 ( .A1(n3327), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4610 ( .A1(n3871), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4611 ( .A1(n3951), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3674)
         );
  NAND2_X1 U4612 ( .A1(n3916), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3673) );
  AND3_X1 U4613 ( .A1(n3674), .A2(n3673), .A3(n3964), .ZN(n3676) );
  AOI22_X1 U4614 ( .A1(n3944), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4615 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3679)
         );
  INV_X1 U4616 ( .A(n3927), .ZN(n3970) );
  NAND2_X1 U4617 ( .A1(n3970), .A2(n3964), .ZN(n3751) );
  OAI21_X1 U4618 ( .B1(n3680), .B2(n3679), .A(n3751), .ZN(n3682) );
  AOI22_X1 U4619 ( .A1(n3975), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3407), .ZN(n3681) );
  NAND2_X1 U4620 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  NAND2_X1 U4621 ( .A1(n3684), .A2(n3683), .ZN(n5363) );
  AOI22_X1 U4622 ( .A1(n3876), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4623 ( .A1(n3871), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4624 ( .A1(n3952), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4625 ( .A1(n3944), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4626 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3696)
         );
  AOI22_X1 U4627 ( .A1(n3941), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3327), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4628 ( .A1(n3940), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4629 ( .A1(n3916), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4630 ( .A1(n3390), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4631 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3695)
         );
  NOR2_X1 U4632 ( .A1(n3696), .A2(n3695), .ZN(n3701) );
  INV_X1 U4633 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4634 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3697)
         );
  OAI211_X1 U4635 ( .C1(n3967), .C2(n3698), .A(n3964), .B(n3697), .ZN(n3699)
         );
  INV_X1 U4636 ( .A(n3699), .ZN(n3700) );
  OAI21_X1 U4637 ( .B1(n3970), .B2(n3701), .A(n3700), .ZN(n3705) );
  OAI21_X1 U4638 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3703), .A(n3723), 
        .ZN(n5969) );
  OR2_X1 U4639 ( .A1(n3964), .A2(n5969), .ZN(n3704) );
  NAND2_X1 U4640 ( .A1(n3705), .A2(n3704), .ZN(n5484) );
  AOI22_X1 U4641 ( .A1(n3943), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4642 ( .A1(n3951), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4643 ( .A1(n3942), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4644 ( .A1(n3876), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4645 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3718)
         );
  AOI22_X1 U4646 ( .A1(n3347), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U4647 ( .A1(n3248), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4648 ( .A1(n3346), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3711)
         );
  AND3_X1 U4649 ( .A1(n3712), .A2(n3711), .A3(n3964), .ZN(n3715) );
  AOI22_X1 U4650 ( .A1(n3871), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4651 ( .A1(n3348), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4652 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  OAI21_X1 U4653 ( .B1(n3718), .B2(n3717), .A(n3751), .ZN(n3720) );
  AOI22_X1 U4654 ( .A1(n3975), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3407), .ZN(n3719) );
  NAND2_X1 U4655 ( .A1(n3720), .A2(n3719), .ZN(n3722) );
  XNOR2_X1 U4656 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3723), .ZN(n5861)
         );
  NAND2_X1 U4657 ( .A1(n5861), .A2(n3885), .ZN(n3721) );
  NAND2_X1 U4658 ( .A1(n3722), .A2(n3721), .ZN(n5475) );
  INV_X1 U4659 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5863) );
  OR2_X1 U4660 ( .A1(n3724), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3725)
         );
  NAND2_X1 U4661 ( .A1(n3725), .A2(n3775), .ZN(n5855) );
  AOI22_X1 U4662 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3943), .B1(n3348), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4663 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3952), .B1(n3942), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4664 ( .A1(n3944), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4665 ( .A1(n3346), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3726) );
  NAND4_X1 U4666 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3735)
         );
  AOI22_X1 U4667 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3916), .B1(n3950), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4668 ( .A1(n3871), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4669 ( .A1(n3347), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4670 ( .A1(n3876), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3730) );
  NAND4_X1 U4671 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3734)
         );
  OAI21_X1 U4672 ( .B1(n3735), .B2(n3734), .A(n3927), .ZN(n3738) );
  NAND2_X1 U4673 ( .A1(n3975), .A2(EAX_REG_20__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4674 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3736)
         );
  NAND4_X1 U4675 ( .A1(n3738), .A2(n3964), .A3(n3737), .A4(n3736), .ZN(n3739)
         );
  OAI21_X1 U4676 ( .B1(n5855), .B2(n3964), .A(n3739), .ZN(n5469) );
  INV_X1 U4677 ( .A(n5469), .ZN(n3740) );
  AOI22_X1 U4678 ( .A1(n3952), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4679 ( .A1(n3940), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4680 ( .A1(n3871), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4681 ( .A1(n3942), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4682 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3753)
         );
  AOI22_X1 U4683 ( .A1(n3944), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4684 ( .A1(n3354), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3749) );
  NAND2_X1 U4685 ( .A1(n3346), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3746)
         );
  NAND2_X1 U4686 ( .A1(n3943), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3745)
         );
  AND3_X1 U4687 ( .A1(n3746), .A2(n3745), .A3(n3964), .ZN(n3748) );
  AOI22_X1 U4688 ( .A1(n3440), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4689 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3752)
         );
  OAI21_X1 U4690 ( .B1(n3753), .B2(n3752), .A(n3751), .ZN(n3756) );
  NAND2_X1 U4691 ( .A1(n3975), .A2(EAX_REG_21__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4692 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3754)
         );
  NAND3_X1 U4693 ( .A1(n3756), .A2(n3755), .A3(n3754), .ZN(n3758) );
  XNOR2_X1 U4694 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3775), .ZN(n5843)
         );
  NAND2_X1 U4695 ( .A1(n5843), .A2(n3885), .ZN(n3757) );
  NAND2_X1 U4696 ( .A1(n3758), .A2(n3757), .ZN(n5459) );
  AOI22_X1 U4697 ( .A1(n3346), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4698 ( .A1(n3952), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4699 ( .A1(n3944), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4700 ( .A1(n3354), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4701 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3769)
         );
  AOI22_X1 U4702 ( .A1(n3871), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4703 ( .A1(n3943), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4704 ( .A1(n3916), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4705 ( .A1(n3347), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4706 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  NOR2_X1 U4707 ( .A1(n3769), .A2(n3768), .ZN(n3774) );
  INV_X1 U4708 ( .A(EAX_REG_22__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4709 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3770)
         );
  OAI211_X1 U4710 ( .C1(n3967), .C2(n3771), .A(n3964), .B(n3770), .ZN(n3772)
         );
  INV_X1 U4711 ( .A(n3772), .ZN(n3773) );
  OAI21_X1 U4712 ( .B1(n3970), .B2(n3774), .A(n3773), .ZN(n3779) );
  OAI21_X1 U4713 ( .B1(n3777), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3821), 
        .ZN(n5593) );
  OR2_X1 U4714 ( .A1(n5593), .A2(n3964), .ZN(n3778) );
  NAND2_X1 U4715 ( .A1(n3779), .A2(n3778), .ZN(n5345) );
  AOI22_X1 U4716 ( .A1(n3943), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4717 ( .A1(n3951), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4718 ( .A1(n3941), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4719 ( .A1(n3871), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4720 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4721 ( .A1(n3876), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4722 ( .A1(n3327), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4723 ( .A1(n3944), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4724 ( .A1(n3916), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4725 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  NOR2_X1 U4726 ( .A1(n3789), .A2(n3788), .ZN(n3807) );
  AOI22_X1 U4727 ( .A1(n3327), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4728 ( .A1(n3943), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4729 ( .A1(n3916), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4730 ( .A1(n3876), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4731 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3799)
         );
  AOI22_X1 U4732 ( .A1(n3871), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4733 ( .A1(n3952), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4734 ( .A1(n3944), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4735 ( .A1(n3941), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4736 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3798)
         );
  NOR2_X1 U4737 ( .A1(n3799), .A2(n3798), .ZN(n3808) );
  XOR2_X1 U4738 ( .A(n3807), .B(n3808), .Z(n3800) );
  NAND2_X1 U4739 ( .A1(n3800), .A2(n3927), .ZN(n3806) );
  INV_X1 U4740 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3802) );
  NAND2_X1 U4741 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3801)
         );
  OAI211_X1 U4742 ( .C1(n3967), .C2(n3802), .A(n3964), .B(n3801), .ZN(n3803)
         );
  INV_X1 U4743 ( .A(n3803), .ZN(n3805) );
  XNOR2_X1 U4744 ( .A(n3821), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5337)
         );
  AOI21_X1 U4745 ( .B1(n3806), .B2(n3805), .A(n3804), .ZN(n5332) );
  NOR2_X1 U4746 ( .A1(n3808), .A2(n3807), .ZN(n3838) );
  AOI22_X1 U4747 ( .A1(n3871), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4748 ( .A1(n3952), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4749 ( .A1(n3951), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4750 ( .A1(n3876), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4751 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3818)
         );
  AOI22_X1 U4752 ( .A1(n3346), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4753 ( .A1(n3916), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4754 ( .A1(n3347), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4755 ( .A1(n3944), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3813) );
  NAND4_X1 U4756 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3817)
         );
  OR2_X1 U4757 ( .A1(n3818), .A2(n3817), .ZN(n3837) );
  INV_X1 U4758 ( .A(n3837), .ZN(n3819) );
  XNOR2_X1 U4759 ( .A(n3838), .B(n3819), .ZN(n3820) );
  NAND2_X1 U4760 ( .A1(n3820), .A2(n3927), .ZN(n3826) );
  INV_X1 U4761 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3823) );
  INV_X1 U4762 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5336) );
  XNOR2_X1 U4763 ( .A(n3843), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5578)
         );
  AOI22_X1 U4764 ( .A1(n5578), .A2(n3885), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3822) );
  OAI21_X1 U4765 ( .B1(n3967), .B2(n3823), .A(n3822), .ZN(n3824) );
  INV_X1 U4766 ( .A(n3824), .ZN(n3825) );
  NAND2_X1 U4767 ( .A1(n3826), .A2(n3825), .ZN(n5322) );
  AOI22_X1 U4768 ( .A1(n3941), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4769 ( .A1(n3916), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4770 ( .A1(n3327), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4771 ( .A1(n3944), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3827) );
  NAND4_X1 U4772 ( .A1(n3830), .A2(n3829), .A3(n3828), .A4(n3827), .ZN(n3836)
         );
  AOI22_X1 U4773 ( .A1(n3871), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4774 ( .A1(n3952), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4775 ( .A1(n3951), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4776 ( .A1(n3354), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4777 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3835)
         );
  NOR2_X1 U4778 ( .A1(n3836), .A2(n3835), .ZN(n3851) );
  NAND2_X1 U4779 ( .A1(n3838), .A2(n3837), .ZN(n3850) );
  XOR2_X1 U4780 ( .A(n3851), .B(n3850), .Z(n3839) );
  NAND2_X1 U4781 ( .A1(n3839), .A2(n3927), .ZN(n3842) );
  INV_X1 U4782 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6704) );
  OAI21_X1 U4783 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6704), .A(n3964), .ZN(
        n3840) );
  AOI21_X1 U4784 ( .B1(n3975), .B2(EAX_REG_25__SCAN_IN), .A(n3840), .ZN(n3841)
         );
  NAND2_X1 U4785 ( .A1(n3842), .A2(n3841), .ZN(n3847) );
  NOR2_X1 U4786 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n3844), .ZN(n3845)
         );
  NOR2_X1 U4787 ( .A1(n3866), .A2(n3845), .ZN(n5833) );
  NAND2_X1 U4788 ( .A1(n5833), .A2(n3885), .ZN(n3846) );
  NAND2_X1 U4789 ( .A1(n3847), .A2(n3846), .ZN(n5444) );
  NOR2_X1 U4790 ( .A1(n3851), .A2(n3850), .ZN(n3870) );
  AOI22_X1 U4791 ( .A1(n3871), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4792 ( .A1(n3952), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4793 ( .A1(n3951), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4794 ( .A1(n3876), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4795 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3861)
         );
  AOI22_X1 U4796 ( .A1(n3346), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4797 ( .A1(n3916), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4798 ( .A1(n3347), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4799 ( .A1(n3944), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4800 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3860)
         );
  OR2_X1 U4801 ( .A1(n3861), .A2(n3860), .ZN(n3869) );
  INV_X1 U4802 ( .A(n3869), .ZN(n3862) );
  XNOR2_X1 U4803 ( .A(n3870), .B(n3862), .ZN(n3865) );
  NAND2_X1 U4804 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3863)
         );
  OAI211_X1 U4805 ( .C1(n3967), .C2(n6706), .A(n3964), .B(n3863), .ZN(n3864)
         );
  AOI21_X1 U4806 ( .B1(n3865), .B2(n3927), .A(n3864), .ZN(n3868) );
  OAI21_X1 U4807 ( .B1(n3866), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n3906), 
        .ZN(n5823) );
  NOR2_X1 U4808 ( .A1(n5823), .A2(n3964), .ZN(n3867) );
  NAND2_X1 U4809 ( .A1(n3870), .A2(n3869), .ZN(n3889) );
  AOI22_X1 U4810 ( .A1(n3941), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4811 ( .A1(n3327), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4812 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3952), .B1(n3871), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4813 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3951), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4814 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3882)
         );
  AOI22_X1 U4815 ( .A1(n3943), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4816 ( .A1(n3945), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4817 ( .A1(n3876), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4818 ( .A1(n3944), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4819 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  NOR2_X1 U4820 ( .A1(n3882), .A2(n3881), .ZN(n3890) );
  XOR2_X1 U4821 ( .A(n3889), .B(n3890), .Z(n3883) );
  NAND2_X1 U4822 ( .A1(n3883), .A2(n3927), .ZN(n3888) );
  INV_X1 U4823 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5552) );
  OAI21_X1 U4824 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5552), .A(n3964), .ZN(
        n3884) );
  AOI21_X1 U4825 ( .B1(n3975), .B2(EAX_REG_27__SCAN_IN), .A(n3884), .ZN(n3887)
         );
  XNOR2_X1 U4826 ( .A(n3906), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5815)
         );
  AOI21_X1 U4827 ( .B1(n3888), .B2(n3887), .A(n3886), .ZN(n5257) );
  NOR2_X1 U4828 ( .A1(n3890), .A2(n3889), .ZN(n3915) );
  AOI22_X1 U4829 ( .A1(n3871), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4830 ( .A1(n3952), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4831 ( .A1(n3951), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4832 ( .A1(n3354), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4833 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3900)
         );
  AOI22_X1 U4834 ( .A1(n3346), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4835 ( .A1(n3916), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4836 ( .A1(n3347), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4837 ( .A1(n3944), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3895) );
  NAND4_X1 U4838 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3899)
         );
  OR2_X1 U4839 ( .A1(n3900), .A2(n3899), .ZN(n3914) );
  INV_X1 U4840 ( .A(n3914), .ZN(n3901) );
  XNOR2_X1 U4841 ( .A(n3915), .B(n3901), .ZN(n3902) );
  NAND2_X1 U4842 ( .A1(n3902), .A2(n3927), .ZN(n3913) );
  INV_X1 U4843 ( .A(EAX_REG_28__SCAN_IN), .ZN(n3904) );
  NAND2_X1 U4844 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3903)
         );
  OAI211_X1 U4845 ( .C1(n3967), .C2(n3904), .A(n3964), .B(n3903), .ZN(n3905)
         );
  INV_X1 U4846 ( .A(n3905), .ZN(n3912) );
  NAND2_X1 U4847 ( .A1(n3907), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3935)
         );
  INV_X1 U4848 ( .A(n3907), .ZN(n3909) );
  INV_X1 U4849 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3908) );
  NAND2_X1 U4850 ( .A1(n3909), .A2(n3908), .ZN(n3910) );
  NAND2_X1 U4851 ( .A1(n3935), .A2(n3910), .ZN(n5545) );
  NOR2_X1 U4852 ( .A1(n5545), .A2(n3964), .ZN(n3911) );
  NAND2_X1 U4853 ( .A1(n3915), .A2(n3914), .ZN(n3960) );
  AOI22_X1 U4854 ( .A1(n3944), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4855 ( .A1(n3941), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4856 ( .A1(n3354), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4857 ( .A1(n3942), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4858 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3926)
         );
  AOI22_X1 U4859 ( .A1(n3943), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4860 ( .A1(n3952), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4861 ( .A1(n3945), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4862 ( .A1(n3871), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4863 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  NOR2_X1 U4864 ( .A1(n3926), .A2(n3925), .ZN(n3961) );
  XOR2_X1 U4865 ( .A(n3960), .B(n3961), .Z(n3928) );
  NAND2_X1 U4866 ( .A1(n3928), .A2(n3927), .ZN(n3933) );
  INV_X1 U4867 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3930) );
  NAND2_X1 U4868 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3929)
         );
  OAI211_X1 U4869 ( .C1(n3967), .C2(n3930), .A(n3964), .B(n3929), .ZN(n3931)
         );
  INV_X1 U4870 ( .A(n3931), .ZN(n3932) );
  NAND2_X1 U4871 ( .A1(n3933), .A2(n3932), .ZN(n3938) );
  INV_X1 U4872 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U4873 ( .A1(n3935), .A2(n3934), .ZN(n3936) );
  NAND2_X1 U4874 ( .A1(n5534), .A2(n3885), .ZN(n3937) );
  NAND2_X1 U4875 ( .A1(n3938), .A2(n3937), .ZN(n5298) );
  AOI22_X1 U4876 ( .A1(n3941), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4877 ( .A1(n3943), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4878 ( .A1(n3944), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4879 ( .A1(n3916), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4880 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3959)
         );
  AOI22_X1 U4881 ( .A1(n3327), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4882 ( .A1(n3952), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4883 ( .A1(n3354), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4884 ( .A1(n3871), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4885 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3958)
         );
  NOR2_X1 U4886 ( .A1(n3959), .A2(n3958), .ZN(n3963) );
  NOR2_X1 U4887 ( .A1(n3961), .A2(n3960), .ZN(n3962) );
  XOR2_X1 U4888 ( .A(n3963), .B(n3962), .Z(n3971) );
  INV_X1 U4889 ( .A(EAX_REG_30__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4890 ( .A1(n3407), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3965)
         );
  OAI211_X1 U4891 ( .C1(n3967), .C2(n3966), .A(n3965), .B(n3964), .ZN(n3968)
         );
  INV_X1 U4892 ( .A(n3968), .ZN(n3969) );
  OAI21_X1 U4893 ( .B1(n3971), .B2(n3970), .A(n3969), .ZN(n3973) );
  XNOR2_X1 U4894 ( .A(n4129), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5287)
         );
  NAND2_X1 U4895 ( .A1(n5287), .A2(n3885), .ZN(n3972) );
  NAND2_X1 U4896 ( .A1(n3973), .A2(n3972), .ZN(n5275) );
  AOI22_X1 U4897 ( .A1(n3975), .A2(EAX_REG_31__SCAN_IN), .B1(n3974), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3976) );
  NAND3_X1 U4898 ( .A1(n6493), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U4899 ( .A1(n4285), .A2(n5894), .ZN(n4136) );
  INV_X1 U4900 ( .A(n3281), .ZN(n6614) );
  NAND2_X1 U4901 ( .A1(n4491), .A2(n4529), .ZN(n3990) );
  OAI21_X1 U4902 ( .B1(n6614), .B2(n3983), .A(n3990), .ZN(n3977) );
  INV_X1 U4903 ( .A(n3977), .ZN(n3978) );
  NAND2_X1 U4904 ( .A1(n4311), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3979)
         );
  INV_X1 U4905 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U4906 ( .A1(n3979), .A2(n4673), .ZN(n3981) );
  AND2_X1 U4907 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3980) );
  NAND2_X1 U4908 ( .A1(n4311), .A2(n3980), .ZN(n3987) );
  AND2_X1 U4909 ( .A1(n3981), .A2(n3987), .ZN(n4480) );
  NAND2_X1 U4910 ( .A1(n3982), .A2(n3983), .ZN(n4001) );
  OAI21_X1 U4911 ( .B1(n3983), .B2(n3982), .A(n4001), .ZN(n3984) );
  OAI211_X1 U4912 ( .C1(n3984), .C2(n6614), .A(n4338), .B(n3263), .ZN(n3985)
         );
  INV_X1 U4913 ( .A(n3985), .ZN(n3986) );
  NAND2_X1 U4914 ( .A1(n4480), .A2(n4481), .ZN(n3988) );
  NAND2_X1 U4915 ( .A1(n6197), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3993)
         );
  XNOR2_X1 U4916 ( .A(n4001), .B(n3999), .ZN(n3991) );
  OAI21_X1 U4917 ( .B1(n3991), .B2(n6614), .A(n3990), .ZN(n3992) );
  NAND2_X1 U4918 ( .A1(n3993), .A2(n6196), .ZN(n3997) );
  INV_X1 U4919 ( .A(n6197), .ZN(n3995) );
  INV_X1 U4920 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4921 ( .A1(n3995), .A2(n3994), .ZN(n3996) );
  AND2_X1 U4922 ( .A1(n3997), .A2(n3996), .ZN(n4738) );
  NAND2_X1 U4923 ( .A1(n3998), .A2(n4085), .ZN(n4005) );
  INV_X1 U4924 ( .A(n3999), .ZN(n4000) );
  NAND2_X1 U4925 ( .A1(n4001), .A2(n4000), .ZN(n4010) );
  INV_X1 U4926 ( .A(n4009), .ZN(n4002) );
  XNOR2_X1 U4927 ( .A(n4010), .B(n4002), .ZN(n4003) );
  NAND2_X1 U4928 ( .A1(n4003), .A2(n3281), .ZN(n4004) );
  INV_X1 U4929 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U4930 ( .A1(n4738), .A2(n4737), .ZN(n4739) );
  NAND2_X1 U4931 ( .A1(n4006), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4007)
         );
  NAND2_X1 U4932 ( .A1(n4739), .A2(n4007), .ZN(n6187) );
  NAND2_X1 U4933 ( .A1(n4008), .A2(n4085), .ZN(n4013) );
  NAND2_X1 U4934 ( .A1(n4010), .A2(n4009), .ZN(n4019) );
  XNOR2_X1 U4935 ( .A(n4019), .B(n4017), .ZN(n4011) );
  NAND2_X1 U4936 ( .A1(n4011), .A2(n3281), .ZN(n4012) );
  NAND2_X1 U4937 ( .A1(n4013), .A2(n4012), .ZN(n4014) );
  INV_X1 U4938 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6271) );
  XNOR2_X1 U4939 ( .A(n4014), .B(n6271), .ZN(n6186) );
  NAND2_X1 U4940 ( .A1(n6187), .A2(n6186), .ZN(n6185) );
  NAND2_X1 U4941 ( .A1(n4014), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4015)
         );
  NAND2_X1 U4942 ( .A1(n6185), .A2(n4015), .ZN(n4871) );
  NAND2_X1 U4943 ( .A1(n4016), .A2(n4085), .ZN(n4022) );
  INV_X1 U4944 ( .A(n4017), .ZN(n4018) );
  OR2_X1 U4945 ( .A1(n4019), .A2(n4018), .ZN(n4027) );
  XNOR2_X1 U4946 ( .A(n4027), .B(n4028), .ZN(n4020) );
  NAND2_X1 U4947 ( .A1(n4020), .A2(n3281), .ZN(n4021) );
  NAND2_X1 U4948 ( .A1(n4022), .A2(n4021), .ZN(n4024) );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4023) );
  XNOR2_X1 U4950 ( .A(n4024), .B(n4023), .ZN(n4870) );
  NAND2_X1 U4951 ( .A1(n4871), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U4952 ( .A1(n4024), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4025)
         );
  NAND3_X1 U4953 ( .A1(n4047), .A2(n4085), .A3(n4026), .ZN(n4032) );
  INV_X1 U4954 ( .A(n4027), .ZN(n4029) );
  NAND2_X1 U4955 ( .A1(n4029), .A2(n4028), .ZN(n4036) );
  XNOR2_X1 U4956 ( .A(n4036), .B(n4037), .ZN(n4030) );
  NAND2_X1 U4957 ( .A1(n4030), .A2(n3281), .ZN(n4031) );
  NAND2_X1 U4958 ( .A1(n4032), .A2(n4031), .ZN(n4033) );
  INV_X1 U4959 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6218) );
  XNOR2_X1 U4960 ( .A(n4033), .B(n6218), .ZN(n4669) );
  NAND2_X1 U4961 ( .A1(n4033), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4034)
         );
  NAND2_X1 U4962 ( .A1(n4035), .A2(n4085), .ZN(n4041) );
  INV_X1 U4963 ( .A(n4036), .ZN(n4038) );
  NAND2_X1 U4964 ( .A1(n4038), .A2(n4037), .ZN(n4050) );
  XNOR2_X1 U4965 ( .A(n4050), .B(n4048), .ZN(n4039) );
  NAND2_X1 U4966 ( .A1(n4039), .A2(n3281), .ZN(n4040) );
  NAND2_X1 U4967 ( .A1(n4041), .A2(n4040), .ZN(n4043) );
  INV_X1 U4968 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4042) );
  XNOR2_X1 U4969 ( .A(n4043), .B(n4042), .ZN(n4951) );
  NAND2_X1 U4970 ( .A1(n4043), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4044)
         );
  NOR2_X1 U4971 ( .A1(n3029), .A2(n4104), .ZN(n4046) );
  NAND2_X1 U4972 ( .A1(n3281), .A2(n4048), .ZN(n4049) );
  OR2_X1 U4973 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NAND2_X1 U4974 ( .A1(n6169), .A2(n4051), .ZN(n4052) );
  INV_X1 U4975 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4185) );
  XNOR2_X1 U4976 ( .A(n4052), .B(n4185), .ZN(n5074) );
  NAND2_X1 U4977 ( .A1(n4052), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4053)
         );
  INV_X4 U4978 ( .A(n3004), .ZN(n6169) );
  INV_X1 U4979 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U4980 ( .A1(n6169), .A2(n6236), .ZN(n5114) );
  OR2_X1 U4981 ( .A1(n6169), .A2(n6236), .ZN(n5115) );
  INV_X1 U4982 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4054) );
  NAND2_X1 U4983 ( .A1(n6169), .A2(n4054), .ZN(n5208) );
  AND2_X1 U4984 ( .A1(n6169), .A2(n6214), .ZN(n4058) );
  INV_X1 U4985 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5242) );
  NOR2_X1 U4986 ( .A1(n6169), .A2(n5242), .ZN(n5233) );
  NAND2_X1 U4987 ( .A1(n6169), .A2(n5242), .ZN(n5231) );
  XNOR2_X1 U4988 ( .A(n6169), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5893)
         );
  NAND2_X1 U4989 ( .A1(n6169), .A2(n5792), .ZN(n4059) );
  INV_X1 U4990 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5920) );
  INV_X1 U4991 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U4992 ( .A1(n6169), .A2(n5928), .ZN(n4061) );
  INV_X1 U4993 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U4994 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5771) );
  INV_X1 U4995 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5910) );
  INV_X1 U4996 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5900) );
  AND3_X1 U4997 ( .A1(n5910), .A2(n5900), .A3(n5921), .ZN(n4062) );
  NOR2_X1 U4998 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5738) );
  INV_X1 U4999 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5774) );
  INV_X1 U5000 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6716) );
  INV_X1 U5001 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5756) );
  NAND4_X1 U5002 ( .A1(n5738), .A2(n5774), .A3(n6716), .A4(n5756), .ZN(n4065)
         );
  AND2_X1 U5003 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5773) );
  AND2_X1 U5004 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U5005 ( .A1(n5773), .A2(n5659), .ZN(n5736) );
  NAND2_X1 U5006 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5669) );
  NOR2_X1 U5007 ( .A1(n5736), .A2(n5669), .ZN(n5673) );
  NAND2_X1 U5008 ( .A1(n5610), .A2(n5673), .ZN(n4066) );
  XOR2_X1 U5009 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n6169), .Z(n5564) );
  INV_X1 U5010 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5732) );
  INV_X1 U5011 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5541) );
  NOR2_X1 U5012 ( .A1(n3004), .A2(n5541), .ZN(n5557) );
  NAND2_X1 U5013 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5707) );
  INV_X1 U5014 ( .A(n5563), .ZN(n4070) );
  NOR2_X1 U5015 ( .A1(n6169), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5556)
         );
  NOR2_X1 U5016 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5706) );
  INV_X1 U5017 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5686) );
  INV_X1 U5018 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5683) );
  NAND4_X1 U5019 ( .A1(n5556), .A2(n5706), .A3(n5686), .A4(n5683), .ZN(n4069)
         );
  NAND2_X1 U5020 ( .A1(n4071), .A2(n3109), .ZN(n4072) );
  AND2_X1 U5021 ( .A1(n3298), .A2(n3263), .ZN(n4073) );
  NAND2_X1 U5022 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6460), .ZN(n4080) );
  OAI21_X1 U5023 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6460), .A(n4080), 
        .ZN(n4081) );
  OAI21_X1 U5024 ( .B1(n3242), .B2(n4081), .A(n4074), .ZN(n4075) );
  NAND2_X1 U5025 ( .A1(n4106), .A2(n4075), .ZN(n4083) );
  INV_X1 U5026 ( .A(n4083), .ZN(n4087) );
  NAND2_X1 U5027 ( .A1(n4775), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U5028 ( .A1(n4076), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U5029 ( .A1(n4091), .A2(n4077), .ZN(n4079) );
  INV_X1 U5030 ( .A(n4092), .ZN(n4078) );
  AOI21_X1 U5031 ( .B1(n4080), .B2(n4079), .A(n4078), .ZN(n4138) );
  INV_X1 U5032 ( .A(n4118), .ZN(n4082) );
  NOR2_X1 U5033 ( .A1(n4082), .A2(n4081), .ZN(n4084) );
  OAI211_X1 U5034 ( .C1(n4088), .C2(n4138), .A(n4084), .B(n4083), .ZN(n4086)
         );
  AOI22_X1 U5035 ( .A1(n4087), .A2(n4138), .B1(n4086), .B2(n4119), .ZN(n4097)
         );
  INV_X1 U5036 ( .A(n4088), .ZN(n4090) );
  INV_X1 U5037 ( .A(n4138), .ZN(n4089) );
  NOR3_X1 U5038 ( .A1(n4090), .A2(n6493), .A3(n4089), .ZN(n4096) );
  NAND2_X1 U5039 ( .A1(n4092), .A2(n4091), .ZN(n4101) );
  NAND2_X1 U5040 ( .A1(n4395), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4093) );
  NAND2_X1 U5041 ( .A1(n4102), .A2(n4093), .ZN(n4099) );
  XNOR2_X1 U5042 ( .A(n4101), .B(n4099), .ZN(n4139) );
  NAND2_X1 U5043 ( .A1(n4118), .A2(n4139), .ZN(n4105) );
  OAI211_X1 U5044 ( .C1(n4094), .C2(n4139), .A(n4106), .B(n4105), .ZN(n4095)
         );
  OAI21_X1 U5045 ( .B1(n4097), .B2(n4096), .A(n4095), .ZN(n4098) );
  INV_X1 U5046 ( .A(n4098), .ZN(n4108) );
  INV_X1 U5047 ( .A(n4099), .ZN(n4100) );
  NAND2_X1 U5048 ( .A1(n4101), .A2(n4100), .ZN(n4103) );
  XNOR2_X1 U5049 ( .A(n3450), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4110)
         );
  XNOR2_X1 U5050 ( .A(n4109), .B(n4110), .ZN(n4140) );
  OAI22_X1 U5051 ( .A1(n4106), .A2(n4105), .B1(n4140), .B2(n4104), .ZN(n4107)
         );
  NAND3_X1 U5052 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4117), .A3(n4470), .ZN(n4137) );
  NOR2_X1 U5053 ( .A1(n4137), .A2(n4113), .ZN(n4114) );
  INV_X1 U5054 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6297) );
  NOR2_X1 U5055 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6297), .ZN(n4116)
         );
  INV_X1 U5056 ( .A(n4119), .ZN(n4120) );
  NAND2_X1 U5057 ( .A1(n4142), .A2(n4120), .ZN(n4121) );
  NAND2_X1 U5058 ( .A1(n4122), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U5059 ( .A1(n4123), .A2(n4124), .ZN(n6476) );
  NAND2_X1 U5060 ( .A1(n4125), .A2(n6400), .ZN(n6611) );
  NAND2_X1 U5061 ( .A1(n6611), .A2(n6493), .ZN(n4126) );
  AND2_X2 U5062 ( .A1(n6178), .A2(n4126), .ZN(n6194) );
  NAND2_X1 U5063 ( .A1(n6493), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4128) );
  INV_X1 U5064 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5002) );
  NAND2_X1 U5065 ( .A1(n5002), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4127) );
  AND2_X1 U5066 ( .A1(n4128), .A2(n4127), .ZN(n4407) );
  INV_X1 U5067 ( .A(n4129), .ZN(n4130) );
  NAND2_X1 U5068 ( .A1(n4130), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4132)
         );
  INV_X1 U5069 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4131) );
  NAND2_X1 U5070 ( .A1(n6493), .A2(n3407), .ZN(n6509) );
  INV_X1 U5071 ( .A(n6509), .ZN(n6502) );
  AND2_X1 U5072 ( .A1(n6206), .A2(REIP_REG_31__SCAN_IN), .ZN(n5676) );
  AOI21_X1 U5073 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5676), 
        .ZN(n4133) );
  OAI21_X1 U5074 ( .B1(n6204), .B2(n5034), .A(n4133), .ZN(n4134) );
  INV_X1 U5075 ( .A(n4134), .ZN(n4135) );
  AND4_X1 U5076 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4141)
         );
  NOR2_X1 U5077 ( .A1(n4142), .A2(n4141), .ZN(n4297) );
  NAND2_X1 U5078 ( .A1(n4297), .A2(n4143), .ZN(n4291) );
  NAND2_X1 U5079 ( .A1(n3407), .A2(n6501), .ZN(n6508) );
  NOR3_X1 U5080 ( .A1(n6493), .A2(n6591), .A3(n6508), .ZN(n6484) );
  NOR3_X1 U5081 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6509), .A3(n6501), .ZN(
        n6504) );
  NOR2_X1 U5082 ( .A1(n5034), .A2(n6501), .ZN(n4146) );
  NAND2_X1 U5083 ( .A1(n5042), .A2(n4146), .ZN(n5977) );
  INV_X1 U5084 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6569) );
  INV_X1 U5085 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6560) );
  NAND3_X1 U5086 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n4149) );
  NAND2_X1 U5087 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5126) );
  INV_X1 U5088 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U5089 ( .A1(n4147), .A2(n6522), .ZN(n6517) );
  INV_X1 U5090 ( .A(n6517), .ZN(n4489) );
  OR2_X1 U5091 ( .A1(n3288), .A2(n4489), .ZN(n4324) );
  NOR2_X1 U5092 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5036) );
  INV_X1 U5093 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6533) );
  NAND4_X1 U5094 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .A4(n5042), .ZN(n5063) );
  INV_X1 U5095 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U5096 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5980), .ZN(n5429) );
  NAND3_X1 U5097 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        n5397), .ZN(n5372) );
  INV_X1 U5098 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U5099 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5868) );
  INV_X1 U5100 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U5101 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5835) );
  INV_X1 U5102 ( .A(n5835), .ZN(n4151) );
  NOR2_X2 U5103 ( .A1(n6569), .A2(n5830), .ZN(n5819) );
  NAND2_X1 U5104 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5819), .ZN(n5315) );
  INV_X1 U5105 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6570) );
  INV_X1 U5106 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6547) );
  AND2_X1 U5107 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4152), .ZN(n5033) );
  NAND4_X1 U5108 ( .A1(n5033), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5131) );
  NOR3_X1 U5109 ( .A1(n6547), .A2(n5131), .A3(n5126), .ZN(n5218) );
  NAND4_X1 U5110 ( .A1(n5218), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U5111 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4153) );
  NOR3_X1 U5112 ( .A1(n6667), .A2(n5378), .A3(n4153), .ZN(n5369) );
  NAND4_X1 U5113 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5369), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U5114 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5346) );
  NOR2_X1 U5115 ( .A1(n5347), .A2(n5346), .ZN(n4154) );
  NAND2_X1 U5116 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5831), .ZN(n5820) );
  OAI21_X1 U5117 ( .B1(n5820), .B2(n6570), .A(n5379), .ZN(n4155) );
  INV_X1 U5118 ( .A(n4155), .ZN(n5318) );
  NOR2_X1 U5119 ( .A1(n5302), .A2(n5318), .ZN(n5294) );
  NAND2_X1 U5120 ( .A1(n5294), .A2(n3110), .ZN(n4272) );
  INV_X1 U5121 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4158) );
  NAND2_X1 U5122 ( .A1(n5477), .A2(n4158), .ZN(n4164) );
  NAND2_X1 U5123 ( .A1(n4423), .A2(n4158), .ZN(n4162) );
  NAND2_X1 U5124 ( .A1(n4159), .A2(n3271), .ZN(n4231) );
  NAND2_X1 U5125 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4160)
         );
  NAND2_X1 U5126 ( .A1(n4231), .A2(n4160), .ZN(n4161) );
  NAND2_X1 U5127 ( .A1(n4162), .A2(n4161), .ZN(n4163) );
  NAND2_X1 U5128 ( .A1(n4231), .A2(EBX_REG_0__SCAN_IN), .ZN(n4166) );
  INV_X1 U5129 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U5130 ( .A1(n4157), .A2(n4434), .ZN(n4165) );
  NAND2_X1 U5131 ( .A1(n4166), .A2(n4165), .ZN(n4353) );
  INV_X1 U5132 ( .A(n4431), .ZN(n4172) );
  NAND2_X1 U5133 ( .A1(n4231), .A2(n3994), .ZN(n4168) );
  INV_X1 U5134 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U5135 ( .A1(n4423), .A2(n6729), .ZN(n4167) );
  NAND3_X1 U5136 ( .A1(n4168), .A2(n4157), .A3(n4167), .ZN(n4170) );
  NAND2_X1 U5137 ( .A1(n5477), .A2(n6729), .ZN(n4169) );
  AND2_X1 U5138 ( .A1(n4170), .A2(n4169), .ZN(n4432) );
  NAND2_X1 U5139 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4173)
         );
  OAI211_X1 U5140 ( .C1(n4294), .C2(EBX_REG_3__SCAN_IN), .A(n4231), .B(n4173), 
        .ZN(n4174) );
  OAI21_X1 U5141 ( .B1(n4258), .B2(EBX_REG_3__SCAN_IN), .A(n4174), .ZN(n4440)
         );
  NAND2_X1 U5142 ( .A1(n4231), .A2(n6271), .ZN(n4176) );
  INV_X1 U5143 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U5144 ( .A1(n4423), .A2(n6662), .ZN(n4175) );
  NAND3_X1 U5145 ( .A1(n4176), .A2(n4157), .A3(n4175), .ZN(n4178) );
  NAND2_X1 U5146 ( .A1(n5477), .A2(n6662), .ZN(n4177) );
  NAND2_X1 U5147 ( .A1(n4178), .A2(n4177), .ZN(n4554) );
  NAND2_X1 U5148 ( .A1(n4555), .A2(n4554), .ZN(n4557) );
  MUX2_X1 U5149 ( .A(n4258), .B(n4157), .S(EBX_REG_5__SCAN_IN), .Z(n4179) );
  OAI21_X1 U5150 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4340), .A(n4179), 
        .ZN(n4513) );
  NAND2_X1 U5151 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4180)
         );
  NAND2_X1 U5152 ( .A1(n4231), .A2(n4180), .ZN(n4182) );
  INV_X1 U5153 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5154 ( .A1(n4423), .A2(n4863), .ZN(n4181) );
  AOI22_X1 U5155 ( .A1(n4182), .A2(n4181), .B1(n5477), .B2(n4863), .ZN(n4671)
         );
  NAND2_X1 U5156 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4183)
         );
  OAI211_X1 U5157 ( .C1(n4294), .C2(EBX_REG_7__SCAN_IN), .A(n4231), .B(n4183), 
        .ZN(n4184) );
  OAI21_X1 U5158 ( .B1(n4258), .B2(EBX_REG_7__SCAN_IN), .A(n4184), .ZN(n4867)
         );
  NAND2_X1 U5159 ( .A1(n4231), .A2(n4185), .ZN(n4187) );
  INV_X1 U5160 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4188) );
  NAND2_X1 U5161 ( .A1(n4423), .A2(n4188), .ZN(n4186) );
  NAND3_X1 U5162 ( .A1(n4187), .A2(n4157), .A3(n4186), .ZN(n4190) );
  NAND2_X1 U5163 ( .A1(n5477), .A2(n4188), .ZN(n4189) );
  NAND2_X1 U5164 ( .A1(n4190), .A2(n4189), .ZN(n4945) );
  MUX2_X1 U5165 ( .A(n4258), .B(n4157), .S(EBX_REG_9__SCAN_IN), .Z(n4192) );
  OR2_X1 U5166 ( .A1(n4340), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4191)
         );
  NAND2_X1 U5167 ( .A1(n4192), .A2(n4191), .ZN(n5990) );
  INV_X1 U5168 ( .A(n5990), .ZN(n4193) );
  NAND2_X1 U5169 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U5170 ( .A1(n4231), .A2(n4194), .ZN(n4197) );
  INV_X1 U5171 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U5172 ( .A1(n4423), .A2(n4195), .ZN(n4196) );
  AOI22_X1 U5173 ( .A1(n4197), .A2(n4196), .B1(n5477), .B2(n4195), .ZN(n5125)
         );
  MUX2_X1 U5174 ( .A(n4258), .B(n4157), .S(EBX_REG_11__SCAN_IN), .Z(n4198) );
  OAI21_X1 U5175 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n4340), .A(n4198), 
        .ZN(n5205) );
  NAND2_X1 U5176 ( .A1(n4231), .A2(n5242), .ZN(n4200) );
  INV_X1 U5177 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U5178 ( .A1(n4423), .A2(n4201), .ZN(n4199) );
  NAND3_X1 U5179 ( .A1(n4200), .A2(n4157), .A3(n4199), .ZN(n4203) );
  NAND2_X1 U5180 ( .A1(n5477), .A2(n4201), .ZN(n4202) );
  NAND2_X1 U5181 ( .A1(n4203), .A2(n4202), .ZN(n5219) );
  NAND2_X1 U5182 ( .A1(n5220), .A2(n5219), .ZN(n5420) );
  NAND2_X1 U5183 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4204) );
  OAI211_X1 U5184 ( .C1(n4294), .C2(EBX_REG_13__SCAN_IN), .A(n4231), .B(n4204), 
        .ZN(n4205) );
  OAI21_X1 U5185 ( .B1(n4258), .B2(EBX_REG_13__SCAN_IN), .A(n4205), .ZN(n5421)
         );
  NAND2_X1 U5186 ( .A1(n4231), .A2(n5920), .ZN(n4209) );
  INV_X1 U5187 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U5188 ( .A1(n4423), .A2(n5498), .ZN(n4208) );
  NAND3_X1 U5189 ( .A1(n4209), .A2(n4157), .A3(n4208), .ZN(n4211) );
  NAND2_X1 U5190 ( .A1(n5477), .A2(n5498), .ZN(n4210) );
  AND2_X1 U5191 ( .A1(n4211), .A2(n4210), .ZN(n5404) );
  MUX2_X1 U5192 ( .A(n4258), .B(n4157), .S(EBX_REG_15__SCAN_IN), .Z(n4212) );
  OAI21_X1 U5193 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4340), .A(n4212), 
        .ZN(n5393) );
  NAND2_X1 U5194 ( .A1(n4231), .A2(n5921), .ZN(n4214) );
  INV_X1 U5195 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U5196 ( .A1(n4423), .A2(n5493), .ZN(n4213) );
  NAND3_X1 U5197 ( .A1(n4214), .A2(n4157), .A3(n4213), .ZN(n4216) );
  NAND2_X1 U5198 ( .A1(n5477), .A2(n5493), .ZN(n4215) );
  NAND2_X1 U5199 ( .A1(n4216), .A2(n4215), .ZN(n5381) );
  MUX2_X1 U5200 ( .A(n4258), .B(n4157), .S(EBX_REG_17__SCAN_IN), .Z(n4217) );
  OAI21_X1 U5201 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4340), .A(n4217), 
        .ZN(n5366) );
  NAND2_X1 U5202 ( .A1(n4231), .A2(n4064), .ZN(n4219) );
  INV_X1 U5203 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U5204 ( .A1(n4423), .A2(n6687), .ZN(n4218) );
  NAND3_X1 U5205 ( .A1(n4219), .A2(n4157), .A3(n4218), .ZN(n4221) );
  NAND2_X1 U5206 ( .A1(n5477), .A2(n6687), .ZN(n4220) );
  AND2_X1 U5207 ( .A1(n4221), .A2(n4220), .ZN(n5481) );
  INV_X1 U5208 ( .A(n4340), .ZN(n4355) );
  NOR2_X1 U5209 ( .A1(n4294), .A2(EBX_REG_20__SCAN_IN), .ZN(n4223) );
  AOI21_X1 U5210 ( .B1(n4355), .B2(n5774), .A(n4223), .ZN(n5470) );
  OR2_X1 U5211 ( .A1(n4340), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4224)
         );
  INV_X1 U5212 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U5213 ( .A1(n4423), .A2(n5490), .ZN(n5478) );
  NAND2_X1 U5214 ( .A1(n4224), .A2(n5478), .ZN(n5479) );
  NAND2_X1 U5215 ( .A1(n5477), .A2(EBX_REG_20__SCAN_IN), .ZN(n4226) );
  NAND2_X1 U5216 ( .A1(n5479), .A2(n4157), .ZN(n4225) );
  OAI211_X1 U5217 ( .C1(n5470), .C2(n5479), .A(n4226), .B(n4225), .ZN(n4227)
         );
  INV_X1 U5218 ( .A(n4227), .ZN(n4228) );
  INV_X1 U5219 ( .A(n4258), .ZN(n4229) );
  INV_X1 U5220 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U5221 ( .A1(n4229), .A2(n5845), .ZN(n4233) );
  NAND2_X1 U5222 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4230) );
  OAI211_X1 U5223 ( .C1(n4294), .C2(EBX_REG_21__SCAN_IN), .A(n4231), .B(n4230), 
        .ZN(n4232) );
  AND2_X1 U5224 ( .A1(n4233), .A2(n4232), .ZN(n5461) );
  NAND2_X1 U5225 ( .A1(n4231), .A2(n6716), .ZN(n4235) );
  INV_X1 U5226 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U5227 ( .A1(n4423), .A2(n5454), .ZN(n4234) );
  NAND3_X1 U5228 ( .A1(n4235), .A2(n4157), .A3(n4234), .ZN(n4237) );
  NAND2_X1 U5229 ( .A1(n5477), .A2(n5454), .ZN(n4236) );
  AND2_X1 U5230 ( .A1(n4237), .A2(n4236), .ZN(n5349) );
  NAND2_X1 U5231 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4238) );
  OAI211_X1 U5232 ( .C1(n4294), .C2(EBX_REG_23__SCAN_IN), .A(n4231), .B(n4238), 
        .ZN(n4239) );
  OAI21_X1 U5233 ( .B1(n4258), .B2(EBX_REG_23__SCAN_IN), .A(n4239), .ZN(n5333)
         );
  INV_X1 U5234 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U5235 ( .A1(n4231), .A2(n6648), .ZN(n4241) );
  INV_X1 U5236 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U5237 ( .A1(n4423), .A2(n4242), .ZN(n4240) );
  NAND3_X1 U5238 ( .A1(n4241), .A2(n4157), .A3(n4240), .ZN(n4244) );
  NAND2_X1 U5239 ( .A1(n5477), .A2(n4242), .ZN(n4243) );
  NAND2_X1 U5240 ( .A1(n4244), .A2(n4243), .ZN(n5324) );
  NAND2_X1 U5241 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4245) );
  OAI211_X1 U5242 ( .C1(n4294), .C2(EBX_REG_25__SCAN_IN), .A(n4231), .B(n4245), 
        .ZN(n4246) );
  OAI21_X1 U5243 ( .B1(n4258), .B2(EBX_REG_25__SCAN_IN), .A(n4246), .ZN(n5446)
         );
  NAND2_X1 U5244 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4247) );
  NAND2_X1 U5245 ( .A1(n4231), .A2(n4247), .ZN(n4250) );
  INV_X1 U5246 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4248) );
  NAND2_X1 U5247 ( .A1(n4423), .A2(n4248), .ZN(n4249) );
  AOI22_X1 U5248 ( .A1(n4250), .A2(n4249), .B1(n5477), .B2(n4248), .ZN(n5440)
         );
  NAND2_X1 U5249 ( .A1(n4157), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4251) );
  OAI211_X1 U5250 ( .C1(n4294), .C2(EBX_REG_27__SCAN_IN), .A(n4231), .B(n4251), 
        .ZN(n4252) );
  OAI21_X1 U5251 ( .B1(n4258), .B2(EBX_REG_27__SCAN_IN), .A(n4252), .ZN(n5262)
         );
  INV_X1 U5252 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5253 ( .A1(n4231), .A2(n4253), .ZN(n4255) );
  INV_X1 U5254 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U5255 ( .A1(n4423), .A2(n5312), .ZN(n4254) );
  NAND3_X1 U5256 ( .A1(n4255), .A2(n4157), .A3(n4254), .ZN(n4257) );
  NAND2_X1 U5257 ( .A1(n5477), .A2(n5312), .ZN(n4256) );
  NAND2_X1 U5258 ( .A1(n4257), .A2(n4256), .ZN(n5310) );
  MUX2_X1 U5259 ( .A(EBX_REG_29__SCAN_IN), .B(n3116), .S(n4157), .Z(n4260) );
  NOR2_X1 U5260 ( .A1(n4258), .A2(EBX_REG_29__SCAN_IN), .ZN(n4259) );
  NOR2_X1 U5261 ( .A1(n4260), .A2(n4259), .ZN(n5299) );
  AND2_X1 U5262 ( .A1(n4294), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4261)
         );
  AOI21_X1 U5263 ( .B1(n4340), .B2(EBX_REG_30__SCAN_IN), .A(n4261), .ZN(n5277)
         );
  NAND2_X1 U5264 ( .A1(n5299), .A2(n5277), .ZN(n4264) );
  OAI22_X1 U5265 ( .A1(n4340), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4294), .ZN(n4265) );
  NOR2_X1 U5266 ( .A1(n3051), .A2(n5036), .ZN(n4267) );
  NAND2_X1 U5267 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4270)
         );
  NAND2_X1 U5268 ( .A1(n4489), .A2(n5036), .ZN(n6491) );
  NAND4_X1 U5269 ( .A1(n3281), .A2(n5052), .A3(EBX_REG_31__SCAN_IN), .A4(n6491), .ZN(n4269) );
  INV_X1 U5270 ( .A(n5315), .ZN(n4271) );
  NAND3_X1 U5271 ( .A1(n4271), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5289) );
  INV_X1 U5272 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U5273 ( .A1(n4338), .A2(n5053), .ZN(n4273) );
  NOR2_X1 U5274 ( .A1(n4273), .A2(n5267), .ZN(n4298) );
  NAND2_X1 U5275 ( .A1(n4382), .A2(n4298), .ZN(n4278) );
  INV_X1 U5276 ( .A(n4297), .ZN(n4275) );
  NOR2_X1 U5277 ( .A1(READY_N), .A2(n4275), .ZN(n4319) );
  INV_X1 U5278 ( .A(n4319), .ZN(n4276) );
  OR2_X1 U5279 ( .A1(n4274), .A2(n4276), .ZN(n4277) );
  NAND2_X1 U5280 ( .A1(n4278), .A2(n4277), .ZN(n4366) );
  AND3_X1 U5281 ( .A1(n3044), .A2(n4421), .A3(n3267), .ZN(n4412) );
  AND2_X1 U5282 ( .A1(n4279), .A2(n4412), .ZN(n4280) );
  NAND2_X1 U5283 ( .A1(n4338), .A2(n3155), .ZN(n4282) );
  NAND2_X1 U5284 ( .A1(n4371), .A2(n4423), .ZN(n4358) );
  AND2_X1 U5285 ( .A1(n6074), .A2(n4421), .ZN(n4284) );
  NOR2_X2 U5286 ( .A1(n6067), .A2(n4325), .ZN(n6065) );
  AOI22_X1 U5287 ( .A1(n6065), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6067), .ZN(n4286) );
  NAND2_X1 U5288 ( .A1(n4287), .A2(n4286), .ZN(U2860) );
  NOR2_X1 U5289 ( .A1(n6400), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5043) );
  INV_X1 U5290 ( .A(n4288), .ZN(n4307) );
  AOI211_X1 U5291 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4289), .A(n5043), .B(
        n4307), .ZN(n4290) );
  INV_X1 U5292 ( .A(n4290), .ZN(U2788) );
  OR2_X1 U5293 ( .A1(n4382), .A2(n5053), .ZN(n4293) );
  NAND2_X1 U5294 ( .A1(n4291), .A2(n4299), .ZN(n4292) );
  NAND2_X1 U5295 ( .A1(n4293), .A2(n4292), .ZN(n5944) );
  INV_X1 U5296 ( .A(n5053), .ZN(n4295) );
  NAND3_X1 U5297 ( .A1(n4295), .A2(n6517), .A3(n4294), .ZN(n4296) );
  INV_X1 U5298 ( .A(READY_N), .ZN(n6612) );
  AND2_X1 U5299 ( .A1(n4296), .A2(n6612), .ZN(n6613) );
  NOR2_X1 U5300 ( .A1(n5944), .A2(n6613), .ZN(n6474) );
  OR2_X1 U5301 ( .A1(n6474), .A2(n6499), .ZN(n4302) );
  INV_X1 U5302 ( .A(n4302), .ZN(n5950) );
  INV_X1 U5303 ( .A(MORE_REG_SCAN_IN), .ZN(n4304) );
  INV_X1 U5304 ( .A(n5267), .ZN(n4314) );
  NAND3_X1 U5305 ( .A1(n4123), .A2(n4314), .A3(n3288), .ZN(n4386) );
  INV_X1 U5306 ( .A(n4386), .ZN(n4345) );
  NOR2_X1 U5307 ( .A1(n4297), .A2(n4347), .ZN(n4301) );
  INV_X1 U5308 ( .A(n4298), .ZN(n4387) );
  AND2_X1 U5309 ( .A1(n4387), .A2(n6476), .ZN(n4332) );
  AOI21_X1 U5310 ( .B1(n4332), .B2(n4299), .A(n4382), .ZN(n4300) );
  AOI211_X1 U5311 ( .C1(n4345), .C2(n4382), .A(n4301), .B(n4300), .ZN(n6477)
         );
  OR2_X1 U5312 ( .A1(n6477), .A2(n4302), .ZN(n4303) );
  OAI21_X1 U5313 ( .B1(n5950), .B2(n4304), .A(n4303), .ZN(U3471) );
  NOR2_X1 U5314 ( .A1(n5043), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4306) );
  OAI21_X1 U5315 ( .B1(n5053), .B2(n4423), .A(n6610), .ZN(n4305) );
  OAI21_X1 U5316 ( .B1(n4306), .B2(n6610), .A(n4305), .ZN(U3474) );
  INV_X1 U5317 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U5318 ( .A1(n4371), .A2(n3281), .ZN(n6490) );
  INV_X1 U5319 ( .A(n6166), .ZN(n4309) );
  INV_X1 U5320 ( .A(DATAI_9_), .ZN(n4308) );
  NOR2_X1 U5321 ( .A1(n6124), .A2(n4308), .ZN(n6148) );
  AOI21_X1 U5322 ( .B1(n4309), .B2(EAX_REG_25__SCAN_IN), .A(n6148), .ZN(n4310)
         );
  OAI21_X1 U5323 ( .B1(n6113), .B2(n6659), .A(n4310), .ZN(U2933) );
  XNOR2_X1 U5324 ( .A(n4311), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4406)
         );
  NAND2_X1 U5325 ( .A1(n4314), .A2(n3288), .ZN(n4322) );
  NAND2_X1 U5326 ( .A1(n4281), .A2(n3271), .ZN(n4313) );
  INV_X1 U5327 ( .A(n3272), .ZN(n4312) );
  MUX2_X1 U5328 ( .A(n4313), .B(n6614), .S(n4312), .Z(n4343) );
  INV_X1 U5329 ( .A(n4123), .ZN(n4316) );
  NAND2_X1 U5330 ( .A1(n4314), .A2(n4338), .ZN(n4315) );
  AOI21_X1 U5331 ( .B1(n4316), .B2(n4315), .A(n4334), .ZN(n4317) );
  NAND2_X1 U5332 ( .A1(n4343), .A2(n4317), .ZN(n4318) );
  NAND2_X1 U5333 ( .A1(n4318), .A2(n4347), .ZN(n4362) );
  NAND2_X1 U5334 ( .A1(n3288), .A2(n6517), .ZN(n4320) );
  NAND3_X1 U5335 ( .A1(n4320), .A2(n4319), .A3(n4533), .ZN(n4321) );
  OAI211_X1 U5336 ( .C1(n4382), .C2(n4322), .A(n4362), .B(n4321), .ZN(n4323)
         );
  NAND2_X1 U5337 ( .A1(n4323), .A2(n4416), .ZN(n4330) );
  NAND3_X1 U5338 ( .A1(n4371), .A2(n4324), .A3(n6612), .ZN(n4326) );
  NAND3_X1 U5339 ( .A1(n4326), .A2(n3271), .A3(n4325), .ZN(n4327) );
  NAND2_X1 U5340 ( .A1(n4327), .A2(n3278), .ZN(n4328) );
  OR2_X1 U5341 ( .A1(n4350), .A2(n3044), .ZN(n4331) );
  NAND4_X1 U5342 ( .A1(n4332), .A2(n4274), .A3(n4358), .A4(n4331), .ZN(n4333)
         );
  NAND2_X1 U5343 ( .A1(n4334), .A2(n5477), .ZN(n4336) );
  OAI211_X1 U5344 ( .C1(n3278), .C2(n3300), .A(n4336), .B(n4335), .ZN(n4337)
         );
  INV_X1 U5345 ( .A(n4337), .ZN(n4342) );
  NOR2_X1 U5346 ( .A1(n5057), .A2(n4533), .ZN(n4360) );
  INV_X1 U5347 ( .A(n4338), .ZN(n4339) );
  OAI21_X1 U5348 ( .B1(n4360), .B2(n4340), .A(n4339), .ZN(n4341) );
  AND4_X1 U5349 ( .A1(n4343), .A2(n4342), .A3(n3277), .A4(n4341), .ZN(n4376)
         );
  OAI211_X1 U5350 ( .C1(n4374), .C2(n3271), .A(n4376), .B(n4450), .ZN(n4344)
         );
  INV_X1 U5351 ( .A(n5794), .ZN(n4346) );
  AND2_X1 U5352 ( .A1(n4346), .A2(n6288), .ZN(n5790) );
  OR2_X1 U5353 ( .A1(n4352), .A2(n6206), .ZN(n4675) );
  INV_X1 U5354 ( .A(n4675), .ZN(n4348) );
  NOR2_X1 U5355 ( .A1(n4347), .A2(n3298), .ZN(n4456) );
  NOR2_X1 U5356 ( .A1(n4348), .A2(n5788), .ZN(n4349) );
  MUX2_X1 U5357 ( .A(n5790), .B(n4349), .S(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .Z(n4357) );
  OAI21_X1 U5358 ( .B1(n4350), .B2(n3244), .A(n6490), .ZN(n4351) );
  INV_X1 U5359 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4674) );
  INV_X1 U5360 ( .A(n4353), .ZN(n4354) );
  AOI21_X1 U5361 ( .B1(n4355), .B2(n4674), .A(n4354), .ZN(n5103) );
  AOI22_X1 U5362 ( .A1(n6286), .A2(n5103), .B1(n6258), .B2(REIP_REG_0__SCAN_IN), .ZN(n4356) );
  OAI211_X1 U5363 ( .C1(n4406), .C2(n6208), .A(n4357), .B(n4356), .ZN(U3018)
         );
  NOR2_X1 U5364 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6591), .ZN(n6587) );
  OAI21_X1 U5365 ( .B1(n4456), .B2(n4371), .A(n4489), .ZN(n4359) );
  AOI21_X1 U5366 ( .B1(n4359), .B2(n4358), .A(READY_N), .ZN(n4364) );
  INV_X1 U5367 ( .A(n4360), .ZN(n4361) );
  NAND2_X1 U5368 ( .A1(n4362), .A2(n4361), .ZN(n4363) );
  AOI21_X1 U5369 ( .B1(n4382), .B2(n4364), .A(n4363), .ZN(n4365) );
  OR2_X1 U5370 ( .A1(n4382), .A2(n4386), .ZN(n4415) );
  AND2_X1 U5371 ( .A1(n4365), .A2(n4415), .ZN(n4368) );
  INV_X1 U5372 ( .A(n4366), .ZN(n4367) );
  NAND2_X1 U5373 ( .A1(n4368), .A2(n4367), .ZN(n6464) );
  INV_X1 U5374 ( .A(n6464), .ZN(n4369) );
  NOR2_X1 U5375 ( .A1(n3407), .A2(n6501), .ZN(n5803) );
  NAND2_X1 U5376 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5803), .ZN(n6588) );
  INV_X1 U5377 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5949) );
  OAI22_X1 U5378 ( .A1(n4369), .A2(n6499), .B1(n6588), .B2(n5949), .ZN(n5940)
         );
  NOR2_X1 U5379 ( .A1(n6587), .A2(n5940), .ZN(n6598) );
  INV_X1 U5380 ( .A(n4279), .ZN(n4373) );
  INV_X1 U5381 ( .A(n4371), .ZN(n4372) );
  AND4_X1 U5382 ( .A1(n4374), .A2(n4274), .A3(n4373), .A4(n4372), .ZN(n4375)
         );
  NAND2_X1 U5383 ( .A1(n4376), .A2(n4375), .ZN(n4446) );
  INV_X1 U5384 ( .A(n4446), .ZN(n5268) );
  NOR3_X1 U5385 ( .A1(n5267), .A2(n4377), .A3(n4378), .ZN(n4379) );
  AOI21_X1 U5386 ( .B1(n4456), .B2(n4076), .A(n4379), .ZN(n4380) );
  OAI21_X1 U5387 ( .B1(n6049), .B2(n5268), .A(n4380), .ZN(n6463) );
  INV_X1 U5388 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U5389 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4381), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4673), .ZN(n4398) );
  NAND2_X1 U5390 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4397) );
  INV_X1 U5391 ( .A(n4397), .ZN(n5269) );
  INV_X1 U5392 ( .A(n4377), .ZN(n4466) );
  NOR2_X1 U5393 ( .A1(n4378), .A2(n6595), .ZN(n4400) );
  AOI222_X1 U5394 ( .A1(n6463), .A2(n6593), .B1(n4398), .B2(n5269), .C1(n4466), 
        .C2(n4400), .ZN(n4384) );
  NAND2_X1 U5395 ( .A1(n6598), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U5396 ( .B1(n6598), .B2(n4384), .A(n4383), .ZN(U3460) );
  INV_X1 U5397 ( .A(n4456), .ZN(n5271) );
  XNOR2_X1 U5398 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5399 ( .A1(n4385), .A2(n4446), .ZN(n4393) );
  NAND2_X1 U5400 ( .A1(n4387), .A2(n4386), .ZN(n4453) );
  INV_X1 U5401 ( .A(n4378), .ZN(n4388) );
  NAND2_X1 U5402 ( .A1(n4388), .A2(n4395), .ZN(n4447) );
  NAND2_X1 U5403 ( .A1(n4378), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U5404 ( .A1(n4447), .A2(n4389), .ZN(n4391) );
  NOR2_X1 U5405 ( .A1(n4450), .A2(n4391), .ZN(n4390) );
  AOI21_X1 U5406 ( .B1(n4453), .B2(n4391), .A(n4390), .ZN(n4392) );
  OAI211_X1 U5407 ( .C1(n5271), .C2(n4394), .A(n4393), .B(n4392), .ZN(n4444)
         );
  INV_X1 U5408 ( .A(n6595), .ZN(n6492) );
  NAND3_X1 U5409 ( .A1(n4378), .A2(n4395), .A3(n6492), .ZN(n4396) );
  OAI21_X1 U5410 ( .B1(n4398), .B2(n4397), .A(n4396), .ZN(n4399) );
  AOI21_X1 U5411 ( .B1(n4444), .B2(n6593), .A(n4399), .ZN(n4402) );
  OAI21_X1 U5412 ( .B1(n6598), .B2(n4400), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4401) );
  OAI21_X1 U5413 ( .B1(n6598), .B2(n4402), .A(n4401), .ZN(U3459) );
  XNOR2_X1 U5414 ( .A(n4404), .B(n4403), .ZN(n5109) );
  INV_X1 U5415 ( .A(n5109), .ZN(n4410) );
  INV_X1 U5416 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4405) );
  OAI22_X1 U5417 ( .A1(n6178), .A2(n4406), .B1(n5907), .B2(n4405), .ZN(n4409)
         );
  INV_X1 U5418 ( .A(n6194), .ZN(n5652) );
  AOI21_X1 U5419 ( .B1(n5652), .B2(n4407), .A(n5105), .ZN(n4408) );
  AOI211_X1 U5420 ( .C1(n5894), .C2(n4410), .A(n4409), .B(n4408), .ZN(n4411)
         );
  INV_X1 U5421 ( .A(n4411), .ZN(U2986) );
  NAND3_X1 U5422 ( .A1(n4413), .A2(n4412), .A3(n4423), .ZN(n4414) );
  NAND2_X1 U5423 ( .A1(n4415), .A2(n4414), .ZN(n4417) );
  OR2_X2 U5424 ( .A1(n6625), .A2(n4421), .ZN(n5460) );
  OAI21_X1 U5425 ( .B1(n4420), .B2(n4419), .A(n4418), .ZN(n6055) );
  OAI21_X1 U5426 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(n6046) );
  AOI22_X1 U5427 ( .A1(n6622), .A2(n6046), .B1(n6625), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4425) );
  OAI21_X1 U5428 ( .B1(n5460), .B2(n6055), .A(n4425), .ZN(U2858) );
  NAND3_X1 U5429 ( .A1(n4428), .A2(n4427), .A3(n4418), .ZN(n4429) );
  NAND2_X1 U5430 ( .A1(n4426), .A2(n4429), .ZN(n6195) );
  INV_X1 U5431 ( .A(n4441), .ZN(n4430) );
  AOI21_X1 U5432 ( .B1(n4432), .B2(n4431), .A(n4430), .ZN(n6285) );
  AOI22_X1 U5433 ( .A1(n6622), .A2(n6285), .B1(n6625), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4433) );
  OAI21_X1 U5434 ( .B1(n6195), .B2(n5460), .A(n4433), .ZN(U2857) );
  INV_X1 U5435 ( .A(n5103), .ZN(n4435) );
  OAI222_X1 U5436 ( .A1(n5499), .A2(n4435), .B1(n4434), .B2(n5497), .C1(n5460), 
        .C2(n5109), .ZN(U2859) );
  NAND2_X1 U5437 ( .A1(n3272), .A2(n5258), .ZN(n4436) );
  INV_X1 U5438 ( .A(DATAI_2_), .ZN(n4532) );
  OAI222_X1 U5439 ( .A1(n6195), .A2(n5871), .B1(n5521), .B2(n4532), .C1(n6074), 
        .C2(n3423), .ZN(U2889) );
  INV_X1 U5440 ( .A(DATAI_0_), .ZN(n4540) );
  OAI222_X1 U5441 ( .A1(n5871), .A2(n5109), .B1(n5521), .B2(n4540), .C1(n6074), 
        .C2(n3419), .ZN(U2891) );
  INV_X1 U5442 ( .A(DATAI_1_), .ZN(n6098) );
  OAI222_X1 U5443 ( .A1(n6055), .A2(n5871), .B1(n6074), .B2(n4437), .C1(n5521), 
        .C2(n6098), .ZN(U2890) );
  INV_X1 U5444 ( .A(n4426), .ZN(n4439) );
  AND2_X1 U5445 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  OR2_X1 U5446 ( .A1(n4555), .A2(n4442), .ZN(n6273) );
  INV_X1 U5447 ( .A(n6273), .ZN(n5065) );
  AOI22_X1 U5448 ( .A1(n6622), .A2(n5065), .B1(n6625), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4443) );
  OAI21_X1 U5449 ( .B1(n5072), .B2(n5460), .A(n4443), .ZN(U2856) );
  MUX2_X1 U5450 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4444), .S(n6464), 
        .Z(n6467) );
  NAND2_X1 U5451 ( .A1(n6344), .A2(n4446), .ZN(n4460) );
  XNOR2_X1 U5452 ( .A(n4447), .B(n3043), .ZN(n4452) );
  INV_X1 U5453 ( .A(n4448), .ZN(n4449) );
  OAI211_X1 U5454 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n4378), .A(n3315), .B(n4449), .ZN(n6594) );
  NOR2_X1 U5455 ( .A1(n4450), .A2(n6594), .ZN(n4451) );
  AOI21_X1 U5456 ( .B1(n4453), .B2(n4452), .A(n4451), .ZN(n4458) );
  NAND2_X1 U5457 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4454) );
  XNOR2_X1 U5458 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4454), .ZN(n4455)
         );
  NAND2_X1 U5459 ( .A1(n4456), .A2(n4455), .ZN(n4457) );
  AND2_X1 U5460 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND2_X1 U5461 ( .A1(n4460), .A2(n4459), .ZN(n6592) );
  NAND2_X1 U5462 ( .A1(n6464), .A2(n6592), .ZN(n4461) );
  OAI21_X1 U5463 ( .B1(n6464), .B2(n3450), .A(n4461), .ZN(n6470) );
  NAND3_X1 U5464 ( .A1(n6467), .A2(n6501), .A3(n6470), .ZN(n4465) );
  NAND2_X1 U5465 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5949), .ZN(n4471) );
  INV_X1 U5466 ( .A(n4471), .ZN(n4462) );
  NAND2_X1 U5467 ( .A1(n4463), .A2(n4462), .ZN(n4464) );
  NAND2_X1 U5468 ( .A1(n4465), .A2(n4464), .ZN(n6480) );
  NAND2_X1 U5469 ( .A1(n6480), .A2(n4466), .ZN(n4474) );
  INV_X1 U5470 ( .A(n4467), .ZN(n5006) );
  NOR2_X1 U5471 ( .A1(n4468), .A2(n5006), .ZN(n4469) );
  XNOR2_X1 U5472 ( .A(n4469), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6036)
         );
  OAI22_X1 U5473 ( .A1(n6464), .A2(n4470), .B1(n6036), .B2(n4274), .ZN(n4473)
         );
  NOR2_X1 U5474 ( .A1(n4470), .A2(n4471), .ZN(n4472) );
  AOI21_X1 U5475 ( .B1(n4473), .B2(n6501), .A(n4472), .ZN(n6478) );
  NAND2_X1 U5476 ( .A1(n4474), .A2(n6478), .ZN(n6483) );
  NOR2_X1 U5477 ( .A1(n6483), .A2(FLUSH_REG_SCAN_IN), .ZN(n4475) );
  INV_X1 U5478 ( .A(n6508), .ZN(n6615) );
  OAI21_X1 U5479 ( .B1(n4475), .B2(n6588), .A(n4543), .ZN(n6296) );
  NOR2_X1 U5480 ( .A1(n4476), .A2(n5002), .ZN(n6299) );
  AOI211_X1 U5481 ( .C1(n5002), .C2(n4476), .A(n6400), .B(n6299), .ZN(n4478)
         );
  AND2_X1 U5482 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6591), .ZN(n5811) );
  NOR2_X1 U5483 ( .A1(n6049), .A2(n5811), .ZN(n4477) );
  OAI21_X1 U5484 ( .B1(n4478), .B2(n4477), .A(n6296), .ZN(n4479) );
  OAI21_X1 U5485 ( .B1(n6296), .B2(n4775), .A(n4479), .ZN(U3464) );
  INV_X1 U5486 ( .A(DATAI_3_), .ZN(n4528) );
  INV_X1 U5487 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6134) );
  OAI222_X1 U5488 ( .A1(n5072), .A2(n5871), .B1(n5521), .B2(n4528), .C1(n6074), 
        .C2(n6134), .ZN(U2888) );
  XNOR2_X1 U5489 ( .A(n4481), .B(n4480), .ZN(n4687) );
  OAI21_X1 U5490 ( .B1(n5790), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4675), 
        .ZN(n4482) );
  NAND2_X1 U5491 ( .A1(n4482), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4486)
         );
  INV_X1 U5492 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6600) );
  NOR2_X1 U5493 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5788), .ZN(n4678)
         );
  NAND2_X1 U5494 ( .A1(n5238), .A2(n6288), .ZN(n6222) );
  INV_X1 U5495 ( .A(n6222), .ZN(n6220) );
  OR3_X1 U5496 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4678), .A3(n6220), 
        .ZN(n4483) );
  OAI21_X1 U5497 ( .B1(n5907), .B2(n6600), .A(n4483), .ZN(n4484) );
  AOI21_X1 U5498 ( .B1(n6286), .B2(n6046), .A(n4484), .ZN(n4485) );
  OAI211_X1 U5499 ( .C1(n4687), .C2(n6208), .A(n4486), .B(n4485), .ZN(U3017)
         );
  NAND2_X1 U5500 ( .A1(n5803), .A2(n6493), .ZN(n6487) );
  INV_X2 U5501 ( .A(n6487), .ZN(n6094) );
  NOR2_X4 U5502 ( .A1(n4492), .A2(n6094), .ZN(n6090) );
  AOI22_X1 U5503 ( .A1(DATAO_REG_22__SCAN_IN), .A2(n6090), .B1(n6094), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4493) );
  OAI21_X1 U5504 ( .B1(n3771), .B2(n6075), .A(n4493), .ZN(U2901) );
  INV_X1 U5505 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6103) );
  AOI22_X1 U5506 ( .A1(DATAO_REG_19__SCAN_IN), .A2(n6090), .B1(n6094), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4494) );
  OAI21_X1 U5507 ( .B1(n6103), .B2(n6075), .A(n4494), .ZN(U2904) );
  AOI22_X1 U5508 ( .A1(n6094), .A2(UWORD_REG_12__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4495) );
  OAI21_X1 U5509 ( .B1(n3904), .B2(n6075), .A(n4495), .ZN(U2895) );
  AOI22_X1 U5510 ( .A1(n6094), .A2(UWORD_REG_13__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4496) );
  OAI21_X1 U5511 ( .B1(n3930), .B2(n6075), .A(n4496), .ZN(U2894) );
  INV_X1 U5512 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U5513 ( .A1(n6094), .A2(UWORD_REG_10__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4497) );
  OAI21_X1 U5514 ( .B1(n6706), .B2(n6075), .A(n4497), .ZN(U2897) );
  INV_X1 U5515 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6701) );
  AOI22_X1 U5516 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6094), .B1(n6090), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4498) );
  OAI21_X1 U5517 ( .B1(n6701), .B2(n6075), .A(n4498), .ZN(U2902) );
  AOI22_X1 U5518 ( .A1(n6094), .A2(UWORD_REG_7__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4499) );
  OAI21_X1 U5519 ( .B1(n3802), .B2(n6075), .A(n4499), .ZN(U2900) );
  AOI22_X1 U5520 ( .A1(n6094), .A2(UWORD_REG_8__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4500) );
  OAI21_X1 U5521 ( .B1(n3823), .B2(n6075), .A(n4500), .ZN(U2899) );
  AOI22_X1 U5522 ( .A1(n6094), .A2(UWORD_REG_14__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4501) );
  OAI21_X1 U5523 ( .B1(n3966), .B2(n6075), .A(n4501), .ZN(U2893) );
  AOI22_X1 U5524 ( .A1(n6094), .A2(UWORD_REG_0__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5525 ( .B1(n3664), .B2(n6075), .A(n4502), .ZN(U2907) );
  INV_X1 U5526 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U5527 ( .A1(n6094), .A2(UWORD_REG_1__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4503) );
  OAI21_X1 U5528 ( .B1(n6100), .B2(n6075), .A(n4503), .ZN(U2906) );
  AOI22_X1 U5529 ( .A1(n6094), .A2(UWORD_REG_2__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4504) );
  OAI21_X1 U5530 ( .B1(n3698), .B2(n6075), .A(n4504), .ZN(U2905) );
  INV_X1 U5531 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6105) );
  AOI22_X1 U5532 ( .A1(n6094), .A2(UWORD_REG_4__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4505) );
  OAI21_X1 U5533 ( .B1(n6105), .B2(n6075), .A(n4505), .ZN(U2903) );
  INV_X1 U5534 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6118) );
  AOI22_X1 U5535 ( .A1(n6094), .A2(UWORD_REG_11__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4506) );
  OAI21_X1 U5536 ( .B1(n6118), .B2(n6075), .A(n4506), .ZN(U2896) );
  OAI21_X1 U5537 ( .B1(n4507), .B2(n4510), .A(n4509), .ZN(n6025) );
  INV_X1 U5538 ( .A(n4511), .ZN(n4512) );
  AOI21_X1 U5539 ( .B1(n4513), .B2(n4557), .A(n4512), .ZN(n6256) );
  AOI22_X1 U5540 ( .A1(n6622), .A2(n6256), .B1(n6625), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4514) );
  OAI21_X1 U5541 ( .B1(n6025), .B2(n5460), .A(n4514), .ZN(U2854) );
  NAND2_X1 U5542 ( .A1(n5894), .A2(DATAI_20_), .ZN(n6434) );
  AND2_X1 U5543 ( .A1(n4476), .A2(n4559), .ZN(n4516) );
  AOI21_X1 U5544 ( .B1(n4525), .B2(STATEBS16_REG_SCAN_IN), .A(n6400), .ZN(
        n4519) );
  AND2_X1 U5545 ( .A1(n6344), .A2(n3418), .ZN(n4707) );
  NAND2_X1 U5546 ( .A1(n4385), .A2(n6049), .ZN(n4817) );
  INV_X1 U5547 ( .A(n4817), .ZN(n5005) );
  NOR2_X1 U5548 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6469), .ZN(n4561)
         );
  NAND2_X1 U5549 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4561), .ZN(n4812) );
  NOR2_X1 U5550 ( .A1(n6460), .A2(n4812), .ZN(n4549) );
  AOI21_X1 U5551 ( .B1(n4707), .B2(n5005), .A(n4549), .ZN(n4523) );
  AOI22_X1 U5552 ( .A1(n4519), .A2(n4523), .B1(n6400), .B2(n4812), .ZN(n4518)
         );
  NAND2_X1 U5553 ( .A1(n6402), .A2(n4518), .ZN(n4547) );
  INV_X1 U5554 ( .A(DATAI_4_), .ZN(n4598) );
  NOR2_X1 U5555 ( .A1(n4598), .A2(n4543), .ZN(n6431) );
  INV_X1 U5556 ( .A(n4519), .ZN(n4522) );
  INV_X1 U5557 ( .A(n4561), .ZN(n4521) );
  NAND2_X1 U5558 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4520) );
  OAI22_X1 U5559 ( .A1(n4523), .A2(n4522), .B1(n4521), .B2(n4520), .ZN(n4546)
         );
  AOI22_X1 U5560 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4547), .B1(n6431), 
        .B2(n4546), .ZN(n4527) );
  NAND2_X1 U5561 ( .A1(n4548), .A2(n3244), .ZN(n5198) );
  INV_X1 U5562 ( .A(n5198), .ZN(n6429) );
  NAND2_X1 U5563 ( .A1(n5894), .A2(DATAI_28_), .ZN(n6369) );
  INV_X1 U5564 ( .A(n6369), .ZN(n6430) );
  AOI22_X1 U5565 ( .A1(n6429), .A2(n4549), .B1(n6430), .B2(n4859), .ZN(n4526)
         );
  OAI211_X1 U5566 ( .C1(n6434), .C2(n4602), .A(n4527), .B(n4526), .ZN(U3128)
         );
  NAND2_X1 U5567 ( .A1(n5894), .A2(DATAI_19_), .ZN(n6363) );
  NOR2_X1 U5568 ( .A1(n4528), .A2(n4543), .ZN(n6425) );
  AOI22_X1 U5569 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4547), .B1(n6425), 
        .B2(n4546), .ZN(n4531) );
  NAND2_X1 U5570 ( .A1(n4548), .A2(n4529), .ZN(n5177) );
  NAND2_X1 U5571 ( .A1(n5894), .A2(DATAI_27_), .ZN(n6428) );
  INV_X1 U5572 ( .A(n6428), .ZN(n6360) );
  AOI22_X1 U5573 ( .A1(n6423), .A2(n4549), .B1(n6360), .B2(n4859), .ZN(n4530)
         );
  OAI211_X1 U5574 ( .C1(n6363), .C2(n4602), .A(n4531), .B(n4530), .ZN(U3127)
         );
  NAND2_X1 U5575 ( .A1(n5894), .A2(DATAI_18_), .ZN(n6315) );
  NOR2_X1 U5576 ( .A1(n4532), .A2(n4543), .ZN(n6419) );
  AOI22_X1 U5577 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4547), .B1(n6419), 
        .B2(n4546), .ZN(n4535) );
  NAND2_X1 U5578 ( .A1(n4548), .A2(n4533), .ZN(n5171) );
  INV_X1 U5579 ( .A(n5171), .ZN(n6417) );
  NAND2_X1 U5580 ( .A1(n5894), .A2(DATAI_26_), .ZN(n6422) );
  INV_X1 U5581 ( .A(n6422), .ZN(n6312) );
  AOI22_X1 U5582 ( .A1(n6417), .A2(n4549), .B1(n6312), .B2(n4859), .ZN(n4534)
         );
  OAI211_X1 U5583 ( .C1(n6315), .C2(n4602), .A(n4535), .B(n4534), .ZN(U3126)
         );
  NAND2_X1 U5584 ( .A1(n5894), .A2(DATAI_22_), .ZN(n6375) );
  AOI22_X1 U5585 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4547), .B1(n6444), 
        .B2(n4546), .ZN(n4537) );
  NAND2_X1 U5586 ( .A1(n4548), .A2(n3267), .ZN(n4982) );
  NAND2_X1 U5587 ( .A1(n5894), .A2(DATAI_30_), .ZN(n6448) );
  INV_X1 U5588 ( .A(n6448), .ZN(n6372) );
  AOI22_X1 U5589 ( .A1(n6441), .A2(n4549), .B1(n6372), .B2(n4859), .ZN(n4536)
         );
  OAI211_X1 U5590 ( .C1(n6375), .C2(n4602), .A(n4537), .B(n4536), .ZN(U3130)
         );
  NAND2_X1 U5591 ( .A1(n5894), .A2(DATAI_23_), .ZN(n6459) );
  AOI22_X1 U5592 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4547), .B1(n6454), 
        .B2(n4546), .ZN(n4539) );
  NAND2_X1 U5593 ( .A1(n4548), .A2(n5258), .ZN(n4965) );
  AOI22_X1 U5594 ( .A1(n6450), .A2(n4549), .B1(n6451), .B2(n4859), .ZN(n4538)
         );
  OAI211_X1 U5595 ( .C1(n6459), .C2(n4602), .A(n4539), .B(n4538), .ZN(U3131)
         );
  NAND2_X1 U5596 ( .A1(n5894), .A2(DATAI_16_), .ZN(n6410) );
  NOR2_X1 U5597 ( .A1(n4540), .A2(n4543), .ZN(n6407) );
  AOI22_X1 U5598 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4547), .B1(n6407), 
        .B2(n4546), .ZN(n4542) );
  NAND2_X1 U5599 ( .A1(n4548), .A2(n3271), .ZN(n5183) );
  NAND2_X1 U5600 ( .A1(n5894), .A2(DATAI_24_), .ZN(n6309) );
  INV_X1 U5601 ( .A(n6309), .ZN(n6394) );
  AOI22_X1 U5602 ( .A1(n6393), .A2(n4549), .B1(n6394), .B2(n4859), .ZN(n4541)
         );
  OAI211_X1 U5603 ( .C1(n6410), .C2(n4602), .A(n4542), .B(n4541), .ZN(U3124)
         );
  NAND2_X1 U5604 ( .A1(n5894), .A2(DATAI_21_), .ZN(n6440) );
  INV_X1 U5605 ( .A(DATAI_5_), .ZN(n4624) );
  NOR2_X1 U5606 ( .A1(n4624), .A2(n4543), .ZN(n6437) );
  AOI22_X1 U5607 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4547), .B1(n6437), 
        .B2(n4546), .ZN(n4545) );
  NAND2_X1 U5608 ( .A1(n4548), .A2(n3263), .ZN(n5189) );
  INV_X1 U5609 ( .A(n5189), .ZN(n6435) );
  NAND2_X1 U5610 ( .A1(n5894), .A2(DATAI_29_), .ZN(n6324) );
  INV_X1 U5611 ( .A(n6324), .ZN(n6436) );
  AOI22_X1 U5612 ( .A1(n6435), .A2(n4549), .B1(n6436), .B2(n4859), .ZN(n4544)
         );
  OAI211_X1 U5613 ( .C1(n6440), .C2(n4602), .A(n4545), .B(n4544), .ZN(U3129)
         );
  NAND2_X1 U5614 ( .A1(n5894), .A2(DATAI_17_), .ZN(n6416) );
  AOI22_X1 U5615 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4547), .B1(n6413), 
        .B2(n4546), .ZN(n4551) );
  NAND2_X1 U5616 ( .A1(n4548), .A2(n3288), .ZN(n4972) );
  NAND2_X1 U5617 ( .A1(n5894), .A2(DATAI_25_), .ZN(n6357) );
  INV_X1 U5618 ( .A(n6357), .ZN(n6412) );
  AOI22_X1 U5619 ( .A1(n6411), .A2(n4549), .B1(n6412), .B2(n4859), .ZN(n4550)
         );
  OAI211_X1 U5620 ( .C1(n6416), .C2(n4602), .A(n4551), .B(n4550), .ZN(U3125)
         );
  INV_X1 U5621 ( .A(n4552), .ZN(n4553) );
  XNOR2_X1 U5622 ( .A(n4553), .B(n4438), .ZN(n6189) );
  INV_X1 U5623 ( .A(n6189), .ZN(n4599) );
  OR2_X1 U5624 ( .A1(n4555), .A2(n4554), .ZN(n4556) );
  AND2_X1 U5625 ( .A1(n4557), .A2(n4556), .ZN(n6265) );
  AOI22_X1 U5626 ( .A1(n6622), .A2(n6265), .B1(n6625), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4558) );
  OAI21_X1 U5627 ( .B1(n4599), .B2(n5460), .A(n4558), .ZN(U2855) );
  INV_X1 U5628 ( .A(n4559), .ZN(n4600) );
  AND2_X1 U5629 ( .A1(n5809), .A2(n4476), .ZN(n4568) );
  INV_X1 U5630 ( .A(n4568), .ZN(n4560) );
  INV_X1 U5631 ( .A(n6400), .ZN(n6396) );
  OAI21_X1 U5632 ( .B1(n4560), .B2(n5002), .A(n6396), .ZN(n4567) );
  INV_X1 U5633 ( .A(n4567), .ZN(n4564) );
  NAND2_X1 U5634 ( .A1(n3418), .A2(n5006), .ZN(n4562) );
  NAND2_X1 U5635 ( .A1(n4561), .A2(n6391), .ZN(n5001) );
  OR2_X1 U5636 ( .A1(n6460), .A2(n5001), .ZN(n4592) );
  OAI21_X1 U5637 ( .B1(n4817), .B2(n4562), .A(n4592), .ZN(n4566) );
  INV_X1 U5638 ( .A(n5001), .ZN(n4563) );
  AOI22_X1 U5639 ( .A1(n4564), .A2(n4566), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4563), .ZN(n4597) );
  INV_X1 U5640 ( .A(n6419), .ZN(n5170) );
  NAND2_X1 U5641 ( .A1(n5001), .A2(n6400), .ZN(n4565) );
  OAI211_X1 U5642 ( .C1(n4567), .C2(n4566), .A(n6402), .B(n4565), .ZN(n4591)
         );
  NAND2_X1 U5643 ( .A1(n4591), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U5644 ( .A1(n4568), .A2(n4517), .ZN(n5003) );
  AND2_X1 U5645 ( .A1(n4476), .A2(n4773), .ZN(n4569) );
  OAI22_X1 U5646 ( .A1(n6315), .A2(n4593), .B1(n5171), .B2(n4592), .ZN(n4570)
         );
  AOI21_X1 U5647 ( .B1(n6312), .B2(n5100), .A(n4570), .ZN(n4571) );
  OAI211_X1 U5648 ( .C1(n4597), .C2(n5170), .A(n4572), .B(n4571), .ZN(U3062)
         );
  INV_X1 U5649 ( .A(n6413), .ZN(n5012) );
  NAND2_X1 U5650 ( .A1(n4591), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4575) );
  OAI22_X1 U5651 ( .A1(n6416), .A2(n4593), .B1(n4972), .B2(n4592), .ZN(n4573)
         );
  AOI21_X1 U5652 ( .B1(n6412), .B2(n5100), .A(n4573), .ZN(n4574) );
  OAI211_X1 U5653 ( .C1(n4597), .C2(n5012), .A(n4575), .B(n4574), .ZN(U3061)
         );
  INV_X1 U5654 ( .A(n6454), .ZN(n5015) );
  NAND2_X1 U5655 ( .A1(n4591), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4578) );
  OAI22_X1 U5656 ( .A1(n6459), .A2(n4593), .B1(n4965), .B2(n4592), .ZN(n4576)
         );
  AOI21_X1 U5657 ( .B1(n6451), .B2(n5100), .A(n4576), .ZN(n4577) );
  OAI211_X1 U5658 ( .C1(n4597), .C2(n5015), .A(n4578), .B(n4577), .ZN(U3067)
         );
  INV_X1 U5659 ( .A(n6407), .ZN(n5182) );
  NAND2_X1 U5660 ( .A1(n4591), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4581) );
  OAI22_X1 U5661 ( .A1(n6410), .A2(n4593), .B1(n5183), .B2(n4592), .ZN(n4579)
         );
  AOI21_X1 U5662 ( .B1(n6394), .B2(n5100), .A(n4579), .ZN(n4580) );
  OAI211_X1 U5663 ( .C1(n4597), .C2(n5182), .A(n4581), .B(n4580), .ZN(U3060)
         );
  INV_X1 U5664 ( .A(n6431), .ZN(n5195) );
  NAND2_X1 U5665 ( .A1(n4591), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4584) );
  OAI22_X1 U5666 ( .A1(n6434), .A2(n4593), .B1(n5198), .B2(n4592), .ZN(n4582)
         );
  AOI21_X1 U5667 ( .B1(n6430), .B2(n5100), .A(n4582), .ZN(n4583) );
  OAI211_X1 U5668 ( .C1(n4597), .C2(n5195), .A(n4584), .B(n4583), .ZN(U3064)
         );
  INV_X1 U5669 ( .A(n6425), .ZN(n5176) );
  NAND2_X1 U5670 ( .A1(n4591), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4587) );
  OAI22_X1 U5671 ( .A1(n6363), .A2(n4593), .B1(n5177), .B2(n4592), .ZN(n4585)
         );
  AOI21_X1 U5672 ( .B1(n6360), .B2(n5100), .A(n4585), .ZN(n4586) );
  OAI211_X1 U5673 ( .C1(n4597), .C2(n5176), .A(n4587), .B(n4586), .ZN(U3063)
         );
  INV_X1 U5674 ( .A(n6444), .ZN(n5018) );
  NAND2_X1 U5675 ( .A1(n4591), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4590) );
  OAI22_X1 U5676 ( .A1(n6375), .A2(n4593), .B1(n4982), .B2(n4592), .ZN(n4588)
         );
  AOI21_X1 U5677 ( .B1(n6372), .B2(n5100), .A(n4588), .ZN(n4589) );
  OAI211_X1 U5678 ( .C1(n4597), .C2(n5018), .A(n4590), .B(n4589), .ZN(U3066)
         );
  INV_X1 U5679 ( .A(n6437), .ZN(n5188) );
  NAND2_X1 U5680 ( .A1(n4591), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4596) );
  OAI22_X1 U5681 ( .A1(n6440), .A2(n4593), .B1(n5189), .B2(n4592), .ZN(n4594)
         );
  AOI21_X1 U5682 ( .B1(n6436), .B2(n5100), .A(n4594), .ZN(n4595) );
  OAI211_X1 U5683 ( .C1(n4597), .C2(n5188), .A(n4596), .B(n4595), .ZN(U3065)
         );
  INV_X1 U5684 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6137) );
  OAI222_X1 U5685 ( .A1(n5871), .A2(n4599), .B1(n5521), .B2(n4598), .C1(n6074), 
        .C2(n6137), .ZN(U2887) );
  NOR2_X1 U5686 ( .A1(n4476), .A2(n4600), .ZN(n4601) );
  NAND2_X1 U5687 ( .A1(n4515), .A2(n4601), .ZN(n4697) );
  NOR2_X2 U5688 ( .A1(n4697), .A2(n4773), .ZN(n4938) );
  INV_X1 U5689 ( .A(n4938), .ZN(n4623) );
  NOR2_X1 U5690 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4695), .ZN(n4651)
         );
  OAI21_X1 U5691 ( .B1(n4880), .B2(n3407), .A(n4881), .ZN(n4960) );
  NOR2_X1 U5692 ( .A1(n4606), .A2(n3407), .ZN(n5147) );
  NOR3_X1 U5693 ( .A1(n4960), .A2(n6391), .A3(n5147), .ZN(n4605) );
  INV_X1 U5694 ( .A(n6049), .ZN(n4706) );
  NAND2_X1 U5695 ( .A1(n4385), .A2(n4706), .ZN(n6345) );
  OAI21_X1 U5696 ( .B1(n4650), .B2(n4938), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4603) );
  NAND3_X1 U5697 ( .A1(n6345), .A2(n6396), .A3(n4603), .ZN(n4604) );
  OAI211_X1 U5698 ( .C1(n4651), .C2(n6591), .A(n4605), .B(n4604), .ZN(n4642)
         );
  NAND2_X1 U5699 ( .A1(n4642), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4609)
         );
  INV_X1 U5700 ( .A(n4651), .ZN(n4619) );
  NOR2_X1 U5701 ( .A1(n6345), .A2(n6400), .ZN(n4628) );
  AND2_X1 U5702 ( .A1(n4606), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4996) );
  INV_X1 U5703 ( .A(n4880), .ZN(n4744) );
  NOR2_X1 U5704 ( .A1(n4744), .A2(n6391), .ZN(n4959) );
  AOI22_X1 U5705 ( .A1(n4628), .A2(n6344), .B1(n4996), .B2(n4959), .ZN(n4643)
         );
  OAI22_X1 U5706 ( .A1(n5198), .A2(n4619), .B1(n4643), .B2(n5195), .ZN(n4607)
         );
  AOI21_X1 U5707 ( .B1(n6430), .B2(n4650), .A(n4607), .ZN(n4608) );
  OAI211_X1 U5708 ( .C1(n4623), .C2(n6434), .A(n4609), .B(n4608), .ZN(U3136)
         );
  NAND2_X1 U5709 ( .A1(n4642), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4612)
         );
  OAI22_X1 U5710 ( .A1(n5183), .A2(n4619), .B1(n4643), .B2(n5182), .ZN(n4610)
         );
  AOI21_X1 U5711 ( .B1(n6394), .B2(n4650), .A(n4610), .ZN(n4611) );
  OAI211_X1 U5712 ( .C1(n4623), .C2(n6410), .A(n4612), .B(n4611), .ZN(U3132)
         );
  NAND2_X1 U5713 ( .A1(n4642), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4615)
         );
  OAI22_X1 U5714 ( .A1(n5177), .A2(n4619), .B1(n4643), .B2(n5176), .ZN(n4613)
         );
  AOI21_X1 U5715 ( .B1(n6360), .B2(n4650), .A(n4613), .ZN(n4614) );
  OAI211_X1 U5716 ( .C1(n4623), .C2(n6363), .A(n4615), .B(n4614), .ZN(U3135)
         );
  NAND2_X1 U5717 ( .A1(n4642), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4618)
         );
  OAI22_X1 U5718 ( .A1(n5189), .A2(n4619), .B1(n4643), .B2(n5188), .ZN(n4616)
         );
  AOI21_X1 U5719 ( .B1(n6436), .B2(n4650), .A(n4616), .ZN(n4617) );
  OAI211_X1 U5720 ( .C1(n4623), .C2(n6440), .A(n4618), .B(n4617), .ZN(U3137)
         );
  NAND2_X1 U5721 ( .A1(n4642), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4622)
         );
  OAI22_X1 U5722 ( .A1(n5171), .A2(n4619), .B1(n4643), .B2(n5170), .ZN(n4620)
         );
  AOI21_X1 U5723 ( .B1(n6312), .B2(n4650), .A(n4620), .ZN(n4621) );
  OAI211_X1 U5724 ( .C1(n4623), .C2(n6315), .A(n4622), .B(n4621), .ZN(U3134)
         );
  INV_X1 U5725 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6140) );
  OAI222_X1 U5726 ( .A1(n6025), .A2(n5871), .B1(n5521), .B2(n4624), .C1(n6074), 
        .C2(n6140), .ZN(U2886) );
  NAND2_X1 U5727 ( .A1(n5809), .A2(n5137), .ZN(n6368) );
  OAI21_X1 U5728 ( .B1(n6376), .B2(n6337), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4625) );
  NAND3_X1 U5729 ( .A1(n6345), .A2(n6396), .A3(n4625), .ZN(n4627) );
  NOR2_X1 U5730 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6349), .ZN(n6336)
         );
  INV_X1 U5731 ( .A(n6336), .ZN(n4638) );
  AOI211_X1 U5732 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4638), .A(n5147), .B(
        n4960), .ZN(n4626) );
  NAND3_X1 U5733 ( .A1(n6391), .A2(n4627), .A3(n4626), .ZN(n6338) );
  NAND2_X1 U5734 ( .A1(n6338), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4631) );
  AND2_X1 U5735 ( .A1(n4880), .A2(n6391), .ZN(n5146) );
  AOI22_X1 U5736 ( .A1(n4628), .A2(n5812), .B1(n5146), .B2(n4996), .ZN(n4657)
         );
  OAI22_X1 U5737 ( .A1(n5189), .A2(n4638), .B1(n4657), .B2(n5188), .ZN(n4629)
         );
  AOI21_X1 U5738 ( .B1(n6436), .B2(n6337), .A(n4629), .ZN(n4630) );
  OAI211_X1 U5739 ( .C1(n6368), .C2(n6440), .A(n4631), .B(n4630), .ZN(U3073)
         );
  NAND2_X1 U5740 ( .A1(n6338), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4634) );
  OAI22_X1 U5741 ( .A1(n5198), .A2(n4638), .B1(n4657), .B2(n5195), .ZN(n4632)
         );
  AOI21_X1 U5742 ( .B1(n6430), .B2(n6337), .A(n4632), .ZN(n4633) );
  OAI211_X1 U5743 ( .C1(n6368), .C2(n6434), .A(n4634), .B(n4633), .ZN(U3072)
         );
  NAND2_X1 U5744 ( .A1(n6338), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4637) );
  OAI22_X1 U5745 ( .A1(n5171), .A2(n4638), .B1(n4657), .B2(n5170), .ZN(n4635)
         );
  AOI21_X1 U5746 ( .B1(n6312), .B2(n6337), .A(n4635), .ZN(n4636) );
  OAI211_X1 U5747 ( .C1(n6368), .C2(n6315), .A(n4637), .B(n4636), .ZN(U3070)
         );
  NAND2_X1 U5748 ( .A1(n6338), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4641) );
  OAI22_X1 U5749 ( .A1(n5177), .A2(n4638), .B1(n4657), .B2(n5176), .ZN(n4639)
         );
  AOI21_X1 U5750 ( .B1(n6360), .B2(n6337), .A(n4639), .ZN(n4640) );
  OAI211_X1 U5751 ( .C1(n6368), .C2(n6363), .A(n4641), .B(n4640), .ZN(U3071)
         );
  INV_X1 U5752 ( .A(n4642), .ZN(n4656) );
  INV_X1 U5753 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5754 ( .A1(n6450), .A2(n4651), .B1(n6451), .B2(n4650), .ZN(n4645)
         );
  INV_X1 U5755 ( .A(n4643), .ZN(n4652) );
  INV_X1 U5756 ( .A(n6459), .ZN(n5150) );
  AOI22_X1 U5757 ( .A1(n6454), .A2(n4652), .B1(n5150), .B2(n4938), .ZN(n4644)
         );
  OAI211_X1 U5758 ( .C1(n4656), .C2(n4646), .A(n4645), .B(n4644), .ZN(U3139)
         );
  INV_X1 U5759 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5760 ( .A1(n6411), .A2(n4651), .B1(n6412), .B2(n4650), .ZN(n4648)
         );
  INV_X1 U5761 ( .A(n6416), .ZN(n6354) );
  AOI22_X1 U5762 ( .A1(n6413), .A2(n4652), .B1(n6354), .B2(n4938), .ZN(n4647)
         );
  OAI211_X1 U5763 ( .C1(n4656), .C2(n4649), .A(n4648), .B(n4647), .ZN(U3133)
         );
  INV_X1 U5764 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5765 ( .A1(n6441), .A2(n4651), .B1(n6372), .B2(n4650), .ZN(n4654)
         );
  INV_X1 U5766 ( .A(n6375), .ZN(n6443) );
  AOI22_X1 U5767 ( .A1(n6444), .A2(n4652), .B1(n6443), .B2(n4938), .ZN(n4653)
         );
  OAI211_X1 U5768 ( .C1(n4656), .C2(n4655), .A(n4654), .B(n4653), .ZN(U3138)
         );
  INV_X1 U5769 ( .A(n6338), .ZN(n4667) );
  INV_X1 U5770 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5771 ( .A1(n6441), .A2(n6336), .B1(n6372), .B2(n6337), .ZN(n4659)
         );
  INV_X1 U5772 ( .A(n4657), .ZN(n6335) );
  AOI22_X1 U5773 ( .A1(n6444), .A2(n6335), .B1(n6443), .B2(n6376), .ZN(n4658)
         );
  OAI211_X1 U5774 ( .C1(n4667), .C2(n4660), .A(n4659), .B(n4658), .ZN(U3074)
         );
  INV_X1 U5775 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5776 ( .A1(n6450), .A2(n6336), .B1(n6451), .B2(n6337), .ZN(n4662)
         );
  AOI22_X1 U5777 ( .A1(n6454), .A2(n6335), .B1(n5150), .B2(n6376), .ZN(n4661)
         );
  OAI211_X1 U5778 ( .C1(n4667), .C2(n4663), .A(n4662), .B(n4661), .ZN(U3075)
         );
  INV_X1 U5779 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5780 ( .A1(n6411), .A2(n6336), .B1(n6412), .B2(n6337), .ZN(n4665)
         );
  AOI22_X1 U5781 ( .A1(n6413), .A2(n6335), .B1(n6354), .B2(n6376), .ZN(n4664)
         );
  OAI211_X1 U5782 ( .C1(n4667), .C2(n4666), .A(n4665), .B(n4664), .ZN(U3069)
         );
  OAI21_X1 U5783 ( .B1(n4670), .B2(n4669), .A(n4668), .ZN(n6179) );
  NAND2_X1 U5784 ( .A1(n4511), .A2(n4671), .ZN(n4672) );
  NAND2_X1 U5785 ( .A1(n4866), .A2(n4672), .ZN(n6015) );
  NOR2_X1 U5786 ( .A1(n6274), .A2(n6015), .ZN(n4682) );
  AOI21_X1 U5788 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6283) );
  NOR2_X1 U5789 ( .A1(n6271), .A2(n6279), .ZN(n6263) );
  NAND2_X1 U5790 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6263), .ZN(n6217)
         );
  NOR2_X1 U5791 ( .A1(n6283), .A2(n6217), .ZN(n5237) );
  INV_X1 U5792 ( .A(n5237), .ZN(n4677) );
  NOR2_X1 U5793 ( .A1(n3994), .A2(n4673), .ZN(n6284) );
  NAND2_X1 U5794 ( .A1(n5794), .A2(n4674), .ZN(n4676) );
  OAI21_X1 U5795 ( .B1(n5238), .B2(n6284), .A(n6219), .ZN(n6282) );
  AOI21_X1 U5796 ( .B1(n4677), .B2(n6222), .A(n6282), .ZN(n6262) );
  INV_X1 U5797 ( .A(n4678), .ZN(n4679) );
  NAND2_X1 U5798 ( .A1(n6281), .A2(n6284), .ZN(n6253) );
  AOI21_X1 U5799 ( .B1(n6288), .B2(n6253), .A(n6283), .ZN(n6225) );
  INV_X1 U5800 ( .A(n6225), .ZN(n6280) );
  OAI33_X1 U5801 ( .A1(1'b0), .A2(n6262), .A3(n6218), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6217), .B3(n6280), .ZN(n4681) );
  AOI211_X1 U5802 ( .C1(n6206), .C2(REIP_REG_6__SCAN_IN), .A(n4682), .B(n4681), 
        .ZN(n4683) );
  OAI21_X1 U5803 ( .B1(n6208), .B2(n6179), .A(n4683), .ZN(U3012) );
  INV_X1 U5804 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6050) );
  AOI22_X1 U5805 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6258), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4684) );
  OAI21_X1 U5806 ( .B1(n6055), .B2(n6173), .A(n4684), .ZN(n4685) );
  AOI21_X1 U5807 ( .B1(n5657), .B2(n6050), .A(n4685), .ZN(n4686) );
  OAI21_X1 U5808 ( .B1(n4687), .B2(n6178), .A(n4686), .ZN(U2985) );
  INV_X1 U5809 ( .A(n4697), .ZN(n4689) );
  NOR2_X1 U5810 ( .A1(n6400), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5142) );
  INV_X1 U5811 ( .A(n5142), .ZN(n4688) );
  OAI21_X1 U5812 ( .B1(n4689), .B2(n6173), .A(n4688), .ZN(n4694) );
  INV_X1 U5813 ( .A(n6345), .ZN(n4691) );
  INV_X1 U5814 ( .A(n4690), .ZN(n4934) );
  AOI21_X1 U5815 ( .B1(n4707), .B2(n4691), .A(n4934), .ZN(n4696) );
  OAI21_X1 U5816 ( .B1(n6396), .B2(n4692), .A(n6402), .ZN(n4693) );
  AOI21_X1 U5817 ( .B1(n4694), .B2(n4696), .A(n4693), .ZN(n4941) );
  INV_X1 U5818 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4700) );
  OAI22_X1 U5819 ( .A1(n4696), .A2(n6400), .B1(n4695), .B2(n3407), .ZN(n4933)
         );
  AOI22_X1 U5820 ( .A1(n6444), .A2(n4933), .B1(n6372), .B2(n4938), .ZN(n4699)
         );
  NOR2_X2 U5821 ( .A1(n4697), .A2(n4517), .ZN(n5024) );
  AOI22_X1 U5822 ( .A1(n6441), .A2(n4934), .B1(n6443), .B2(n5024), .ZN(n4698)
         );
  OAI211_X1 U5823 ( .C1(n4941), .C2(n4700), .A(n4699), .B(n4698), .ZN(U3146)
         );
  INV_X1 U5824 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5825 ( .A1(n6454), .A2(n4933), .B1(n6451), .B2(n4938), .ZN(n4702)
         );
  AOI22_X1 U5826 ( .A1(n6450), .A2(n4934), .B1(n5150), .B2(n5024), .ZN(n4701)
         );
  OAI211_X1 U5827 ( .C1(n4941), .C2(n4703), .A(n4702), .B(n4701), .ZN(U3147)
         );
  AOI22_X1 U5828 ( .A1(n6413), .A2(n4933), .B1(n6412), .B2(n4938), .ZN(n4705)
         );
  AOI22_X1 U5829 ( .A1(n6411), .A2(n4934), .B1(n6354), .B2(n5024), .ZN(n4704)
         );
  OAI211_X1 U5830 ( .C1(n4941), .C2(n3199), .A(n4705), .B(n4704), .ZN(U3141)
         );
  NOR2_X1 U5831 ( .A1(n4385), .A2(n4706), .ZN(n4774) );
  NAND3_X1 U5832 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6469), .A3(n4775), .ZN(n4743) );
  NOR2_X1 U5833 ( .A1(n6460), .A2(n4743), .ZN(n4730) );
  AOI21_X1 U5834 ( .B1(n4707), .B2(n4774), .A(n4730), .ZN(n4710) );
  AOI21_X1 U5835 ( .B1(n4712), .B2(STATEBS16_REG_SCAN_IN), .A(n6400), .ZN(
        n4709) );
  AOI22_X1 U5836 ( .A1(n4710), .A2(n4709), .B1(n6400), .B2(n4743), .ZN(n4708)
         );
  NAND2_X1 U5837 ( .A1(n6402), .A2(n4708), .ZN(n4729) );
  INV_X1 U5838 ( .A(n4709), .ZN(n4711) );
  OAI22_X1 U5839 ( .A1(n4711), .A2(n4710), .B1(n3407), .B2(n4743), .ZN(n4728)
         );
  AOI22_X1 U5840 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4729), .B1(n6407), 
        .B2(n4728), .ZN(n4715) );
  INV_X1 U5841 ( .A(n4712), .ZN(n4713) );
  AOI22_X1 U5842 ( .A1(n6386), .A2(n6394), .B1(n6393), .B2(n4730), .ZN(n4714)
         );
  OAI211_X1 U5843 ( .C1(n4964), .C2(n6410), .A(n4715), .B(n4714), .ZN(U3092)
         );
  AOI22_X1 U5844 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4729), .B1(n6413), 
        .B2(n4728), .ZN(n4717) );
  AOI22_X1 U5845 ( .A1(n6386), .A2(n6412), .B1(n6411), .B2(n4730), .ZN(n4716)
         );
  OAI211_X1 U5846 ( .C1(n4964), .C2(n6416), .A(n4717), .B(n4716), .ZN(U3093)
         );
  AOI22_X1 U5847 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4729), .B1(n6454), 
        .B2(n4728), .ZN(n4719) );
  AOI22_X1 U5848 ( .A1(n6386), .A2(n6451), .B1(n6450), .B2(n4730), .ZN(n4718)
         );
  OAI211_X1 U5849 ( .C1(n4964), .C2(n6459), .A(n4719), .B(n4718), .ZN(U3099)
         );
  AOI22_X1 U5850 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4729), .B1(n6444), 
        .B2(n4728), .ZN(n4721) );
  AOI22_X1 U5851 ( .A1(n6386), .A2(n6372), .B1(n6441), .B2(n4730), .ZN(n4720)
         );
  OAI211_X1 U5852 ( .C1(n4964), .C2(n6375), .A(n4721), .B(n4720), .ZN(U3098)
         );
  AOI22_X1 U5853 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4729), .B1(n6437), 
        .B2(n4728), .ZN(n4723) );
  AOI22_X1 U5854 ( .A1(n6386), .A2(n6436), .B1(n6435), .B2(n4730), .ZN(n4722)
         );
  OAI211_X1 U5855 ( .C1(n4964), .C2(n6440), .A(n4723), .B(n4722), .ZN(U3097)
         );
  AOI22_X1 U5856 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4729), .B1(n6431), 
        .B2(n4728), .ZN(n4725) );
  AOI22_X1 U5857 ( .A1(n6386), .A2(n6430), .B1(n6429), .B2(n4730), .ZN(n4724)
         );
  OAI211_X1 U5858 ( .C1(n4964), .C2(n6434), .A(n4725), .B(n4724), .ZN(U3096)
         );
  AOI22_X1 U5859 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4729), .B1(n6425), 
        .B2(n4728), .ZN(n4727) );
  AOI22_X1 U5860 ( .A1(n6386), .A2(n6360), .B1(n6423), .B2(n4730), .ZN(n4726)
         );
  OAI211_X1 U5861 ( .C1(n4964), .C2(n6363), .A(n4727), .B(n4726), .ZN(U3095)
         );
  AOI22_X1 U5862 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4729), .B1(n6419), 
        .B2(n4728), .ZN(n4732) );
  AOI22_X1 U5863 ( .A1(n6386), .A2(n6312), .B1(n6417), .B2(n4730), .ZN(n4731)
         );
  OAI211_X1 U5864 ( .C1(n4964), .C2(n6315), .A(n4732), .B(n4731), .ZN(U3094)
         );
  INV_X1 U5865 ( .A(n5068), .ZN(n4736) );
  INV_X1 U5866 ( .A(n6206), .ZN(n5907) );
  INV_X1 U5867 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4733) );
  OAI22_X1 U5868 ( .A1(n5652), .A2(n4734), .B1(n5907), .B2(n4733), .ZN(n4735)
         );
  AOI21_X1 U5869 ( .B1(n4736), .B2(n5657), .A(n4735), .ZN(n4741) );
  OR2_X1 U5870 ( .A1(n4738), .A2(n4737), .ZN(n6272) );
  NAND3_X1 U5871 ( .A1(n6272), .A2(n4739), .A3(n6199), .ZN(n4740) );
  OAI211_X1 U5872 ( .C1(n5072), .C2(n6173), .A(n4741), .B(n4740), .ZN(U2983)
         );
  INV_X1 U5873 ( .A(n6386), .ZN(n4769) );
  NOR2_X1 U5874 ( .A1(n4476), .A2(n4517), .ZN(n4999) );
  NAND2_X1 U5875 ( .A1(n5809), .A2(n4999), .ZN(n6390) );
  OAI21_X1 U5876 ( .B1(n6386), .B2(n6364), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4742) );
  NAND2_X1 U5877 ( .A1(n4774), .A2(n6344), .ZN(n4747) );
  NAND3_X1 U5878 ( .A1(n4742), .A2(n6396), .A3(n4747), .ZN(n4746) );
  NOR2_X1 U5879 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4743), .ZN(n6384)
         );
  INV_X1 U5880 ( .A(n6384), .ZN(n4765) );
  AND2_X1 U5881 ( .A1(n4744), .A2(n4879), .ZN(n4818) );
  OAI21_X1 U5882 ( .B1(n4818), .B2(n3407), .A(n4881), .ZN(n4813) );
  AOI211_X1 U5883 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4765), .A(n4996), .B(
        n4813), .ZN(n4745) );
  NAND2_X1 U5884 ( .A1(n4746), .A2(n4745), .ZN(n6387) );
  NAND2_X1 U5885 ( .A1(n6387), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4751) );
  INV_X1 U5886 ( .A(n4747), .ZN(n4748) );
  AOI22_X1 U5887 ( .A1(n4748), .A2(n6396), .B1(n5147), .B2(n4818), .ZN(n4764)
         );
  OAI22_X1 U5888 ( .A1(n5189), .A2(n4765), .B1(n4764), .B2(n5188), .ZN(n4749)
         );
  AOI21_X1 U5889 ( .B1(n6436), .B2(n6364), .A(n4749), .ZN(n4750) );
  OAI211_X1 U5890 ( .C1(n4769), .C2(n6440), .A(n4751), .B(n4750), .ZN(U3089)
         );
  NAND2_X1 U5891 ( .A1(n6387), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4754) );
  OAI22_X1 U5892 ( .A1(n5171), .A2(n4765), .B1(n4764), .B2(n5170), .ZN(n4752)
         );
  AOI21_X1 U5893 ( .B1(n6312), .B2(n6364), .A(n4752), .ZN(n4753) );
  OAI211_X1 U5894 ( .C1(n4769), .C2(n6315), .A(n4754), .B(n4753), .ZN(U3086)
         );
  NAND2_X1 U5895 ( .A1(n6387), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4757) );
  INV_X1 U5896 ( .A(n4764), .ZN(n6385) );
  OAI22_X1 U5897 ( .A1(n4972), .A2(n4765), .B1(n6357), .B2(n6390), .ZN(n4755)
         );
  AOI21_X1 U5898 ( .B1(n6413), .B2(n6385), .A(n4755), .ZN(n4756) );
  OAI211_X1 U5899 ( .C1(n4769), .C2(n6416), .A(n4757), .B(n4756), .ZN(U3085)
         );
  NAND2_X1 U5900 ( .A1(n6387), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4760) );
  OAI22_X1 U5901 ( .A1(n5183), .A2(n4765), .B1(n4764), .B2(n5182), .ZN(n4758)
         );
  AOI21_X1 U5902 ( .B1(n6394), .B2(n6364), .A(n4758), .ZN(n4759) );
  OAI211_X1 U5903 ( .C1(n4769), .C2(n6410), .A(n4760), .B(n4759), .ZN(U3084)
         );
  NAND2_X1 U5904 ( .A1(n6387), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4763) );
  INV_X1 U5905 ( .A(n6451), .ZN(n5153) );
  OAI22_X1 U5906 ( .A1(n4965), .A2(n4765), .B1(n5153), .B2(n6390), .ZN(n4761)
         );
  AOI21_X1 U5907 ( .B1(n6454), .B2(n6385), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5908 ( .C1(n4769), .C2(n6459), .A(n4763), .B(n4762), .ZN(U3091)
         );
  NAND2_X1 U5909 ( .A1(n6387), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4768) );
  OAI22_X1 U5910 ( .A1(n5198), .A2(n4765), .B1(n4764), .B2(n5195), .ZN(n4766)
         );
  AOI21_X1 U5911 ( .B1(n6430), .B2(n6364), .A(n4766), .ZN(n4767) );
  OAI211_X1 U5912 ( .C1(n4769), .C2(n6434), .A(n4768), .B(n4767), .ZN(U3088)
         );
  INV_X1 U5913 ( .A(n3998), .ZN(n4771) );
  INV_X1 U5914 ( .A(n6300), .ZN(n4772) );
  NAND2_X1 U5915 ( .A1(n4772), .A2(n4476), .ZN(n4781) );
  NAND2_X1 U5916 ( .A1(n4774), .A2(n5812), .ZN(n4876) );
  INV_X1 U5917 ( .A(n4876), .ZN(n4884) );
  NAND3_X1 U5918 ( .A1(n6391), .A2(n6469), .A3(n4775), .ZN(n4878) );
  NOR2_X1 U5919 ( .A1(n6460), .A2(n4878), .ZN(n4782) );
  AOI21_X1 U5920 ( .B1(n4884), .B2(n3418), .A(n4782), .ZN(n4780) );
  OR2_X1 U5921 ( .A1(n4781), .A2(n5002), .ZN(n4776) );
  AOI22_X1 U5922 ( .A1(n4780), .A2(n4778), .B1(n6400), .B2(n4878), .ZN(n4777)
         );
  NAND2_X1 U5923 ( .A1(n6402), .A2(n4777), .ZN(n4805) );
  INV_X1 U5924 ( .A(n4778), .ZN(n4779) );
  OAI22_X1 U5925 ( .A1(n4780), .A2(n4779), .B1(n3407), .B2(n4878), .ZN(n4804)
         );
  AOI22_X1 U5926 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4805), .B1(n6407), 
        .B2(n4804), .ZN(n4785) );
  INV_X1 U5927 ( .A(n4782), .ZN(n4806) );
  OAI22_X1 U5928 ( .A1(n5203), .A2(n6410), .B1(n5183), .B2(n4806), .ZN(n4783)
         );
  INV_X1 U5929 ( .A(n4783), .ZN(n4784) );
  OAI211_X1 U5930 ( .C1(n6309), .C2(n5029), .A(n4785), .B(n4784), .ZN(U3028)
         );
  AOI22_X1 U5931 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4805), .B1(n6413), 
        .B2(n4804), .ZN(n4788) );
  OAI22_X1 U5932 ( .A1(n5203), .A2(n6416), .B1(n4972), .B2(n4806), .ZN(n4786)
         );
  INV_X1 U5933 ( .A(n4786), .ZN(n4787) );
  OAI211_X1 U5934 ( .C1(n6357), .C2(n5029), .A(n4788), .B(n4787), .ZN(U3029)
         );
  AOI22_X1 U5935 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4805), .B1(n6425), 
        .B2(n4804), .ZN(n4791) );
  OAI22_X1 U5936 ( .A1(n5203), .A2(n6363), .B1(n5177), .B2(n4806), .ZN(n4789)
         );
  INV_X1 U5937 ( .A(n4789), .ZN(n4790) );
  OAI211_X1 U5938 ( .C1(n6428), .C2(n5029), .A(n4791), .B(n4790), .ZN(U3031)
         );
  AOI22_X1 U5939 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4805), .B1(n6431), 
        .B2(n4804), .ZN(n4794) );
  OAI22_X1 U5940 ( .A1(n5203), .A2(n6434), .B1(n5198), .B2(n4806), .ZN(n4792)
         );
  INV_X1 U5941 ( .A(n4792), .ZN(n4793) );
  OAI211_X1 U5942 ( .C1(n6369), .C2(n5029), .A(n4794), .B(n4793), .ZN(U3032)
         );
  AOI22_X1 U5943 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4805), .B1(n6444), 
        .B2(n4804), .ZN(n4797) );
  OAI22_X1 U5944 ( .A1(n5203), .A2(n6375), .B1(n4982), .B2(n4806), .ZN(n4795)
         );
  INV_X1 U5945 ( .A(n4795), .ZN(n4796) );
  OAI211_X1 U5946 ( .C1(n6448), .C2(n5029), .A(n4797), .B(n4796), .ZN(U3034)
         );
  AOI22_X1 U5947 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4805), .B1(n6454), 
        .B2(n4804), .ZN(n4800) );
  OAI22_X1 U5948 ( .A1(n5203), .A2(n6459), .B1(n4965), .B2(n4806), .ZN(n4798)
         );
  INV_X1 U5949 ( .A(n4798), .ZN(n4799) );
  OAI211_X1 U5950 ( .C1(n5153), .C2(n5029), .A(n4800), .B(n4799), .ZN(U3035)
         );
  AOI22_X1 U5951 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4805), .B1(n6419), 
        .B2(n4804), .ZN(n4803) );
  OAI22_X1 U5952 ( .A1(n5203), .A2(n6315), .B1(n5171), .B2(n4806), .ZN(n4801)
         );
  INV_X1 U5953 ( .A(n4801), .ZN(n4802) );
  OAI211_X1 U5954 ( .C1(n6422), .C2(n5029), .A(n4803), .B(n4802), .ZN(U3030)
         );
  AOI22_X1 U5955 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4805), .B1(n6437), 
        .B2(n4804), .ZN(n4809) );
  OAI22_X1 U5956 ( .A1(n5203), .A2(n6440), .B1(n5189), .B2(n4806), .ZN(n4807)
         );
  INV_X1 U5957 ( .A(n4807), .ZN(n4808) );
  OAI211_X1 U5958 ( .C1(n6324), .C2(n5029), .A(n4809), .B(n4808), .ZN(U3033)
         );
  INV_X1 U5959 ( .A(DATAI_6_), .ZN(n6107) );
  XOR2_X1 U5960 ( .A(n4509), .B(n4810), .Z(n6180) );
  INV_X1 U5961 ( .A(n6180), .ZN(n4862) );
  OAI222_X1 U5962 ( .A1(n6107), .A2(n5521), .B1(n5871), .B2(n4862), .C1(n4811), 
        .C2(n6074), .ZN(U2885) );
  NOR2_X1 U5963 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4812), .ZN(n4844)
         );
  INV_X1 U5964 ( .A(n4844), .ZN(n4857) );
  AOI211_X1 U5965 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4857), .A(n5147), .B(
        n4813), .ZN(n4816) );
  NAND2_X1 U5966 ( .A1(n6395), .A2(n4999), .ZN(n6458) );
  INV_X1 U5967 ( .A(n6458), .ZN(n6442) );
  NOR3_X1 U5968 ( .A1(n6442), .A2(n4859), .A3(n6400), .ZN(n4814) );
  OAI22_X1 U5969 ( .A1(n4814), .A2(n5142), .B1(n5006), .B2(n4817), .ZN(n4815)
         );
  NAND2_X1 U5970 ( .A1(n4816), .A2(n4815), .ZN(n4855) );
  NOR2_X1 U5971 ( .A1(n4817), .A2(n6400), .ZN(n4998) );
  NAND2_X1 U5972 ( .A1(n4998), .A2(n6344), .ZN(n4820) );
  NAND2_X1 U5973 ( .A1(n4818), .A2(n4996), .ZN(n4819) );
  AND2_X1 U5974 ( .A1(n4820), .A2(n4819), .ZN(n4856) );
  OAI22_X1 U5975 ( .A1(n5171), .A2(n4857), .B1(n4856), .B2(n5170), .ZN(n4821)
         );
  INV_X1 U5976 ( .A(n4821), .ZN(n4823) );
  INV_X1 U5977 ( .A(n6315), .ZN(n6418) );
  NAND2_X1 U5978 ( .A1(n4859), .A2(n6418), .ZN(n4822) );
  OAI211_X1 U5979 ( .C1(n6458), .C2(n6422), .A(n4823), .B(n4822), .ZN(n4824)
         );
  AOI21_X1 U5980 ( .B1(n4855), .B2(INSTQUEUE_REG_12__2__SCAN_IN), .A(n4824), 
        .ZN(n4825) );
  INV_X1 U5981 ( .A(n4825), .ZN(U3118) );
  OAI22_X1 U5982 ( .A1(n5198), .A2(n4857), .B1(n4856), .B2(n5195), .ZN(n4826)
         );
  INV_X1 U5983 ( .A(n4826), .ZN(n4828) );
  INV_X1 U5984 ( .A(n6434), .ZN(n6365) );
  NAND2_X1 U5985 ( .A1(n4859), .A2(n6365), .ZN(n4827) );
  OAI211_X1 U5986 ( .C1(n6458), .C2(n6369), .A(n4828), .B(n4827), .ZN(n4829)
         );
  AOI21_X1 U5987 ( .B1(n4855), .B2(INSTQUEUE_REG_12__4__SCAN_IN), .A(n4829), 
        .ZN(n4830) );
  INV_X1 U5988 ( .A(n4830), .ZN(U3120) );
  AOI22_X1 U5989 ( .A1(n6441), .A2(n4844), .B1(n6443), .B2(n4859), .ZN(n4832)
         );
  INV_X1 U5990 ( .A(n4856), .ZN(n4845) );
  NAND2_X1 U5991 ( .A1(n6444), .A2(n4845), .ZN(n4831) );
  OAI211_X1 U5992 ( .C1(n6458), .C2(n6448), .A(n4832), .B(n4831), .ZN(n4833)
         );
  AOI21_X1 U5993 ( .B1(n4855), .B2(INSTQUEUE_REG_12__6__SCAN_IN), .A(n4833), 
        .ZN(n4834) );
  INV_X1 U5994 ( .A(n4834), .ZN(U3122) );
  AOI22_X1 U5995 ( .A1(n6411), .A2(n4844), .B1(n6354), .B2(n4859), .ZN(n4836)
         );
  NAND2_X1 U5996 ( .A1(n6413), .A2(n4845), .ZN(n4835) );
  OAI211_X1 U5997 ( .C1(n6458), .C2(n6357), .A(n4836), .B(n4835), .ZN(n4837)
         );
  AOI21_X1 U5998 ( .B1(n4855), .B2(INSTQUEUE_REG_12__1__SCAN_IN), .A(n4837), 
        .ZN(n4838) );
  INV_X1 U5999 ( .A(n4838), .ZN(U3117) );
  OAI22_X1 U6000 ( .A1(n5189), .A2(n4857), .B1(n4856), .B2(n5188), .ZN(n4839)
         );
  INV_X1 U6001 ( .A(n4839), .ZN(n4841) );
  INV_X1 U6002 ( .A(n6440), .ZN(n6320) );
  NAND2_X1 U6003 ( .A1(n4859), .A2(n6320), .ZN(n4840) );
  OAI211_X1 U6004 ( .C1(n6458), .C2(n6324), .A(n4841), .B(n4840), .ZN(n4842)
         );
  AOI21_X1 U6005 ( .B1(n4855), .B2(INSTQUEUE_REG_12__5__SCAN_IN), .A(n4842), 
        .ZN(n4843) );
  INV_X1 U6006 ( .A(n4843), .ZN(U3121) );
  AOI22_X1 U6007 ( .A1(n6450), .A2(n4844), .B1(n5150), .B2(n4859), .ZN(n4847)
         );
  NAND2_X1 U6008 ( .A1(n6454), .A2(n4845), .ZN(n4846) );
  OAI211_X1 U6009 ( .C1(n6458), .C2(n5153), .A(n4847), .B(n4846), .ZN(n4848)
         );
  AOI21_X1 U6010 ( .B1(n4855), .B2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n4848), 
        .ZN(n4849) );
  INV_X1 U6011 ( .A(n4849), .ZN(U3123) );
  OAI22_X1 U6012 ( .A1(n5177), .A2(n4857), .B1(n4856), .B2(n5176), .ZN(n4850)
         );
  INV_X1 U6013 ( .A(n4850), .ZN(n4852) );
  INV_X1 U6014 ( .A(n6363), .ZN(n6424) );
  NAND2_X1 U6015 ( .A1(n4859), .A2(n6424), .ZN(n4851) );
  OAI211_X1 U6016 ( .C1(n6458), .C2(n6428), .A(n4852), .B(n4851), .ZN(n4853)
         );
  AOI21_X1 U6017 ( .B1(n4855), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n4853), 
        .ZN(n4854) );
  INV_X1 U6018 ( .A(n4854), .ZN(U3119) );
  NAND2_X1 U6019 ( .A1(n4855), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4861)
         );
  INV_X1 U6020 ( .A(n6410), .ZN(n6298) );
  OAI22_X1 U6021 ( .A1(n5183), .A2(n4857), .B1(n4856), .B2(n5182), .ZN(n4858)
         );
  AOI21_X1 U6022 ( .B1(n6298), .B2(n4859), .A(n4858), .ZN(n4860) );
  OAI211_X1 U6023 ( .C1(n6458), .C2(n6309), .A(n4861), .B(n4860), .ZN(U3116)
         );
  OAI222_X1 U6024 ( .A1(n6015), .A2(n5499), .B1(n4863), .B2(n5497), .C1(n5460), 
        .C2(n4862), .ZN(U2853) );
  XNOR2_X1 U6025 ( .A(n4864), .B(n4865), .ZN(n5051) );
  AOI21_X1 U6026 ( .B1(n4867), .B2(n4866), .A(n4946), .ZN(n6246) );
  AOI22_X1 U6027 ( .A1(n6622), .A2(n6246), .B1(n6625), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4868) );
  OAI21_X1 U6028 ( .B1(n5051), .B2(n5460), .A(n4868), .ZN(U2852) );
  OAI21_X1 U6029 ( .B1(n4871), .B2(n4870), .A(n4869), .ZN(n6255) );
  OAI22_X1 U6030 ( .A1(n5652), .A2(n4872), .B1(n5907), .B2(n6535), .ZN(n4874)
         );
  NOR2_X1 U6031 ( .A1(n6025), .A2(n6173), .ZN(n4873) );
  AOI211_X1 U6032 ( .C1(n5657), .C2(n6028), .A(n4874), .B(n4873), .ZN(n4875)
         );
  OAI21_X1 U6033 ( .B1(n6178), .B2(n6255), .A(n4875), .ZN(U2981) );
  OAI21_X1 U6034 ( .B1(n4916), .B2(n5024), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4877) );
  NAND3_X1 U6035 ( .A1(n4877), .A2(n6396), .A3(n4876), .ZN(n4883) );
  NOR2_X1 U6036 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4878), .ZN(n5025)
         );
  INV_X1 U6037 ( .A(n5025), .ZN(n4914) );
  NOR2_X1 U6038 ( .A1(n4880), .A2(n4879), .ZN(n4997) );
  OAI21_X1 U6039 ( .B1(n4997), .B2(n3407), .A(n4881), .ZN(n5007) );
  AOI211_X1 U6040 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4914), .A(n4996), .B(
        n5007), .ZN(n4882) );
  AOI22_X1 U6041 ( .A1(n6411), .A2(n5025), .B1(n6412), .B2(n5024), .ZN(n4888)
         );
  NAND2_X1 U6042 ( .A1(n4884), .A2(n6396), .ZN(n4886) );
  NAND2_X1 U6043 ( .A1(n5147), .A2(n4997), .ZN(n4885) );
  NAND2_X1 U6044 ( .A1(n4886), .A2(n4885), .ZN(n5026) );
  NAND2_X1 U6045 ( .A1(n6413), .A2(n5026), .ZN(n4887) );
  OAI211_X1 U6046 ( .C1(n5029), .C2(n6416), .A(n4888), .B(n4887), .ZN(n4889)
         );
  INV_X1 U6047 ( .A(n4889), .ZN(n4890) );
  OAI21_X1 U6048 ( .B1(n5019), .B2(n4891), .A(n4890), .ZN(U3021) );
  NAND2_X1 U6049 ( .A1(n5024), .A2(n6312), .ZN(n4893) );
  NAND2_X1 U6050 ( .A1(n5026), .A2(n6419), .ZN(n4892) );
  OAI211_X1 U6051 ( .C1(n5171), .C2(n4914), .A(n4893), .B(n4892), .ZN(n4894)
         );
  AOI21_X1 U6052 ( .B1(n4916), .B2(n6418), .A(n4894), .ZN(n4895) );
  OAI21_X1 U6053 ( .B1(n5019), .B2(n4896), .A(n4895), .ZN(U3022) );
  NAND2_X1 U6054 ( .A1(n5024), .A2(n6394), .ZN(n4898) );
  NAND2_X1 U6055 ( .A1(n5026), .A2(n6407), .ZN(n4897) );
  OAI211_X1 U6056 ( .C1(n5183), .C2(n4914), .A(n4898), .B(n4897), .ZN(n4899)
         );
  AOI21_X1 U6057 ( .B1(n4916), .B2(n6298), .A(n4899), .ZN(n4900) );
  OAI21_X1 U6058 ( .B1(n5019), .B2(n4901), .A(n4900), .ZN(U3020) );
  NAND2_X1 U6059 ( .A1(n5024), .A2(n6430), .ZN(n4903) );
  NAND2_X1 U6060 ( .A1(n5026), .A2(n6431), .ZN(n4902) );
  OAI211_X1 U6061 ( .C1(n5198), .C2(n4914), .A(n4903), .B(n4902), .ZN(n4904)
         );
  AOI21_X1 U6062 ( .B1(n4916), .B2(n6365), .A(n4904), .ZN(n4905) );
  OAI21_X1 U6063 ( .B1(n5019), .B2(n4906), .A(n4905), .ZN(U3024) );
  NAND2_X1 U6064 ( .A1(n5024), .A2(n6436), .ZN(n4908) );
  NAND2_X1 U6065 ( .A1(n5026), .A2(n6437), .ZN(n4907) );
  OAI211_X1 U6066 ( .C1(n5189), .C2(n4914), .A(n4908), .B(n4907), .ZN(n4909)
         );
  AOI21_X1 U6067 ( .B1(n4916), .B2(n6320), .A(n4909), .ZN(n4910) );
  OAI21_X1 U6068 ( .B1(n5019), .B2(n4911), .A(n4910), .ZN(U3025) );
  INV_X1 U6069 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6070 ( .A1(n5024), .A2(n6360), .ZN(n4913) );
  NAND2_X1 U6071 ( .A1(n5026), .A2(n6425), .ZN(n4912) );
  OAI211_X1 U6072 ( .C1(n5177), .C2(n4914), .A(n4913), .B(n4912), .ZN(n4915)
         );
  AOI21_X1 U6073 ( .B1(n4916), .B2(n6424), .A(n4915), .ZN(n4917) );
  OAI21_X1 U6074 ( .B1(n5019), .B2(n4918), .A(n4917), .ZN(U3023) );
  INV_X1 U6075 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4922) );
  INV_X1 U6076 ( .A(n5024), .ZN(n4936) );
  AOI22_X1 U6077 ( .A1(n6417), .A2(n4934), .B1(n6419), .B2(n4933), .ZN(n4919)
         );
  OAI21_X1 U6078 ( .B1(n6315), .B2(n4936), .A(n4919), .ZN(n4920) );
  AOI21_X1 U6079 ( .B1(n6312), .B2(n4938), .A(n4920), .ZN(n4921) );
  OAI21_X1 U6080 ( .B1(n4941), .B2(n4922), .A(n4921), .ZN(U3142) );
  AOI22_X1 U6081 ( .A1(n6393), .A2(n4934), .B1(n6407), .B2(n4933), .ZN(n4923)
         );
  OAI21_X1 U6082 ( .B1(n6410), .B2(n4936), .A(n4923), .ZN(n4924) );
  AOI21_X1 U6083 ( .B1(n6394), .B2(n4938), .A(n4924), .ZN(n4925) );
  OAI21_X1 U6084 ( .B1(n4941), .B2(n6632), .A(n4925), .ZN(U3140) );
  AOI22_X1 U6085 ( .A1(n6429), .A2(n4934), .B1(n6431), .B2(n4933), .ZN(n4926)
         );
  OAI21_X1 U6086 ( .B1(n6434), .B2(n4936), .A(n4926), .ZN(n4927) );
  AOI21_X1 U6087 ( .B1(n6430), .B2(n4938), .A(n4927), .ZN(n4928) );
  OAI21_X1 U6088 ( .B1(n4941), .B2(n3160), .A(n4928), .ZN(U3144) );
  INV_X1 U6089 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4932) );
  AOI22_X1 U6090 ( .A1(n6423), .A2(n4934), .B1(n6425), .B2(n4933), .ZN(n4929)
         );
  OAI21_X1 U6091 ( .B1(n6363), .B2(n4936), .A(n4929), .ZN(n4930) );
  AOI21_X1 U6092 ( .B1(n6360), .B2(n4938), .A(n4930), .ZN(n4931) );
  OAI21_X1 U6093 ( .B1(n4941), .B2(n4932), .A(n4931), .ZN(U3143) );
  INV_X1 U6094 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4940) );
  AOI22_X1 U6095 ( .A1(n6435), .A2(n4934), .B1(n6437), .B2(n4933), .ZN(n4935)
         );
  OAI21_X1 U6096 ( .B1(n6440), .B2(n4936), .A(n4935), .ZN(n4937) );
  AOI21_X1 U6097 ( .B1(n6436), .B2(n4938), .A(n4937), .ZN(n4939) );
  OAI21_X1 U6098 ( .B1(n4941), .B2(n4940), .A(n4939), .ZN(U3145) );
  OAI21_X1 U6099 ( .B1(n4942), .B2(n4944), .A(n4943), .ZN(n6004) );
  NOR2_X1 U6100 ( .A1(n4946), .A2(n4945), .ZN(n4947) );
  OR2_X1 U6101 ( .A1(n5986), .A2(n4947), .ZN(n6002) );
  INV_X1 U6102 ( .A(n6002), .ZN(n6240) );
  AOI22_X1 U6103 ( .A1(n6622), .A2(n6240), .B1(n6625), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4948) );
  OAI21_X1 U6104 ( .B1(n6004), .B2(n5460), .A(n4948), .ZN(U2851) );
  AOI22_X1 U6105 ( .A1(n6071), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6067), .ZN(n4949) );
  OAI21_X1 U6106 ( .B1(n6004), .B2(n5871), .A(n4949), .ZN(U2883) );
  OAI21_X1 U6107 ( .B1(n4952), .B2(n4951), .A(n4950), .ZN(n4953) );
  INV_X1 U6108 ( .A(n4953), .ZN(n6248) );
  NAND2_X1 U6109 ( .A1(n6248), .A2(n6199), .ZN(n4956) );
  AND2_X1 U6110 ( .A1(n6206), .A2(REIP_REG_7__SCAN_IN), .ZN(n6245) );
  NOR2_X1 U6111 ( .A1(n6204), .A2(n5048), .ZN(n4954) );
  AOI211_X1 U6112 ( .C1(n6194), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6245), 
        .B(n4954), .ZN(n4955) );
  OAI211_X1 U6113 ( .C1(n5051), .C2(n6173), .A(n4956), .B(n4955), .ZN(U2979)
         );
  INV_X1 U6114 ( .A(DATAI_7_), .ZN(n6109) );
  OAI222_X1 U6115 ( .A1(n5521), .A2(n6109), .B1(n5871), .B2(n5051), .C1(n4957), 
        .C2(n6074), .ZN(U2884) );
  NAND2_X1 U6116 ( .A1(n4964), .A2(n6447), .ZN(n4958) );
  AOI21_X1 U6117 ( .B1(n4958), .B2(STATEBS16_REG_SCAN_IN), .A(n6400), .ZN(
        n4962) );
  NOR2_X1 U6118 ( .A1(n4385), .A2(n6049), .ZN(n5140) );
  AND2_X1 U6119 ( .A1(n5140), .A2(n6344), .ZN(n6399) );
  AOI22_X1 U6120 ( .A1(n4962), .A2(n6399), .B1(n5147), .B2(n4959), .ZN(n4995)
         );
  NOR2_X1 U6121 ( .A1(n4996), .A2(n4960), .ZN(n5144) );
  INV_X1 U6122 ( .A(n6399), .ZN(n4961) );
  NAND3_X1 U6123 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6469), .ZN(n6404) );
  OR2_X1 U6124 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6404), .ZN(n4990)
         );
  AOI22_X1 U6125 ( .A1(n4962), .A2(n4961), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4990), .ZN(n4963) );
  OAI211_X1 U6126 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n3407), .A(n5144), .B(n4963), .ZN(n4989) );
  NAND2_X1 U6127 ( .A1(n4989), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4968)
         );
  OAI22_X1 U6128 ( .A1(n6447), .A2(n6459), .B1(n4965), .B2(n4990), .ZN(n4966)
         );
  AOI21_X1 U6129 ( .B1(n4992), .B2(n6451), .A(n4966), .ZN(n4967) );
  OAI211_X1 U6130 ( .C1(n4995), .C2(n5015), .A(n4968), .B(n4967), .ZN(U3107)
         );
  NAND2_X1 U6131 ( .A1(n4989), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4971)
         );
  OAI22_X1 U6132 ( .A1(n6447), .A2(n6440), .B1(n5189), .B2(n4990), .ZN(n4969)
         );
  AOI21_X1 U6133 ( .B1(n4992), .B2(n6436), .A(n4969), .ZN(n4970) );
  OAI211_X1 U6134 ( .C1(n4995), .C2(n5188), .A(n4971), .B(n4970), .ZN(U3105)
         );
  NAND2_X1 U6135 ( .A1(n4989), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4975)
         );
  OAI22_X1 U6136 ( .A1(n6447), .A2(n6416), .B1(n4972), .B2(n4990), .ZN(n4973)
         );
  AOI21_X1 U6137 ( .B1(n4992), .B2(n6412), .A(n4973), .ZN(n4974) );
  OAI211_X1 U6138 ( .C1(n4995), .C2(n5012), .A(n4975), .B(n4974), .ZN(U3101)
         );
  NAND2_X1 U6139 ( .A1(n4989), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4978)
         );
  OAI22_X1 U6140 ( .A1(n6447), .A2(n6363), .B1(n5177), .B2(n4990), .ZN(n4976)
         );
  AOI21_X1 U6141 ( .B1(n4992), .B2(n6360), .A(n4976), .ZN(n4977) );
  OAI211_X1 U6142 ( .C1(n4995), .C2(n5176), .A(n4978), .B(n4977), .ZN(U3103)
         );
  NAND2_X1 U6143 ( .A1(n4989), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4981)
         );
  OAI22_X1 U6144 ( .A1(n6447), .A2(n6434), .B1(n5198), .B2(n4990), .ZN(n4979)
         );
  AOI21_X1 U6145 ( .B1(n4992), .B2(n6430), .A(n4979), .ZN(n4980) );
  OAI211_X1 U6146 ( .C1(n4995), .C2(n5195), .A(n4981), .B(n4980), .ZN(U3104)
         );
  NAND2_X1 U6147 ( .A1(n4989), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4985)
         );
  OAI22_X1 U6148 ( .A1(n6447), .A2(n6375), .B1(n4982), .B2(n4990), .ZN(n4983)
         );
  AOI21_X1 U6149 ( .B1(n4992), .B2(n6372), .A(n4983), .ZN(n4984) );
  OAI211_X1 U6150 ( .C1(n4995), .C2(n5018), .A(n4985), .B(n4984), .ZN(U3106)
         );
  NAND2_X1 U6151 ( .A1(n4989), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4988)
         );
  OAI22_X1 U6152 ( .A1(n6447), .A2(n6315), .B1(n5171), .B2(n4990), .ZN(n4986)
         );
  AOI21_X1 U6153 ( .B1(n4992), .B2(n6312), .A(n4986), .ZN(n4987) );
  OAI211_X1 U6154 ( .C1(n4995), .C2(n5170), .A(n4988), .B(n4987), .ZN(U3102)
         );
  NAND2_X1 U6155 ( .A1(n4989), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4994)
         );
  OAI22_X1 U6156 ( .A1(n6447), .A2(n6410), .B1(n5183), .B2(n4990), .ZN(n4991)
         );
  AOI21_X1 U6157 ( .B1(n4992), .B2(n6394), .A(n4991), .ZN(n4993) );
  OAI211_X1 U6158 ( .C1(n4995), .C2(n5182), .A(n4994), .B(n4993), .ZN(U3100)
         );
  AOI22_X1 U6159 ( .A1(n4998), .A2(n5812), .B1(n4997), .B2(n4996), .ZN(n5082)
         );
  INV_X1 U6160 ( .A(n4999), .ZN(n5000) );
  INV_X1 U6161 ( .A(n6334), .ZN(n6321) );
  AOI22_X1 U6162 ( .A1(n6321), .A2(n6412), .B1(n5100), .B2(n6354), .ZN(n5011)
         );
  NOR2_X1 U6163 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5001), .ZN(n5081)
         );
  AOI21_X1 U6164 ( .B1(n5003), .B2(n6334), .A(n5002), .ZN(n5004) );
  AOI211_X1 U6165 ( .C1(n5006), .C2(n5005), .A(n5004), .B(n6400), .ZN(n5008)
         );
  NOR3_X1 U6166 ( .A1(n5147), .A2(n5008), .A3(n5007), .ZN(n5009) );
  AOI22_X1 U6167 ( .A1(n6411), .A2(n5081), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5095), .ZN(n5010) );
  OAI211_X1 U6168 ( .C1(n5082), .C2(n5012), .A(n5011), .B(n5010), .ZN(U3053)
         );
  AOI22_X1 U6169 ( .A1(n6321), .A2(n6451), .B1(n5100), .B2(n5150), .ZN(n5014)
         );
  AOI22_X1 U6170 ( .A1(n6450), .A2(n5081), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5095), .ZN(n5013) );
  OAI211_X1 U6171 ( .C1(n5082), .C2(n5015), .A(n5014), .B(n5013), .ZN(U3059)
         );
  AOI22_X1 U6172 ( .A1(n6321), .A2(n6372), .B1(n5100), .B2(n6443), .ZN(n5017)
         );
  AOI22_X1 U6173 ( .A1(n6441), .A2(n5081), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5095), .ZN(n5016) );
  OAI211_X1 U6174 ( .C1(n5082), .C2(n5018), .A(n5017), .B(n5016), .ZN(U3058)
         );
  INV_X1 U6175 ( .A(n5019), .ZN(n5031) );
  AOI22_X1 U6176 ( .A1(n6450), .A2(n5025), .B1(n6451), .B2(n5024), .ZN(n5021)
         );
  NAND2_X1 U6177 ( .A1(n6454), .A2(n5026), .ZN(n5020) );
  OAI211_X1 U6178 ( .C1(n5029), .C2(n6459), .A(n5021), .B(n5020), .ZN(n5022)
         );
  AOI21_X1 U6179 ( .B1(n5031), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n5022), 
        .ZN(n5023) );
  INV_X1 U6180 ( .A(n5023), .ZN(U3027) );
  AOI22_X1 U6181 ( .A1(n6441), .A2(n5025), .B1(n6372), .B2(n5024), .ZN(n5028)
         );
  NAND2_X1 U6182 ( .A1(n6444), .A2(n5026), .ZN(n5027) );
  OAI211_X1 U6183 ( .C1(n5029), .C2(n6375), .A(n5028), .B(n5027), .ZN(n5030)
         );
  AOI21_X1 U6184 ( .B1(n5031), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n5030), 
        .ZN(n5032) );
  INV_X1 U6185 ( .A(n5032), .ZN(U3026) );
  NOR2_X1 U6186 ( .A1(n5370), .A2(n5033), .ZN(n6023) );
  AND2_X1 U6187 ( .A1(n5034), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6188 ( .A1(n3281), .A2(n6491), .ZN(n5039) );
  NOR2_X1 U6189 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5036), .ZN(n5037) );
  NAND2_X1 U6190 ( .A1(n3271), .A2(n5037), .ZN(n5038) );
  NAND2_X1 U6191 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  AND2_X2 U6192 ( .A1(n5040), .A2(n5052), .ZN(n6056) );
  INV_X1 U6193 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5045) );
  INV_X1 U6194 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6540) );
  INV_X1 U6195 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U6196 ( .A1(n6540), .A2(n6537), .ZN(n6000) );
  AOI21_X1 U6197 ( .B1(n6540), .B2(n6537), .A(n6000), .ZN(n5041) );
  AOI22_X1 U6198 ( .A1(n6045), .A2(n6246), .B1(n6017), .B2(n5041), .ZN(n5044)
         );
  NAND2_X1 U6199 ( .A1(n5043), .A2(n5042), .ZN(n6030) );
  OAI211_X1 U6200 ( .C1(n6051), .C2(n5045), .A(n5044), .B(n6030), .ZN(n5046)
         );
  AOI21_X1 U6201 ( .B1(n6056), .B2(EBX_REG_7__SCAN_IN), .A(n5046), .ZN(n5047)
         );
  OAI21_X1 U6202 ( .B1(n6061), .B2(n5048), .A(n5047), .ZN(n5049) );
  AOI21_X1 U6203 ( .B1(n6023), .B2(REIP_REG_7__SCAN_IN), .A(n5049), .ZN(n5050)
         );
  OAI21_X1 U6204 ( .B1(n5051), .B2(n5977), .A(n5050), .ZN(U2820) );
  NAND2_X1 U6205 ( .A1(n5053), .A2(n5052), .ZN(n5054) );
  INV_X1 U6206 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6530) );
  AOI211_X1 U6207 ( .C1(n6044), .C2(n6600), .A(n6054), .B(n6530), .ZN(n5064)
         );
  AOI221_X1 U6208 ( .B1(n6600), .B2(n6530), .C1(n5055), .C2(n6530), .A(n5064), 
        .ZN(n5056) );
  INV_X1 U6209 ( .A(n5056), .ZN(n5062) );
  AOI22_X1 U6210 ( .A1(n6285), .A2(n6045), .B1(n6056), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5059) );
  NOR2_X1 U6211 ( .A1(n5057), .A2(n3051), .ZN(n5102) );
  NAND2_X1 U6212 ( .A1(n4385), .A2(n5102), .ZN(n5058) );
  OAI211_X1 U6213 ( .C1(n6061), .C2(n6203), .A(n5059), .B(n5058), .ZN(n5060)
         );
  AOI21_X1 U6214 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6024), .A(n5060), 
        .ZN(n5061) );
  OAI211_X1 U6215 ( .C1(n6026), .C2(n6195), .A(n5062), .B(n5061), .ZN(U2825)
         );
  AND2_X1 U6216 ( .A1(n5379), .A2(n5063), .ZN(n6034) );
  OAI21_X1 U6217 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5064), .A(n6034), .ZN(n5071)
         );
  AOI22_X1 U6218 ( .A1(n5065), .A2(n6045), .B1(n6056), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5067) );
  NAND2_X1 U6219 ( .A1(n6344), .A2(n5102), .ZN(n5066) );
  OAI211_X1 U6220 ( .C1(n6061), .C2(n5068), .A(n5067), .B(n5066), .ZN(n5069)
         );
  AOI21_X1 U6221 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6024), .A(n5069), 
        .ZN(n5070) );
  OAI211_X1 U6222 ( .C1(n6026), .C2(n5072), .A(n5071), .B(n5070), .ZN(U2824)
         );
  OAI21_X1 U6223 ( .B1(n5075), .B2(n5074), .A(n5073), .ZN(n5076) );
  INV_X1 U6224 ( .A(n5076), .ZN(n6241) );
  NAND2_X1 U6225 ( .A1(n6241), .A2(n6199), .ZN(n5080) );
  INV_X1 U6226 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5077) );
  NOR2_X1 U6227 ( .A1(n5907), .A2(n5077), .ZN(n6239) );
  NOR2_X1 U6228 ( .A1(n6204), .A2(n6005), .ZN(n5078) );
  AOI211_X1 U6229 ( .C1(n6194), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6239), 
        .B(n5078), .ZN(n5079) );
  OAI211_X1 U6230 ( .C1(n6173), .C2(n6004), .A(n5080), .B(n5079), .ZN(U2978)
         );
  INV_X1 U6231 ( .A(n5081), .ZN(n5098) );
  INV_X1 U6232 ( .A(n5082), .ZN(n5096) );
  AOI22_X1 U6233 ( .A1(n5096), .A2(n6425), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5095), .ZN(n5083) );
  OAI21_X1 U6234 ( .B1(n5177), .B2(n5098), .A(n5083), .ZN(n5084) );
  AOI21_X1 U6235 ( .B1(n6424), .B2(n5100), .A(n5084), .ZN(n5085) );
  OAI21_X1 U6236 ( .B1(n6428), .B2(n6334), .A(n5085), .ZN(U3055) );
  AOI22_X1 U6237 ( .A1(n5096), .A2(n6407), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5095), .ZN(n5086) );
  OAI21_X1 U6238 ( .B1(n5183), .B2(n5098), .A(n5086), .ZN(n5087) );
  AOI21_X1 U6239 ( .B1(n6298), .B2(n5100), .A(n5087), .ZN(n5088) );
  OAI21_X1 U6240 ( .B1(n6309), .B2(n6334), .A(n5088), .ZN(U3052) );
  AOI22_X1 U6241 ( .A1(n5096), .A2(n6419), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5095), .ZN(n5089) );
  OAI21_X1 U6242 ( .B1(n5171), .B2(n5098), .A(n5089), .ZN(n5090) );
  AOI21_X1 U6243 ( .B1(n6418), .B2(n5100), .A(n5090), .ZN(n5091) );
  OAI21_X1 U6244 ( .B1(n6422), .B2(n6334), .A(n5091), .ZN(U3054) );
  AOI22_X1 U6245 ( .A1(n5096), .A2(n6431), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5095), .ZN(n5092) );
  OAI21_X1 U6246 ( .B1(n5198), .B2(n5098), .A(n5092), .ZN(n5093) );
  AOI21_X1 U6247 ( .B1(n6365), .B2(n5100), .A(n5093), .ZN(n5094) );
  OAI21_X1 U6248 ( .B1(n6369), .B2(n6334), .A(n5094), .ZN(U3056) );
  AOI22_X1 U6249 ( .A1(n5096), .A2(n6437), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5095), .ZN(n5097) );
  OAI21_X1 U6250 ( .B1(n5189), .B2(n5098), .A(n5097), .ZN(n5099) );
  AOI21_X1 U6251 ( .B1(n6320), .B2(n5100), .A(n5099), .ZN(n5101) );
  OAI21_X1 U6252 ( .B1(n6324), .B2(n6334), .A(n5101), .ZN(U3057) );
  INV_X1 U6253 ( .A(n5102), .ZN(n6048) );
  AOI22_X1 U6254 ( .A1(n5103), .A2(n6045), .B1(n6056), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5104) );
  OAI21_X1 U6255 ( .B1(n6343), .B2(n6048), .A(n5104), .ZN(n5107) );
  AOI21_X1 U6256 ( .B1(n6051), .B2(n6061), .A(n5105), .ZN(n5106) );
  AOI211_X1 U6257 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5379), .A(n5107), .B(n5106), 
        .ZN(n5108) );
  OAI21_X1 U6258 ( .B1(n6026), .B2(n5109), .A(n5108), .ZN(U2827) );
  INV_X1 U6259 ( .A(n4943), .ZN(n5112) );
  INV_X1 U6260 ( .A(n5110), .ZN(n5111) );
  OAI21_X1 U6261 ( .B1(n5112), .B2(n5111), .A(n3018), .ZN(n5995) );
  NAND2_X1 U6262 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  XNOR2_X1 U6263 ( .A(n5113), .B(n5116), .ZN(n6233) );
  NAND2_X1 U6264 ( .A1(n6233), .A2(n6199), .ZN(n5119) );
  NAND2_X1 U6265 ( .A1(n6258), .A2(REIP_REG_9__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U6266 ( .B1(n5652), .B2(n5992), .A(n6230), .ZN(n5117) );
  AOI21_X1 U6267 ( .B1(n5657), .B2(n5996), .A(n5117), .ZN(n5118) );
  OAI211_X1 U6268 ( .C1(n6173), .C2(n5995), .A(n5119), .B(n5118), .ZN(U2977)
         );
  AND2_X1 U6269 ( .A1(n3018), .A2(n5120), .ZN(n5122) );
  OR2_X1 U6270 ( .A1(n5122), .A2(n5121), .ZN(n5210) );
  AOI22_X1 U6271 ( .A1(n6071), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6067), .ZN(n5123) );
  OAI21_X1 U6272 ( .B1(n5210), .B2(n5871), .A(n5123), .ZN(U2881) );
  INV_X1 U6273 ( .A(n5212), .ZN(n5134) );
  INV_X1 U6274 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5130) );
  INV_X1 U6275 ( .A(n5204), .ZN(n5124) );
  AOI21_X1 U6276 ( .B1(n5125), .B2(n5987), .A(n5124), .ZN(n6223) );
  OAI21_X1 U6277 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .A(
        n5126), .ZN(n5127) );
  OAI21_X1 U6278 ( .B1(n5127), .B2(n5991), .A(n6030), .ZN(n5128) );
  AOI21_X1 U6279 ( .B1(n6223), .B2(n6045), .A(n5128), .ZN(n5129) );
  OAI21_X1 U6280 ( .B1(n6051), .B2(n5130), .A(n5129), .ZN(n5133) );
  INV_X1 U6281 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U6282 ( .A1(n5379), .A2(n5131), .ZN(n6010) );
  OAI22_X1 U6283 ( .A1(n5846), .A2(n4195), .B1(n6545), .B2(n6010), .ZN(n5132)
         );
  AOI211_X1 U6284 ( .C1(n6027), .C2(n5134), .A(n5133), .B(n5132), .ZN(n5135)
         );
  OAI21_X1 U6285 ( .B1(n5977), .B2(n5210), .A(n5135), .ZN(U2817) );
  INV_X1 U6286 ( .A(n6223), .ZN(n5136) );
  OAI222_X1 U6287 ( .A1(n5210), .A2(n5460), .B1(n5497), .B2(n4195), .C1(n5136), 
        .C2(n5499), .ZN(U2849) );
  NAND3_X1 U6288 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6391), .A3(n6469), .ZN(n6304) );
  NOR2_X1 U6289 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6304), .ZN(n5169)
         );
  INV_X1 U6290 ( .A(n5203), .ZN(n5139) );
  INV_X1 U6291 ( .A(n5137), .ZN(n5138) );
  NOR2_X1 U6292 ( .A1(n5139), .A2(n6329), .ZN(n5143) );
  INV_X1 U6293 ( .A(n6301), .ZN(n5141) );
  OAI21_X1 U6294 ( .B1(n5143), .B2(n5142), .A(n5141), .ZN(n5145) );
  OAI221_X1 U6295 ( .B1(n5169), .B2(n6591), .C1(n5169), .C2(n5145), .A(n5144), 
        .ZN(n5194) );
  NAND2_X1 U6296 ( .A1(n6301), .A2(n6396), .ZN(n5149) );
  NAND2_X1 U6297 ( .A1(n5147), .A2(n5146), .ZN(n5148) );
  AND2_X1 U6298 ( .A1(n5149), .A2(n5148), .ZN(n5196) );
  INV_X1 U6299 ( .A(n5196), .ZN(n5160) );
  AOI22_X1 U6300 ( .A1(n6454), .A2(n5160), .B1(n6450), .B2(n5169), .ZN(n5152)
         );
  NAND2_X1 U6301 ( .A1(n6329), .A2(n5150), .ZN(n5151) );
  OAI211_X1 U6302 ( .C1(n5203), .C2(n5153), .A(n5152), .B(n5151), .ZN(n5154)
         );
  AOI21_X1 U6303 ( .B1(n5194), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n5154), 
        .ZN(n5155) );
  INV_X1 U6304 ( .A(n5155), .ZN(U3043) );
  AOI22_X1 U6305 ( .A1(n6413), .A2(n5160), .B1(n6411), .B2(n5169), .ZN(n5157)
         );
  NAND2_X1 U6306 ( .A1(n6329), .A2(n6354), .ZN(n5156) );
  OAI211_X1 U6307 ( .C1(n5203), .C2(n6357), .A(n5157), .B(n5156), .ZN(n5158)
         );
  AOI21_X1 U6308 ( .B1(n5194), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n5158), 
        .ZN(n5159) );
  INV_X1 U6309 ( .A(n5159), .ZN(U3037) );
  AOI22_X1 U6310 ( .A1(n6444), .A2(n5160), .B1(n6441), .B2(n5169), .ZN(n5162)
         );
  NAND2_X1 U6311 ( .A1(n6329), .A2(n6443), .ZN(n5161) );
  OAI211_X1 U6312 ( .C1(n5203), .C2(n6448), .A(n5162), .B(n5161), .ZN(n5163)
         );
  AOI21_X1 U6313 ( .B1(n5194), .B2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n5163), 
        .ZN(n5164) );
  INV_X1 U6314 ( .A(n5164), .ZN(U3042) );
  NOR2_X1 U6315 ( .A1(n5121), .A2(n5166), .ZN(n5167) );
  OR2_X1 U6316 ( .A1(n5165), .A2(n5167), .ZN(n6174) );
  AOI22_X1 U6317 ( .A1(n6071), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6067), .ZN(n5168) );
  OAI21_X1 U6318 ( .B1(n6174), .B2(n5871), .A(n5168), .ZN(U2880) );
  NAND2_X1 U6319 ( .A1(n5194), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5175) );
  NOR2_X1 U6320 ( .A1(n6325), .A2(n6315), .ZN(n5173) );
  INV_X1 U6321 ( .A(n5169), .ZN(n5197) );
  OAI22_X1 U6322 ( .A1(n5171), .A2(n5197), .B1(n5196), .B2(n5170), .ZN(n5172)
         );
  NOR2_X1 U6323 ( .A1(n5173), .A2(n5172), .ZN(n5174) );
  OAI211_X1 U6324 ( .C1(n5203), .C2(n6422), .A(n5175), .B(n5174), .ZN(U3038)
         );
  NAND2_X1 U6325 ( .A1(n5194), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5181) );
  NOR2_X1 U6326 ( .A1(n6325), .A2(n6363), .ZN(n5179) );
  OAI22_X1 U6327 ( .A1(n5177), .A2(n5197), .B1(n5196), .B2(n5176), .ZN(n5178)
         );
  NOR2_X1 U6328 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  OAI211_X1 U6329 ( .C1(n5203), .C2(n6428), .A(n5181), .B(n5180), .ZN(U3039)
         );
  NAND2_X1 U6330 ( .A1(n5194), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5187) );
  NOR2_X1 U6331 ( .A1(n6325), .A2(n6410), .ZN(n5185) );
  OAI22_X1 U6332 ( .A1(n5183), .A2(n5197), .B1(n5196), .B2(n5182), .ZN(n5184)
         );
  NOR2_X1 U6333 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  OAI211_X1 U6334 ( .C1(n6309), .C2(n5203), .A(n5187), .B(n5186), .ZN(U3036)
         );
  NAND2_X1 U6335 ( .A1(n5194), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5193) );
  NOR2_X1 U6336 ( .A1(n6325), .A2(n6440), .ZN(n5191) );
  OAI22_X1 U6337 ( .A1(n5189), .A2(n5197), .B1(n5196), .B2(n5188), .ZN(n5190)
         );
  NOR2_X1 U6338 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  OAI211_X1 U6339 ( .C1(n5203), .C2(n6324), .A(n5193), .B(n5192), .ZN(U3041)
         );
  NAND2_X1 U6340 ( .A1(n5194), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5202) );
  NOR2_X1 U6341 ( .A1(n6325), .A2(n6434), .ZN(n5200) );
  OAI22_X1 U6342 ( .A1(n5198), .A2(n5197), .B1(n5196), .B2(n5195), .ZN(n5199)
         );
  NOR2_X1 U6343 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  OAI211_X1 U6344 ( .C1(n5203), .C2(n6369), .A(n5202), .B(n5201), .ZN(U3040)
         );
  INV_X1 U6345 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5206) );
  AOI21_X1 U6346 ( .B1(n5205), .B2(n5204), .A(n5220), .ZN(n5975) );
  INV_X1 U6347 ( .A(n5975), .ZN(n6207) );
  OAI222_X1 U6348 ( .A1(n6174), .A2(n5460), .B1(n5206), .B2(n5497), .C1(n5499), 
        .C2(n6207), .ZN(U2848) );
  NAND2_X1 U6349 ( .A1(n6167), .A2(n5208), .ZN(n5209) );
  XNOR2_X1 U6350 ( .A(n5207), .B(n5209), .ZN(n6224) );
  INV_X1 U6351 ( .A(n6224), .ZN(n5216) );
  INV_X1 U6352 ( .A(n5210), .ZN(n5214) );
  AOI22_X1 U6353 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6206), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5211) );
  OAI21_X1 U6354 ( .B1(n6204), .B2(n5212), .A(n5211), .ZN(n5213) );
  AOI21_X1 U6355 ( .B1(n5214), .B2(n5894), .A(n5213), .ZN(n5215) );
  OAI21_X1 U6356 ( .B1(n5216), .B2(n6178), .A(n5215), .ZN(U2976) );
  XOR2_X1 U6357 ( .A(n5217), .B(n5165), .Z(n5252) );
  NOR2_X1 U6358 ( .A1(n5370), .A2(n5218), .ZN(n5979) );
  OR2_X1 U6359 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  NAND2_X1 U6360 ( .A1(n5420), .A2(n5221), .ZN(n5243) );
  INV_X1 U6361 ( .A(n6030), .ZN(n6038) );
  AOI21_X1 U6362 ( .B1(n6056), .B2(EBX_REG_12__SCAN_IN), .A(n6038), .ZN(n5222)
         );
  OAI21_X1 U6363 ( .B1(n5243), .B2(n6014), .A(n5222), .ZN(n5223) );
  AOI21_X1 U6364 ( .B1(n6024), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5223), 
        .ZN(n5224) );
  OAI21_X1 U6365 ( .B1(n6061), .B2(n5250), .A(n5224), .ZN(n5225) );
  NOR2_X1 U6366 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5429), .ZN(n5426) );
  AOI211_X1 U6367 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5979), .A(n5225), .B(n5426), .ZN(n5226) );
  OAI21_X1 U6368 ( .B1(n5230), .B2(n5977), .A(n5226), .ZN(U2815) );
  INV_X1 U6369 ( .A(n5243), .ZN(n5227) );
  AOI22_X1 U6370 ( .A1(n6622), .A2(n5227), .B1(n6625), .B2(EBX_REG_12__SCAN_IN), .ZN(n5228) );
  OAI21_X1 U6371 ( .B1(n5230), .B2(n5460), .A(n5228), .ZN(U2847) );
  INV_X1 U6372 ( .A(DATAI_12_), .ZN(n6119) );
  OAI222_X1 U6373 ( .A1(n5521), .A2(n6119), .B1(n5871), .B2(n5230), .C1(n5229), 
        .C2(n6074), .ZN(U2879) );
  INV_X1 U6374 ( .A(n5231), .ZN(n5232) );
  NOR2_X1 U6375 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  XNOR2_X1 U6376 ( .A(n5235), .B(n5234), .ZN(n5254) );
  INV_X1 U6377 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6214) );
  NOR2_X1 U6378 ( .A1(n6214), .A2(n5242), .ZN(n5791) );
  INV_X1 U6379 ( .A(n6288), .ZN(n6216) );
  INV_X1 U6380 ( .A(n6217), .ZN(n6226) );
  NAND2_X1 U6381 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U6382 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6227) );
  NOR3_X1 U6383 ( .A1(n6218), .A2(n6238), .A3(n6227), .ZN(n5236) );
  AND3_X1 U6384 ( .A1(n6226), .A2(n5236), .A3(n6284), .ZN(n5660) );
  NOR2_X1 U6385 ( .A1(n6216), .A2(n5241), .ZN(n5240) );
  NAND2_X1 U6386 ( .A1(n5237), .A2(n5236), .ZN(n5665) );
  OAI21_X1 U6387 ( .B1(n5238), .B2(n5660), .A(n6219), .ZN(n5239) );
  AOI21_X1 U6388 ( .B1(n6216), .B2(n5665), .A(n5239), .ZN(n6215) );
  OAI21_X1 U6389 ( .B1(n5791), .B2(n5240), .A(n6215), .ZN(n5246) );
  NOR2_X1 U6390 ( .A1(n6288), .A2(n5665), .ZN(n5795) );
  OAI21_X1 U6391 ( .B1(n6205), .B2(n6214), .A(n5242), .ZN(n5245) );
  NAND2_X1 U6392 ( .A1(n6258), .A2(REIP_REG_12__SCAN_IN), .ZN(n5249) );
  OAI21_X1 U6393 ( .B1(n6274), .B2(n5243), .A(n5249), .ZN(n5244) );
  AOI21_X1 U6394 ( .B1(n5246), .B2(n5245), .A(n5244), .ZN(n5247) );
  OAI21_X1 U6395 ( .B1(n5254), .B2(n6208), .A(n5247), .ZN(U3006) );
  NAND2_X1 U6396 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5248)
         );
  OAI211_X1 U6397 ( .C1(n6204), .C2(n5250), .A(n5249), .B(n5248), .ZN(n5251)
         );
  AOI21_X1 U6398 ( .B1(n5252), .B2(n5894), .A(n5251), .ZN(n5253) );
  OAI21_X1 U6399 ( .B1(n5254), .B2(n6178), .A(n5253), .ZN(U2974) );
  INV_X1 U6400 ( .A(n5256), .ZN(n5307) );
  AND2_X1 U6401 ( .A1(n3155), .A2(n5258), .ZN(n5259) );
  AOI22_X1 U6402 ( .A1(n6068), .A2(DATAI_11_), .B1(n6067), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6403 ( .A1(n6065), .A2(DATAI_27_), .ZN(n5260) );
  OAI211_X1 U6404 ( .C1(n5818), .C2(n5871), .A(n5261), .B(n5260), .ZN(U2864)
         );
  AND2_X1 U6405 ( .A1(n5442), .A2(n5262), .ZN(n5263) );
  NOR2_X1 U6406 ( .A1(n5311), .A2(n5263), .ZN(n5816) );
  INV_X1 U6407 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U6408 ( .A1(n5497), .A2(n5822), .ZN(n5264) );
  AOI21_X1 U6409 ( .B1(n5816), .B2(n6622), .A(n5264), .ZN(n5265) );
  OAI21_X1 U6410 ( .B1(n5818), .B2(n5460), .A(n5265), .ZN(U2832) );
  INV_X1 U6411 ( .A(n6598), .ZN(n5942) );
  OAI22_X1 U6412 ( .A1(n6343), .A2(n5268), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5267), .ZN(n6461) );
  AOI21_X1 U6413 ( .B1(n6461), .B2(n6591), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n5270) );
  OAI22_X1 U6414 ( .A1(n5270), .A2(n5269), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6595), .ZN(n5272) );
  NOR2_X1 U6415 ( .A1(n5271), .A2(n5266), .ZN(n6462) );
  AOI22_X1 U6416 ( .A1(n5942), .A2(n5272), .B1(n6593), .B2(n6462), .ZN(n5273)
         );
  OAI21_X1 U6417 ( .B1(n5266), .B2(n5942), .A(n5273), .ZN(U3461) );
  INV_X1 U6418 ( .A(n5528), .ZN(n5286) );
  AOI21_X1 U6419 ( .B1(n5279), .B2(n5276), .A(n5277), .ZN(n5282) );
  INV_X1 U6420 ( .A(n5277), .ZN(n5278) );
  AOI21_X1 U6421 ( .B1(n5309), .B2(n5477), .A(n5278), .ZN(n5280) );
  AOI22_X1 U6422 ( .A1(n5282), .A2(n5281), .B1(n5280), .B2(n5279), .ZN(n5690)
         );
  AOI22_X1 U6423 ( .A1(n5690), .A2(n6622), .B1(EBX_REG_30__SCAN_IN), .B2(n6625), .ZN(n5283) );
  OAI21_X1 U6424 ( .B1(n5286), .B2(n5460), .A(n5283), .ZN(U2829) );
  AOI22_X1 U6425 ( .A1(n6065), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6067), .ZN(n5285) );
  NAND2_X1 U6426 ( .A1(n6068), .A2(DATAI_14_), .ZN(n5284) );
  OAI211_X1 U6427 ( .C1(n5286), .C2(n5871), .A(n5285), .B(n5284), .ZN(U2861)
         );
  NAND2_X1 U6428 ( .A1(n5528), .A2(n6018), .ZN(n5293) );
  INV_X1 U6429 ( .A(n5287), .ZN(n5526) );
  AOI22_X1 U6430 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n6056), .ZN(n5288) );
  OAI21_X1 U6431 ( .B1(n6061), .B2(n5526), .A(n5288), .ZN(n5291) );
  NOR2_X1 U6432 ( .A1(n5289), .A2(REIP_REG_30__SCAN_IN), .ZN(n5290) );
  AOI211_X1 U6433 ( .C1(n6045), .C2(n5690), .A(n5291), .B(n5290), .ZN(n5292)
         );
  OAI211_X1 U6434 ( .C1(n5294), .C2(n6580), .A(n5293), .B(n5292), .ZN(U2797)
         );
  INV_X1 U6435 ( .A(n5296), .ZN(n5297) );
  INV_X1 U6436 ( .A(n5538), .ZN(n5505) );
  XNOR2_X1 U6437 ( .A(n5276), .B(n5299), .ZN(n5693) );
  AOI22_X1 U6438 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .B1(n6056), 
        .B2(EBX_REG_29__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6439 ( .A1(n6027), .A2(n5534), .ZN(n5300) );
  OAI211_X1 U6440 ( .C1(n5693), .C2(n6014), .A(n5301), .B(n5300), .ZN(n5303)
         );
  AOI211_X1 U6441 ( .C1(n5318), .C2(REIP_REG_29__SCAN_IN), .A(n5303), .B(n5302), .ZN(n5304) );
  OAI21_X1 U6442 ( .B1(n5505), .B2(n5977), .A(n5304), .ZN(U2798) );
  INV_X1 U6443 ( .A(n5305), .ZN(n5308) );
  OAI21_X1 U6444 ( .B1(n5311), .B2(n5310), .A(n5309), .ZN(n5702) );
  OAI22_X1 U6445 ( .A1(n5846), .A2(n5312), .B1(n5545), .B2(n6061), .ZN(n5313)
         );
  AOI21_X1 U6446 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6024), .A(n5313), 
        .ZN(n5314) );
  OAI21_X1 U6447 ( .B1(n5702), .B2(n6014), .A(n5314), .ZN(n5317) );
  NOR2_X1 U6448 ( .A1(n5315), .A2(REIP_REG_28__SCAN_IN), .ZN(n5316) );
  AOI211_X1 U6449 ( .C1(n5318), .C2(REIP_REG_28__SCAN_IN), .A(n5317), .B(n5316), .ZN(n5319) );
  OAI21_X1 U6450 ( .B1(n5508), .B2(n5977), .A(n5319), .ZN(U2799) );
  OAI21_X1 U6451 ( .B1(n5320), .B2(n5322), .A(n5443), .ZN(n5576) );
  OAI21_X1 U6452 ( .B1(n5335), .B2(n5324), .A(n5323), .ZN(n5449) );
  INV_X1 U6453 ( .A(n5578), .ZN(n5325) );
  AOI22_X1 U6454 ( .A1(n6027), .A2(n5325), .B1(n6056), .B2(EBX_REG_24__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6455 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5326)
         );
  OAI211_X1 U6456 ( .C1(n5449), .C2(n6014), .A(n5327), .B(n5326), .ZN(n5328)
         );
  AOI21_X1 U6457 ( .B1(n5832), .B2(REIP_REG_24__SCAN_IN), .A(n5328), .ZN(n5330) );
  INV_X1 U6458 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U6459 ( .A1(n5836), .A2(n6688), .ZN(n5329) );
  OAI211_X1 U6460 ( .C1(n5576), .C2(n5977), .A(n5330), .B(n5329), .ZN(U2803)
         );
  XOR2_X1 U6461 ( .A(n5332), .B(n5331), .Z(n5587) );
  INV_X1 U6462 ( .A(n5587), .ZN(n5513) );
  AND2_X1 U6463 ( .A1(n5351), .A2(n5333), .ZN(n5334) );
  NOR2_X1 U6464 ( .A1(n5335), .A2(n5334), .ZN(n5750) );
  INV_X1 U6465 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5451) );
  OAI22_X1 U6466 ( .A1(n5846), .A2(n5451), .B1(n5336), .B2(n6051), .ZN(n5339)
         );
  INV_X1 U6467 ( .A(n5337), .ZN(n5585) );
  NOR2_X1 U6468 ( .A1(n6061), .A2(n5585), .ZN(n5338) );
  AOI211_X1 U6469 ( .C1(n5750), .C2(n6045), .A(n5339), .B(n5338), .ZN(n5343)
         );
  NAND2_X1 U6470 ( .A1(n6565), .A2(n5340), .ZN(n5341) );
  NAND2_X1 U6471 ( .A1(n5341), .A2(n5832), .ZN(n5342) );
  OAI211_X1 U6472 ( .C1(n5513), .C2(n5977), .A(n5343), .B(n5342), .ZN(U2804)
         );
  AOI21_X1 U6473 ( .B1(n5345), .B2(n5344), .A(n5331), .ZN(n5878) );
  INV_X1 U6474 ( .A(n5878), .ZN(n5457) );
  OAI211_X1 U6475 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5848), .B(n5346), .ZN(n5359) );
  NAND2_X1 U6476 ( .A1(n5379), .A2(n5347), .ZN(n5853) );
  INV_X1 U6477 ( .A(n5853), .ZN(n5849) );
  NAND2_X1 U6478 ( .A1(n5348), .A2(n5349), .ZN(n5350) );
  AND2_X1 U6479 ( .A1(n5351), .A2(n5350), .ZN(n5755) );
  INV_X1 U6480 ( .A(n5755), .ZN(n5356) );
  INV_X1 U6481 ( .A(n5593), .ZN(n5354) );
  INV_X1 U6482 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5352) );
  OAI22_X1 U6483 ( .A1(n6051), .A2(n5352), .B1(n5454), .B2(n5846), .ZN(n5353)
         );
  AOI21_X1 U6484 ( .B1(n5354), .B2(n6027), .A(n5353), .ZN(n5355) );
  OAI21_X1 U6485 ( .B1(n5356), .B2(n6014), .A(n5355), .ZN(n5357) );
  AOI21_X1 U6486 ( .B1(n5849), .B2(REIP_REG_22__SCAN_IN), .A(n5357), .ZN(n5358) );
  OAI211_X1 U6487 ( .C1(n5457), .C2(n5977), .A(n5359), .B(n5358), .ZN(U2805)
         );
  INV_X1 U6488 ( .A(n5361), .ZN(n5362) );
  AOI21_X1 U6489 ( .B1(n5363), .B2(n5360), .A(n5362), .ZN(n5624) );
  INV_X1 U6490 ( .A(n5624), .ZN(n5518) );
  INV_X1 U6491 ( .A(n5364), .ZN(n5365) );
  AOI21_X1 U6492 ( .B1(n5366), .B2(n5383), .A(n5364), .ZN(n5905) );
  AOI22_X1 U6493 ( .A1(EBX_REG_17__SCAN_IN), .A2(n6056), .B1(n5620), .B2(n6027), .ZN(n5367) );
  OAI211_X1 U6494 ( .C1(n6051), .C2(n5368), .A(n6030), .B(n5367), .ZN(n5374)
         );
  NOR2_X1 U6495 ( .A1(n5370), .A2(n5369), .ZN(n5967) );
  INV_X1 U6496 ( .A(n5967), .ZN(n5371) );
  AOI21_X1 U6497 ( .B1(n6667), .B2(n5372), .A(n5371), .ZN(n5373) );
  AOI211_X1 U6498 ( .C1(n5905), .C2(n6045), .A(n5374), .B(n5373), .ZN(n5375)
         );
  OAI21_X1 U6499 ( .B1(n5518), .B2(n5977), .A(n5375), .ZN(U2810) );
  OAI21_X1 U6500 ( .B1(n5376), .B2(n5377), .A(n5360), .ZN(n5633) );
  AND2_X1 U6501 ( .A1(n5379), .A2(n5378), .ZN(n5411) );
  INV_X1 U6502 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U6503 ( .A(REIP_REG_16__SCAN_IN), .B(n6554), .ZN(n5380) );
  AOI22_X1 U6504 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5411), .B1(n5397), .B2(
        n5380), .ZN(n5388) );
  OR2_X1 U6505 ( .A1(n5392), .A2(n5381), .ZN(n5382) );
  NAND2_X1 U6506 ( .A1(n5383), .A2(n5382), .ZN(n5915) );
  AOI21_X1 U6507 ( .B1(n6056), .B2(EBX_REG_16__SCAN_IN), .A(n6038), .ZN(n5385)
         );
  AOI22_X1 U6508 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6024), .B1(n6027), 
        .B2(n5636), .ZN(n5384) );
  OAI211_X1 U6509 ( .C1(n5915), .C2(n6014), .A(n5385), .B(n5384), .ZN(n5386)
         );
  INV_X1 U6510 ( .A(n5386), .ZN(n5387) );
  OAI211_X1 U6511 ( .C1(n5633), .C2(n5977), .A(n5388), .B(n5387), .ZN(U2811)
         );
  AND2_X1 U6512 ( .A1(n5389), .A2(n5390), .ZN(n5391) );
  OR2_X1 U6513 ( .A1(n5391), .A2(n5376), .ZN(n5641) );
  AOI21_X1 U6514 ( .B1(n5393), .B2(n5406), .A(n5392), .ZN(n5924) );
  AOI22_X1 U6515 ( .A1(n5924), .A2(n6045), .B1(n6056), .B2(EBX_REG_15__SCAN_IN), .ZN(n5394) );
  OAI211_X1 U6516 ( .C1(n6051), .C2(n5395), .A(n5394), .B(n6030), .ZN(n5396)
         );
  AOI21_X1 U6517 ( .B1(n5397), .B2(n6554), .A(n5396), .ZN(n5400) );
  INV_X1 U6518 ( .A(n5643), .ZN(n5398) );
  AOI22_X1 U6519 ( .A1(n5411), .A2(REIP_REG_15__SCAN_IN), .B1(n6027), .B2(
        n5398), .ZN(n5399) );
  OAI211_X1 U6520 ( .C1(n5641), .C2(n5977), .A(n5400), .B(n5399), .ZN(U2812)
         );
  OAI21_X1 U6521 ( .B1(n5401), .B2(n5402), .A(n5389), .ZN(n5653) );
  NAND2_X1 U6522 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5403) );
  INV_X1 U6523 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6552) );
  OAI21_X1 U6524 ( .B1(n5403), .B2(n5429), .A(n6552), .ZN(n5412) );
  INV_X1 U6525 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5651) );
  OAI21_X1 U6526 ( .B1(n5846), .B2(n5498), .A(n6030), .ZN(n5408) );
  NAND2_X1 U6527 ( .A1(n5418), .A2(n5404), .ZN(n5405) );
  NAND2_X1 U6528 ( .A1(n5406), .A2(n5405), .ZN(n5787) );
  NOR2_X1 U6529 ( .A1(n5787), .A2(n6014), .ZN(n5407) );
  AOI211_X1 U6530 ( .C1(n5656), .C2(n6027), .A(n5408), .B(n5407), .ZN(n5409)
         );
  OAI21_X1 U6531 ( .B1(n5651), .B2(n6051), .A(n5409), .ZN(n5410) );
  AOI21_X1 U6532 ( .B1(n5412), .B2(n5411), .A(n5410), .ZN(n5413) );
  OAI21_X1 U6533 ( .B1(n5653), .B2(n5977), .A(n5413), .ZN(U2813) );
  AOI21_X1 U6534 ( .B1(n5417), .B2(n5414), .A(n5416), .ZN(n5895) );
  INV_X1 U6535 ( .A(n5895), .ZN(n5523) );
  INV_X1 U6536 ( .A(n5898), .ZN(n5422) );
  INV_X1 U6537 ( .A(n5418), .ZN(n5419) );
  AOI21_X1 U6538 ( .B1(n5421), .B2(n5420), .A(n5419), .ZN(n5932) );
  AOI22_X1 U6539 ( .A1(n5422), .A2(n6027), .B1(n6045), .B2(n5932), .ZN(n5423)
         );
  OAI211_X1 U6540 ( .C1(n6051), .C2(n5424), .A(n5423), .B(n6030), .ZN(n5425)
         );
  INV_X1 U6541 ( .A(n5425), .ZN(n5428) );
  OAI21_X1 U6542 ( .B1(n5979), .B2(n5426), .A(REIP_REG_13__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6543 ( .A1(n5428), .A2(n5427), .ZN(n5431) );
  INV_X1 U6544 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6549) );
  NOR3_X1 U6545 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6549), .A3(n5429), .ZN(n5430) );
  AOI211_X1 U6546 ( .C1(EBX_REG_13__SCAN_IN), .C2(n6056), .A(n5431), .B(n5430), 
        .ZN(n5432) );
  OAI21_X1 U6547 ( .B1(n5523), .B2(n5977), .A(n5432), .ZN(U2814) );
  INV_X1 U6548 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5433) );
  OAI22_X1 U6549 ( .A1(n5678), .A2(n5499), .B1(n5497), .B2(n5433), .ZN(U2828)
         );
  INV_X1 U6550 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5434) );
  OAI222_X1 U6551 ( .A1(n5460), .A2(n5505), .B1(n5434), .B2(n5497), .C1(n5693), 
        .C2(n5499), .ZN(U2830) );
  INV_X1 U6552 ( .A(n5702), .ZN(n5435) );
  AOI22_X1 U6553 ( .A1(n5435), .A2(n6622), .B1(EBX_REG_28__SCAN_IN), .B2(n6625), .ZN(n5436) );
  OAI21_X1 U6554 ( .B1(n5508), .B2(n5460), .A(n5436), .ZN(U2831) );
  AND2_X1 U6555 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  NAND2_X1 U6556 ( .A1(n5445), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U6557 ( .A1(n5442), .A2(n5441), .ZN(n5825) );
  OAI222_X1 U6558 ( .A1(n5460), .A2(n5826), .B1(n5497), .B2(n4248), .C1(n5825), 
        .C2(n5499), .ZN(U2833) );
  XOR2_X1 U6559 ( .A(n5444), .B(n5443), .Z(n5875) );
  INV_X1 U6560 ( .A(n5875), .ZN(n5448) );
  AOI21_X1 U6561 ( .B1(n5446), .B2(n5323), .A(n3067), .ZN(n5834) );
  AOI22_X1 U6562 ( .A1(n5834), .A2(n6622), .B1(EBX_REG_25__SCAN_IN), .B2(n6625), .ZN(n5447) );
  OAI21_X1 U6563 ( .B1(n5448), .B2(n5460), .A(n5447), .ZN(U2834) );
  INV_X1 U6564 ( .A(n5449), .ZN(n5742) );
  AOI22_X1 U6565 ( .A1(n5742), .A2(n6622), .B1(EBX_REG_24__SCAN_IN), .B2(n6625), .ZN(n5450) );
  OAI21_X1 U6566 ( .B1(n5576), .B2(n5460), .A(n5450), .ZN(U2835) );
  NOR2_X1 U6567 ( .A1(n5497), .A2(n5451), .ZN(n5452) );
  AOI21_X1 U6568 ( .B1(n5750), .B2(n6622), .A(n5452), .ZN(n5453) );
  OAI21_X1 U6569 ( .B1(n5513), .B2(n5460), .A(n5453), .ZN(U2836) );
  NOR2_X1 U6570 ( .A1(n5497), .A2(n5454), .ZN(n5455) );
  AOI21_X1 U6571 ( .B1(n5755), .B2(n6622), .A(n5455), .ZN(n5456) );
  OAI21_X1 U6572 ( .B1(n5457), .B2(n5460), .A(n5456), .ZN(U2837) );
  XOR2_X1 U6573 ( .A(n5459), .B(n5458), .Z(n5881) );
  INV_X1 U6574 ( .A(n5460), .ZN(n6624) );
  OR2_X1 U6575 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  NAND2_X1 U6576 ( .A1(n5348), .A2(n5463), .ZN(n5841) );
  OAI22_X1 U6577 ( .A1(n5841), .A2(n5499), .B1(n5845), .B2(n5497), .ZN(n5464)
         );
  AOI21_X1 U6578 ( .B1(n5881), .B2(n6624), .A(n5464), .ZN(n5465) );
  INV_X1 U6579 ( .A(n5465), .ZN(U2838) );
  INV_X1 U6580 ( .A(n5466), .ZN(n5468) );
  INV_X1 U6581 ( .A(n5458), .ZN(n5467) );
  AOI21_X1 U6582 ( .B1(n5469), .B2(n5468), .A(n5467), .ZN(n5884) );
  INV_X1 U6583 ( .A(n5884), .ZN(n5473) );
  MUX2_X1 U6584 ( .A(n4157), .B(n5479), .S(n3118), .Z(n5471) );
  XNOR2_X1 U6585 ( .A(n5471), .B(n5470), .ZN(n5852) );
  AOI22_X1 U6586 ( .A1(n5852), .A2(n6622), .B1(EBX_REG_20__SCAN_IN), .B2(n6625), .ZN(n5472) );
  OAI21_X1 U6587 ( .B1(n5473), .B2(n5460), .A(n5472), .ZN(U2839) );
  AND2_X1 U6588 ( .A1(n5474), .A2(n5475), .ZN(n5476) );
  NOR2_X1 U6589 ( .A1(n5466), .A2(n5476), .ZN(n5614) );
  MUX2_X1 U6590 ( .A(n5479), .B(n5478), .S(n5477), .Z(n5486) );
  INV_X1 U6591 ( .A(n5486), .ZN(n5480) );
  NAND2_X1 U6592 ( .A1(n5364), .A2(n5480), .ZN(n5488) );
  XNOR2_X1 U6593 ( .A(n5488), .B(n5481), .ZN(n5864) );
  OAI22_X1 U6594 ( .A1(n5864), .A2(n5499), .B1(n6687), .B2(n5497), .ZN(n5482)
         );
  AOI21_X1 U6595 ( .B1(n5614), .B2(n6624), .A(n5482), .ZN(n5483) );
  INV_X1 U6596 ( .A(n5483), .ZN(U2840) );
  NAND2_X1 U6597 ( .A1(n5361), .A2(n5484), .ZN(n5485) );
  AND2_X1 U6598 ( .A1(n5474), .A2(n5485), .ZN(n6062) );
  INV_X1 U6599 ( .A(n6062), .ZN(n5491) );
  NAND2_X1 U6600 ( .A1(n5365), .A2(n5486), .ZN(n5487) );
  INV_X1 U6601 ( .A(n5971), .ZN(n5489) );
  OAI222_X1 U6602 ( .A1(n5460), .A2(n5491), .B1(n5490), .B2(n5497), .C1(n5489), 
        .C2(n5499), .ZN(U2841) );
  AOI22_X1 U6603 ( .A1(n5905), .A2(n6622), .B1(EBX_REG_17__SCAN_IN), .B2(n6625), .ZN(n5492) );
  OAI21_X1 U6604 ( .B1(n5518), .B2(n5460), .A(n5492), .ZN(U2842) );
  INV_X1 U6605 ( .A(n5633), .ZN(n6066) );
  OAI22_X1 U6606 ( .A1(n5915), .A2(n5499), .B1(n5493), .B2(n5497), .ZN(n5494)
         );
  AOI21_X1 U6607 ( .B1(n6066), .B2(n6624), .A(n5494), .ZN(n5495) );
  INV_X1 U6608 ( .A(n5495), .ZN(U2843) );
  AOI22_X1 U6609 ( .A1(n5924), .A2(n6622), .B1(EBX_REG_15__SCAN_IN), .B2(n6625), .ZN(n5496) );
  OAI21_X1 U6610 ( .B1(n5641), .B2(n5460), .A(n5496), .ZN(U2844) );
  OAI22_X1 U6611 ( .A1(n5787), .A2(n5499), .B1(n5498), .B2(n5497), .ZN(n5500)
         );
  INV_X1 U6612 ( .A(n5500), .ZN(n5501) );
  OAI21_X1 U6613 ( .B1(n5653), .B2(n5460), .A(n5501), .ZN(U2845) );
  AOI22_X1 U6614 ( .A1(n5932), .A2(n6622), .B1(EBX_REG_13__SCAN_IN), .B2(n6625), .ZN(n5502) );
  OAI21_X1 U6615 ( .B1(n5523), .B2(n5460), .A(n5502), .ZN(U2846) );
  AOI22_X1 U6616 ( .A1(n6065), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6067), .ZN(n5504) );
  NAND2_X1 U6617 ( .A1(n6068), .A2(DATAI_13_), .ZN(n5503) );
  OAI211_X1 U6618 ( .C1(n5505), .C2(n5871), .A(n5504), .B(n5503), .ZN(U2862)
         );
  AOI22_X1 U6619 ( .A1(n6065), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6067), .ZN(n5507) );
  NAND2_X1 U6620 ( .A1(n6068), .A2(DATAI_12_), .ZN(n5506) );
  OAI211_X1 U6621 ( .C1(n5508), .C2(n5871), .A(n5507), .B(n5506), .ZN(U2863)
         );
  AOI22_X1 U6622 ( .A1(n6065), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6067), .ZN(n5510) );
  NAND2_X1 U6623 ( .A1(n6068), .A2(DATAI_8_), .ZN(n5509) );
  OAI211_X1 U6624 ( .C1(n5576), .C2(n5871), .A(n5510), .B(n5509), .ZN(U2867)
         );
  AOI22_X1 U6625 ( .A1(n6065), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6067), .ZN(n5512) );
  NAND2_X1 U6626 ( .A1(n6068), .A2(DATAI_7_), .ZN(n5511) );
  OAI211_X1 U6627 ( .C1(n5513), .C2(n5871), .A(n5512), .B(n5511), .ZN(U2868)
         );
  INV_X1 U6628 ( .A(n5614), .ZN(n5865) );
  AOI22_X1 U6629 ( .A1(n6068), .A2(DATAI_3_), .B1(n6067), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U6630 ( .A1(n6065), .A2(DATAI_19_), .ZN(n5514) );
  OAI211_X1 U6631 ( .C1(n5865), .C2(n5871), .A(n5515), .B(n5514), .ZN(U2872)
         );
  AOI22_X1 U6632 ( .A1(n6065), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6067), .ZN(n5517) );
  NAND2_X1 U6633 ( .A1(n6068), .A2(DATAI_1_), .ZN(n5516) );
  OAI211_X1 U6634 ( .C1(n5518), .C2(n5871), .A(n5517), .B(n5516), .ZN(U2874)
         );
  AOI22_X1 U6635 ( .A1(n6071), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6067), .ZN(n5519) );
  OAI21_X1 U6636 ( .B1(n5641), .B2(n5871), .A(n5519), .ZN(U2876) );
  INV_X1 U6637 ( .A(DATAI_14_), .ZN(n6123) );
  OAI222_X1 U6638 ( .A1(n5653), .A2(n5871), .B1(n6074), .B2(n5520), .C1(n6123), 
        .C2(n5521), .ZN(U2877) );
  INV_X1 U6639 ( .A(DATAI_13_), .ZN(n6121) );
  OAI222_X1 U6640 ( .A1(n5523), .A2(n5871), .B1(n6074), .B2(n5522), .C1(n6121), 
        .C2(n5521), .ZN(U2878) );
  XNOR2_X1 U6641 ( .A(n5524), .B(n5686), .ZN(n5692) );
  AND2_X1 U6642 ( .A1(n6206), .A2(REIP_REG_30__SCAN_IN), .ZN(n5684) );
  AOI21_X1 U6643 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5684), 
        .ZN(n5525) );
  OAI21_X1 U6644 ( .B1(n6204), .B2(n5526), .A(n5525), .ZN(n5527) );
  AOI21_X1 U6645 ( .B1(n5528), .B2(n5894), .A(n5527), .ZN(n5529) );
  OAI21_X1 U6646 ( .B1(n5692), .B2(n6178), .A(n5529), .ZN(U2956) );
  INV_X1 U6647 ( .A(n5530), .ZN(n5531) );
  OAI21_X1 U6648 ( .B1(n5531), .B2(n3006), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n5533) );
  AOI22_X1 U6649 ( .A1(n5533), .A2(n5532), .B1(n3006), .B2(n5683), .ZN(n5701)
         );
  INV_X1 U6650 ( .A(n5534), .ZN(n5536) );
  AND2_X1 U6651 ( .A1(n6206), .A2(REIP_REG_29__SCAN_IN), .ZN(n5694) );
  AOI21_X1 U6652 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5694), 
        .ZN(n5535) );
  OAI21_X1 U6653 ( .B1(n6204), .B2(n5536), .A(n5535), .ZN(n5537) );
  AOI21_X1 U6654 ( .B1(n5538), .B2(n5894), .A(n5537), .ZN(n5539) );
  OAI21_X1 U6655 ( .B1(n5701), .B2(n6178), .A(n5539), .ZN(U2957) );
  NAND3_X1 U6656 ( .A1(n2986), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n6169), .ZN(n5542) );
  NAND2_X1 U6657 ( .A1(n5732), .A2(n5541), .ZN(n5723) );
  AOI22_X1 U6658 ( .A1(n5542), .A2(n5549), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5541), .ZN(n5543) );
  XNOR2_X1 U6659 ( .A(n5543), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5711)
         );
  AND2_X1 U6660 ( .A1(n6206), .A2(REIP_REG_28__SCAN_IN), .ZN(n5704) );
  AOI21_X1 U6661 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5704), 
        .ZN(n5544) );
  OAI21_X1 U6662 ( .B1(n6204), .B2(n5545), .A(n5544), .ZN(n5546) );
  AOI21_X1 U6663 ( .B1(n5547), .B2(n5894), .A(n5546), .ZN(n5548) );
  OAI21_X1 U6664 ( .B1(n6178), .B2(n5711), .A(n5548), .ZN(U2958) );
  NAND2_X1 U6665 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  XNOR2_X1 U6666 ( .A(n5551), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5719)
         );
  NAND2_X1 U6667 ( .A1(n6206), .A2(REIP_REG_27__SCAN_IN), .ZN(n5712) );
  OAI21_X1 U6668 ( .B1(n5652), .B2(n5552), .A(n5712), .ZN(n5554) );
  NOR2_X1 U6669 ( .A1(n5818), .A2(n6173), .ZN(n5553) );
  AOI211_X1 U6670 ( .C1(n5657), .C2(n5815), .A(n5554), .B(n5553), .ZN(n5555)
         );
  OAI21_X1 U6671 ( .B1(n5719), .B2(n6178), .A(n5555), .ZN(U2959) );
  NOR2_X1 U6672 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  XNOR2_X1 U6673 ( .A(n5559), .B(n5558), .ZN(n5727) );
  INV_X1 U6674 ( .A(n5826), .ZN(n5872) );
  AND2_X1 U6675 ( .A1(n6206), .A2(REIP_REG_26__SCAN_IN), .ZN(n5721) );
  AOI21_X1 U6676 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5721), 
        .ZN(n5560) );
  OAI21_X1 U6677 ( .B1(n6204), .B2(n5823), .A(n5560), .ZN(n5561) );
  AOI21_X1 U6678 ( .B1(n5872), .B2(n5894), .A(n5561), .ZN(n5562) );
  OAI21_X1 U6679 ( .B1(n5727), .B2(n6178), .A(n5562), .ZN(U2960) );
  AOI21_X1 U6680 ( .B1(n5540), .B2(n5564), .A(n5563), .ZN(n5735) );
  NAND2_X1 U6681 ( .A1(n5657), .A2(n5833), .ZN(n5565) );
  NAND2_X1 U6682 ( .A1(n6258), .A2(REIP_REG_25__SCAN_IN), .ZN(n5729) );
  OAI211_X1 U6683 ( .C1(n5652), .C2(n6704), .A(n5565), .B(n5729), .ZN(n5566)
         );
  AOI21_X1 U6684 ( .B1(n5875), .B2(n5894), .A(n5566), .ZN(n5567) );
  OAI21_X1 U6685 ( .B1(n5735), .B2(n6178), .A(n5567), .ZN(U2961) );
  NAND2_X1 U6686 ( .A1(n5568), .A2(n3004), .ZN(n5571) );
  XNOR2_X1 U6687 ( .A(n6169), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5604)
         );
  OR2_X1 U6688 ( .A1(n6169), .A2(n5774), .ZN(n5572) );
  XNOR2_X1 U6689 ( .A(n6169), .B(n5756), .ZN(n5598) );
  NOR2_X1 U6690 ( .A1(n6169), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5589)
         );
  NAND2_X1 U6691 ( .A1(n5596), .A2(n5589), .ZN(n5582) );
  NAND2_X1 U6692 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  XNOR2_X1 U6693 ( .A(n5575), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5744)
         );
  INV_X1 U6694 ( .A(n5576), .ZN(n5580) );
  AND2_X1 U6695 ( .A1(n6206), .A2(REIP_REG_24__SCAN_IN), .ZN(n5741) );
  AOI21_X1 U6696 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5741), 
        .ZN(n5577) );
  OAI21_X1 U6697 ( .B1(n6204), .B2(n5578), .A(n5577), .ZN(n5579) );
  AOI21_X1 U6698 ( .B1(n5580), .B2(n5894), .A(n5579), .ZN(n5581) );
  OAI21_X1 U6699 ( .B1(n5744), .B2(n6178), .A(n5581), .ZN(U2962) );
  OAI21_X1 U6700 ( .B1(n5603), .B2(n5736), .A(n5582), .ZN(n5583) );
  XNOR2_X1 U6701 ( .A(n5583), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5752)
         );
  NAND2_X1 U6702 ( .A1(n6206), .A2(REIP_REG_23__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U6703 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5584)
         );
  OAI211_X1 U6704 ( .C1(n6204), .C2(n5585), .A(n5745), .B(n5584), .ZN(n5586)
         );
  AOI21_X1 U6705 ( .B1(n5587), .B2(n5894), .A(n5586), .ZN(n5588) );
  OAI21_X1 U6706 ( .B1(n5752), .B2(n6178), .A(n5588), .ZN(U2963) );
  AOI21_X1 U6707 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6169), .A(n5589), 
        .ZN(n5591) );
  XOR2_X1 U6708 ( .A(n5591), .B(n5590), .Z(n5760) );
  AND2_X1 U6709 ( .A1(n6206), .A2(REIP_REG_22__SCAN_IN), .ZN(n5754) );
  AOI21_X1 U6710 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5754), 
        .ZN(n5592) );
  OAI21_X1 U6711 ( .B1(n6204), .B2(n5593), .A(n5592), .ZN(n5594) );
  AOI21_X1 U6712 ( .B1(n5878), .B2(n5894), .A(n5594), .ZN(n5595) );
  OAI21_X1 U6713 ( .B1(n5760), .B2(n6178), .A(n5595), .ZN(U2964) );
  AOI21_X1 U6714 ( .B1(n5598), .B2(n5597), .A(n5596), .ZN(n5768) );
  INV_X1 U6715 ( .A(n5843), .ZN(n5600) );
  NAND2_X1 U6716 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5599)
         );
  NAND2_X1 U6717 ( .A1(n6258), .A2(REIP_REG_21__SCAN_IN), .ZN(n5761) );
  OAI211_X1 U6718 ( .C1(n6204), .C2(n5600), .A(n5599), .B(n5761), .ZN(n5601)
         );
  AOI21_X1 U6719 ( .B1(n5881), .B2(n5894), .A(n5601), .ZN(n5602) );
  OAI21_X1 U6720 ( .B1(n5768), .B2(n6178), .A(n5602), .ZN(U2965) );
  OAI21_X1 U6721 ( .B1(n5605), .B2(n5604), .A(n5603), .ZN(n5778) );
  AOI22_X1 U6722 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n6206), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U6723 ( .B1(n6204), .B2(n5855), .A(n5606), .ZN(n5607) );
  AOI21_X1 U6724 ( .B1(n5884), .B2(n5894), .A(n5607), .ZN(n5608) );
  OAI21_X1 U6725 ( .B1(n5778), .B2(n6178), .A(n5608), .ZN(U2966) );
  XNOR2_X1 U6726 ( .A(n3004), .B(n4064), .ZN(n5609) );
  XNOR2_X1 U6727 ( .A(n5610), .B(n5609), .ZN(n5785) );
  INV_X1 U6728 ( .A(n5861), .ZN(n5612) );
  AOI22_X1 U6729 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6206), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5611) );
  OAI21_X1 U6730 ( .B1(n6204), .B2(n5612), .A(n5611), .ZN(n5613) );
  AOI21_X1 U6731 ( .B1(n5614), .B2(n5894), .A(n5613), .ZN(n5615) );
  OAI21_X1 U6732 ( .B1(n5785), .B2(n6178), .A(n5615), .ZN(U2967) );
  NAND2_X1 U6733 ( .A1(n3004), .A2(n5921), .ZN(n5628) );
  AOI21_X1 U6734 ( .B1(n3004), .B2(n5910), .A(n3005), .ZN(n5616) );
  AOI21_X1 U6735 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5628), .A(n5616), 
        .ZN(n5619) );
  NOR3_X1 U6736 ( .A1(n3005), .A2(n3004), .A3(n5910), .ZN(n5888) );
  NOR3_X1 U6737 ( .A1(n2990), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5628), 
        .ZN(n5887) );
  INV_X1 U6738 ( .A(n5887), .ZN(n5618) );
  OAI21_X1 U6739 ( .B1(n5619), .B2(n5888), .A(n5618), .ZN(n5906) );
  INV_X1 U6740 ( .A(n5906), .ZN(n5626) );
  INV_X1 U6741 ( .A(n5620), .ZN(n5622) );
  AOI22_X1 U6742 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n6206), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5621) );
  OAI21_X1 U6743 ( .B1(n6204), .B2(n5622), .A(n5621), .ZN(n5623) );
  AOI21_X1 U6744 ( .B1(n5624), .B2(n5894), .A(n5623), .ZN(n5625) );
  OAI21_X1 U6745 ( .B1(n5626), .B2(n6178), .A(n5625), .ZN(U2969) );
  OAI21_X1 U6746 ( .B1(n3004), .B2(n5921), .A(n5628), .ZN(n5629) );
  XNOR2_X1 U6747 ( .A(n5630), .B(n5629), .ZN(n5916) );
  INV_X1 U6748 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5631) );
  OAI22_X1 U6749 ( .A1(n5652), .A2(n5632), .B1(n5907), .B2(n5631), .ZN(n5635)
         );
  NOR2_X1 U6750 ( .A1(n5633), .A2(n6173), .ZN(n5634) );
  AOI211_X1 U6751 ( .C1(n5657), .C2(n5636), .A(n5635), .B(n5634), .ZN(n5637)
         );
  OAI21_X1 U6752 ( .B1(n5916), .B2(n6178), .A(n5637), .ZN(U2970) );
  XNOR2_X1 U6753 ( .A(n6169), .B(n5928), .ZN(n5639) );
  XNOR2_X1 U6754 ( .A(n5640), .B(n5639), .ZN(n5925) );
  INV_X1 U6755 ( .A(n5925), .ZN(n5647) );
  INV_X1 U6756 ( .A(n5641), .ZN(n5645) );
  AOI22_X1 U6757 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6206), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5642) );
  OAI21_X1 U6758 ( .B1(n6204), .B2(n5643), .A(n5642), .ZN(n5644) );
  AOI21_X1 U6759 ( .B1(n5645), .B2(n5894), .A(n5644), .ZN(n5646) );
  OAI21_X1 U6760 ( .B1(n5647), .B2(n6178), .A(n5646), .ZN(U2971) );
  NAND2_X1 U6761 ( .A1(n3021), .A2(n5649), .ZN(n5650) );
  XNOR2_X1 U6762 ( .A(n5648), .B(n5650), .ZN(n5802) );
  NAND2_X1 U6763 ( .A1(n6258), .A2(REIP_REG_14__SCAN_IN), .ZN(n5786) );
  OAI21_X1 U6764 ( .B1(n5652), .B2(n5651), .A(n5786), .ZN(n5655) );
  NOR2_X1 U6765 ( .A1(n5653), .A2(n6173), .ZN(n5654) );
  AOI211_X1 U6766 ( .C1(n5657), .C2(n5656), .A(n5655), .B(n5654), .ZN(n5658)
         );
  OAI21_X1 U6767 ( .B1(n6178), .B2(n5802), .A(n5658), .ZN(U2972) );
  INV_X1 U6768 ( .A(n5707), .ZN(n5674) );
  NAND2_X1 U6769 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5724) );
  INV_X1 U6770 ( .A(n5659), .ZN(n5668) );
  NAND2_X1 U6771 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5791), .ZN(n5919) );
  NOR2_X1 U6772 ( .A1(n5920), .A2(n5919), .ZN(n5914) );
  NAND3_X1 U6773 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5914), .ZN(n5671) );
  INV_X1 U6774 ( .A(n5671), .ZN(n5661) );
  NAND2_X1 U6775 ( .A1(n5661), .A2(n5660), .ZN(n5662) );
  NAND2_X1 U6776 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  AND2_X1 U6777 ( .A1(n6219), .A2(n5664), .ZN(n5769) );
  NOR2_X1 U6778 ( .A1(n5665), .A2(n5671), .ZN(n5770) );
  INV_X1 U6779 ( .A(n5771), .ZN(n5672) );
  NAND3_X1 U6780 ( .A1(n5770), .A2(n5672), .A3(n5773), .ZN(n5666) );
  NAND2_X1 U6781 ( .A1(n6222), .A2(n5666), .ZN(n5667) );
  NAND2_X1 U6782 ( .A1(n5769), .A2(n5667), .ZN(n5763) );
  AOI21_X1 U6783 ( .B1(n5668), .B2(n6222), .A(n5763), .ZN(n5746) );
  OAI21_X1 U6784 ( .B1(n6281), .B2(n6216), .A(n5669), .ZN(n5670) );
  NAND2_X1 U6785 ( .A1(n5746), .A2(n5670), .ZN(n5728) );
  AOI21_X1 U6786 ( .B1(n5724), .B2(n6222), .A(n5728), .ZN(n5714) );
  OAI21_X1 U6787 ( .B1(n5674), .B2(n6220), .A(n5714), .ZN(n5695) );
  AOI21_X1 U6788 ( .B1(n5683), .B2(n6222), .A(n5695), .ZN(n5687) );
  OAI21_X1 U6789 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n6220), .A(n5687), 
        .ZN(n5677) );
  NOR2_X1 U6790 ( .A1(n6205), .A2(n5671), .ZN(n5911) );
  NAND2_X1 U6791 ( .A1(n5783), .A2(n5673), .ZN(n5722) );
  NOR2_X1 U6792 ( .A1(n5722), .A2(n5724), .ZN(n5717) );
  NAND2_X1 U6793 ( .A1(n5717), .A2(n5674), .ZN(n5697) );
  NOR4_X1 U6794 ( .A1(n5697), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5686), 
        .A4(n5683), .ZN(n5675) );
  AOI211_X1 U6795 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n5677), .A(n5676), .B(n5675), .ZN(n5681) );
  INV_X1 U6796 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U6797 ( .A1(n5679), .A2(n6286), .ZN(n5680) );
  OAI211_X1 U6798 ( .C1(n5682), .C2(n6208), .A(n5681), .B(n5680), .ZN(U2987)
         );
  NOR3_X1 U6799 ( .A1(n5697), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5683), 
        .ZN(n5689) );
  INV_X1 U6800 ( .A(n5684), .ZN(n5685) );
  OAI21_X1 U6801 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5688) );
  AOI211_X1 U6802 ( .C1(n5690), .C2(n6286), .A(n5689), .B(n5688), .ZN(n5691)
         );
  OAI21_X1 U6803 ( .B1(n5692), .B2(n6208), .A(n5691), .ZN(U2988) );
  INV_X1 U6804 ( .A(n5693), .ZN(n5699) );
  AOI21_X1 U6805 ( .B1(n5695), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5694), 
        .ZN(n5696) );
  OAI21_X1 U6806 ( .B1(n5697), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5696), 
        .ZN(n5698) );
  AOI21_X1 U6807 ( .B1(n5699), .B2(n6286), .A(n5698), .ZN(n5700) );
  OAI21_X1 U6808 ( .B1(n5701), .B2(n6208), .A(n5700), .ZN(U2989) );
  INV_X1 U6809 ( .A(n5714), .ZN(n5705) );
  NOR2_X1 U6810 ( .A1(n5702), .A2(n6274), .ZN(n5703) );
  AOI211_X1 U6811 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5705), .A(n5704), .B(n5703), .ZN(n5710) );
  INV_X1 U6812 ( .A(n5706), .ZN(n5708) );
  NAND3_X1 U6813 ( .A1(n5717), .A2(n5708), .A3(n5707), .ZN(n5709) );
  OAI211_X1 U6814 ( .C1(n5711), .C2(n6208), .A(n5710), .B(n5709), .ZN(U2990)
         );
  INV_X1 U6815 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U6816 ( .A1(n5816), .A2(n6286), .ZN(n5713) );
  OAI211_X1 U6817 ( .C1(n5714), .C2(n5716), .A(n5713), .B(n5712), .ZN(n5715)
         );
  AOI21_X1 U6818 ( .B1(n5717), .B2(n5716), .A(n5715), .ZN(n5718) );
  OAI21_X1 U6819 ( .B1(n5719), .B2(n6208), .A(n5718), .ZN(U2991) );
  NOR2_X1 U6820 ( .A1(n5825), .A2(n6274), .ZN(n5720) );
  AOI211_X1 U6821 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5728), .A(n5721), .B(n5720), .ZN(n5726) );
  INV_X1 U6822 ( .A(n5722), .ZN(n5733) );
  NAND3_X1 U6823 ( .A1(n5733), .A2(n5724), .A3(n5723), .ZN(n5725) );
  OAI211_X1 U6824 ( .C1(n5727), .C2(n6208), .A(n5726), .B(n5725), .ZN(U2992)
         );
  INV_X1 U6825 ( .A(n5728), .ZN(n5739) );
  NAND2_X1 U6826 ( .A1(n5834), .A2(n6286), .ZN(n5730) );
  OAI211_X1 U6827 ( .C1(n5739), .C2(n5732), .A(n5730), .B(n5729), .ZN(n5731)
         );
  AOI21_X1 U6828 ( .B1(n5733), .B2(n5732), .A(n5731), .ZN(n5734) );
  OAI21_X1 U6829 ( .B1(n5735), .B2(n6208), .A(n5734), .ZN(U2993) );
  INV_X1 U6830 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U6831 ( .A1(n5783), .A2(n5737), .ZN(n5747) );
  AOI211_X1 U6832 ( .C1(n5747), .C2(n6648), .A(n5739), .B(n5738), .ZN(n5740)
         );
  AOI211_X1 U6833 ( .C1(n6286), .C2(n5742), .A(n5741), .B(n5740), .ZN(n5743)
         );
  OAI21_X1 U6834 ( .B1(n5744), .B2(n6208), .A(n5743), .ZN(U2994) );
  INV_X1 U6835 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6707) );
  OAI21_X1 U6836 ( .B1(n5746), .B2(n6707), .A(n5745), .ZN(n5749) );
  NOR2_X1 U6837 ( .A1(n5747), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5748)
         );
  AOI211_X1 U6838 ( .C1(n6286), .C2(n5750), .A(n5749), .B(n5748), .ZN(n5751)
         );
  OAI21_X1 U6839 ( .B1(n5752), .B2(n6208), .A(n5751), .ZN(U2995) );
  AND4_X1 U6840 ( .A1(n5783), .A2(n5773), .A3(INSTADDRPOINTER_REG_21__SCAN_IN), 
        .A4(n6716), .ZN(n5753) );
  AOI211_X1 U6841 ( .C1(n6286), .C2(n5755), .A(n5754), .B(n5753), .ZN(n5759)
         );
  AND2_X1 U6842 ( .A1(n5773), .A2(n5756), .ZN(n5757) );
  AND2_X1 U6843 ( .A1(n5783), .A2(n5757), .ZN(n5766) );
  OAI21_X1 U6844 ( .B1(n5766), .B2(n5763), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5758) );
  OAI211_X1 U6845 ( .C1(n5760), .C2(n6208), .A(n5759), .B(n5758), .ZN(U2996)
         );
  INV_X1 U6846 ( .A(n5761), .ZN(n5762) );
  AOI21_X1 U6847 ( .B1(n5763), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5762), 
        .ZN(n5764) );
  OAI21_X1 U6848 ( .B1(n5841), .B2(n6274), .A(n5764), .ZN(n5765) );
  NOR2_X1 U6849 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  OAI21_X1 U6850 ( .B1(n5768), .B2(n6208), .A(n5767), .ZN(U2997) );
  OAI221_X1 U6851 ( .B1(n6288), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n6288), .C2(n5770), .A(n5769), .ZN(n5909) );
  AOI21_X1 U6852 ( .B1(n5771), .B2(n6222), .A(n5909), .ZN(n5780) );
  OAI22_X1 U6853 ( .A1(n5780), .A2(n5774), .B1(n6560), .B2(n5907), .ZN(n5776)
         );
  INV_X1 U6854 ( .A(n5783), .ZN(n5772) );
  AOI211_X1 U6855 ( .C1(n4064), .C2(n5774), .A(n5773), .B(n5772), .ZN(n5775)
         );
  AOI211_X1 U6856 ( .C1(n6286), .C2(n5852), .A(n5776), .B(n5775), .ZN(n5777)
         );
  OAI21_X1 U6857 ( .B1(n5778), .B2(n6208), .A(n5777), .ZN(U2998) );
  NAND2_X1 U6858 ( .A1(n6258), .A2(REIP_REG_19__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U6859 ( .B1(n5864), .B2(n6274), .A(n5779), .ZN(n5782) );
  NOR2_X1 U6860 ( .A1(n5780), .A2(n4064), .ZN(n5781) );
  AOI211_X1 U6861 ( .C1(n5783), .C2(n4064), .A(n5782), .B(n5781), .ZN(n5784)
         );
  OAI21_X1 U6862 ( .B1(n5785), .B2(n6208), .A(n5784), .ZN(U2999) );
  NOR2_X1 U6863 ( .A1(n6205), .A2(n5919), .ZN(n5800) );
  OAI21_X1 U6864 ( .B1(n6274), .B2(n5787), .A(n5786), .ZN(n5799) );
  NAND2_X1 U6865 ( .A1(n5788), .A2(n5919), .ZN(n5789) );
  OAI211_X1 U6866 ( .C1(n5791), .C2(n5790), .A(n6215), .B(n5789), .ZN(n5933)
         );
  INV_X1 U6867 ( .A(n5933), .ZN(n5797) );
  INV_X1 U6868 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6869 ( .A1(n5792), .A2(n5791), .ZN(n5937) );
  INV_X1 U6870 ( .A(n5937), .ZN(n5793) );
  OAI21_X1 U6871 ( .B1(n5795), .B2(n5794), .A(n5793), .ZN(n5796) );
  AOI21_X1 U6872 ( .B1(n5797), .B2(n5796), .A(n5920), .ZN(n5798) );
  AOI211_X1 U6873 ( .C1(n5800), .C2(n5920), .A(n5799), .B(n5798), .ZN(n5801)
         );
  OAI21_X1 U6874 ( .B1(n5802), .B2(n6208), .A(n5801), .ZN(U3004) );
  INV_X1 U6875 ( .A(n5803), .ZN(n5804) );
  OAI222_X1 U6876 ( .A1(n4517), .A2(n6400), .B1(n5811), .B2(n6343), .C1(n6483), 
        .C2(n5804), .ZN(n5805) );
  MUX2_X1 U6877 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n5805), .S(n6296), 
        .Z(U3465) );
  INV_X1 U6878 ( .A(n4385), .ZN(n5807) );
  NAND2_X1 U6879 ( .A1(n4515), .A2(n6299), .ZN(n5810) );
  OAI211_X1 U6880 ( .C1(n4515), .C2(n6299), .A(n5810), .B(n6396), .ZN(n5806)
         );
  OAI21_X1 U6881 ( .B1(n5811), .B2(n5807), .A(n5806), .ZN(n5808) );
  MUX2_X1 U6882 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5808), .S(n6296), 
        .Z(U3463) );
  AND2_X1 U6883 ( .A1(n5809), .A2(n6299), .ZN(n6342) );
  AOI21_X1 U6884 ( .B1(n3998), .B2(n5810), .A(n6342), .ZN(n5813) );
  OAI22_X1 U6885 ( .A1(n5813), .A2(n6400), .B1(n5812), .B2(n5811), .ZN(n5814)
         );
  MUX2_X1 U6886 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5814), .S(n6296), 
        .Z(U3462) );
  AND2_X1 U6887 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6090), .ZN(U2892) );
  AOI22_X1 U6888 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6024), .B1(n5815), 
        .B2(n6027), .ZN(n5821) );
  INV_X1 U6889 ( .A(n5816), .ZN(n5817) );
  INV_X1 U6890 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5824) );
  OAI22_X1 U6891 ( .A1(n5824), .A2(n6051), .B1(n5823), .B2(n6061), .ZN(n5828)
         );
  OAI22_X1 U6892 ( .A1(n5826), .A2(n5977), .B1(n5825), .B2(n6014), .ZN(n5827)
         );
  AOI211_X1 U6893 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6056), .A(n5828), .B(n5827), 
        .ZN(n5829) );
  OAI221_X1 U6894 ( .B1(n5831), .B2(n6569), .C1(n5831), .C2(n5830), .A(n5829), 
        .ZN(U2801) );
  AOI22_X1 U6895 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6056), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6024), .ZN(n5840) );
  AOI22_X1 U6896 ( .A1(n5833), .A2(n6027), .B1(n5832), .B2(
        REIP_REG_25__SCAN_IN), .ZN(n5839) );
  AOI22_X1 U6897 ( .A1(n5875), .A2(n6018), .B1(n6045), .B2(n5834), .ZN(n5838)
         );
  OAI211_X1 U6898 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5836), .B(n5835), .ZN(n5837) );
  NAND4_X1 U6899 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(U2802)
         );
  INV_X1 U6900 ( .A(n5841), .ZN(n5842) );
  AOI22_X1 U6901 ( .A1(n5881), .A2(n6018), .B1(n5842), .B2(n6045), .ZN(n5851)
         );
  INV_X1 U6902 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6562) );
  AOI22_X1 U6903 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6024), .B1(n5843), 
        .B2(n6027), .ZN(n5844) );
  OAI21_X1 U6904 ( .B1(n5846), .B2(n5845), .A(n5844), .ZN(n5847) );
  AOI221_X1 U6905 ( .B1(n5849), .B2(REIP_REG_21__SCAN_IN), .C1(n5848), .C2(
        n6562), .A(n5847), .ZN(n5850) );
  NAND2_X1 U6906 ( .A1(n5851), .A2(n5850), .ZN(U2806) );
  AOI22_X1 U6907 ( .A1(n5884), .A2(n6018), .B1(n6045), .B2(n5852), .ZN(n5860)
         );
  AOI21_X1 U6908 ( .B1(n6560), .B2(n5854), .A(n5853), .ZN(n5858) );
  INV_X1 U6909 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5856) );
  OAI22_X1 U6910 ( .A1(n5856), .A2(n6051), .B1(n5855), .B2(n6061), .ZN(n5857)
         );
  AOI211_X1 U6911 ( .C1(EBX_REG_20__SCAN_IN), .C2(n6056), .A(n5858), .B(n5857), 
        .ZN(n5859) );
  NAND2_X1 U6912 ( .A1(n5860), .A2(n5859), .ZN(U2807) );
  AOI22_X1 U6913 ( .A1(n5861), .A2(n6027), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5967), .ZN(n5862) );
  OAI211_X1 U6914 ( .C1(n6051), .C2(n5863), .A(n5862), .B(n6030), .ZN(n5867)
         );
  OAI22_X1 U6915 ( .A1(n5865), .A2(n5977), .B1(n5864), .B2(n6014), .ZN(n5866)
         );
  AOI211_X1 U6916 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6056), .A(n5867), .B(n5866), 
        .ZN(n5870) );
  OAI211_X1 U6917 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5966), .B(n5868), .ZN(n5869) );
  NAND2_X1 U6918 ( .A1(n5870), .A2(n5869), .ZN(U2808) );
  AOI22_X1 U6919 ( .A1(n5872), .A2(n6072), .B1(n6065), .B2(DATAI_26_), .ZN(
        n5874) );
  AOI22_X1 U6920 ( .A1(n6068), .A2(DATAI_10_), .B1(n6067), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U6921 ( .A1(n5874), .A2(n5873), .ZN(U2865) );
  AOI22_X1 U6922 ( .A1(n5875), .A2(n6072), .B1(n6065), .B2(DATAI_25_), .ZN(
        n5877) );
  AOI22_X1 U6923 ( .A1(n6068), .A2(DATAI_9_), .B1(n6067), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U6924 ( .A1(n5877), .A2(n5876), .ZN(U2866) );
  AOI22_X1 U6925 ( .A1(n5878), .A2(n6072), .B1(n6065), .B2(DATAI_22_), .ZN(
        n5880) );
  AOI22_X1 U6926 ( .A1(n6068), .A2(DATAI_6_), .B1(n6067), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U6927 ( .A1(n5880), .A2(n5879), .ZN(U2869) );
  AOI22_X1 U6928 ( .A1(n5881), .A2(n6072), .B1(n6065), .B2(DATAI_21_), .ZN(
        n5883) );
  AOI22_X1 U6929 ( .A1(n6068), .A2(DATAI_5_), .B1(n6067), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U6930 ( .A1(n5883), .A2(n5882), .ZN(U2870) );
  AOI22_X1 U6931 ( .A1(n5884), .A2(n6072), .B1(n6065), .B2(DATAI_20_), .ZN(
        n5886) );
  AOI22_X1 U6932 ( .A1(n6068), .A2(DATAI_4_), .B1(n6067), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U6933 ( .A1(n5886), .A2(n5885), .ZN(U2871) );
  AOI22_X1 U6934 ( .A1(n6206), .A2(REIP_REG_18__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5891) );
  NOR2_X1 U6935 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  XNOR2_X1 U6936 ( .A(n5889), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5899)
         );
  AOI22_X1 U6937 ( .A1(n5899), .A2(n6199), .B1(n5894), .B2(n6062), .ZN(n5890)
         );
  OAI211_X1 U6938 ( .C1(n6204), .C2(n5969), .A(n5891), .B(n5890), .ZN(U2968)
         );
  AOI22_X1 U6939 ( .A1(n6258), .A2(REIP_REG_13__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5897) );
  XNOR2_X1 U6940 ( .A(n5892), .B(n5893), .ZN(n5934) );
  AOI22_X1 U6941 ( .A1(n6199), .A2(n5934), .B1(n5895), .B2(n5894), .ZN(n5896)
         );
  OAI211_X1 U6942 ( .C1(n6204), .C2(n5898), .A(n5897), .B(n5896), .ZN(U2973)
         );
  AOI22_X1 U6943 ( .A1(n5899), .A2(n6292), .B1(n6286), .B2(n5971), .ZN(n5904)
         );
  NAND2_X1 U6944 ( .A1(n6258), .A2(REIP_REG_18__SCAN_IN), .ZN(n5903) );
  NAND3_X1 U6945 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5911), .A3(n5900), .ZN(n5902) );
  OAI221_X1 U6946 ( .B1(n5909), .B2(n6281), .C1(n5909), .C2(n5910), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5901) );
  NAND4_X1 U6947 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(U3000)
         );
  AOI22_X1 U6948 ( .A1(n5906), .A2(n6292), .B1(n6286), .B2(n5905), .ZN(n5913)
         );
  NOR2_X1 U6949 ( .A1(n5907), .A2(n6667), .ZN(n5908) );
  AOI221_X1 U6950 ( .B1(n5911), .B2(n5910), .C1(n5909), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5908), .ZN(n5912) );
  NAND2_X1 U6951 ( .A1(n5913), .A2(n5912), .ZN(U3001) );
  OAI21_X1 U6952 ( .B1(n5914), .B2(n6220), .A(n6215), .ZN(n5927) );
  NOR2_X1 U6953 ( .A1(n5907), .A2(n5631), .ZN(n5918) );
  OAI22_X1 U6954 ( .A1(n5916), .A2(n6208), .B1(n6274), .B2(n5915), .ZN(n5917)
         );
  AOI211_X1 U6955 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5927), .A(n5918), .B(n5917), .ZN(n5923) );
  NOR3_X1 U6956 ( .A1(n6205), .A2(n5920), .A3(n5919), .ZN(n5929) );
  OAI221_X1 U6957 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5928), .C2(n5921), .A(n5929), 
        .ZN(n5922) );
  NAND2_X1 U6958 ( .A1(n5923), .A2(n5922), .ZN(U3002) );
  AOI22_X1 U6959 ( .A1(n5925), .A2(n6292), .B1(n6286), .B2(n5924), .ZN(n5931)
         );
  NOR2_X1 U6960 ( .A1(n5907), .A2(n6554), .ZN(n5926) );
  AOI221_X1 U6961 ( .B1(n5929), .B2(n5928), .C1(n5927), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5926), .ZN(n5930) );
  NAND2_X1 U6962 ( .A1(n5931), .A2(n5930), .ZN(U3003) );
  AOI22_X1 U6963 ( .A1(n5932), .A2(n6286), .B1(n6258), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5936) );
  AOI22_X1 U6964 ( .A1(n5934), .A2(n6292), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5933), .ZN(n5935) );
  OAI211_X1 U6965 ( .C1(n6205), .C2(n5937), .A(n5936), .B(n5935), .ZN(U3005)
         );
  INV_X1 U6966 ( .A(n4274), .ZN(n5939) );
  INV_X1 U6967 ( .A(n6036), .ZN(n5938) );
  NAND4_X1 U6968 ( .A1(n5940), .A2(n5939), .A3(n6593), .A4(n5938), .ZN(n5941)
         );
  OAI21_X1 U6969 ( .B1(n5942), .B2(n4470), .A(n5941), .ZN(U3455) );
  AOI21_X1 U6970 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6528), .A(n6522), .ZN(n5947) );
  INV_X1 U6971 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5943) );
  INV_X1 U6972 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6518) );
  NOR2_X2 U6973 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6518), .ZN(n6620) );
  AOI21_X1 U6974 ( .B1(n5947), .B2(n5943), .A(n6620), .ZN(U2789) );
  OAI21_X1 U6975 ( .B1(n5944), .B2(n6499), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5945) );
  OAI21_X1 U6976 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6500), .A(n5945), .ZN(
        U2790) );
  NOR2_X1 U6977 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5948) );
  OAI21_X1 U6978 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5948), .A(n6609), .ZN(n5946)
         );
  OAI21_X1 U6979 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6609), .A(n5946), .ZN(
        U2791) );
  NOR2_X1 U6980 ( .A1(n6620), .A2(n5947), .ZN(n6586) );
  OAI21_X1 U6981 ( .B1(n5948), .B2(BS16_N), .A(n6586), .ZN(n6584) );
  OAI21_X1 U6982 ( .B1(n6586), .B2(n5002), .A(n6584), .ZN(U2792) );
  OAI21_X1 U6983 ( .B1(n5950), .B2(n5949), .A(n6178), .ZN(U2793) );
  NOR4_X1 U6984 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5954) );
  NOR4_X1 U6985 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5953) );
  NOR4_X1 U6986 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5952) );
  NOR4_X1 U6987 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5951) );
  NAND4_X1 U6988 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n5960)
         );
  NOR4_X1 U6989 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n5958) );
  AOI211_X1 U6990 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n5957) );
  NOR4_X1 U6991 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5956)
         );
  NOR4_X1 U6992 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5955) );
  NAND4_X1 U6993 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n5959)
         );
  NOR2_X1 U6994 ( .A1(n5960), .A2(n5959), .ZN(n6604) );
  INV_X1 U6995 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5962) );
  NOR3_X1 U6996 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5963) );
  OAI21_X1 U6997 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5963), .A(n6604), .ZN(n5961)
         );
  OAI21_X1 U6998 ( .B1(n6604), .B2(n5962), .A(n5961), .ZN(U2794) );
  INV_X1 U6999 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6585) );
  AOI21_X1 U7000 ( .B1(n6600), .B2(n6585), .A(n5963), .ZN(n5965) );
  INV_X1 U7001 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5964) );
  INV_X1 U7002 ( .A(n6604), .ZN(n6606) );
  AOI22_X1 U7003 ( .A1(n6604), .A2(n5965), .B1(n5964), .B2(n6606), .ZN(U2795)
         );
  INV_X1 U7004 ( .A(n5966), .ZN(n5974) );
  AOI22_X1 U7005 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6056), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5967), .ZN(n5968) );
  OAI21_X1 U7006 ( .B1(n5969), .B2(n6061), .A(n5968), .ZN(n5970) );
  AOI211_X1 U7007 ( .C1(n6024), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6038), 
        .B(n5970), .ZN(n5973) );
  AOI22_X1 U7008 ( .A1(n6062), .A2(n6018), .B1(n6045), .B2(n5971), .ZN(n5972)
         );
  OAI211_X1 U7009 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5974), .A(n5973), .B(n5972), .ZN(U2809) );
  AOI22_X1 U7010 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6045), 
        .B2(n5975), .ZN(n5984) );
  AOI21_X1 U7011 ( .B1(EBX_REG_11__SCAN_IN), .B2(n6056), .A(n6038), .ZN(n5983)
         );
  INV_X1 U7012 ( .A(n5976), .ZN(n6172) );
  OAI22_X1 U7013 ( .A1(n6174), .A2(n5977), .B1(n6061), .B2(n6172), .ZN(n5978)
         );
  INV_X1 U7014 ( .A(n5978), .ZN(n5982) );
  OAI21_X1 U7015 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5980), .A(n5979), .ZN(n5981) );
  NAND4_X1 U7016 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(U2816)
         );
  INV_X1 U7017 ( .A(n6010), .ZN(n5985) );
  AOI22_X1 U7018 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6056), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5985), .ZN(n5999) );
  INV_X1 U7019 ( .A(n5986), .ZN(n5989) );
  INV_X1 U7020 ( .A(n5987), .ZN(n5988) );
  AOI21_X1 U7021 ( .B1(n5990), .B2(n5989), .A(n5988), .ZN(n6621) );
  OAI21_X1 U7022 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5991), .A(n6030), .ZN(n5994)
         );
  NOR2_X1 U7023 ( .A1(n6051), .A2(n5992), .ZN(n5993) );
  AOI211_X1 U7024 ( .C1(n6621), .C2(n6045), .A(n5994), .B(n5993), .ZN(n5998)
         );
  INV_X1 U7025 ( .A(n5995), .ZN(n6623) );
  AOI22_X1 U7026 ( .A1(n6623), .A2(n6018), .B1(n6027), .B2(n5996), .ZN(n5997)
         );
  NAND3_X1 U7027 ( .A1(n5999), .A2(n5998), .A3(n5997), .ZN(U2818) );
  AOI21_X1 U7028 ( .B1(n6000), .B2(n6017), .A(REIP_REG_8__SCAN_IN), .ZN(n6011)
         );
  AOI21_X1 U7029 ( .B1(n6056), .B2(EBX_REG_8__SCAN_IN), .A(n6038), .ZN(n6001)
         );
  OAI21_X1 U7030 ( .B1(n6002), .B2(n6014), .A(n6001), .ZN(n6003) );
  AOI21_X1 U7031 ( .B1(n6024), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6003), 
        .ZN(n6009) );
  INV_X1 U7032 ( .A(n6004), .ZN(n6007) );
  INV_X1 U7033 ( .A(n6005), .ZN(n6006) );
  AOI22_X1 U7034 ( .A1(n6007), .A2(n6018), .B1(n6006), .B2(n6027), .ZN(n6008)
         );
  OAI211_X1 U7035 ( .C1(n6011), .C2(n6010), .A(n6009), .B(n6008), .ZN(U2819)
         );
  NAND2_X1 U7036 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6013)
         );
  AOI21_X1 U7037 ( .B1(n6056), .B2(EBX_REG_6__SCAN_IN), .A(n6038), .ZN(n6012)
         );
  OAI211_X1 U7038 ( .C1(n6015), .C2(n6014), .A(n6013), .B(n6012), .ZN(n6016)
         );
  AOI221_X1 U7039 ( .B1(n6023), .B2(REIP_REG_6__SCAN_IN), .C1(n6017), .C2(
        n6537), .A(n6016), .ZN(n6020) );
  NAND2_X1 U7040 ( .A1(n6180), .A2(n6018), .ZN(n6019) );
  OAI211_X1 U7041 ( .C1(n6061), .C2(n6184), .A(n6020), .B(n6019), .ZN(U2821)
         );
  NAND2_X1 U7042 ( .A1(n6535), .A2(n6021), .ZN(n6022) );
  AOI22_X1 U7043 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6056), .B1(n6023), .B2(n6022), 
        .ZN(n6033) );
  AOI22_X1 U7044 ( .A1(n6024), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6045), 
        .B2(n6256), .ZN(n6032) );
  INV_X1 U7045 ( .A(n6025), .ZN(n6029) );
  INV_X1 U7046 ( .A(n6026), .ZN(n6058) );
  AOI22_X1 U7047 ( .A1(n6029), .A2(n6058), .B1(n6028), .B2(n6027), .ZN(n6031)
         );
  NAND4_X1 U7048 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(U2822)
         );
  AOI22_X1 U7049 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6056), .B1(
        REIP_REG_4__SCAN_IN), .B2(n6034), .ZN(n6043) );
  INV_X1 U7050 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6685) );
  NOR3_X1 U7051 ( .A1(n6600), .A2(n4733), .A3(n6530), .ZN(n6035) );
  NAND3_X1 U7052 ( .A1(n6044), .A2(n6035), .A3(n6533), .ZN(n6040) );
  NOR2_X1 U7053 ( .A1(n6036), .A2(n6048), .ZN(n6037) );
  AOI211_X1 U7054 ( .C1(n6045), .C2(n6265), .A(n6038), .B(n6037), .ZN(n6039)
         );
  OAI211_X1 U7055 ( .C1(n6685), .C2(n6051), .A(n6040), .B(n6039), .ZN(n6041)
         );
  AOI21_X1 U7056 ( .B1(n6058), .B2(n6189), .A(n6041), .ZN(n6042) );
  OAI211_X1 U7057 ( .C1(n6193), .C2(n6061), .A(n6043), .B(n6042), .ZN(U2823)
         );
  AOI22_X1 U7058 ( .A1(n6046), .A2(n6045), .B1(n6044), .B2(n6600), .ZN(n6047)
         );
  OAI21_X1 U7059 ( .B1(n6049), .B2(n6048), .A(n6047), .ZN(n6053) );
  NOR2_X1 U7060 ( .A1(n6051), .A2(n6050), .ZN(n6052) );
  AOI211_X1 U7061 ( .C1(n6054), .C2(REIP_REG_1__SCAN_IN), .A(n6053), .B(n6052), 
        .ZN(n6060) );
  INV_X1 U7062 ( .A(n6055), .ZN(n6057) );
  AOI22_X1 U7063 ( .A1(n6058), .A2(n6057), .B1(n6056), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n6059) );
  OAI211_X1 U7064 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6061), .A(n6060), 
        .B(n6059), .ZN(U2826) );
  AOI22_X1 U7065 ( .A1(n6062), .A2(n6072), .B1(n6065), .B2(DATAI_18_), .ZN(
        n6064) );
  AOI22_X1 U7066 ( .A1(n6068), .A2(DATAI_2_), .B1(n6067), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7067 ( .A1(n6064), .A2(n6063), .ZN(U2873) );
  AOI22_X1 U7068 ( .A1(n6066), .A2(n6072), .B1(n6065), .B2(DATAI_16_), .ZN(
        n6070) );
  AOI22_X1 U7069 ( .A1(n6068), .A2(DATAI_0_), .B1(n6067), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7070 ( .A1(n6070), .A2(n6069), .ZN(U2875) );
  INV_X1 U7071 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7072 ( .A1(n6623), .A2(n6072), .B1(n6071), .B2(DATAI_9_), .ZN(
        n6073) );
  OAI21_X1 U7073 ( .B1(n6654), .B2(n6074), .A(n6073), .ZN(U2882) );
  INV_X1 U7074 ( .A(n6075), .ZN(n6076) );
  AOI22_X1 U7075 ( .A1(n6090), .A2(DATAO_REG_25__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6076), .ZN(n6077) );
  OAI21_X1 U7076 ( .B1(n6659), .B2(n6487), .A(n6077), .ZN(U2898) );
  AOI22_X1 U7077 ( .A1(n6094), .A2(LWORD_REG_15__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6078) );
  OAI21_X1 U7078 ( .B1(n3636), .B2(n6096), .A(n6078), .ZN(U2908) );
  AOI22_X1 U7079 ( .A1(n6094), .A2(LWORD_REG_14__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U7080 ( .B1(n5520), .B2(n6096), .A(n6079), .ZN(U2909) );
  AOI22_X1 U7081 ( .A1(n6094), .A2(LWORD_REG_13__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7082 ( .B1(n5522), .B2(n6096), .A(n6080), .ZN(U2910) );
  AOI22_X1 U7083 ( .A1(n6094), .A2(LWORD_REG_12__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U7084 ( .B1(n5229), .B2(n6096), .A(n6081), .ZN(U2911) );
  INV_X1 U7085 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6156) );
  AOI22_X1 U7086 ( .A1(n6094), .A2(LWORD_REG_11__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7087 ( .B1(n6156), .B2(n6096), .A(n6082), .ZN(U2912) );
  INV_X1 U7088 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6153) );
  AOI22_X1 U7089 ( .A1(n6094), .A2(LWORD_REG_10__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6083) );
  OAI21_X1 U7090 ( .B1(n6153), .B2(n6096), .A(n6083), .ZN(U2913) );
  AOI22_X1 U7091 ( .A1(n6094), .A2(LWORD_REG_9__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7092 ( .B1(n6654), .B2(n6096), .A(n6084), .ZN(U2914) );
  INV_X1 U7093 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6147) );
  AOI22_X1 U7094 ( .A1(n6094), .A2(LWORD_REG_8__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6085) );
  OAI21_X1 U7095 ( .B1(n6147), .B2(n6096), .A(n6085), .ZN(U2915) );
  AOI22_X1 U7096 ( .A1(n6094), .A2(LWORD_REG_7__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U7097 ( .B1(n4957), .B2(n6096), .A(n6086), .ZN(U2916) );
  AOI22_X1 U7098 ( .A1(n6094), .A2(LWORD_REG_6__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7099 ( .B1(n4811), .B2(n6096), .A(n6087), .ZN(U2917) );
  AOI22_X1 U7100 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6094), .B1(
        DATAO_REG_5__SCAN_IN), .B2(n6090), .ZN(n6088) );
  OAI21_X1 U7101 ( .B1(n6140), .B2(n6096), .A(n6088), .ZN(U2918) );
  AOI22_X1 U7102 ( .A1(n6094), .A2(LWORD_REG_4__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7103 ( .B1(n6137), .B2(n6096), .A(n6089), .ZN(U2919) );
  AOI22_X1 U7104 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6094), .B1(n6090), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7105 ( .B1(n6134), .B2(n6096), .A(n6091), .ZN(U2920) );
  AOI22_X1 U7106 ( .A1(n6094), .A2(LWORD_REG_2__SCAN_IN), .B1(n6090), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6092) );
  OAI21_X1 U7107 ( .B1(n3423), .B2(n6096), .A(n6092), .ZN(U2921) );
  AOI22_X1 U7108 ( .A1(DATAO_REG_1__SCAN_IN), .A2(n6090), .B1(n6094), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7109 ( .B1(n4437), .B2(n6096), .A(n6093), .ZN(U2922) );
  AOI22_X1 U7110 ( .A1(DATAO_REG_0__SCAN_IN), .A2(n6090), .B1(n6094), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7111 ( .B1(n3419), .B2(n6096), .A(n6095), .ZN(U2923) );
  INV_X1 U7112 ( .A(n6124), .ZN(n6164) );
  AND2_X1 U7113 ( .A1(n6164), .A2(DATAI_0_), .ZN(n6126) );
  AOI21_X1 U7114 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6162), .A(n6126), .ZN(n6097) );
  OAI21_X1 U7115 ( .B1(n3664), .B2(n6166), .A(n6097), .ZN(U2924) );
  NOR2_X1 U7116 ( .A1(n6124), .A2(n6098), .ZN(n6128) );
  AOI21_X1 U7117 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6149), .A(n6128), .ZN(n6099) );
  OAI21_X1 U7118 ( .B1(n6100), .B2(n6166), .A(n6099), .ZN(U2925) );
  AND2_X1 U7119 ( .A1(n6164), .A2(DATAI_2_), .ZN(n6130) );
  AOI21_X1 U7120 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6162), .A(n6130), .ZN(n6101) );
  OAI21_X1 U7121 ( .B1(n3698), .B2(n6166), .A(n6101), .ZN(U2926) );
  AND2_X1 U7122 ( .A1(n6164), .A2(DATAI_3_), .ZN(n6132) );
  AOI21_X1 U7123 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6162), .A(n6132), .ZN(n6102) );
  OAI21_X1 U7124 ( .B1(n6103), .B2(n6166), .A(n6102), .ZN(U2927) );
  AND2_X1 U7125 ( .A1(n6164), .A2(DATAI_4_), .ZN(n6135) );
  AOI21_X1 U7126 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6162), .A(n6135), .ZN(n6104) );
  OAI21_X1 U7127 ( .B1(n6105), .B2(n6166), .A(n6104), .ZN(U2928) );
  AND2_X1 U7128 ( .A1(n6164), .A2(DATAI_5_), .ZN(n6138) );
  AOI21_X1 U7129 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6162), .A(n6138), .ZN(n6106) );
  OAI21_X1 U7130 ( .B1(n6701), .B2(n6166), .A(n6106), .ZN(U2929) );
  NOR2_X1 U7131 ( .A1(n6124), .A2(n6107), .ZN(n6141) );
  AOI21_X1 U7132 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6149), .A(n6141), .ZN(n6108) );
  OAI21_X1 U7133 ( .B1(n3771), .B2(n6166), .A(n6108), .ZN(U2930) );
  NOR2_X1 U7134 ( .A1(n6124), .A2(n6109), .ZN(n6143) );
  AOI21_X1 U7135 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6149), .A(n6143), .ZN(n6110) );
  OAI21_X1 U7136 ( .B1(n3802), .B2(n6166), .A(n6110), .ZN(U2931) );
  INV_X1 U7137 ( .A(DATAI_8_), .ZN(n6111) );
  NOR2_X1 U7138 ( .A1(n6124), .A2(n6111), .ZN(n6145) );
  AOI21_X1 U7139 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6149), .A(n6145), .ZN(n6112) );
  OAI21_X1 U7140 ( .B1(n3823), .B2(n6166), .A(n6112), .ZN(U2932) );
  INV_X1 U7141 ( .A(DATAI_10_), .ZN(n6114) );
  NOR2_X1 U7142 ( .A1(n6124), .A2(n6114), .ZN(n6151) );
  AOI21_X1 U7143 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6162), .A(n6151), .ZN(
        n6115) );
  OAI21_X1 U7144 ( .B1(n6706), .B2(n6166), .A(n6115), .ZN(U2934) );
  INV_X1 U7145 ( .A(DATAI_11_), .ZN(n6116) );
  NOR2_X1 U7146 ( .A1(n6124), .A2(n6116), .ZN(n6154) );
  AOI21_X1 U7147 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6162), .A(n6154), .ZN(
        n6117) );
  OAI21_X1 U7148 ( .B1(n6118), .B2(n6166), .A(n6117), .ZN(U2935) );
  NOR2_X1 U7149 ( .A1(n6124), .A2(n6119), .ZN(n6157) );
  AOI21_X1 U7150 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6162), .A(n6157), .ZN(
        n6120) );
  OAI21_X1 U7151 ( .B1(n3904), .B2(n6166), .A(n6120), .ZN(U2936) );
  NOR2_X1 U7152 ( .A1(n6124), .A2(n6121), .ZN(n6159) );
  AOI21_X1 U7153 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6162), .A(n6159), .ZN(
        n6122) );
  OAI21_X1 U7154 ( .B1(n3930), .B2(n6166), .A(n6122), .ZN(U2937) );
  NOR2_X1 U7155 ( .A1(n6124), .A2(n6123), .ZN(n6161) );
  AOI21_X1 U7156 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6162), .A(n6161), .ZN(
        n6125) );
  OAI21_X1 U7157 ( .B1(n3966), .B2(n6166), .A(n6125), .ZN(U2938) );
  AOI21_X1 U7158 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6162), .A(n6126), .ZN(n6127) );
  OAI21_X1 U7159 ( .B1(n3419), .B2(n6166), .A(n6127), .ZN(U2939) );
  AOI21_X1 U7160 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6162), .A(n6128), .ZN(n6129) );
  OAI21_X1 U7161 ( .B1(n4437), .B2(n6166), .A(n6129), .ZN(U2940) );
  AOI21_X1 U7162 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6162), .A(n6130), .ZN(n6131) );
  OAI21_X1 U7163 ( .B1(n3423), .B2(n6166), .A(n6131), .ZN(U2941) );
  AOI21_X1 U7164 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6162), .A(n6132), .ZN(n6133) );
  OAI21_X1 U7165 ( .B1(n6134), .B2(n6166), .A(n6133), .ZN(U2942) );
  AOI21_X1 U7166 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6149), .A(n6135), .ZN(n6136) );
  OAI21_X1 U7167 ( .B1(n6137), .B2(n6166), .A(n6136), .ZN(U2943) );
  AOI21_X1 U7168 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6149), .A(n6138), .ZN(n6139) );
  OAI21_X1 U7169 ( .B1(n6140), .B2(n6166), .A(n6139), .ZN(U2944) );
  AOI21_X1 U7170 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6149), .A(n6141), .ZN(n6142) );
  OAI21_X1 U7171 ( .B1(n4811), .B2(n6166), .A(n6142), .ZN(U2945) );
  AOI21_X1 U7172 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6149), .A(n6143), .ZN(n6144) );
  OAI21_X1 U7173 ( .B1(n4957), .B2(n6166), .A(n6144), .ZN(U2946) );
  AOI21_X1 U7174 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6162), .A(n6145), .ZN(n6146) );
  OAI21_X1 U7175 ( .B1(n6147), .B2(n6166), .A(n6146), .ZN(U2947) );
  AOI21_X1 U7176 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6149), .A(n6148), .ZN(n6150) );
  OAI21_X1 U7177 ( .B1(n6654), .B2(n6166), .A(n6150), .ZN(U2948) );
  AOI21_X1 U7178 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6162), .A(n6151), .ZN(
        n6152) );
  OAI21_X1 U7179 ( .B1(n6153), .B2(n6166), .A(n6152), .ZN(U2949) );
  AOI21_X1 U7180 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6162), .A(n6154), .ZN(
        n6155) );
  OAI21_X1 U7181 ( .B1(n6156), .B2(n6166), .A(n6155), .ZN(U2950) );
  AOI21_X1 U7182 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6162), .A(n6157), .ZN(
        n6158) );
  OAI21_X1 U7183 ( .B1(n5229), .B2(n6166), .A(n6158), .ZN(U2951) );
  AOI21_X1 U7184 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6162), .A(n6159), .ZN(
        n6160) );
  OAI21_X1 U7185 ( .B1(n5522), .B2(n6166), .A(n6160), .ZN(U2952) );
  AOI21_X1 U7186 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6162), .A(n6161), .ZN(
        n6163) );
  OAI21_X1 U7187 ( .B1(n5520), .B2(n6166), .A(n6163), .ZN(U2953) );
  AOI22_X1 U7188 ( .A1(n6149), .A2(LWORD_REG_15__SCAN_IN), .B1(n6164), .B2(
        DATAI_15_), .ZN(n6165) );
  OAI21_X1 U7189 ( .B1(n3636), .B2(n6166), .A(n6165), .ZN(U2954) );
  NAND2_X1 U7190 ( .A1(n6168), .A2(n6167), .ZN(n6171) );
  XNOR2_X1 U7191 ( .A(n6169), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6170)
         );
  XNOR2_X1 U7192 ( .A(n6171), .B(n6170), .ZN(n6209) );
  AOI22_X1 U7193 ( .A1(n6258), .A2(REIP_REG_11__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6177) );
  OAI22_X1 U7194 ( .A1(n6174), .A2(n6173), .B1(n6204), .B2(n6172), .ZN(n6175)
         );
  INV_X1 U7195 ( .A(n6175), .ZN(n6176) );
  OAI211_X1 U7196 ( .C1(n6209), .C2(n6178), .A(n6177), .B(n6176), .ZN(U2975)
         );
  AOI22_X1 U7197 ( .A1(n6258), .A2(REIP_REG_6__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6183) );
  INV_X1 U7198 ( .A(n6179), .ZN(n6181) );
  AOI22_X1 U7199 ( .A1(n6181), .A2(n6199), .B1(n5894), .B2(n6180), .ZN(n6182)
         );
  OAI211_X1 U7200 ( .C1(n6204), .C2(n6184), .A(n6183), .B(n6182), .ZN(U2980)
         );
  AOI22_X1 U7201 ( .A1(n6206), .A2(REIP_REG_4__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7202 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  NAND2_X1 U7203 ( .A1(n6185), .A2(n6188), .ZN(n6264) );
  INV_X1 U7204 ( .A(n6264), .ZN(n6190) );
  AOI22_X1 U7205 ( .A1(n6190), .A2(n6199), .B1(n5894), .B2(n6189), .ZN(n6191)
         );
  OAI211_X1 U7206 ( .C1(n6204), .C2(n6193), .A(n6192), .B(n6191), .ZN(U2982)
         );
  AOI22_X1 U7207 ( .A1(n6206), .A2(REIP_REG_2__SCAN_IN), .B1(n6194), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6202) );
  INV_X1 U7208 ( .A(n6195), .ZN(n6200) );
  XNOR2_X1 U7209 ( .A(n6197), .B(n3994), .ZN(n6198) );
  XNOR2_X1 U7210 ( .A(n6196), .B(n6198), .ZN(n6291) );
  AOI22_X1 U7211 ( .A1(n5894), .A2(n6200), .B1(n6291), .B2(n6199), .ZN(n6201)
         );
  OAI211_X1 U7212 ( .C1(n6204), .C2(n6203), .A(n6202), .B(n6201), .ZN(U2984)
         );
  INV_X1 U7213 ( .A(n6205), .ZN(n6212) );
  OAI22_X1 U7214 ( .A1(n6274), .A2(n6207), .B1(n6547), .B2(n5907), .ZN(n6211)
         );
  NOR2_X1 U7215 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  AOI211_X1 U7216 ( .C1(n6214), .C2(n6212), .A(n6211), .B(n6210), .ZN(n6213)
         );
  OAI21_X1 U7217 ( .B1(n6215), .B2(n6214), .A(n6213), .ZN(U3007) );
  AOI21_X1 U7218 ( .B1(n6216), .B2(n6283), .A(n6282), .ZN(n6278) );
  NOR2_X1 U7219 ( .A1(n6218), .A2(n6217), .ZN(n6221) );
  AOI22_X1 U7220 ( .A1(n6278), .A2(n6221), .B1(n6220), .B2(n6219), .ZN(n6247)
         );
  AOI21_X1 U7221 ( .B1(n6238), .B2(n6222), .A(n6247), .ZN(n6237) );
  AOI222_X1 U7222 ( .A1(n6224), .A2(n6292), .B1(n6286), .B2(n6223), .C1(
        REIP_REG_10__SCAN_IN), .C2(n6258), .ZN(n6229) );
  NAND3_X1 U7223 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6226), .A3(n6225), 
        .ZN(n6251) );
  NOR2_X1 U7224 ( .A1(n6238), .A2(n6251), .ZN(n6232) );
  OAI211_X1 U7225 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6232), .B(n6227), .ZN(n6228) );
  OAI211_X1 U7226 ( .C1(n6237), .C2(n4054), .A(n6229), .B(n6228), .ZN(U3008)
         );
  INV_X1 U7227 ( .A(n6230), .ZN(n6231) );
  AOI21_X1 U7228 ( .B1(n6286), .B2(n6621), .A(n6231), .ZN(n6235) );
  AOI22_X1 U7229 ( .A1(n6233), .A2(n6292), .B1(n6232), .B2(n6236), .ZN(n6234)
         );
  OAI211_X1 U7230 ( .C1(n6237), .C2(n6236), .A(n6235), .B(n6234), .ZN(U3009)
         );
  OAI21_X1 U7231 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6238), .ZN(n6244) );
  AOI21_X1 U7232 ( .B1(n6286), .B2(n6240), .A(n6239), .ZN(n6243) );
  AOI22_X1 U7233 ( .A1(n6241), .A2(n6292), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6247), .ZN(n6242) );
  OAI211_X1 U7234 ( .C1(n6251), .C2(n6244), .A(n6243), .B(n6242), .ZN(U3010)
         );
  AOI21_X1 U7235 ( .B1(n6286), .B2(n6246), .A(n6245), .ZN(n6250) );
  AOI22_X1 U7236 ( .A1(n6248), .A2(n6292), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6247), .ZN(n6249) );
  OAI211_X1 U7237 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6251), .A(n6250), 
        .B(n6249), .ZN(U3011) );
  INV_X1 U7238 ( .A(n6263), .ZN(n6252) );
  AOI211_X1 U7239 ( .C1(n6253), .C2(n6288), .A(n6283), .B(n6252), .ZN(n6254)
         );
  NOR2_X1 U7240 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6254), .ZN(n6261)
         );
  INV_X1 U7241 ( .A(n6255), .ZN(n6257) );
  AOI22_X1 U7242 ( .A1(n6257), .A2(n6292), .B1(n6286), .B2(n6256), .ZN(n6260)
         );
  NAND2_X1 U7243 ( .A1(n6258), .A2(REIP_REG_5__SCAN_IN), .ZN(n6259) );
  OAI211_X1 U7244 ( .C1(n6262), .C2(n6261), .A(n6260), .B(n6259), .ZN(U3013)
         );
  AOI211_X1 U7245 ( .C1(n6271), .C2(n6279), .A(n6263), .B(n6280), .ZN(n6269)
         );
  NOR2_X1 U7246 ( .A1(n6264), .A2(n6208), .ZN(n6268) );
  NAND2_X1 U7247 ( .A1(n6286), .A2(n6265), .ZN(n6266) );
  OAI21_X1 U7248 ( .B1(n6533), .B2(n5907), .A(n6266), .ZN(n6267) );
  NOR3_X1 U7249 ( .A1(n6269), .A2(n6268), .A3(n6267), .ZN(n6270) );
  OAI21_X1 U7250 ( .B1(n6278), .B2(n6271), .A(n6270), .ZN(U3014) );
  AND3_X1 U7251 ( .A1(n4739), .A2(n6272), .A3(n6292), .ZN(n6276) );
  OAI22_X1 U7252 ( .A1(n6274), .A2(n6273), .B1(n4733), .B2(n5907), .ZN(n6275)
         );
  NOR2_X1 U7253 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  OAI221_X1 U7254 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6280), .C1(n6279), .C2(n6278), .A(n6277), .ZN(U3015) );
  NAND2_X1 U7255 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6281), .ZN(n6295)
         );
  INV_X1 U7256 ( .A(n6282), .ZN(n6294) );
  AOI21_X1 U7257 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6284), .A(n6283), 
        .ZN(n6289) );
  AOI22_X1 U7258 ( .A1(n6286), .A2(n6285), .B1(n6206), .B2(REIP_REG_2__SCAN_IN), .ZN(n6287) );
  OAI21_X1 U7259 ( .B1(n6289), .B2(n6288), .A(n6287), .ZN(n6290) );
  AOI21_X1 U7260 ( .B1(n6292), .B2(n6291), .A(n6290), .ZN(n6293) );
  OAI221_X1 U7261 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6295), .C1(n3994), .C2(n6294), .A(n6293), .ZN(U3016) );
  NOR2_X1 U7262 ( .A1(n6297), .A2(n6296), .ZN(U3019) );
  NOR2_X1 U7263 ( .A1(n6392), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6328)
         );
  AOI22_X1 U7264 ( .A1(n6321), .A2(n6298), .B1(n6393), .B2(n6328), .ZN(n6308)
         );
  INV_X1 U7265 ( .A(n6299), .ZN(n6397) );
  OAI21_X1 U7266 ( .B1(n6300), .B2(n6397), .A(n6396), .ZN(n6306) );
  AOI21_X1 U7267 ( .B1(n6301), .B2(n3418), .A(n6328), .ZN(n6305) );
  INV_X1 U7268 ( .A(n6305), .ZN(n6303) );
  NAND2_X1 U7269 ( .A1(n6400), .A2(n6304), .ZN(n6302) );
  OAI211_X1 U7270 ( .C1(n6306), .C2(n6303), .A(n6402), .B(n6302), .ZN(n6331)
         );
  OAI22_X1 U7271 ( .A1(n6306), .A2(n6305), .B1(n6304), .B2(n3407), .ZN(n6330)
         );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6331), .B1(n6407), 
        .B2(n6330), .ZN(n6307) );
  OAI211_X1 U7273 ( .C1(n6309), .C2(n6325), .A(n6308), .B(n6307), .ZN(U3044)
         );
  AOI22_X1 U7274 ( .A1(n6329), .A2(n6412), .B1(n6411), .B2(n6328), .ZN(n6311)
         );
  AOI22_X1 U7275 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6331), .B1(n6413), 
        .B2(n6330), .ZN(n6310) );
  OAI211_X1 U7276 ( .C1(n6416), .C2(n6334), .A(n6311), .B(n6310), .ZN(U3045)
         );
  AOI22_X1 U7277 ( .A1(n6329), .A2(n6312), .B1(n6417), .B2(n6328), .ZN(n6314)
         );
  AOI22_X1 U7278 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6331), .B1(n6419), 
        .B2(n6330), .ZN(n6313) );
  OAI211_X1 U7279 ( .C1(n6315), .C2(n6334), .A(n6314), .B(n6313), .ZN(U3046)
         );
  AOI22_X1 U7280 ( .A1(n6329), .A2(n6360), .B1(n6423), .B2(n6328), .ZN(n6317)
         );
  AOI22_X1 U7281 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6331), .B1(n6425), 
        .B2(n6330), .ZN(n6316) );
  OAI211_X1 U7282 ( .C1(n6363), .C2(n6334), .A(n6317), .B(n6316), .ZN(U3047)
         );
  AOI22_X1 U7283 ( .A1(n6329), .A2(n6430), .B1(n6429), .B2(n6328), .ZN(n6319)
         );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6331), .B1(n6431), 
        .B2(n6330), .ZN(n6318) );
  OAI211_X1 U7285 ( .C1(n6434), .C2(n6334), .A(n6319), .B(n6318), .ZN(U3048)
         );
  AOI22_X1 U7286 ( .A1(n6321), .A2(n6320), .B1(n6435), .B2(n6328), .ZN(n6323)
         );
  AOI22_X1 U7287 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6331), .B1(n6437), 
        .B2(n6330), .ZN(n6322) );
  OAI211_X1 U7288 ( .C1(n6325), .C2(n6324), .A(n6323), .B(n6322), .ZN(U3049)
         );
  AOI22_X1 U7289 ( .A1(n6329), .A2(n6372), .B1(n6441), .B2(n6328), .ZN(n6327)
         );
  AOI22_X1 U7290 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6331), .B1(n6444), 
        .B2(n6330), .ZN(n6326) );
  OAI211_X1 U7291 ( .C1(n6375), .C2(n6334), .A(n6327), .B(n6326), .ZN(U3050)
         );
  AOI22_X1 U7292 ( .A1(n6329), .A2(n6451), .B1(n6450), .B2(n6328), .ZN(n6333)
         );
  AOI22_X1 U7293 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6331), .B1(n6454), 
        .B2(n6330), .ZN(n6332) );
  OAI211_X1 U7294 ( .C1(n6459), .C2(n6334), .A(n6333), .B(n6332), .ZN(U3051)
         );
  AOI22_X1 U7295 ( .A1(n6393), .A2(n6336), .B1(n6407), .B2(n6335), .ZN(n6340)
         );
  AOI22_X1 U7296 ( .A1(n6338), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6394), 
        .B2(n6337), .ZN(n6339) );
  OAI211_X1 U7297 ( .C1(n6410), .C2(n6368), .A(n6340), .B(n6339), .ZN(U3068)
         );
  INV_X1 U7298 ( .A(n6341), .ZN(n6377) );
  AOI22_X1 U7299 ( .A1(n6393), .A2(n6377), .B1(n6394), .B2(n6376), .ZN(n6353)
         );
  NOR2_X1 U7300 ( .A1(n6342), .A2(n6400), .ZN(n6348) );
  NOR3_X1 U7301 ( .A1(n6345), .A2(n6344), .A3(n6343), .ZN(n6346) );
  NOR2_X1 U7302 ( .A1(n6346), .A2(n6377), .ZN(n6351) );
  AOI22_X1 U7303 ( .A1(n6348), .A2(n6351), .B1(n6349), .B2(n6400), .ZN(n6347)
         );
  NAND2_X1 U7304 ( .A1(n6402), .A2(n6347), .ZN(n6379) );
  INV_X1 U7305 ( .A(n6348), .ZN(n6350) );
  OAI22_X1 U7306 ( .A1(n6351), .A2(n6350), .B1(n3407), .B2(n6349), .ZN(n6378)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6379), .B1(n6407), 
        .B2(n6378), .ZN(n6352) );
  OAI211_X1 U7308 ( .C1(n6410), .C2(n6390), .A(n6353), .B(n6352), .ZN(U3076)
         );
  AOI22_X1 U7309 ( .A1(n6411), .A2(n6377), .B1(n6354), .B2(n6364), .ZN(n6356)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6379), .B1(n6413), 
        .B2(n6378), .ZN(n6355) );
  OAI211_X1 U7311 ( .C1(n6357), .C2(n6368), .A(n6356), .B(n6355), .ZN(U3077)
         );
  AOI22_X1 U7312 ( .A1(n6417), .A2(n6377), .B1(n6418), .B2(n6364), .ZN(n6359)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6379), .B1(n6419), 
        .B2(n6378), .ZN(n6358) );
  OAI211_X1 U7314 ( .C1(n6422), .C2(n6368), .A(n6359), .B(n6358), .ZN(U3078)
         );
  AOI22_X1 U7315 ( .A1(n6423), .A2(n6377), .B1(n6360), .B2(n6376), .ZN(n6362)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6379), .B1(n6425), 
        .B2(n6378), .ZN(n6361) );
  OAI211_X1 U7317 ( .C1(n6363), .C2(n6390), .A(n6362), .B(n6361), .ZN(U3079)
         );
  AOI22_X1 U7318 ( .A1(n6429), .A2(n6377), .B1(n6365), .B2(n6364), .ZN(n6367)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6379), .B1(n6431), 
        .B2(n6378), .ZN(n6366) );
  OAI211_X1 U7320 ( .C1(n6369), .C2(n6368), .A(n6367), .B(n6366), .ZN(U3080)
         );
  AOI22_X1 U7321 ( .A1(n6435), .A2(n6377), .B1(n6436), .B2(n6376), .ZN(n6371)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6379), .B1(n6437), 
        .B2(n6378), .ZN(n6370) );
  OAI211_X1 U7323 ( .C1(n6440), .C2(n6390), .A(n6371), .B(n6370), .ZN(U3081)
         );
  AOI22_X1 U7324 ( .A1(n6441), .A2(n6377), .B1(n6372), .B2(n6376), .ZN(n6374)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6379), .B1(n6444), 
        .B2(n6378), .ZN(n6373) );
  OAI211_X1 U7326 ( .C1(n6375), .C2(n6390), .A(n6374), .B(n6373), .ZN(U3082)
         );
  AOI22_X1 U7327 ( .A1(n6450), .A2(n6377), .B1(n6451), .B2(n6376), .ZN(n6381)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6379), .B1(n6454), 
        .B2(n6378), .ZN(n6380) );
  OAI211_X1 U7329 ( .C1(n6459), .C2(n6390), .A(n6381), .B(n6380), .ZN(U3083)
         );
  AOI22_X1 U7330 ( .A1(n6423), .A2(n6384), .B1(n6425), .B2(n6385), .ZN(n6383)
         );
  AOI22_X1 U7331 ( .A1(n6387), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6424), 
        .B2(n6386), .ZN(n6382) );
  OAI211_X1 U7332 ( .C1(n6428), .C2(n6390), .A(n6383), .B(n6382), .ZN(U3087)
         );
  AOI22_X1 U7333 ( .A1(n6444), .A2(n6385), .B1(n6441), .B2(n6384), .ZN(n6389)
         );
  AOI22_X1 U7334 ( .A1(n6387), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6443), 
        .B2(n6386), .ZN(n6388) );
  OAI211_X1 U7335 ( .C1(n6448), .C2(n6390), .A(n6389), .B(n6388), .ZN(U3090)
         );
  INV_X1 U7336 ( .A(n6447), .ZN(n6452) );
  NOR2_X1 U7337 ( .A1(n6392), .A2(n6391), .ZN(n6449) );
  AOI22_X1 U7338 ( .A1(n6452), .A2(n6394), .B1(n6393), .B2(n6449), .ZN(n6409)
         );
  INV_X1 U7339 ( .A(n6395), .ZN(n6398) );
  OAI21_X1 U7340 ( .B1(n6398), .B2(n6397), .A(n6396), .ZN(n6406) );
  AOI21_X1 U7341 ( .B1(n6399), .B2(n3418), .A(n6449), .ZN(n6405) );
  INV_X1 U7342 ( .A(n6405), .ZN(n6403) );
  NAND2_X1 U7343 ( .A1(n6400), .A2(n6404), .ZN(n6401) );
  OAI211_X1 U7344 ( .C1(n6406), .C2(n6403), .A(n6402), .B(n6401), .ZN(n6455)
         );
  OAI22_X1 U7345 ( .A1(n6406), .A2(n6405), .B1(n6404), .B2(n3407), .ZN(n6453)
         );
  AOI22_X1 U7346 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6455), .B1(n6407), 
        .B2(n6453), .ZN(n6408) );
  OAI211_X1 U7347 ( .C1(n6410), .C2(n6458), .A(n6409), .B(n6408), .ZN(U3108)
         );
  AOI22_X1 U7348 ( .A1(n6452), .A2(n6412), .B1(n6411), .B2(n6449), .ZN(n6415)
         );
  AOI22_X1 U7349 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6455), .B1(n6413), 
        .B2(n6453), .ZN(n6414) );
  OAI211_X1 U7350 ( .C1(n6416), .C2(n6458), .A(n6415), .B(n6414), .ZN(U3109)
         );
  AOI22_X1 U7351 ( .A1(n6418), .A2(n6442), .B1(n6417), .B2(n6449), .ZN(n6421)
         );
  AOI22_X1 U7352 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6455), .B1(n6419), 
        .B2(n6453), .ZN(n6420) );
  OAI211_X1 U7353 ( .C1(n6422), .C2(n6447), .A(n6421), .B(n6420), .ZN(U3110)
         );
  AOI22_X1 U7354 ( .A1(n6424), .A2(n6442), .B1(n6423), .B2(n6449), .ZN(n6427)
         );
  AOI22_X1 U7355 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6455), .B1(n6425), 
        .B2(n6453), .ZN(n6426) );
  OAI211_X1 U7356 ( .C1(n6428), .C2(n6447), .A(n6427), .B(n6426), .ZN(U3111)
         );
  AOI22_X1 U7357 ( .A1(n6452), .A2(n6430), .B1(n6429), .B2(n6449), .ZN(n6433)
         );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6455), .B1(n6431), 
        .B2(n6453), .ZN(n6432) );
  OAI211_X1 U7359 ( .C1(n6434), .C2(n6458), .A(n6433), .B(n6432), .ZN(U3112)
         );
  AOI22_X1 U7360 ( .A1(n6452), .A2(n6436), .B1(n6435), .B2(n6449), .ZN(n6439)
         );
  AOI22_X1 U7361 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6455), .B1(n6437), 
        .B2(n6453), .ZN(n6438) );
  OAI211_X1 U7362 ( .C1(n6440), .C2(n6458), .A(n6439), .B(n6438), .ZN(U3113)
         );
  AOI22_X1 U7363 ( .A1(n6443), .A2(n6442), .B1(n6441), .B2(n6449), .ZN(n6446)
         );
  AOI22_X1 U7364 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6455), .B1(n6444), 
        .B2(n6453), .ZN(n6445) );
  OAI211_X1 U7365 ( .C1(n6448), .C2(n6447), .A(n6446), .B(n6445), .ZN(U3114)
         );
  AOI22_X1 U7366 ( .A1(n6452), .A2(n6451), .B1(n6450), .B2(n6449), .ZN(n6457)
         );
  AOI22_X1 U7367 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6455), .B1(n6454), 
        .B2(n6453), .ZN(n6456) );
  OAI211_X1 U7368 ( .C1(n6459), .C2(n6458), .A(n6457), .B(n6456), .ZN(U3115)
         );
  NOR3_X1 U7369 ( .A1(n6462), .A2(n6461), .A3(n6460), .ZN(n6466) );
  NAND2_X1 U7370 ( .A1(n6464), .A2(n6463), .ZN(n6465) );
  AOI222_X1 U7371 ( .A1(n6466), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6466), .B2(n6465), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6465), 
        .ZN(n6468) );
  AOI21_X1 U7372 ( .B1(n6468), .B2(n6469), .A(n6467), .ZN(n6472) );
  NOR2_X1 U7373 ( .A1(n6469), .A2(n6468), .ZN(n6471) );
  INV_X1 U7374 ( .A(n6470), .ZN(n6473) );
  OAI22_X1 U7375 ( .A1(n6472), .A2(n6471), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6473), .ZN(n6482) );
  AOI21_X1 U7376 ( .B1(n6473), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U7377 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6474), 
        .ZN(n6475) );
  NAND4_X1 U7378 ( .A1(n6478), .A2(n6477), .A3(n6476), .A4(n6475), .ZN(n6479)
         );
  AOI211_X1 U7379 ( .C1(n6482), .C2(n6481), .A(n6480), .B(n6479), .ZN(n6498)
         );
  INV_X1 U7380 ( .A(n6483), .ZN(n6486) );
  INV_X1 U7381 ( .A(n6588), .ZN(n6485) );
  AOI21_X1 U7382 ( .B1(n6486), .B2(n6485), .A(n6484), .ZN(n6497) );
  INV_X1 U7383 ( .A(n6498), .ZN(n6488) );
  OAI22_X1 U7384 ( .A1(n6488), .A2(n6499), .B1(n6487), .B2(n6612), .ZN(n6489)
         );
  OAI21_X1 U7385 ( .B1(n6491), .B2(n6490), .A(n6489), .ZN(n6590) );
  AOI21_X1 U7386 ( .B1(n6615), .B2(n6492), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6495) );
  NAND2_X1 U7387 ( .A1(READY_N), .A2(n3407), .ZN(n6507) );
  AOI21_X1 U7388 ( .B1(n6507), .B2(n6590), .A(n6493), .ZN(n6494) );
  AOI21_X1 U7389 ( .B1(n6590), .B2(n6495), .A(n6494), .ZN(n6496) );
  OAI211_X1 U7390 ( .C1(n6498), .C2(n6499), .A(n6497), .B(n6496), .ZN(U3148)
         );
  OAI21_X1 U7391 ( .B1(READY_N), .B2(n6500), .A(n6499), .ZN(n6505) );
  AOI211_X1 U7392 ( .C1(n6590), .C2(n6507), .A(n6502), .B(n6501), .ZN(n6503)
         );
  AOI211_X1 U7393 ( .C1(n6590), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6506)
         );
  INV_X1 U7394 ( .A(n6506), .ZN(U3149) );
  NAND4_X1 U7395 ( .A1(n6509), .A2(n6508), .A3(n6507), .A4(n6588), .ZN(n6510)
         );
  NAND2_X1 U7396 ( .A1(n6511), .A2(n6510), .ZN(U3150) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6582), .ZN(U3151) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6582), .ZN(U3152) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6582), .ZN(U3153) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6582), .ZN(U3154) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6582), .ZN(U3155) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6582), .ZN(U3156) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6582), .ZN(U3157) );
  AND2_X1 U7404 ( .A1(n6582), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U7405 ( .A1(n6582), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6582), .ZN(U3160) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6582), .ZN(U3161) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6582), .ZN(U3162) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6582), .ZN(U3163) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6582), .ZN(U3164) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6582), .ZN(U3165) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6582), .ZN(U3166) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6582), .ZN(U3167) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6582), .ZN(U3168) );
  AND2_X1 U7415 ( .A1(n6582), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6582), .ZN(U3170) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6582), .ZN(U3171) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6582), .ZN(U3172) );
  INV_X1 U7419 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U7420 ( .A1(n6586), .A2(n6628), .ZN(U3173) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6582), .ZN(U3174) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6582), .ZN(U3175) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6582), .ZN(U3176) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6582), .ZN(U3177) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6582), .ZN(U3178) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6582), .ZN(U3179) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6582), .ZN(U3180) );
  NOR2_X1 U7428 ( .A1(n6518), .A2(n6528), .ZN(n6519) );
  AOI22_X1 U7429 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6527) );
  AND2_X1 U7430 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6515) );
  INV_X1 U7431 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6513) );
  INV_X1 U7432 ( .A(NA_N), .ZN(n6520) );
  AOI221_X1 U7433 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6520), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6524) );
  AOI221_X1 U7434 ( .B1(n6515), .B2(n6609), .C1(n6513), .C2(n6609), .A(n6524), 
        .ZN(n6512) );
  OAI21_X1 U7435 ( .B1(n6519), .B2(n6527), .A(n6512), .ZN(U3181) );
  NOR2_X1 U7436 ( .A1(n6522), .A2(n6513), .ZN(n6521) );
  NAND2_X1 U7437 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6514) );
  OAI21_X1 U7438 ( .B1(n6521), .B2(n6515), .A(n6514), .ZN(n6516) );
  OAI211_X1 U7439 ( .C1(n6518), .C2(n6612), .A(n6517), .B(n6516), .ZN(U3182)
         );
  AOI21_X1 U7440 ( .B1(n6521), .B2(n6520), .A(n6519), .ZN(n6526) );
  AOI221_X1 U7441 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6612), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6523) );
  AOI221_X1 U7442 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6523), .C2(HOLD), .A(n6522), .ZN(n6525) );
  OAI22_X1 U7443 ( .A1(n6527), .A2(n6526), .B1(n6525), .B2(n6524), .ZN(U3183)
         );
  NAND2_X1 U7444 ( .A1(n6620), .A2(n6528), .ZN(n6574) );
  INV_X1 U7445 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7446 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6620), .ZN(n6579) );
  OAI222_X1 U7447 ( .A1(n6574), .A2(n6530), .B1(n6529), .B2(n6620), .C1(n6600), 
        .C2(n6579), .ZN(U3184) );
  INV_X1 U7448 ( .A(n6579), .ZN(n6572) );
  AOI22_X1 U7449 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6609), .ZN(n6531) );
  OAI21_X1 U7450 ( .B1(n4733), .B2(n6574), .A(n6531), .ZN(U3185) );
  AOI22_X1 U7451 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6609), .ZN(n6532) );
  OAI21_X1 U7452 ( .B1(n6533), .B2(n6574), .A(n6532), .ZN(U3186) );
  AOI22_X1 U7453 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6609), .ZN(n6534) );
  OAI21_X1 U7454 ( .B1(n6535), .B2(n6574), .A(n6534), .ZN(U3187) );
  INV_X1 U7455 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6536) );
  OAI222_X1 U7456 ( .A1(n6574), .A2(n6537), .B1(n6536), .B2(n6620), .C1(n6535), 
        .C2(n6579), .ZN(U3188) );
  AOI22_X1 U7457 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6609), .ZN(n6538) );
  OAI21_X1 U7458 ( .B1(n6540), .B2(n6574), .A(n6538), .ZN(U3189) );
  INV_X1 U7459 ( .A(n6574), .ZN(n6577) );
  AOI22_X1 U7460 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6609), .ZN(n6539) );
  OAI21_X1 U7461 ( .B1(n6540), .B2(n6579), .A(n6539), .ZN(U3190) );
  INV_X1 U7462 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6542) );
  AOI22_X1 U7463 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6609), .ZN(n6541) );
  OAI21_X1 U7464 ( .B1(n6542), .B2(n6574), .A(n6541), .ZN(U3191) );
  AOI22_X1 U7465 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6609), .ZN(n6543) );
  OAI21_X1 U7466 ( .B1(n6545), .B2(n6574), .A(n6543), .ZN(U3192) );
  INV_X1 U7467 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6544) );
  OAI222_X1 U7468 ( .A1(n6579), .A2(n6545), .B1(n6544), .B2(n6620), .C1(n6547), 
        .C2(n6574), .ZN(U3193) );
  AOI22_X1 U7469 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6609), .ZN(n6546) );
  OAI21_X1 U7470 ( .B1(n6547), .B2(n6579), .A(n6546), .ZN(U3194) );
  AOI22_X1 U7471 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6609), .ZN(n6548) );
  OAI21_X1 U7472 ( .B1(n6549), .B2(n6579), .A(n6548), .ZN(U3195) );
  AOI22_X1 U7473 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6609), .ZN(n6550) );
  OAI21_X1 U7474 ( .B1(n6552), .B2(n6574), .A(n6550), .ZN(U3196) );
  AOI22_X1 U7475 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6609), .ZN(n6551) );
  OAI21_X1 U7476 ( .B1(n6552), .B2(n6579), .A(n6551), .ZN(U3197) );
  AOI22_X1 U7477 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6609), .ZN(n6553) );
  OAI21_X1 U7478 ( .B1(n6554), .B2(n6579), .A(n6553), .ZN(U3198) );
  AOI22_X1 U7479 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6609), .ZN(n6555) );
  OAI21_X1 U7480 ( .B1(n6667), .B2(n6574), .A(n6555), .ZN(U3199) );
  AOI22_X1 U7481 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6609), .ZN(n6556) );
  OAI21_X1 U7482 ( .B1(n6667), .B2(n6579), .A(n6556), .ZN(U3200) );
  INV_X1 U7483 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6722) );
  AOI22_X1 U7484 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6609), .ZN(n6557) );
  OAI21_X1 U7485 ( .B1(n6722), .B2(n6574), .A(n6557), .ZN(U3201) );
  AOI22_X1 U7486 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6609), .ZN(n6558) );
  OAI21_X1 U7487 ( .B1(n6560), .B2(n6574), .A(n6558), .ZN(U3202) );
  INV_X1 U7488 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6559) );
  OAI222_X1 U7489 ( .A1(n6579), .A2(n6560), .B1(n6559), .B2(n6620), .C1(n6562), 
        .C2(n6574), .ZN(U3203) );
  AOI22_X1 U7490 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6609), .ZN(n6561) );
  OAI21_X1 U7491 ( .B1(n6562), .B2(n6579), .A(n6561), .ZN(U3204) );
  AOI22_X1 U7492 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6609), .ZN(n6563) );
  OAI21_X1 U7493 ( .B1(n6565), .B2(n6574), .A(n6563), .ZN(U3205) );
  AOI22_X1 U7494 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6609), .ZN(n6564) );
  OAI21_X1 U7495 ( .B1(n6565), .B2(n6579), .A(n6564), .ZN(U3206) );
  AOI22_X1 U7496 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6609), .ZN(n6566) );
  OAI21_X1 U7497 ( .B1(n6688), .B2(n6579), .A(n6566), .ZN(U3207) );
  INV_X1 U7498 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6672) );
  AOI22_X1 U7499 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6609), .ZN(n6567) );
  OAI21_X1 U7500 ( .B1(n6672), .B2(n6579), .A(n6567), .ZN(U3208) );
  AOI22_X1 U7501 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6609), .ZN(n6568) );
  OAI21_X1 U7502 ( .B1(n6569), .B2(n6579), .A(n6568), .ZN(U3209) );
  INV_X1 U7503 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6571) );
  INV_X1 U7504 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6658) );
  OAI222_X1 U7505 ( .A1(n6579), .A2(n6571), .B1(n6658), .B2(n6620), .C1(n6570), 
        .C2(n6574), .ZN(U3210) );
  INV_X1 U7506 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6576) );
  AOI22_X1 U7507 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6572), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6609), .ZN(n6573) );
  OAI21_X1 U7508 ( .B1(n6576), .B2(n6574), .A(n6573), .ZN(U3211) );
  AOI22_X1 U7509 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6609), .ZN(n6575) );
  OAI21_X1 U7510 ( .B1(n6576), .B2(n6579), .A(n6575), .ZN(U3212) );
  AOI22_X1 U7511 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6609), .ZN(n6578) );
  OAI21_X1 U7512 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(U3213) );
  MUX2_X1 U7513 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6620), .Z(U3445) );
  MUX2_X1 U7514 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6620), .Z(U3446) );
  MUX2_X1 U7515 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6620), .Z(U3447) );
  MUX2_X1 U7516 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6620), .Z(U3448) );
  INV_X1 U7517 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6583) );
  INV_X1 U7518 ( .A(n6584), .ZN(n6581) );
  AOI21_X1 U7519 ( .B1(n6583), .B2(n6582), .A(n6581), .ZN(U3451) );
  OAI21_X1 U7520 ( .B1(n6586), .B2(n6585), .A(n6584), .ZN(U3452) );
  INV_X1 U7521 ( .A(n6587), .ZN(n6589) );
  OAI211_X1 U7522 ( .C1(n6591), .C2(n6590), .A(n6589), .B(n6588), .ZN(U3453)
         );
  INV_X1 U7523 ( .A(n6592), .ZN(n6597) );
  INV_X1 U7524 ( .A(n6593), .ZN(n6596) );
  OAI22_X1 U7525 ( .A1(n6597), .A2(n6596), .B1(n6595), .B2(n6594), .ZN(n6599)
         );
  MUX2_X1 U7526 ( .A(n6599), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6598), 
        .Z(U3456) );
  AOI21_X1 U7527 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7528 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6601), .B2(n6600), .ZN(n6603) );
  INV_X1 U7529 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7530 ( .A1(n6604), .A2(n6603), .B1(n6602), .B2(n6606), .ZN(U3468)
         );
  INV_X1 U7531 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6607) );
  NOR2_X1 U7532 ( .A1(n6606), .A2(REIP_REG_1__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U7533 ( .A1(n6607), .A2(n6606), .B1(n4405), .B2(n6605), .ZN(U3469)
         );
  NAND2_X1 U7534 ( .A1(n6609), .A2(W_R_N_REG_SCAN_IN), .ZN(n6608) );
  OAI21_X1 U7535 ( .B1(n6609), .B2(READREQUEST_REG_SCAN_IN), .A(n6608), .ZN(
        U3470) );
  AOI211_X1 U7536 ( .C1(n6094), .C2(n6612), .A(n6611), .B(n6610), .ZN(n6619)
         );
  OAI211_X1 U7537 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6614), .A(n6613), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6616) );
  AOI21_X1 U7538 ( .B1(n6616), .B2(STATE2_REG_0__SCAN_IN), .A(n6615), .ZN(
        n6618) );
  NAND2_X1 U7539 ( .A1(n6619), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6617) );
  OAI21_X1 U7540 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(U3472) );
  MUX2_X1 U7541 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6620), .Z(U3473) );
  AOI222_X1 U7542 ( .A1(n6625), .A2(EBX_REG_9__SCAN_IN), .B1(n6624), .B2(n6623), .C1(n6622), .C2(n6621), .ZN(n6778) );
  AOI22_X1 U7543 ( .A1(n3930), .A2(keyinput0), .B1(keyinput11), .B2(n5631), 
        .ZN(n6626) );
  OAI221_X1 U7544 ( .B1(n3930), .B2(keyinput0), .C1(n5631), .C2(keyinput11), 
        .A(n6626), .ZN(n6638) );
  INV_X1 U7545 ( .A(keyinput12), .ZN(n6629) );
  AOI22_X1 U7546 ( .A1(n6629), .A2(DATAO_REG_19__SCAN_IN), .B1(keyinput23), 
        .B2(n6628), .ZN(n6627) );
  OAI221_X1 U7547 ( .B1(n6629), .B2(DATAO_REG_19__SCAN_IN), .C1(n6628), .C2(
        keyinput23), .A(n6627), .ZN(n6637) );
  INV_X1 U7548 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6632) );
  INV_X1 U7549 ( .A(keyinput55), .ZN(n6631) );
  AOI22_X1 U7550 ( .A1(n6632), .A2(keyinput57), .B1(ADDRESS_REG_9__SCAN_IN), 
        .B2(n6631), .ZN(n6630) );
  OAI221_X1 U7551 ( .B1(n6632), .B2(keyinput57), .C1(n6631), .C2(
        ADDRESS_REG_9__SCAN_IN), .A(n6630), .ZN(n6636) );
  XNOR2_X1 U7552 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .B(keyinput37), .ZN(n6634)
         );
  XNOR2_X1 U7553 ( .A(keyinput59), .B(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U7554 ( .A1(n6634), .A2(n6633), .ZN(n6635) );
  NOR4_X1 U7555 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6776)
         );
  INV_X1 U7556 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6641) );
  INV_X1 U7557 ( .A(keyinput48), .ZN(n6640) );
  AOI22_X1 U7558 ( .A1(n6641), .A2(keyinput6), .B1(DATAO_REG_0__SCAN_IN), .B2(
        n6640), .ZN(n6639) );
  OAI221_X1 U7559 ( .B1(n6641), .B2(keyinput6), .C1(n6640), .C2(
        DATAO_REG_0__SCAN_IN), .A(n6639), .ZN(n6652) );
  INV_X1 U7560 ( .A(DATAI_20_), .ZN(n6643) );
  AOI22_X1 U7561 ( .A1(n6643), .A2(keyinput22), .B1(n3664), .B2(keyinput19), 
        .ZN(n6642) );
  OAI221_X1 U7562 ( .B1(n6643), .B2(keyinput22), .C1(n3664), .C2(keyinput19), 
        .A(n6642), .ZN(n6651) );
  INV_X1 U7563 ( .A(keyinput13), .ZN(n6645) );
  AOI22_X1 U7564 ( .A1(n4700), .A2(keyinput40), .B1(DATAWIDTH_REG_23__SCAN_IN), 
        .B2(n6645), .ZN(n6644) );
  OAI221_X1 U7565 ( .B1(n4700), .B2(keyinput40), .C1(n6645), .C2(
        DATAWIDTH_REG_23__SCAN_IN), .A(n6644), .ZN(n6650) );
  INV_X1 U7566 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U7567 ( .A1(n6648), .A2(keyinput61), .B1(n6647), .B2(keyinput14), 
        .ZN(n6646) );
  OAI221_X1 U7568 ( .B1(n6648), .B2(keyinput61), .C1(n6647), .C2(keyinput14), 
        .A(n6646), .ZN(n6649) );
  NOR4_X1 U7569 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6775)
         );
  INV_X1 U7570 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7571 ( .A1(n6655), .A2(keyinput30), .B1(keyinput60), .B2(n6654), 
        .ZN(n6653) );
  OAI221_X1 U7572 ( .B1(n6655), .B2(keyinput30), .C1(n6654), .C2(keyinput60), 
        .A(n6653), .ZN(n6746) );
  AOI22_X1 U7573 ( .A1(n4660), .A2(keyinput32), .B1(keyinput38), .B2(n4195), 
        .ZN(n6656) );
  OAI221_X1 U7574 ( .B1(n4660), .B2(keyinput32), .C1(n4195), .C2(keyinput38), 
        .A(n6656), .ZN(n6745) );
  OAI22_X1 U7575 ( .A1(keyinput36), .A2(n6659), .B1(n6658), .B2(keyinput2), 
        .ZN(n6657) );
  AOI221_X1 U7576 ( .B1(n6659), .B2(keyinput36), .C1(n6658), .C2(keyinput2), 
        .A(n6657), .ZN(n6679) );
  INV_X1 U7577 ( .A(keyinput1), .ZN(n6661) );
  OAI22_X1 U7578 ( .A1(n6662), .A2(keyinput42), .B1(n6661), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n6660) );
  AOI221_X1 U7579 ( .B1(n6662), .B2(keyinput42), .C1(ADDRESS_REG_4__SCAN_IN), 
        .C2(n6661), .A(n6660), .ZN(n6678) );
  INV_X1 U7580 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6665) );
  INV_X1 U7581 ( .A(keyinput45), .ZN(n6664) );
  AOI22_X1 U7582 ( .A1(n6665), .A2(keyinput49), .B1(LWORD_REG_3__SCAN_IN), 
        .B2(n6664), .ZN(n6663) );
  OAI221_X1 U7583 ( .B1(n6665), .B2(keyinput49), .C1(n6664), .C2(
        LWORD_REG_3__SCAN_IN), .A(n6663), .ZN(n6676) );
  INV_X1 U7584 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7585 ( .A1(n6668), .A2(keyinput28), .B1(keyinput43), .B2(n6667), 
        .ZN(n6666) );
  OAI221_X1 U7586 ( .B1(n6668), .B2(keyinput28), .C1(n6667), .C2(keyinput43), 
        .A(n6666), .ZN(n6675) );
  AOI22_X1 U7587 ( .A1(n6121), .A2(keyinput29), .B1(n3407), .B2(keyinput10), 
        .ZN(n6669) );
  OAI221_X1 U7588 ( .B1(n6121), .B2(keyinput29), .C1(n3407), .C2(keyinput10), 
        .A(n6669), .ZN(n6674) );
  INV_X1 U7589 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7590 ( .A1(n6672), .A2(keyinput44), .B1(n6671), .B2(keyinput15), 
        .ZN(n6670) );
  OAI221_X1 U7591 ( .B1(n6672), .B2(keyinput44), .C1(n6671), .C2(keyinput15), 
        .A(n6670), .ZN(n6673) );
  NOR4_X1 U7592 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6677)
         );
  NAND3_X1 U7593 ( .A1(n6679), .A2(n6678), .A3(n6677), .ZN(n6744) );
  INV_X1 U7594 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6682) );
  INV_X1 U7595 ( .A(keyinput47), .ZN(n6681) );
  AOI22_X1 U7596 ( .A1(n6682), .A2(keyinput26), .B1(DATAWIDTH_REG_13__SCAN_IN), 
        .B2(n6681), .ZN(n6680) );
  OAI221_X1 U7597 ( .B1(n6682), .B2(keyinput26), .C1(n6681), .C2(
        DATAWIDTH_REG_13__SCAN_IN), .A(n6680), .ZN(n6695) );
  INV_X1 U7598 ( .A(keyinput53), .ZN(n6684) );
  AOI22_X1 U7599 ( .A1(n6685), .A2(keyinput34), .B1(UWORD_REG_5__SCAN_IN), 
        .B2(n6684), .ZN(n6683) );
  OAI221_X1 U7600 ( .B1(n6685), .B2(keyinput34), .C1(n6684), .C2(
        UWORD_REG_5__SCAN_IN), .A(n6683), .ZN(n6694) );
  AOI22_X1 U7601 ( .A1(n6688), .A2(keyinput24), .B1(n6687), .B2(keyinput50), 
        .ZN(n6686) );
  OAI221_X1 U7602 ( .B1(n6688), .B2(keyinput24), .C1(n6687), .C2(keyinput50), 
        .A(n6686), .ZN(n6693) );
  INV_X1 U7603 ( .A(DATAI_31_), .ZN(n6691) );
  INV_X1 U7604 ( .A(keyinput46), .ZN(n6690) );
  AOI22_X1 U7605 ( .A1(n6691), .A2(keyinput35), .B1(ADDRESS_REG_0__SCAN_IN), 
        .B2(n6690), .ZN(n6689) );
  OAI221_X1 U7606 ( .B1(n6691), .B2(keyinput35), .C1(n6690), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n6689), .ZN(n6692) );
  NOR4_X1 U7607 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6742)
         );
  INV_X1 U7608 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6698) );
  INV_X1 U7609 ( .A(keyinput20), .ZN(n6697) );
  AOI22_X1 U7610 ( .A1(n6698), .A2(keyinput31), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n6697), .ZN(n6696) );
  OAI221_X1 U7611 ( .B1(n6698), .B2(keyinput31), .C1(n6697), .C2(
        DATAO_REG_31__SCAN_IN), .A(n6696), .ZN(n6711) );
  AOI22_X1 U7612 ( .A1(n6701), .A2(keyinput41), .B1(n6700), .B2(keyinput39), 
        .ZN(n6699) );
  OAI221_X1 U7613 ( .B1(n6701), .B2(keyinput41), .C1(n6700), .C2(keyinput39), 
        .A(n6699), .ZN(n6710) );
  INV_X1 U7614 ( .A(keyinput17), .ZN(n6703) );
  AOI22_X1 U7615 ( .A1(n6704), .A2(keyinput16), .B1(ADDRESS_REG_6__SCAN_IN), 
        .B2(n6703), .ZN(n6702) );
  OAI221_X1 U7616 ( .B1(n6704), .B2(keyinput16), .C1(n6703), .C2(
        ADDRESS_REG_6__SCAN_IN), .A(n6702), .ZN(n6709) );
  AOI22_X1 U7617 ( .A1(n6707), .A2(keyinput51), .B1(keyinput4), .B2(n6706), 
        .ZN(n6705) );
  OAI221_X1 U7618 ( .B1(n6707), .B2(keyinput51), .C1(n6706), .C2(keyinput4), 
        .A(n6705), .ZN(n6708) );
  NOR4_X1 U7619 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n6741)
         );
  INV_X1 U7620 ( .A(keyinput54), .ZN(n6713) );
  AOI22_X1 U7621 ( .A1(n4703), .A2(keyinput58), .B1(DATAWIDTH_REG_24__SCAN_IN), 
        .B2(n6713), .ZN(n6712) );
  OAI221_X1 U7622 ( .B1(n4703), .B2(keyinput58), .C1(n6713), .C2(
        DATAWIDTH_REG_24__SCAN_IN), .A(n6712), .ZN(n6726) );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U7624 ( .A1(n6716), .A2(keyinput3), .B1(n6715), .B2(keyinput5), 
        .ZN(n6714) );
  OAI221_X1 U7625 ( .B1(n6716), .B2(keyinput3), .C1(n6715), .C2(keyinput5), 
        .A(n6714), .ZN(n6725) );
  INV_X1 U7626 ( .A(keyinput21), .ZN(n6719) );
  INV_X1 U7627 ( .A(keyinput18), .ZN(n6718) );
  AOI22_X1 U7628 ( .A1(n6719), .A2(ADDRESS_REG_19__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n6718), .ZN(n6717) );
  OAI221_X1 U7629 ( .B1(n6719), .B2(ADDRESS_REG_19__SCAN_IN), .C1(n6718), .C2(
        DATAO_REG_1__SCAN_IN), .A(n6717), .ZN(n6724) );
  INV_X1 U7630 ( .A(keyinput62), .ZN(n6721) );
  AOI22_X1 U7631 ( .A1(n6722), .A2(keyinput7), .B1(LWORD_REG_5__SCAN_IN), .B2(
        n6721), .ZN(n6720) );
  OAI221_X1 U7632 ( .B1(n6722), .B2(keyinput7), .C1(n6721), .C2(
        LWORD_REG_5__SCAN_IN), .A(n6720), .ZN(n6723) );
  NOR4_X1 U7633 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6740)
         );
  AOI22_X1 U7634 ( .A1(n3802), .A2(keyinput9), .B1(n3423), .B2(keyinput56), 
        .ZN(n6727) );
  OAI221_X1 U7635 ( .B1(n3802), .B2(keyinput9), .C1(n3423), .C2(keyinput56), 
        .A(n6727), .ZN(n6738) );
  AOI22_X1 U7636 ( .A1(n4666), .A2(keyinput52), .B1(keyinput25), .B2(n6729), 
        .ZN(n6728) );
  OAI221_X1 U7637 ( .B1(n4666), .B2(keyinput52), .C1(n6729), .C2(keyinput25), 
        .A(n6728), .ZN(n6737) );
  INV_X1 U7638 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6731) );
  INV_X1 U7639 ( .A(keyinput63), .ZN(n6758) );
  AOI22_X1 U7640 ( .A1(n6731), .A2(keyinput33), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n6758), .ZN(n6730) );
  OAI221_X1 U7641 ( .B1(n6731), .B2(keyinput33), .C1(n6758), .C2(
        DATAO_REG_22__SCAN_IN), .A(n6730), .ZN(n6736) );
  INV_X1 U7642 ( .A(keyinput27), .ZN(n6732) );
  XOR2_X1 U7643 ( .A(DATAO_REG_5__SCAN_IN), .B(n6732), .Z(n6734) );
  XNOR2_X1 U7644 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput8), .ZN(
        n6733) );
  NAND2_X1 U7645 ( .A1(n6734), .A2(n6733), .ZN(n6735) );
  NOR4_X1 U7646 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .ZN(n6739)
         );
  NAND4_X1 U7647 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6743)
         );
  NOR4_X1 U7648 ( .A1(n6746), .A2(n6745), .A3(n6744), .A4(n6743), .ZN(n6774)
         );
  NAND2_X1 U7649 ( .A1(keyinput26), .A2(keyinput47), .ZN(n6752) );
  NOR2_X1 U7650 ( .A1(keyinput50), .A2(keyinput46), .ZN(n6750) );
  NAND2_X1 U7651 ( .A1(keyinput20), .A2(keyinput41), .ZN(n6748) );
  NAND4_X1 U7652 ( .A1(keyinput17), .A2(keyinput16), .A3(keyinput51), .A4(
        keyinput4), .ZN(n6747) );
  NOR4_X1 U7653 ( .A1(keyinput31), .A2(keyinput39), .A3(n6748), .A4(n6747), 
        .ZN(n6749) );
  NAND4_X1 U7654 ( .A1(keyinput24), .A2(keyinput35), .A3(n6750), .A4(n6749), 
        .ZN(n6751) );
  NOR4_X1 U7655 ( .A1(keyinput34), .A2(keyinput53), .A3(n6752), .A4(n6751), 
        .ZN(n6772) );
  INV_X1 U7656 ( .A(keyinput6), .ZN(n6753) );
  NOR4_X1 U7657 ( .A1(keyinput59), .A2(keyinput30), .A3(keyinput23), .A4(n6753), .ZN(n6771) );
  NAND4_X1 U7658 ( .A1(keyinput57), .A2(keyinput60), .A3(keyinput0), .A4(
        keyinput48), .ZN(n6756) );
  NAND4_X1 U7659 ( .A1(keyinput11), .A2(keyinput55), .A3(keyinput15), .A4(
        keyinput10), .ZN(n6755) );
  NAND4_X1 U7660 ( .A1(keyinput2), .A2(keyinput14), .A3(keyinput22), .A4(
        keyinput19), .ZN(n6754) );
  NOR3_X1 U7661 ( .A1(n6756), .A2(n6755), .A3(n6754), .ZN(n6770) );
  NOR2_X1 U7662 ( .A1(keyinput21), .A2(keyinput62), .ZN(n6757) );
  NAND3_X1 U7663 ( .A1(keyinput18), .A2(keyinput7), .A3(n6757), .ZN(n6768) );
  NAND4_X1 U7664 ( .A1(keyinput33), .A2(keyinput52), .A3(keyinput25), .A4(
        n6758), .ZN(n6767) );
  NOR3_X1 U7665 ( .A1(keyinput54), .A2(keyinput3), .A3(keyinput5), .ZN(n6760)
         );
  NOR3_X1 U7666 ( .A1(keyinput56), .A2(keyinput27), .A3(keyinput8), .ZN(n6759)
         );
  NAND4_X1 U7667 ( .A1(keyinput58), .A2(n6760), .A3(keyinput9), .A4(n6759), 
        .ZN(n6766) );
  NOR4_X1 U7668 ( .A1(keyinput13), .A2(keyinput1), .A3(keyinput29), .A4(
        keyinput37), .ZN(n6764) );
  NOR4_X1 U7669 ( .A1(keyinput45), .A2(keyinput49), .A3(keyinput61), .A4(
        keyinput12), .ZN(n6763) );
  NOR4_X1 U7670 ( .A1(keyinput28), .A2(keyinput36), .A3(keyinput40), .A4(
        keyinput44), .ZN(n6762) );
  NOR4_X1 U7671 ( .A1(keyinput32), .A2(keyinput42), .A3(keyinput43), .A4(
        keyinput38), .ZN(n6761) );
  NAND4_X1 U7672 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6765)
         );
  NOR4_X1 U7673 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6769)
         );
  NAND4_X1 U7674 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6773)
         );
  NAND4_X1 U7675 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6777)
         );
  XOR2_X1 U7676 ( .A(n6778), .B(n6777), .Z(U2850) );
  AND2_X2 U4117 ( .A1(n4377), .A2(n4463), .ZN(n3440) );
  MUX2_X1 U3610 ( .A(n3885), .B(n4404), .S(n4403), .Z(n4420) );
  CLKBUF_X1 U3575 ( .A(n3348), .Z(n3940) );
  CLKBUF_X1 U3648 ( .A(n3373), .Z(n2987) );
  CLKBUF_X1 U3770 ( .A(n5321), .Z(n5443) );
  CLKBUF_X1 U4271 ( .A(n3346), .Z(n3941) );
endmodule

