

module b15_C_SARLock_k_128_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009;

  INV_X1 U3540 ( .A(n3928), .ZN(n5418) );
  CLKBUF_X1 U3542 ( .A(n5397), .Z(n4019) );
  CLKBUF_X2 U3543 ( .A(n3112), .Z(n3093) );
  CLKBUF_X2 U3544 ( .A(n3390), .Z(n5398) );
  CLKBUF_X1 U3545 ( .A(n3345), .Z(n4460) );
  AND2_X2 U3547 ( .A1(n3217), .A2(n4606), .ZN(n3097) );
  AND2_X1 U3548 ( .A1(n3217), .A2(n3218), .ZN(n3446) );
  AND2_X1 U3549 ( .A1(n4606), .A2(n4634), .ZN(n3390) );
  AOI22_X1 U3550 ( .A1(n6849), .A2(keyinput110), .B1(n6848), .B2(keyinput13), 
        .ZN(n6847) );
  AND2_X1 U3551 ( .A1(n3193), .A2(n3377), .ZN(n3388) );
  OAI221_X1 U3552 ( .B1(n6849), .B2(keyinput110), .C1(n6848), .C2(keyinput13), 
        .A(n6847), .ZN(n6854) );
  INV_X1 U3553 ( .A(n6100), .ZN(n6091) );
  INV_X1 U3554 ( .A(n6081), .ZN(n6146) );
  AND2_X1 U3555 ( .A1(n4633), .A2(n4606), .ZN(n3116) );
  OR2_X1 U3556 ( .A1(n5892), .A2(n6360), .ZN(n3091) );
  AND2_X1 U3557 ( .A1(n4428), .A2(n3256), .ZN(n3092) );
  OAI21_X2 U3558 ( .B1(n5434), .B2(n5376), .A(n5375), .ZN(n5377) );
  BUF_X1 U3559 ( .A(n3121), .Z(n3094) );
  BUF_X4 U3560 ( .A(n3121), .Z(n3095) );
  BUF_X2 U3561 ( .A(n3809), .Z(n3121) );
  NAND2_X2 U3562 ( .A1(n4373), .A2(n4355), .ZN(n6137) );
  AND2_X1 U3563 ( .A1(n3217), .A2(n4606), .ZN(n3096) );
  AND2_X2 U3564 ( .A1(n3217), .A2(n4606), .ZN(n4133) );
  NOR2_X1 U3565 ( .A1(n5499), .A2(n5500), .ZN(n4151) );
  BUF_X1 U3566 ( .A(n4461), .Z(n3110) );
  AND2_X1 U3567 ( .A1(n3486), .A2(n3485), .ZN(n4566) );
  INV_X2 U3569 ( .A(n3489), .ZN(n3341) );
  AND4_X1 U3570 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3297)
         );
  AND4_X1 U3571 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  CLKBUF_X2 U3572 ( .A(n3317), .Z(n5395) );
  CLKBUF_X2 U3573 ( .A(n3318), .Z(n5396) );
  BUF_X2 U3574 ( .A(n3446), .Z(n4094) );
  CLKBUF_X1 U3575 ( .A(n3116), .Z(n3118) );
  CLKBUF_X1 U3576 ( .A(n3116), .Z(n3119) );
  AND2_X2 U3577 ( .A1(n3210), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5459)
         );
  OAI22_X1 U3578 ( .A1(n5744), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5755), .B2(n4168), .ZN(n4169) );
  NOR2_X1 U3579 ( .A1(n3635), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5433)
         );
  AND2_X1 U3580 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  AOI211_X1 U3581 ( .C1(n6298), .C2(n5716), .A(n5715), .B(n5714), .ZN(n5717)
         );
  OR2_X1 U3582 ( .A1(n5619), .A2(n6325), .ZN(n4160) );
  INV_X1 U3583 ( .A(n3170), .ZN(n5699) );
  AOI21_X1 U3584 ( .B1(n5771), .B2(n3171), .A(n3174), .ZN(n3170) );
  XNOR2_X1 U3585 ( .A(n3200), .B(n3199), .ZN(n5673) );
  NOR2_X1 U3586 ( .A1(n4151), .A2(n3129), .ZN(n5707) );
  NAND2_X1 U3587 ( .A1(n5509), .A2(n5510), .ZN(n5499) );
  CLKBUF_X1 U3588 ( .A(n5509), .Z(n5525) );
  NOR2_X1 U3589 ( .A1(n5970), .A2(n5593), .ZN(n6178) );
  CLKBUF_X1 U3590 ( .A(n5535), .Z(n5536) );
  NOR2_X1 U3591 ( .A1(n5626), .A2(n5625), .ZN(n5535) );
  CLKBUF_X1 U3592 ( .A(n3621), .Z(n3102) );
  AND2_X1 U3593 ( .A1(n5591), .A2(n5590), .ZN(n5970) );
  NOR2_X1 U3594 ( .A1(n5562), .A2(n3968), .ZN(n5642) );
  NAND2_X2 U3595 ( .A1(n5271), .A2(n3842), .ZN(n5589) );
  NAND2_X1 U3596 ( .A1(n3830), .A2(n3125), .ZN(n5273) );
  AND2_X1 U3597 ( .A1(n5188), .A2(n3842), .ZN(n3828) );
  NAND2_X1 U3598 ( .A1(n6065), .A2(n3201), .ZN(n3842) );
  OAI21_X1 U3599 ( .B1(n5342), .B2(n3169), .A(n3623), .ZN(n3168) );
  INV_X1 U3600 ( .A(n3622), .ZN(n3169) );
  NOR2_X1 U3601 ( .A1(n4781), .A2(n4997), .ZN(n4935) );
  NAND2_X1 U3602 ( .A1(n3186), .A2(n3185), .ZN(n4781) );
  OAI21_X1 U3603 ( .B1(n3610), .B2(n3593), .A(n3592), .ZN(n3594) );
  INV_X1 U3604 ( .A(n4442), .ZN(n3186) );
  OR2_X1 U3605 ( .A1(n3610), .A2(n3609), .ZN(n3619) );
  AND2_X1 U3606 ( .A1(n4809), .A2(n3738), .ZN(n3185) );
  XNOR2_X1 U3607 ( .A(n3600), .B(n3599), .ZN(n3743) );
  NOR2_X1 U3608 ( .A1(n4450), .A2(n4559), .ZN(n4443) );
  AND2_X1 U3609 ( .A1(n3188), .A2(n3187), .ZN(n4559) );
  OR2_X1 U3610 ( .A1(n3563), .A2(n3562), .ZN(n3140) );
  NAND2_X1 U3611 ( .A1(n4386), .A2(n3523), .ZN(n6306) );
  NOR2_X1 U3612 ( .A1(n3126), .A2(n4267), .ZN(n5645) );
  CLKBUF_X1 U3613 ( .A(n4462), .Z(n5906) );
  OR2_X1 U3614 ( .A1(n5608), .A2(n5597), .ZN(n5897) );
  XNOR2_X1 U3615 ( .A(n3513), .B(n3512), .ZN(n4462) );
  NOR2_X1 U3616 ( .A1(n5078), .A2(n3342), .ZN(n4373) );
  OR2_X1 U3617 ( .A1(n5671), .A2(n5610), .ZN(n5608) );
  MUX2_X1 U3618 ( .A(n4436), .B(n4344), .S(n4434), .Z(n4438) );
  INV_X1 U3619 ( .A(n4566), .ZN(n3098) );
  NAND2_X1 U3620 ( .A1(n6092), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U3621 ( .A1(n6186), .A2(n4681), .ZN(n5951) );
  NAND2_X1 U3622 ( .A1(n3418), .A2(n3417), .ZN(n3159) );
  NOR2_X1 U3623 ( .A1(n3145), .A2(n3134), .ZN(n5669) );
  AND2_X1 U3624 ( .A1(n5047), .A2(n4937), .ZN(n6072) );
  OR2_X1 U3625 ( .A1(n3388), .A2(n3387), .ZN(n3389) );
  NOR2_X1 U3626 ( .A1(n5049), .A2(n5048), .ZN(n5047) );
  AND2_X2 U3627 ( .A1(n4622), .A2(n6543), .ZN(n4419) );
  OR2_X2 U3628 ( .A1(n3686), .A2(n3685), .ZN(n4622) );
  NOR2_X1 U3629 ( .A1(n3309), .A2(n3308), .ZN(n3336) );
  OAI211_X1 U3630 ( .C1(n3435), .C2(n3434), .A(n3433), .B(n3453), .ZN(n3510)
         );
  OR2_X1 U3631 ( .A1(n3598), .A2(n4540), .ZN(n3460) );
  CLKBUF_X1 U3632 ( .A(n3361), .Z(n3362) );
  INV_X1 U3633 ( .A(n3683), .ZN(n3667) );
  OR2_X1 U3634 ( .A1(n4601), .A2(n3344), .ZN(n4282) );
  NOR2_X1 U3635 ( .A1(n4673), .A2(n3130), .ZN(n3668) );
  NOR2_X2 U3636 ( .A1(n3474), .A2(n6786), .ZN(n3676) );
  AND2_X2 U3637 ( .A1(n3474), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U3638 ( .A1(n3324), .A2(n3299), .ZN(n3373) );
  NAND2_X1 U3639 ( .A1(n3342), .A2(n3489), .ZN(n5077) );
  NOR2_X1 U3640 ( .A1(n3342), .A2(n3489), .ZN(n3490) );
  OR2_X2 U3641 ( .A1(n3255), .A2(n3254), .ZN(n4678) );
  AND4_X1 U3643 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3245)
         );
  AND4_X1 U3644 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3234)
         );
  AND4_X1 U3645 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3323)
         );
  AND4_X1 U3646 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3225)
         );
  AND4_X1 U3647 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3274)
         );
  NOR2_X1 U3648 ( .A1(n6325), .A2(n4483), .ZN(n6475) );
  AND4_X1 U3649 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3235)
         );
  AND4_X1 U3650 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3244)
         );
  AND4_X1 U3651 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3224)
         );
  AND4_X1 U3652 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3276)
         );
  AND4_X1 U3653 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3275)
         );
  AND4_X1 U3654 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3296)
         );
  AND4_X1 U3655 ( .A1(n3289), .A2(n3288), .A3(n3287), .A4(n3286), .ZN(n3295)
         );
  AND4_X1 U3656 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3294)
         );
  NOR2_X1 U3657 ( .A1(n6325), .A2(n4474), .ZN(n6495) );
  NOR2_X1 U3658 ( .A1(n6325), .A2(n4479), .ZN(n6489) );
  BUF_X2 U3659 ( .A(n3312), .Z(n5404) );
  CLKBUF_X1 U3660 ( .A(n3311), .Z(n4132) );
  BUF_X2 U3661 ( .A(n3444), .Z(n4135) );
  AND2_X2 U3662 ( .A1(n5459), .A2(n3219), .ZN(n5397) );
  AND2_X2 U3663 ( .A1(n3217), .A2(n4645), .ZN(n4134) );
  AND2_X2 U3664 ( .A1(n3217), .A2(n4645), .ZN(n3111) );
  AND2_X1 U3665 ( .A1(n3211), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3218)
         );
  AND2_X1 U3666 ( .A1(n3216), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3219)
         );
  AND2_X2 U3667 ( .A1(n4645), .A2(n4634), .ZN(n3445) );
  AND2_X2 U3668 ( .A1(n3209), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3217)
         );
  INV_X1 U3669 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3209) );
  AND2_X2 U3670 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4634) );
  NAND2_X2 U3671 ( .A1(n3468), .A2(n3099), .ZN(n3549) );
  AND2_X2 U3672 ( .A1(n3495), .A2(n3098), .ZN(n3099) );
  NAND2_X1 U3673 ( .A1(n4428), .A2(n3256), .ZN(n3100) );
  AND2_X1 U3674 ( .A1(n5760), .A2(n5761), .ZN(n3101) );
  AND2_X1 U3675 ( .A1(n5698), .A2(n3203), .ZN(n3635) );
  AOI21_X1 U3676 ( .B1(n3743), .B2(n3901), .A(n3742), .ZN(n4997) );
  AND2_X1 U3677 ( .A1(n3590), .A2(n3140), .ZN(n3724) );
  NAND2_X1 U3678 ( .A1(n3436), .A2(n3439), .ZN(n3103) );
  CLKBUF_X1 U3679 ( .A(n4596), .Z(n3104) );
  CLKBUF_X1 U3680 ( .A(n5199), .Z(n3105) );
  CLKBUF_X1 U3681 ( .A(n4557), .Z(n3106) );
  NAND2_X1 U3682 ( .A1(n3436), .A2(n3439), .ZN(n3437) );
  XNOR2_X1 U3683 ( .A(n3526), .B(n6694), .ZN(n4557) );
  OR2_X1 U3684 ( .A1(n5432), .A2(n6370), .ZN(n3154) );
  CLKBUF_X1 U3685 ( .A(n4443), .Z(n3107) );
  OR2_X1 U3686 ( .A1(n5822), .A2(n6284), .ZN(n3108) );
  NAND2_X1 U3687 ( .A1(n5717), .A2(n3108), .ZN(U2959) );
  NOR2_X1 U3688 ( .A1(n5562), .A2(n3109), .ZN(n5550) );
  OR2_X1 U3689 ( .A1(n3968), .A2(n3138), .ZN(n3109) );
  XNOR2_X1 U3690 ( .A(n3495), .B(n3494), .ZN(n4461) );
  OR2_X1 U3691 ( .A1(n3373), .A2(n4201), .ZN(n3361) );
  AND2_X1 U3692 ( .A1(n3217), .A2(n5459), .ZN(n3312) );
  NAND2_X1 U3693 ( .A1(n5372), .A2(n3633), .ZN(n5698) );
  OAI222_X1 U3694 ( .A1(n6148), .A2(n5713), .B1(n5622), .B2(n6170), .C1(n5815), 
        .C2(n6153), .ZN(U2832) );
  NAND2_X1 U3695 ( .A1(n3493), .A2(n3492), .ZN(n3526) );
  OAI21_X1 U3696 ( .B1(n4151), .B2(n4152), .A(n5465), .ZN(n5619) );
  OR2_X1 U3697 ( .A1(n3378), .A2(n4635), .ZN(n3473) );
  AND2_X1 U3698 ( .A1(n4633), .A2(n4645), .ZN(n3112) );
  AND2_X1 U3699 ( .A1(n4633), .A2(n4645), .ZN(n3424) );
  AND2_X4 U3700 ( .A1(n3218), .A2(n4634), .ZN(n3311) );
  BUF_X4 U3701 ( .A(n3445), .Z(n3114) );
  BUF_X8 U3702 ( .A(n5403), .Z(n3115) );
  AND2_X2 U3703 ( .A1(n4633), .A2(n3218), .ZN(n5403) );
  AND2_X1 U3704 ( .A1(n4633), .A2(n4606), .ZN(n3117) );
  CLKBUF_X1 U3705 ( .A(n3395), .Z(n3120) );
  AND2_X1 U3706 ( .A1(n4633), .A2(n4606), .ZN(n3395) );
  AND2_X1 U3707 ( .A1(n3219), .A2(n4645), .ZN(n3444) );
  OR2_X1 U3708 ( .A1(n5499), .A2(n3194), .ZN(n3200) );
  NOR2_X2 U3709 ( .A1(n5698), .A2(n5719), .ZN(n5709) );
  OAI21_X2 U3710 ( .B1(n3378), .B2(n6513), .A(n3360), .ZN(n3436) );
  AOI21_X2 U3711 ( .B1(n5765), .B2(n5766), .A(n4167), .ZN(n5760) );
  AOI21_X1 U3712 ( .B1(n3372), .B2(n4673), .A(n3375), .ZN(n4296) );
  NAND2_X4 U3713 ( .A1(n3245), .A2(n3244), .ZN(n3310) );
  OR2_X2 U3714 ( .A1(n5499), .A2(n3197), .ZN(n5465) );
  OAI21_X2 U3715 ( .B1(n5199), .B2(n5201), .A(n5200), .ZN(n5210) );
  INV_X4 U3716 ( .A(n3617), .ZN(n5892) );
  OAI21_X2 U3717 ( .B1(n5771), .B2(n3174), .A(n3172), .ZN(n5372) );
  BUF_X4 U3718 ( .A(n3809), .Z(n3122) );
  NAND2_X1 U3719 ( .A1(n3139), .A2(n5643), .ZN(n3138) );
  INV_X1 U3720 ( .A(n5638), .ZN(n3139) );
  INV_X1 U3721 ( .A(n3910), .ZN(n3192) );
  AND2_X1 U3722 ( .A1(n3827), .A2(n5188), .ZN(n3201) );
  NOR2_X2 U3723 ( .A1(n4460), .A2(n6455), .ZN(n3901) );
  NOR2_X1 U3724 ( .A1(n3152), .A2(n4280), .ZN(n3151) );
  INV_X1 U3725 ( .A(n4275), .ZN(n3152) );
  INV_X1 U3726 ( .A(n3516), .ZN(n3457) );
  INV_X1 U3727 ( .A(n4156), .ZN(n3384) );
  AND2_X2 U3728 ( .A1(n3342), .A2(n3341), .ZN(n4673) );
  NAND2_X1 U3729 ( .A1(n4419), .A2(n4624), .ZN(n6239) );
  NAND2_X1 U3730 ( .A1(n5647), .A2(n3151), .ZN(n5539) );
  OR2_X1 U3731 ( .A1(n3453), .A2(n3457), .ZN(n3502) );
  AND2_X1 U3732 ( .A1(n4657), .A2(n4656), .ZN(n4858) );
  AND2_X1 U3733 ( .A1(n4657), .A2(n4821), .ZN(n4690) );
  AND2_X1 U3734 ( .A1(n6186), .A2(n4682), .ZN(n6180) );
  AOI21_X1 U3735 ( .B1(n3384), .B2(n4962), .A(n3352), .ZN(n3355) );
  NAND2_X1 U3736 ( .A1(n3100), .A2(n3277), .ZN(n4188) );
  AND2_X1 U3737 ( .A1(n3347), .A2(n4678), .ZN(n3327) );
  OAI21_X1 U3738 ( .B1(n3666), .B2(n3664), .A(n3642), .ZN(n3672) );
  XNOR2_X1 U3739 ( .A(n4635), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3671)
         );
  OR2_X1 U3740 ( .A1(n3462), .A2(n6786), .ZN(n3609) );
  INV_X1 U3741 ( .A(n3345), .ZN(n3363) );
  NOR3_X1 U3742 ( .A1(n3192), .A2(n5578), .A3(n5563), .ZN(n3191) );
  NOR2_X1 U3743 ( .A1(n5454), .A2(n6786), .ZN(n4146) );
  NAND2_X1 U3744 ( .A1(n5647), .A2(n3149), .ZN(n3153) );
  NOR2_X1 U3745 ( .A1(n5540), .A2(n3150), .ZN(n3149) );
  INV_X1 U3746 ( .A(n3151), .ZN(n3150) );
  NAND2_X1 U3747 ( .A1(n5892), .A2(n3632), .ZN(n3633) );
  NAND2_X1 U3748 ( .A1(n5892), .A2(n3178), .ZN(n3175) );
  NOR2_X1 U3749 ( .A1(n5892), .A2(n3177), .ZN(n3176) );
  NOR2_X1 U3750 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3177)
         );
  INV_X1 U3751 ( .A(n3175), .ZN(n3174) );
  NOR2_X1 U3752 ( .A1(n3169), .A2(n3166), .ZN(n3165) );
  INV_X1 U3753 ( .A(n5275), .ZN(n3166) );
  NAND2_X1 U3754 ( .A1(n6072), .A2(n3141), .ZN(n3145) );
  NOR2_X1 U3755 ( .A1(n3142), .A2(n5216), .ZN(n3141) );
  INV_X1 U3756 ( .A(n3143), .ZN(n3142) );
  CLKBUF_X1 U3757 ( .A(n4201), .Z(n4226) );
  NOR2_X1 U3758 ( .A1(n3364), .A2(n3346), .ZN(n4427) );
  XNOR2_X1 U3759 ( .A(n3469), .B(n5004), .ZN(n4463) );
  NOR2_X1 U3760 ( .A1(n3688), .A2(n3690), .ZN(n4194) );
  AND2_X1 U3761 ( .A1(n3948), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3951)
         );
  INV_X1 U3762 ( .A(n4226), .ZN(n5652) );
  OR2_X1 U3763 ( .A1(n4112), .A2(n6688), .ZN(n4348) );
  OR2_X1 U3764 ( .A1(n4088), .A2(n4087), .ZN(n4108) );
  INV_X1 U3765 ( .A(n5589), .ZN(n3190) );
  AND2_X1 U3766 ( .A1(n3821), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3822)
         );
  NAND2_X1 U3767 ( .A1(n3828), .A2(n6065), .ZN(n3830) );
  AOI21_X1 U3768 ( .B1(n5210), .B2(n5211), .A(n5213), .ZN(n5277) );
  NAND2_X1 U3769 ( .A1(n3731), .A2(n3730), .ZN(n4809) );
  INV_X1 U3770 ( .A(n3729), .ZN(n3730) );
  NAND2_X1 U3771 ( .A1(n3692), .A2(n3824), .ZN(n4452) );
  NAND2_X1 U3772 ( .A1(n4387), .A2(n4388), .ZN(n4386) );
  AND2_X1 U3773 ( .A1(n5840), .A2(n4315), .ZN(n4322) );
  NOR2_X1 U3774 ( .A1(n3161), .A2(n3131), .ZN(n3160) );
  INV_X1 U3775 ( .A(n3127), .ZN(n3161) );
  NAND2_X1 U3776 ( .A1(n3162), .A2(n3127), .ZN(n5881) );
  OR2_X1 U3777 ( .A1(n5864), .A2(n4303), .ZN(n5347) );
  OR2_X1 U3778 ( .A1(n4756), .A2(n4755), .ZN(n4758) );
  AND2_X1 U3779 ( .A1(n3489), .A2(n4490), .ZN(n4382) );
  INV_X1 U3780 ( .A(n4302), .ZN(n4299) );
  INV_X1 U3781 ( .A(n3455), .ZN(n3456) );
  OAI21_X1 U3782 ( .B1(n3454), .B2(n6786), .A(n3502), .ZN(n3455) );
  CLKBUF_X1 U3783 ( .A(n4467), .Z(n4468) );
  INV_X1 U3784 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6513) );
  OR2_X1 U3785 ( .A1(n6449), .A2(n4957), .ZN(n5116) );
  OR2_X1 U3786 ( .A1(n4466), .A2(n5907), .ZN(n6398) );
  CLKBUF_X1 U3787 ( .A(n4463), .Z(n4464) );
  NOR2_X1 U3788 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4471), .ZN(n4689) );
  AND2_X1 U3789 ( .A1(n3110), .A2(n3098), .ZN(n4657) );
  INV_X2 U3790 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6455) );
  AND2_X1 U3791 ( .A1(n5429), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4370) );
  NAND2_X1 U3792 ( .A1(n6092), .A2(n4352), .ZN(n6100) );
  NAND2_X1 U3793 ( .A1(n4375), .A2(n4374), .ZN(n6125) );
  OAI21_X1 U3794 ( .B1(n4676), .B2(n4675), .A(n6543), .ZN(n4677) );
  AND2_X1 U3795 ( .A1(n5539), .A2(n4281), .ZN(n5916) );
  OR2_X1 U3796 ( .A1(n5875), .A2(n5862), .ZN(n5861) );
  INV_X1 U3797 ( .A(n6352), .ZN(n6377) );
  INV_X1 U3798 ( .A(n4468), .ZN(n5907) );
  CLKBUF_X1 U3799 ( .A(n4465), .Z(n4466) );
  INV_X1 U3800 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6532) );
  AND2_X1 U3801 ( .A1(n4858), .A2(n5115), .ZN(n4894) );
  AND2_X1 U3802 ( .A1(n3638), .A2(n3637), .ZN(n3649) );
  OR2_X1 U3803 ( .A1(n3584), .A2(n3583), .ZN(n3602) );
  OR2_X1 U3804 ( .A1(n3559), .A2(n3558), .ZN(n3567) );
  NAND2_X1 U3805 ( .A1(n3364), .A2(n3489), .ZN(n4201) );
  OR2_X1 U3806 ( .A1(n3538), .A2(n3537), .ZN(n3564) );
  OR2_X1 U3807 ( .A1(n3430), .A2(n3429), .ZN(n3612) );
  AND2_X1 U3808 ( .A1(n3324), .A2(n4678), .ZN(n3256) );
  OR2_X1 U3809 ( .A1(n3416), .A2(n3415), .ZN(n3515) );
  INV_X1 U3810 ( .A(n3346), .ZN(n3374) );
  OAI211_X1 U3811 ( .C1(n3329), .C2(n3328), .A(n3327), .B(n3326), .ZN(n3372)
         );
  AOI22_X1 U3812 ( .A1(n5403), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U3813 ( .A1(n3311), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U3814 ( .A1(n5397), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3228) );
  OR2_X1 U3815 ( .A1(n3484), .A2(n3483), .ZN(n3491) );
  NAND2_X1 U3816 ( .A1(n3310), .A2(n4490), .ZN(n3474) );
  AOI21_X1 U3817 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6532), .A(n3644), 
        .ZN(n3645) );
  NOR2_X1 U3818 ( .A1(n3643), .A2(n3671), .ZN(n3644) );
  NAND2_X1 U3819 ( .A1(n4152), .A2(n3198), .ZN(n3197) );
  INV_X1 U3820 ( .A(n5500), .ZN(n3198) );
  INV_X1 U3821 ( .A(n4146), .ZN(n5420) );
  AND2_X1 U3822 ( .A1(n5044), .A2(n5067), .ZN(n3181) );
  INV_X1 U3823 ( .A(n3608), .ZN(n3182) );
  NAND2_X1 U3824 ( .A1(n5787), .A2(n5786), .ZN(n3163) );
  NOR2_X1 U3825 ( .A1(n3144), .A2(n4241), .ZN(n3143) );
  INV_X1 U3826 ( .A(n6071), .ZN(n3144) );
  INV_X1 U3827 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6974) );
  NAND3_X1 U3828 ( .A1(n3146), .A2(n3147), .A3(n3208), .ZN(n5049) );
  INV_X1 U3829 ( .A(n4758), .ZN(n3146) );
  NOR2_X1 U3830 ( .A1(n3148), .A2(n4446), .ZN(n3147) );
  INV_X1 U3831 ( .A(n6108), .ZN(n3148) );
  AND2_X1 U3832 ( .A1(n3299), .A2(n3489), .ZN(n3655) );
  OR2_X1 U3833 ( .A1(n3452), .A2(n3451), .ZN(n3516) );
  NAND2_X1 U3834 ( .A1(n3377), .A2(n3358), .ZN(n3405) );
  AND3_X1 U3835 ( .A1(n3092), .A2(n3348), .A3(n3347), .ZN(n4189) );
  AND3_X1 U3836 ( .A1(n3342), .A2(n4460), .A3(n3346), .ZN(n3348) );
  OR2_X1 U3837 ( .A1(n3378), .A2(n3379), .ZN(n3386) );
  INV_X1 U3838 ( .A(n5906), .ZN(n4656) );
  AOI21_X1 U3839 ( .B1(n6560), .B2(n4652), .A(n5460), .ZN(n4471) );
  INV_X1 U3840 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6526) );
  INV_X1 U3841 ( .A(n3373), .ZN(n3691) );
  AND2_X1 U3842 ( .A1(n3676), .A2(n3655), .ZN(n3684) );
  AOI21_X1 U3843 ( .B1(n3667), .B2(n3655), .A(n4177), .ZN(n3680) );
  INV_X1 U3844 ( .A(n4343), .ZN(n4402) );
  AND2_X1 U3845 ( .A1(n4405), .A2(n4189), .ZN(n4399) );
  INV_X1 U3846 ( .A(n4605), .ZN(n4406) );
  NAND2_X1 U3847 ( .A1(n3341), .A2(n6671), .ZN(n4354) );
  OR2_X1 U3848 ( .A1(n5896), .A2(n3137), .ZN(n3158) );
  AND2_X1 U3849 ( .A1(n4256), .A2(n4255), .ZN(n5597) );
  OR2_X1 U3850 ( .A1(n4618), .A2(n4287), .ZN(n4605) );
  INV_X1 U3851 ( .A(n3716), .ZN(n3187) );
  NAND2_X1 U3852 ( .A1(n4617), .A2(n4616), .ZN(n4676) );
  OR2_X1 U3853 ( .A1(n4428), .A2(n4429), .ZN(n4674) );
  INV_X1 U3854 ( .A(n4673), .ZN(n5076) );
  INV_X1 U3855 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6701) );
  NOR2_X1 U3856 ( .A1(n4678), .A2(n6455), .ZN(n3725) );
  INV_X1 U3857 ( .A(n3824), .ZN(n5425) );
  NAND2_X1 U3858 ( .A1(n3196), .A2(n3195), .ZN(n3194) );
  INV_X1 U3859 ( .A(n5464), .ZN(n3195) );
  INV_X1 U3860 ( .A(n3197), .ZN(n3196) );
  NAND2_X1 U3861 ( .A1(n4107), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4112)
         );
  INV_X1 U3862 ( .A(n4069), .ZN(n4070) );
  NAND2_X1 U3863 ( .A1(n4050), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4069)
         );
  INV_X1 U3864 ( .A(n4000), .ZN(n4001) );
  AND2_X1 U3865 ( .A1(n4002), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4050)
         );
  INV_X1 U3866 ( .A(n5649), .ZN(n3968) );
  NOR2_X1 U3867 ( .A1(n3911), .A2(n6031), .ZN(n3912) );
  AND2_X1 U3868 ( .A1(n3912), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3948)
         );
  NOR2_X1 U3869 ( .A1(n6849), .A2(n3856), .ZN(n3874) );
  NOR2_X1 U3870 ( .A1(n6814), .A2(n3892), .ZN(n3891) );
  NOR2_X1 U3871 ( .A1(n3804), .A2(n3803), .ZN(n3821) );
  INV_X1 U3872 ( .A(n5087), .ZN(n3788) );
  NAND2_X1 U3873 ( .A1(n3758), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3773)
         );
  NOR2_X1 U3874 ( .A1(n3732), .A2(n6107), .ZN(n3739) );
  NOR2_X1 U3875 ( .A1(n3707), .A2(n4451), .ZN(n3189) );
  NAND2_X1 U3876 ( .A1(n4219), .A2(n4226), .ZN(n5390) );
  NOR2_X2 U3877 ( .A1(n3153), .A2(n3136), .ZN(n5516) );
  NOR2_X1 U3878 ( .A1(n5892), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5718)
         );
  AND2_X1 U3879 ( .A1(n5732), .A2(n3173), .ZN(n3172) );
  NAND2_X1 U3880 ( .A1(n3176), .A2(n3175), .ZN(n3173) );
  INV_X1 U3881 ( .A(n3176), .ZN(n3171) );
  AND2_X1 U3882 ( .A1(n4279), .A2(n4278), .ZN(n4280) );
  NAND2_X1 U3883 ( .A1(n5647), .A2(n4275), .ZN(n5555) );
  NAND2_X1 U3884 ( .A1(n5760), .A2(n5761), .ZN(n5759) );
  NOR2_X1 U3885 ( .A1(n5897), .A2(n5896), .ZN(n5898) );
  INV_X1 U3886 ( .A(n3168), .ZN(n3167) );
  NAND2_X1 U3887 ( .A1(n5340), .A2(n5342), .ZN(n5341) );
  NAND2_X1 U3888 ( .A1(n6072), .A2(n3143), .ZN(n5217) );
  NAND2_X1 U3889 ( .A1(n3616), .A2(n3091), .ZN(n3184) );
  NAND2_X1 U3890 ( .A1(n4299), .A2(n4406), .ZN(n5864) );
  XNOR2_X1 U3891 ( .A(n3607), .B(n5057), .ZN(n5044) );
  NAND2_X1 U3892 ( .A1(n3146), .A2(n3147), .ZN(n6110) );
  NOR2_X1 U3893 ( .A1(n4758), .A2(n4446), .ZN(n6109) );
  XNOR2_X1 U3894 ( .A(n3544), .B(n4218), .ZN(n4597) );
  OAI21_X1 U3895 ( .B1(n6306), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6305), 
        .ZN(n3525) );
  INV_X1 U3896 ( .A(n5864), .ZN(n6378) );
  NAND2_X1 U3897 ( .A1(n4214), .A2(n4213), .ZN(n4756) );
  NAND2_X1 U3898 ( .A1(n4193), .A2(n6543), .ZN(n4302) );
  NAND2_X1 U3899 ( .A1(n4192), .A2(n4191), .ZN(n4193) );
  AND2_X1 U3900 ( .A1(n4626), .A2(n4286), .ZN(n4191) );
  XNOR2_X1 U3901 ( .A(n3159), .B(n3510), .ZN(n3513) );
  INV_X1 U3902 ( .A(n3511), .ZN(n3512) );
  OAI22_X1 U3903 ( .A1(n3598), .A2(n4548), .B1(n3497), .B2(n3434), .ZN(n3402)
         );
  NAND2_X1 U3904 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  OR2_X1 U3905 ( .A1(n3368), .A2(n3689), .ZN(n5454) );
  NAND4_X1 U3906 ( .A1(n3697), .A2(n3342), .A3(n4427), .A4(n3310), .ZN(n4632)
         );
  NAND2_X1 U3907 ( .A1(n4189), .A2(n3341), .ZN(n4196) );
  INV_X1 U3908 ( .A(n3110), .ZN(n4823) );
  OR2_X1 U3909 ( .A1(n4466), .A2(n4468), .ZN(n5003) );
  AND2_X1 U3910 ( .A1(n3110), .A2(n4566), .ZN(n4583) );
  AND2_X1 U3911 ( .A1(n5288), .A2(n4464), .ZN(n6450) );
  NAND2_X1 U3912 ( .A1(n4822), .A2(n4823), .ZN(n6449) );
  NOR2_X1 U3913 ( .A1(n6637), .A2(n4471), .ZN(n4500) );
  NAND2_X1 U3914 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4652) );
  AND2_X1 U3915 ( .A1(n6645), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3687) );
  INV_X1 U3916 ( .A(n6554), .ZN(n6543) );
  INV_X1 U3917 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6849) );
  INV_X1 U3918 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6107) );
  INV_X1 U3919 ( .A(n6128), .ZN(n6113) );
  AND2_X1 U3920 ( .A1(n6092), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U3921 ( .A1(n4369), .A2(n4368), .ZN(n6130) );
  INV_X1 U3922 ( .A(n6153), .ZN(n6165) );
  INV_X1 U3923 ( .A(n6170), .ZN(n5663) );
  NAND2_X1 U3924 ( .A1(n6170), .A2(n5672), .ZN(n6153) );
  INV_X1 U3925 ( .A(n5751), .ZN(n5690) );
  INV_X1 U3926 ( .A(n5282), .ZN(n5198) );
  INV_X1 U3927 ( .A(n5951), .ZN(n6184) );
  NAND2_X1 U3928 ( .A1(n4684), .A2(n4683), .ZN(n6183) );
  INV_X1 U3929 ( .A(n6183), .ZN(n5001) );
  AND2_X1 U3930 ( .A1(n4680), .A2(n3344), .ZN(n4681) );
  NOR2_X1 U3931 ( .A1(n4652), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6665) );
  AND2_X1 U3932 ( .A1(n4419), .A2(n4418), .ZN(n6682) );
  NOR2_X1 U3933 ( .A1(n6665), .A2(n6682), .ZN(n6192) );
  NAND2_X2 U3936 ( .A1(n4419), .A2(n6545), .ZN(n6278) );
  OR2_X1 U3937 ( .A1(n5422), .A2(n5467), .ZN(n4351) );
  OAI21_X1 U3938 ( .B1(n5470), .B2(n6318), .A(n5469), .ZN(n5471) );
  AND2_X1 U3939 ( .A1(n3123), .A2(n5580), .ZN(n6171) );
  NAND2_X1 U3940 ( .A1(n5589), .A2(n3910), .ZN(n5579) );
  AND2_X1 U3941 ( .A1(n5667), .A2(n5666), .ZN(n6046) );
  AND2_X1 U3942 ( .A1(n4780), .A2(n4811), .ZN(n6300) );
  NAND2_X1 U3943 ( .A1(n4419), .A2(n6535), .ZN(n6284) );
  NAND2_X1 U3944 ( .A1(n6304), .A2(n6321), .ZN(n6318) );
  INV_X1 U3945 ( .A(n6304), .ZN(n6322) );
  INV_X1 U3946 ( .A(n6284), .ZN(n6320) );
  INV_X1 U3947 ( .A(n3156), .ZN(n3155) );
  AOI21_X1 U3948 ( .B1(n5394), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n3157), 
        .ZN(n3156) );
  INV_X1 U3949 ( .A(n5428), .ZN(n3157) );
  AND2_X1 U3950 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U3951 ( .A1(n4300), .A2(n6327), .ZN(n5994) );
  NAND2_X1 U3952 ( .A1(n5347), .A2(n5863), .ZN(n6327) );
  CLKBUF_X1 U3953 ( .A(n6295), .Z(n6296) );
  NOR2_X1 U3954 ( .A1(n4305), .A2(n4381), .ZN(n6384) );
  NOR2_X1 U3955 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4510), .ZN(n4381)
         );
  INV_X1 U3956 ( .A(n5359), .ZN(n4510) );
  INV_X1 U3957 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6799) );
  NAND2_X2 U3958 ( .A1(n3505), .A2(n3504), .ZN(n4957) );
  BUF_X1 U3959 ( .A(n3436), .Z(n3438) );
  NOR2_X2 U3960 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6447) );
  AND2_X1 U3961 ( .A1(n5906), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6446) );
  INV_X1 U3962 ( .A(n6447), .ZN(n6452) );
  INV_X1 U3963 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6530) );
  INV_X1 U3964 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6645) );
  INV_X1 U3965 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5462) );
  INV_X1 U3966 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3379) );
  INV_X1 U3967 ( .A(n6640), .ZN(n5460) );
  INV_X1 U3968 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6796) );
  CLKBUF_X1 U3969 ( .A(n4196), .Z(n6003) );
  INV_X1 U3970 ( .A(n4748), .ZN(n4665) );
  OAI21_X1 U3971 ( .B1(n4924), .B2(n4903), .A(n5295), .ZN(n4927) );
  INV_X1 U3972 ( .A(n4900), .ZN(n4929) );
  INV_X1 U3973 ( .A(n6441), .ZN(n6396) );
  AND2_X1 U3974 ( .A1(n4583), .A2(n4571), .ZN(n6434) );
  AOI22_X1 U3975 ( .A1(n5293), .A2(n6450), .B1(n5289), .B2(n6400), .ZN(n5338)
         );
  INV_X1 U3976 ( .A(n5128), .ZN(n6490) );
  INV_X1 U3977 ( .A(n6487), .ZN(n6501) );
  INV_X1 U3978 ( .A(n6459), .ZN(n5339) );
  INV_X1 U3979 ( .A(n5143), .ZN(n6464) );
  INV_X1 U3980 ( .A(n6465), .ZN(n5331) );
  INV_X1 U3981 ( .A(n5137), .ZN(n6470) );
  INV_X1 U3982 ( .A(n6477), .ZN(n5313) );
  INV_X1 U3983 ( .A(n5131), .ZN(n6483) );
  INV_X1 U3984 ( .A(n6484), .ZN(n5327) );
  INV_X1 U3985 ( .A(n6491), .ZN(n5319) );
  INV_X1 U3986 ( .A(n6497), .ZN(n5307) );
  INV_X1 U3987 ( .A(n4894), .ZN(n4879) );
  OAI211_X1 U3988 ( .C1(n4719), .C2(n6959), .A(n4693), .B(n4692), .ZN(n4716)
         );
  INV_X1 U3989 ( .A(n5122), .ZN(n6504) );
  INV_X1 U3990 ( .A(n6506), .ZN(n5301) );
  NOR2_X1 U3991 ( .A1(n4870), .A2(n4963), .ZN(n6459) );
  NOR2_X1 U3992 ( .A1(n4785), .A2(n4963), .ZN(n6465) );
  NOR2_X1 U3993 ( .A1(n4788), .A2(n4963), .ZN(n6471) );
  AND2_X1 U3994 ( .A1(DATAI_3_), .A2(n4689), .ZN(n6477) );
  NOR2_X1 U3995 ( .A1(n6962), .A2(n4963), .ZN(n6484) );
  AND2_X1 U3996 ( .A1(DATAI_5_), .A2(n4689), .ZN(n6491) );
  AND2_X1 U3997 ( .A1(DATAI_6_), .A2(n4689), .ZN(n6497) );
  AND2_X1 U3998 ( .A1(n4657), .A2(n4571), .ZN(n4663) );
  INV_X1 U3999 ( .A(n4663), .ZN(n4552) );
  INV_X1 U4000 ( .A(n4690), .ZN(n4717) );
  NAND2_X1 U4001 ( .A1(n6645), .A2(n6455), .ZN(n6560) );
  INV_X1 U4002 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U4003 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4622), .ZN(n6640) );
  INV_X1 U4004 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U4005 ( .A1(n4171), .A2(n6573), .ZN(n6671) );
  INV_X1 U4006 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6601) );
  AND4_X1 U4007 ( .A1(n6143), .A2(n6142), .A3(n6141), .A4(n6140), .ZN(n6144)
         );
  AND2_X1 U4008 ( .A1(n4340), .A2(n3204), .ZN(n4341) );
  AND2_X1 U4009 ( .A1(n4318), .A2(n4317), .ZN(n4319) );
  AND2_X1 U4010 ( .A1(n3219), .A2(n4606), .ZN(n3318) );
  OR3_X1 U4011 ( .A1(n5578), .A2(n3192), .A3(n3190), .ZN(n3123) );
  AND4_X1 U4012 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3124)
         );
  NAND2_X1 U4013 ( .A1(n3368), .A2(n3364), .ZN(n3347) );
  NAND2_X1 U4014 ( .A1(n3842), .A2(n3827), .ZN(n3125) );
  BUF_X1 U4015 ( .A(n4226), .Z(n5384) );
  OR3_X1 U4016 ( .A1(n5897), .A2(n5582), .A3(n3158), .ZN(n3126) );
  AND2_X1 U4017 ( .A1(n3163), .A2(n3626), .ZN(n3127) );
  NAND2_X1 U4018 ( .A1(n3162), .A2(n3160), .ZN(n4163) );
  NAND2_X1 U4019 ( .A1(n5341), .A2(n3622), .ZN(n5797) );
  AND3_X1 U4020 ( .A1(n3300), .A2(n3301), .A3(n3302), .ZN(n3128) );
  AND2_X1 U4021 ( .A1(n5499), .A2(n5500), .ZN(n3129) );
  AND2_X1 U4022 ( .A1(n3299), .A2(n3341), .ZN(n3130) );
  AND2_X1 U4023 ( .A1(n5892), .A2(n4301), .ZN(n3131) );
  NOR2_X1 U4024 ( .A1(n5393), .A2(n3155), .ZN(n3132) );
  AND2_X1 U4025 ( .A1(n3615), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3133)
         );
  NAND2_X1 U4026 ( .A1(n5354), .A2(n5355), .ZN(n3134) );
  NAND2_X1 U4027 ( .A1(n3184), .A2(n3618), .ZN(n5199) );
  NAND2_X1 U4028 ( .A1(n3183), .A2(n3608), .ZN(n5066) );
  NAND2_X1 U4029 ( .A1(n3102), .A2(n5275), .ZN(n5340) );
  NAND2_X1 U4030 ( .A1(n3364), .A2(n3374), .ZN(n4289) );
  OR2_X1 U4031 ( .A1(n5897), .A2(n3158), .ZN(n3135) );
  OR2_X1 U4032 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5416) );
  OR2_X1 U4033 ( .A1(n5513), .A2(n5512), .ZN(n3136) );
  NAND2_X1 U4034 ( .A1(n3186), .A2(n4809), .ZN(n4780) );
  NAND2_X1 U4035 ( .A1(n6072), .A2(n6071), .ZN(n5092) );
  XNOR2_X1 U4036 ( .A(n3571), .B(n6969), .ZN(n6294) );
  OAI21_X1 U4037 ( .B1(n4452), .B2(n3189), .A(n3708), .ZN(n4450) );
  INV_X2 U4038 ( .A(n6325), .ZN(n6314) );
  AND2_X1 U4039 ( .A1(n4262), .A2(n4261), .ZN(n3137) );
  NOR2_X1 U4040 ( .A1(n3346), .A2(n3341), .ZN(n4290) );
  AOI21_X1 U4041 ( .B1(n3333), .B2(n3369), .A(n3341), .ZN(n3370) );
  NAND2_X1 U4042 ( .A1(n5642), .A2(n5643), .ZN(n5637) );
  NAND2_X1 U4043 ( .A1(n5550), .A2(n4036), .ZN(n5626) );
  AND2_X2 U4044 ( .A1(n5086), .A2(n6064), .ZN(n6065) );
  AND2_X2 U4045 ( .A1(n5060), .A2(n3788), .ZN(n5086) );
  NOR2_X2 U4046 ( .A1(n5059), .A2(n3772), .ZN(n5060) );
  NAND3_X2 U4047 ( .A1(n3124), .A2(n3303), .A3(n3128), .ZN(n3364) );
  NAND2_X2 U4048 ( .A1(n3363), .A2(n3299), .ZN(n3368) );
  NOR2_X2 U4049 ( .A1(n3549), .A2(n3548), .ZN(n3563) );
  NAND2_X1 U4050 ( .A1(n3724), .A2(n3901), .ZN(n3731) );
  OAI21_X2 U4051 ( .B1(n5525), .B2(n5510), .A(n5499), .ZN(n5713) );
  INV_X1 U4052 ( .A(n3145), .ZN(n5356) );
  INV_X1 U4053 ( .A(n3153), .ZN(n5538) );
  OAI211_X1 U4054 ( .C1(n5618), .C2(n6352), .A(n3132), .B(n3154), .ZN(U2987)
         );
  XNOR2_X2 U4055 ( .A(n5392), .B(n5391), .ZN(n5618) );
  INV_X1 U4056 ( .A(n3159), .ZN(n3465) );
  NAND2_X1 U4057 ( .A1(n3159), .A2(n3510), .ZN(n3463) );
  NAND2_X1 U4058 ( .A1(n5790), .A2(n5786), .ZN(n3162) );
  OAI21_X1 U4059 ( .B1(n5790), .B2(n5787), .A(n5786), .ZN(n5780) );
  NAND2_X1 U4060 ( .A1(n3164), .A2(n3167), .ZN(n3625) );
  NAND2_X1 U4061 ( .A1(n3621), .A2(n3165), .ZN(n3164) );
  NAND2_X1 U4062 ( .A1(n5771), .A2(n3629), .ZN(n5772) );
  NAND2_X1 U4063 ( .A1(n4337), .A2(n5742), .ZN(n3178) );
  NAND2_X1 U4064 ( .A1(n5043), .A2(n5044), .ZN(n3183) );
  NAND2_X1 U4065 ( .A1(n3180), .A2(n3179), .ZN(n5154) );
  AOI21_X1 U4066 ( .B1(n3182), .B2(n5067), .A(n3133), .ZN(n3179) );
  NAND2_X1 U4067 ( .A1(n5043), .A2(n3181), .ZN(n3180) );
  NAND2_X1 U4068 ( .A1(n4521), .A2(n3901), .ZN(n3188) );
  AND2_X2 U4069 ( .A1(n3549), .A2(n3488), .ZN(n4521) );
  NAND2_X1 U4070 ( .A1(n5589), .A2(n3191), .ZN(n5562) );
  NAND2_X1 U4071 ( .A1(n3437), .A2(n3358), .ZN(n3193) );
  INV_X1 U4072 ( .A(n5426), .ZN(n3199) );
  NAND2_X1 U4073 ( .A1(n3570), .A2(n3569), .ZN(n3571) );
  OAI21_X1 U4074 ( .B1(n5476), .B2(n6325), .A(n5472), .ZN(n5473) );
  CLKBUF_X1 U4075 ( .A(n4521), .Z(n4822) );
  CLKBUF_X1 U4076 ( .A(n4935), .Z(n4999) );
  NAND2_X1 U4077 ( .A1(n4678), .A2(n3345), .ZN(n3344) );
  AND2_X4 U4078 ( .A1(n5459), .A2(n4634), .ZN(n3574) );
  NAND2_X1 U4079 ( .A1(n5709), .A2(n5808), .ZN(n5434) );
  OR2_X1 U4080 ( .A1(n3356), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3202)
         );
  AND2_X1 U4081 ( .A1(n5718), .A2(n5807), .ZN(n3203) );
  INV_X1 U4082 ( .A(n3725), .ZN(n3928) );
  OR2_X1 U4083 ( .A1(n5448), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3204)
         );
  INV_X1 U4084 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4350) );
  AND4_X1 U4085 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3205)
         );
  INV_X1 U4086 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U4087 ( .A1(n4299), .A2(n4199), .ZN(n6370) );
  NAND2_X1 U4088 ( .A1(n5507), .A2(REIP_REG_29__SCAN_IN), .ZN(n3206) );
  OR2_X1 U4089 ( .A1(n5619), .A2(n6100), .ZN(n3207) );
  NAND2_X1 U4090 ( .A1(n4229), .A2(n4228), .ZN(n3208) );
  INV_X1 U4091 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3632) );
  NAND2_X2 U4092 ( .A1(n6170), .A2(n4678), .ZN(n6148) );
  AOI21_X1 U4093 ( .B1(n3649), .B2(n3640), .A(n3639), .ZN(n3666) );
  NAND2_X1 U4094 ( .A1(n3724), .A2(n3655), .ZN(n3570) );
  NOR2_X1 U4095 ( .A1(n6530), .A2(n3646), .ZN(n3647) );
  OR2_X1 U4096 ( .A1(n4048), .A2(n4047), .ZN(n4065) );
  INV_X1 U4097 ( .A(n4289), .ZN(n3332) );
  INV_X1 U4098 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4635) );
  INV_X1 U4099 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6688) );
  AND2_X1 U4100 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4001), .ZN(n4002)
         );
  AND2_X1 U4101 ( .A1(n3586), .A2(n3585), .ZN(n3589) );
  NAND2_X1 U4102 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4103 ( .A1(n3444), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3300) );
  INV_X1 U4104 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3803) );
  AND2_X1 U4105 ( .A1(n4354), .A2(n4353), .ZN(n4355) );
  NAND2_X1 U4106 ( .A1(n4382), .A2(n5384), .ZN(n4332) );
  INV_X1 U4107 ( .A(n5551), .ZN(n4036) );
  OR2_X1 U4108 ( .A1(n6003), .A2(n4615), .ZN(n4616) );
  INV_X1 U4109 ( .A(n6517), .ZN(n4637) );
  INV_X1 U4110 ( .A(n4108), .ZN(n4107) );
  NOR2_X1 U4111 ( .A1(n3773), .A2(n6075), .ZN(n3789) );
  AND2_X1 U4112 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3726), .ZN(n3727)
         );
  INV_X1 U4113 ( .A(n4456), .ZN(n4213) );
  NAND2_X1 U4114 ( .A1(n3473), .A2(n3472), .ZN(n5004) );
  AND2_X1 U4115 ( .A1(n4179), .A2(n3684), .ZN(n3685) );
  INV_X1 U4116 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6031) );
  INV_X1 U4117 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6814) );
  OR2_X1 U4118 ( .A1(n4346), .A2(n6548), .ZN(n4347) );
  NAND2_X1 U4119 ( .A1(n5516), .A2(n5501), .ZN(n5388) );
  AND2_X1 U4120 ( .A1(n4269), .A2(n4268), .ZN(n5644) );
  AND2_X1 U4121 ( .A1(n4170), .A2(n4413), .ZN(n4624) );
  AOI21_X1 U4122 ( .B1(n4637), .B2(n4417), .A(n6671), .ZN(n4418) );
  XNOR2_X1 U4123 ( .A(n4351), .B(n4350), .ZN(n5429) );
  NAND2_X1 U4124 ( .A1(n4070), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4088)
         );
  NAND2_X1 U4125 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3951), .ZN(n4000)
         );
  INV_X1 U4126 ( .A(n5562), .ZN(n5650) );
  AND2_X1 U4127 ( .A1(n4322), .A2(n4321), .ZN(n5816) );
  NAND2_X1 U4128 ( .A1(n3625), .A2(n3624), .ZN(n5790) );
  INV_X1 U4129 ( .A(n5052), .ZN(n4305) );
  NAND2_X1 U4130 ( .A1(n4299), .A2(n6517), .ZN(n5359) );
  AND2_X1 U4131 ( .A1(n4522), .A2(n4823), .ZN(n4731) );
  AND2_X1 U4132 ( .A1(n3351), .A2(n3381), .ZN(n4962) );
  INV_X1 U4133 ( .A(n6434), .ZN(n5262) );
  INV_X1 U4134 ( .A(n5290), .ZN(n5334) );
  INV_X1 U4135 ( .A(n4957), .ZN(n5115) );
  AND2_X1 U4136 ( .A1(n4362), .A2(n5923), .ZN(n5914) );
  NOR2_X1 U4137 ( .A1(n4357), .A2(n5566), .ZN(n5945) );
  NAND2_X1 U4138 ( .A1(n3822), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3892)
         );
  OR2_X1 U4139 ( .A1(n6663), .A2(n4347), .ZN(n6092) );
  AND2_X1 U4140 ( .A1(n3739), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3758)
         );
  AND2_X1 U4141 ( .A1(n6092), .A2(n4370), .ZN(n6081) );
  INV_X1 U4142 ( .A(n6130), .ZN(n6112) );
  INV_X1 U4143 ( .A(n6148), .ZN(n6166) );
  NOR2_X2 U4144 ( .A1(n6179), .A2(n3344), .ZN(n6177) );
  INV_X2 U4145 ( .A(n6186), .ZN(n6179) );
  INV_X1 U4146 ( .A(n6222), .ZN(n6271) );
  INV_X1 U4147 ( .A(n4417), .ZN(n6545) );
  INV_X1 U4148 ( .A(n6318), .ZN(n6298) );
  AND2_X1 U4149 ( .A1(n4439), .A2(n3707), .ZN(n6313) );
  NOR2_X1 U4150 ( .A1(n5839), .A2(n4339), .ZN(n5820) );
  INV_X1 U4151 ( .A(n4322), .ZN(n5836) );
  OR2_X1 U4152 ( .A1(n5901), .A2(n4310), .ZN(n5858) );
  NOR2_X1 U4153 ( .A1(n5994), .A2(n5984), .ZN(n5903) );
  OR2_X1 U4154 ( .A1(n6651), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4156) );
  INV_X1 U4155 ( .A(n6001), .ZN(n6333) );
  OR2_X1 U4156 ( .A1(n5348), .A2(n4510), .ZN(n6339) );
  INV_X1 U4157 ( .A(n6001), .ZN(n6375) );
  INV_X1 U4158 ( .A(n6370), .ZN(n6382) );
  INV_X1 U4159 ( .A(n4689), .ZN(n4963) );
  AND2_X1 U4160 ( .A1(n4731), .A2(n4957), .ZN(n4748) );
  AND2_X1 U4161 ( .A1(n4731), .A2(n5115), .ZN(n4931) );
  OAI21_X1 U4162 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(n4853) );
  OAI21_X1 U4163 ( .B1(n5009), .B2(n5008), .A(n5007), .ZN(n5035) );
  INV_X1 U4164 ( .A(n5037), .ZN(n5031) );
  AND2_X1 U4165 ( .A1(n5906), .A2(n4957), .ZN(n4821) );
  NOR2_X1 U4166 ( .A1(n5116), .A2(n5906), .ZN(n5290) );
  NOR2_X1 U4167 ( .A1(n4526), .A2(n6455), .ZN(n6400) );
  INV_X1 U4168 ( .A(n5119), .ZN(n6476) );
  INV_X1 U4169 ( .A(n5125), .ZN(n6496) );
  INV_X1 U4170 ( .A(n6510), .ZN(n6481) );
  OR2_X1 U4171 ( .A1(n4966), .A2(n4965), .ZN(n4990) );
  INV_X1 U4172 ( .A(n5134), .ZN(n6445) );
  NOR2_X1 U4173 ( .A1(n6217), .A2(n4963), .ZN(n6506) );
  AND2_X1 U4174 ( .A1(n6786), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4345) );
  INV_X1 U4175 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U4176 ( .A1(n4393), .A2(n4394), .ZN(n6663) );
  INV_X1 U4177 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6941) );
  AOI211_X1 U4178 ( .C1(n5496), .C2(REIP_REG_31__SCAN_IN), .A(n5495), .B(n5494), .ZN(n5497) );
  NAND2_X1 U4179 ( .A1(n6092), .A2(n5095), .ZN(n6128) );
  INV_X1 U4180 ( .A(n6126), .ZN(n6106) );
  INV_X1 U4181 ( .A(n6125), .ZN(n6123) );
  AND2_X2 U4182 ( .A1(n4431), .A2(n6543), .ZN(n6170) );
  INV_X1 U4183 ( .A(n6046), .ZN(n5697) );
  INV_X1 U4184 ( .A(DATAI_4_), .ZN(n6962) );
  NAND2_X1 U4185 ( .A1(n4677), .A2(n6239), .ZN(n6186) );
  NAND2_X1 U4186 ( .A1(n6682), .A2(n4490), .ZN(n4779) );
  INV_X1 U4187 ( .A(n6682), .ZN(n6203) );
  INV_X1 U4188 ( .A(n6263), .ZN(n6222) );
  OR2_X1 U4189 ( .A1(n5642), .A2(n5651), .ZN(n5942) );
  NAND2_X1 U4190 ( .A1(n6284), .A2(n4153), .ZN(n6304) );
  OR2_X1 U4191 ( .A1(n6562), .A2(n6452), .ZN(n6325) );
  OR2_X1 U4192 ( .A1(n5861), .A2(n4338), .ZN(n5839) );
  INV_X1 U4193 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5987) );
  OR2_X1 U4194 ( .A1(n4156), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U4195 ( .A1(n4299), .A2(n4283), .ZN(n6352) );
  NAND2_X1 U4196 ( .A1(n6959), .A2(n6645), .ZN(n6651) );
  INV_X1 U4197 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4540) );
  AND2_X1 U4198 ( .A1(n4525), .A2(n4524), .ZN(n4670) );
  INV_X1 U4199 ( .A(n4724), .ZN(n4751) );
  AND2_X1 U4200 ( .A1(n4898), .A2(n4897), .ZN(n4928) );
  AOI22_X1 U4201 ( .A1(n4820), .A2(n4827), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4819), .ZN(n4855) );
  AOI22_X1 U4202 ( .A1(n4587), .A2(n4589), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4586), .ZN(n4808) );
  NAND2_X1 U4203 ( .A1(n4583), .A2(n4821), .ZN(n6441) );
  AOI21_X1 U4204 ( .B1(n5230), .B2(n5228), .A(n5227), .ZN(n5270) );
  INV_X1 U4205 ( .A(n5108), .ZN(n5142) );
  OR2_X1 U4206 ( .A1(n6449), .A2(n5285), .ZN(n6487) );
  NAND2_X1 U4207 ( .A1(n4958), .A2(n5906), .ZN(n6510) );
  INV_X1 U4208 ( .A(n4891), .ZN(n4882) );
  INV_X1 U4209 ( .A(n6471), .ZN(n5323) );
  NAND2_X1 U4210 ( .A1(n4500), .A2(n3364), .ZN(n5119) );
  NAND2_X1 U4211 ( .A1(n3687), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U4212 ( .A1(n6786), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U4213 ( .A1(n6679), .A2(n6012), .ZN(n6635) );
  INV_X1 U4214 ( .A(READY_N), .ZN(n6666) );
  INV_X1 U4215 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6718) );
  INV_X1 U4216 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U4217 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6679), .ZN(n6625) );
  NOR2_X4 U4218 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4633) );
  NOR2_X4 U4219 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4645) );
  AND2_X4 U4220 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4606) );
  AOI22_X1 U4221 ( .A1(n3112), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3215) );
  INV_X1 U4222 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4223 ( .A1(n4134), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3214) );
  INV_X1 U4224 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3211) );
  AND2_X2 U4225 ( .A1(n5459), .A2(n4633), .ZN(n3809) );
  AOI22_X1 U4226 ( .A1(n5403), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3809), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4227 ( .A1(n3446), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3212) );
  INV_X1 U4228 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4229 ( .A1(n3444), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4230 ( .A1(n3311), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3222) );
  AND2_X2 U4231 ( .A1(n3218), .A2(n3219), .ZN(n3317) );
  AOI22_X1 U4232 ( .A1(n4133), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4233 ( .A1(n5397), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3220) );
  NAND2_X4 U4234 ( .A1(n3225), .A2(n3224), .ZN(n3299) );
  INV_X1 U4235 ( .A(n3299), .ZN(n4679) );
  AOI22_X1 U4236 ( .A1(n3112), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4237 ( .A1(n3446), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4238 ( .A1(n4134), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4239 ( .A1(n3094), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4240 ( .A1(n4133), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3231) );
  NAND2_X2 U4241 ( .A1(n3235), .A2(n3234), .ZN(n3345) );
  NAND2_X2 U4242 ( .A1(n4679), .A2(n3345), .ZN(n4428) );
  AOI22_X1 U4243 ( .A1(n5403), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3809), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4244 ( .A1(n3111), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4245 ( .A1(n3424), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4246 ( .A1(n3446), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4247 ( .A1(n3574), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5397), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4248 ( .A1(n3096), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4249 ( .A1(n3311), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4250 ( .A1(n3444), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3240) );
  INV_X2 U4251 ( .A(n3310), .ZN(n3324) );
  AOI22_X1 U4252 ( .A1(n4134), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5403), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4253 ( .A1(n3097), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4254 ( .A1(n3311), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4255 ( .A1(n3444), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4256 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3255)
         );
  AOI22_X1 U4257 ( .A1(n5397), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4258 ( .A1(n3312), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3424), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4259 ( .A1(n3122), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4260 ( .A1(n3446), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3250) );
  NAND4_X1 U4261 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3254)
         );
  NAND2_X1 U4262 ( .A1(n3446), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3260) );
  NAND2_X1 U4263 ( .A1(n3312), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4264 ( .A1(n3574), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3258)
         );
  NAND2_X1 U4265 ( .A1(n3113), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3257)
         );
  NAND2_X1 U4266 ( .A1(n5397), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3264) );
  NAND2_X1 U4267 ( .A1(n4133), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4268 ( .A1(n3317), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3262)
         );
  NAND2_X1 U4269 ( .A1(n3311), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3261)
         );
  NAND2_X1 U4270 ( .A1(n3122), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4271 ( .A1(n3318), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3267)
         );
  NAND2_X1 U4272 ( .A1(n3444), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4273 ( .A1(n3390), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3265)
         );
  NAND2_X1 U4274 ( .A1(n4134), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4275 ( .A1(n3115), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4276 ( .A1(n3424), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4277 ( .A1(n3118), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3269) );
  AND2_X1 U4278 ( .A1(n3340), .A2(n3368), .ZN(n3277) );
  NAND2_X1 U4279 ( .A1(n3446), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4280 ( .A1(n3115), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4281 ( .A1(n3122), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4282 ( .A1(n3113), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3278)
         );
  NAND2_X1 U4283 ( .A1(n3311), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4284 ( .A1(n4133), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4285 ( .A1(n3317), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4286 ( .A1(n3318), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3282)
         );
  NAND2_X1 U4287 ( .A1(n3444), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4288 ( .A1(n5397), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4289 ( .A1(n3574), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3287)
         );
  NAND2_X1 U4290 ( .A1(n3390), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3286)
         );
  NAND2_X1 U4291 ( .A1(n4134), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4292 ( .A1(n3312), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U4293 ( .A1(n3118), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4294 ( .A1(n3112), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3290) );
  NAND4_X4 U4295 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3489)
         );
  NAND2_X1 U4296 ( .A1(n3100), .A2(n3490), .ZN(n3298) );
  NAND2_X1 U4297 ( .A1(n4188), .A2(n3298), .ZN(n3309) );
  XNOR2_X1 U4298 ( .A(n6564), .B(STATE_REG_1__SCAN_IN), .ZN(n4171) );
  NOR2_X1 U4299 ( .A1(n3489), .A2(n4171), .ZN(n3349) );
  AOI22_X1 U4300 ( .A1(n3311), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4301 ( .A1(n4133), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4302 ( .A1(n5397), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4303 ( .A1(n3115), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4304 ( .A1(n4134), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4305 ( .A1(n3424), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4306 ( .A1(n3446), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3304) );
  INV_X2 U4307 ( .A(n3340), .ZN(n3342) );
  OAI211_X1 U4308 ( .C1(n3349), .C2(n3299), .A(n3361), .B(n5077), .ZN(n3308)
         );
  AOI22_X1 U4309 ( .A1(n3115), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4310 ( .A1(n3311), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4311 ( .A1(n3312), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4312 ( .A1(n3446), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4313 ( .A1(n4133), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4314 ( .A1(n5397), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4315 ( .A1(n4134), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3112), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4316 ( .A1(n3444), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3319) );
  NAND2_X2 U4317 ( .A1(n3323), .A2(n3205), .ZN(n3346) );
  MUX2_X1 U4318 ( .A(n3310), .B(n3346), .S(n3345), .Z(n3329) );
  INV_X1 U4319 ( .A(n4428), .ZN(n3328) );
  NAND2_X1 U4320 ( .A1(n4428), .A2(n3324), .ZN(n3325) );
  NAND2_X1 U4321 ( .A1(n3325), .A2(n3346), .ZN(n3326) );
  NAND2_X1 U4322 ( .A1(n3372), .A2(n3342), .ZN(n3335) );
  NAND2_X1 U4323 ( .A1(n3373), .A2(n4678), .ZN(n3330) );
  NAND2_X1 U4324 ( .A1(n3330), .A2(n3344), .ZN(n3331) );
  NAND2_X1 U4325 ( .A1(n3331), .A2(n4428), .ZN(n3367) );
  INV_X1 U4326 ( .A(n3367), .ZN(n3333) );
  NAND2_X1 U4327 ( .A1(n3333), .A2(n3332), .ZN(n3688) );
  INV_X1 U4328 ( .A(n3688), .ZN(n3334) );
  NAND3_X1 U4329 ( .A1(n3336), .A2(n3335), .A3(n3334), .ZN(n3337) );
  NAND2_X2 U4330 ( .A1(n3337), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3378) );
  INV_X1 U4331 ( .A(n3378), .ZN(n3338) );
  NAND2_X1 U4332 ( .A1(n3338), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3353) );
  NOR2_X1 U4333 ( .A1(n4289), .A2(n3299), .ZN(n3339) );
  AND2_X2 U4334 ( .A1(n3092), .A2(n3339), .ZN(n4170) );
  NAND2_X1 U4335 ( .A1(n4170), .A2(n4490), .ZN(n4343) );
  NOR2_X1 U4336 ( .A1(n3299), .A2(n3364), .ZN(n3343) );
  NAND3_X1 U4337 ( .A1(n3343), .A2(n3374), .A3(n4673), .ZN(n4601) );
  OAI211_X1 U4338 ( .C1(n4343), .C2(n3349), .A(n4282), .B(n4196), .ZN(n3350)
         );
  NAND2_X1 U4339 ( .A1(n3350), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4340 ( .A1(n6799), .A2(n6701), .ZN(n3351) );
  NAND2_X1 U4341 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3381) );
  INV_X1 U4342 ( .A(n3687), .ZN(n3383) );
  AND2_X1 U4343 ( .A1(n3383), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3352)
         );
  NAND3_X1 U4344 ( .A1(n3353), .A2(n3354), .A3(n3355), .ZN(n3377) );
  INV_X1 U4345 ( .A(n3354), .ZN(n3357) );
  INV_X1 U4346 ( .A(n3355), .ZN(n3356) );
  NAND2_X1 U4347 ( .A1(n3357), .A2(n3202), .ZN(n3358) );
  MUX2_X1 U4348 ( .A(n3383), .B(n3384), .S(n6799), .Z(n3359) );
  INV_X1 U4349 ( .A(n3359), .ZN(n3360) );
  OAI21_X1 U4350 ( .B1(n3100), .B2(n3347), .A(n3490), .ZN(n3366) );
  OR2_X1 U4351 ( .A1(n6651), .A2(n6786), .ZN(n6555) );
  INV_X1 U4352 ( .A(n6555), .ZN(n3365) );
  AND2_X1 U4353 ( .A1(n3363), .A2(n4678), .ZN(n3697) );
  NAND4_X1 U4354 ( .A1(n3366), .A2(n3365), .A3(n3362), .A4(n4632), .ZN(n3371)
         );
  INV_X1 U4355 ( .A(n3364), .ZN(n4200) );
  AOI21_X1 U4356 ( .B1(n3368), .B2(n3310), .A(n4200), .ZN(n3369) );
  NOR2_X1 U4357 ( .A1(n3371), .A2(n3370), .ZN(n3376) );
  OAI22_X1 U4358 ( .A1(n3691), .A2(n5077), .B1(n3342), .B2(n3374), .ZN(n3375)
         );
  NAND2_X1 U4359 ( .A1(n3376), .A2(n4296), .ZN(n3439) );
  INV_X1 U4360 ( .A(n3381), .ZN(n3380) );
  NAND2_X1 U4361 ( .A1(n3380), .A2(n6526), .ZN(n6443) );
  NAND2_X1 U4362 ( .A1(n3381), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4363 ( .A1(n6443), .A2(n3382), .ZN(n4526) );
  AOI22_X1 U4364 ( .A1(n3384), .A2(n4526), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3383), .ZN(n3385) );
  NAND2_X1 U4365 ( .A1(n3386), .A2(n3385), .ZN(n3387) );
  NAND2_X1 U4366 ( .A1(n3388), .A2(n3387), .ZN(n3469) );
  NAND2_X1 U4367 ( .A1(n3389), .A2(n3469), .ZN(n4465) );
  AOI22_X1 U4368 ( .A1(n5397), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4369 ( .A1(n4133), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4370 ( .A1(n3311), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4371 ( .A1(n4135), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4372 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3401)
         );
  AOI22_X1 U4373 ( .A1(n4134), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4374 ( .A1(n3115), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4375 ( .A1(n3093), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4376 ( .A1(n4094), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3396) );
  NAND4_X1 U4377 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3400)
         );
  NOR2_X1 U4378 ( .A1(n3401), .A2(n3400), .ZN(n3497) );
  NAND2_X1 U4379 ( .A1(n3324), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3406) );
  OAI22_X1 U4380 ( .A1(n4465), .A2(STATE2_REG_0__SCAN_IN), .B1(n3497), .B2(
        n3406), .ZN(n3403) );
  INV_X1 U4381 ( .A(n3676), .ZN(n3598) );
  INV_X1 U4382 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4548) );
  NAND2_X1 U4383 ( .A1(n3342), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3434) );
  XNOR2_X1 U4384 ( .A(n3403), .B(n3402), .ZN(n3494) );
  INV_X1 U4385 ( .A(n3494), .ZN(n3468) );
  INV_X1 U4386 ( .A(n3437), .ZN(n3404) );
  XNOR2_X1 U4387 ( .A(n3405), .B(n3404), .ZN(n4467) );
  NAND2_X1 U4388 ( .A1(n4467), .A2(n6786), .ZN(n3418) );
  INV_X1 U4389 ( .A(n3406), .ZN(n3432) );
  AOI22_X1 U4390 ( .A1(n4135), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4391 ( .A1(n4133), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4392 ( .A1(n5397), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4393 ( .A1(n4134), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3407) );
  NAND4_X1 U4394 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3416)
         );
  AOI22_X1 U4395 ( .A1(n3115), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4396 ( .A1(n5404), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4397 ( .A1(n4094), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4398 ( .A1(n3311), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3411) );
  NAND4_X1 U4399 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n3415)
         );
  NAND2_X1 U4400 ( .A1(n3432), .A2(n3515), .ZN(n3417) );
  INV_X1 U4401 ( .A(n3515), .ZN(n3435) );
  INV_X1 U4402 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4556) );
  OR2_X1 U4403 ( .A1(n3598), .A2(n4556), .ZN(n3433) );
  AOI22_X1 U4404 ( .A1(n5397), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4405 ( .A1(n4133), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4406 ( .A1(n3311), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3421) );
  INV_X1 U4407 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4408 ( .A1(n4135), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3420) );
  NAND4_X1 U4409 ( .A1(n3423), .A2(n3422), .A3(n3421), .A4(n3420), .ZN(n3430)
         );
  AOI22_X1 U4410 ( .A1(n4134), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4411 ( .A1(n3115), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4412 ( .A1(n3093), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4413 ( .A1(n4094), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3425) );
  NAND4_X1 U4414 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3429)
         );
  INV_X1 U4415 ( .A(n3612), .ZN(n3431) );
  NAND2_X1 U4416 ( .A1(n3432), .A2(n3431), .ZN(n3453) );
  OAI21_X2 U4417 ( .B1(n3439), .B2(n3438), .A(n3103), .ZN(n3698) );
  NAND2_X1 U4418 ( .A1(n3324), .A2(n3612), .ZN(n3462) );
  AOI22_X1 U4419 ( .A1(n4134), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4420 ( .A1(n3097), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4421 ( .A1(n3095), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4422 ( .A1(n3115), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3440) );
  NAND4_X1 U4423 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3452)
         );
  AOI22_X1 U4424 ( .A1(n3311), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4425 ( .A1(n4135), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4426 ( .A1(n3395), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4427 ( .A1(n4094), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4428 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3451)
         );
  OR2_X1 U4429 ( .A1(n3462), .A2(n3516), .ZN(n3454) );
  OAI21_X1 U4430 ( .B1(n3698), .B2(STATE2_REG_0__SCAN_IN), .A(n3456), .ZN(
        n3461) );
  OAI211_X1 U4431 ( .C1(n3457), .C2(n4490), .A(n3462), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3458) );
  INV_X1 U4432 ( .A(n3458), .ZN(n3459) );
  NAND2_X1 U4433 ( .A1(n3460), .A2(n3459), .ZN(n3501) );
  NAND2_X1 U4434 ( .A1(n3461), .A2(n3501), .ZN(n3505) );
  AND2_X2 U4435 ( .A1(n3505), .A2(n3609), .ZN(n3511) );
  NAND2_X1 U4436 ( .A1(n3463), .A2(n3511), .ZN(n3467) );
  INV_X1 U4437 ( .A(n3510), .ZN(n3464) );
  AND2_X2 U4438 ( .A1(n3467), .A2(n3466), .ZN(n3495) );
  NAND2_X1 U4439 ( .A1(n3468), .A2(n3495), .ZN(n3487) );
  NOR3_X1 U4440 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6526), .A3(n6701), 
        .ZN(n4568) );
  NAND2_X1 U4441 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4568), .ZN(n4582) );
  NAND2_X1 U4442 ( .A1(n6532), .A2(n4582), .ZN(n3470) );
  NAND3_X1 U4443 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4688) );
  INV_X1 U4444 ( .A(n4688), .ZN(n4473) );
  NAND2_X1 U4445 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4473), .ZN(n4507) );
  NAND2_X1 U4446 ( .A1(n3470), .A2(n4507), .ZN(n4961) );
  OAI22_X1 U4447 ( .A1(n4156), .A2(n4961), .B1(n3687), .B2(n6532), .ZN(n3471)
         );
  INV_X1 U4448 ( .A(n3471), .ZN(n3472) );
  NAND2_X1 U4449 ( .A1(n4463), .A2(n6786), .ZN(n3486) );
  AOI22_X1 U4450 ( .A1(n4019), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4451 ( .A1(n3097), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4452 ( .A1(n4132), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4453 ( .A1(n4135), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3475) );
  NAND4_X1 U4454 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3484)
         );
  AOI22_X1 U4455 ( .A1(n4134), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4456 ( .A1(n3115), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4457 ( .A1(n3093), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4458 ( .A1(n4094), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4459 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3483)
         );
  AOI22_X1 U4460 ( .A1(n3676), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3683), 
        .B2(n3491), .ZN(n3485) );
  NAND2_X1 U4461 ( .A1(n3487), .A2(n4566), .ZN(n3488) );
  NAND2_X1 U4462 ( .A1(n4521), .A2(n3655), .ZN(n3493) );
  NAND2_X1 U4463 ( .A1(n3515), .A2(n3516), .ZN(n3514) );
  NAND2_X1 U4464 ( .A1(n3514), .A2(n3497), .ZN(n3496) );
  NAND2_X1 U4465 ( .A1(n3496), .A2(n3491), .ZN(n3566) );
  OAI211_X1 U4466 ( .C1(n3491), .C2(n3496), .A(n3566), .B(n6668), .ZN(n3492)
         );
  INV_X1 U4467 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U4468 ( .A1(n4461), .A2(n3655), .ZN(n3500) );
  OAI21_X1 U4469 ( .B1(n3497), .B2(n3514), .A(n3496), .ZN(n3498) );
  AND2_X1 U4470 ( .A1(n3342), .A2(n3364), .ZN(n3506) );
  AOI21_X1 U4471 ( .B1(n3498), .B2(n6668), .A(n3506), .ZN(n3499) );
  NAND2_X1 U4472 ( .A1(n3500), .A2(n3499), .ZN(n6305) );
  INV_X1 U4473 ( .A(n3501), .ZN(n3503) );
  NAND2_X1 U4474 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  INV_X1 U4475 ( .A(n3655), .ZN(n3673) );
  INV_X1 U4476 ( .A(n6668), .ZN(n3517) );
  INV_X1 U4477 ( .A(n3506), .ZN(n3507) );
  OAI21_X1 U4478 ( .B1(n3517), .B2(n3516), .A(n3507), .ZN(n3508) );
  INV_X1 U4479 ( .A(n3508), .ZN(n3509) );
  OAI21_X2 U4480 ( .B1(n4957), .B2(n3673), .A(n3509), .ZN(n4511) );
  NAND2_X1 U4481 ( .A1(n4511), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3522)
         );
  XNOR2_X1 U4482 ( .A(n3522), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4388)
         );
  NAND2_X1 U4483 ( .A1(n4462), .A2(n3655), .ZN(n3521) );
  OAI21_X1 U4484 ( .B1(n3516), .B2(n3515), .A(n3514), .ZN(n3518) );
  OAI211_X1 U4485 ( .C1(n3518), .C2(n3517), .A(n3332), .B(n3299), .ZN(n3519)
         );
  INV_X1 U4486 ( .A(n3519), .ZN(n3520) );
  NAND2_X1 U4487 ( .A1(n3521), .A2(n3520), .ZN(n4387) );
  INV_X1 U4488 ( .A(n3522), .ZN(n4512) );
  NAND2_X1 U4489 ( .A1(n4512), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3523)
         );
  NAND2_X1 U4490 ( .A1(n6306), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3524)
         );
  NAND2_X1 U4491 ( .A1(n3525), .A2(n3524), .ZN(n4558) );
  NAND2_X1 U4492 ( .A1(n4557), .A2(n4558), .ZN(n3528) );
  NAND2_X1 U4493 ( .A1(n3526), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3527)
         );
  NAND2_X1 U4494 ( .A1(n3528), .A2(n3527), .ZN(n4596) );
  NAND2_X1 U4495 ( .A1(n3676), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4496 ( .A1(n4019), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4497 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4133), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4498 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3311), .B1(n5396), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4499 ( .A1(n4135), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4500 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3538)
         );
  AOI22_X1 U4501 ( .A1(n3111), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4502 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3115), .B1(n3095), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4503 ( .A1(n3093), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4504 ( .A1(n4094), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3533) );
  NAND4_X1 U4505 ( .A1(n3536), .A2(n3535), .A3(n3534), .A4(n3533), .ZN(n3537)
         );
  NAND2_X1 U4506 ( .A1(n3683), .A2(n3564), .ZN(n3539) );
  NAND2_X1 U4507 ( .A1(n3540), .A2(n3539), .ZN(n3547) );
  XNOR2_X1 U4508 ( .A(n3549), .B(n3547), .ZN(n3717) );
  NAND2_X1 U4509 ( .A1(n3717), .A2(n3655), .ZN(n3543) );
  XNOR2_X1 U4510 ( .A(n3566), .B(n3564), .ZN(n3541) );
  NAND2_X1 U4511 ( .A1(n3541), .A2(n6668), .ZN(n3542) );
  NAND2_X1 U4512 ( .A1(n3543), .A2(n3542), .ZN(n3544) );
  INV_X1 U4513 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U4514 ( .A1(n4596), .A2(n4597), .ZN(n3546) );
  NAND2_X1 U4515 ( .A1(n3544), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3545)
         );
  NAND2_X1 U4516 ( .A1(n3546), .A2(n3545), .ZN(n6295) );
  INV_X1 U4517 ( .A(n3547), .ZN(n3548) );
  NAND2_X1 U4518 ( .A1(n3676), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4519 ( .A1(n4019), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4520 ( .A1(n3097), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4521 ( .A1(n4132), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4522 ( .A1(n4135), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3550) );
  NAND4_X1 U4523 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(n3559)
         );
  AOI22_X1 U4524 ( .A1(n4134), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4525 ( .A1(n3115), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4526 ( .A1(n3093), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4527 ( .A1(n4094), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3554) );
  NAND4_X1 U4528 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3558)
         );
  NAND2_X1 U4529 ( .A1(n3683), .A2(n3567), .ZN(n3560) );
  NAND2_X1 U4530 ( .A1(n3561), .A2(n3560), .ZN(n3562) );
  NAND2_X1 U4531 ( .A1(n3563), .A2(n3562), .ZN(n3590) );
  INV_X1 U4532 ( .A(n3564), .ZN(n3565) );
  NOR2_X1 U4533 ( .A1(n3566), .A2(n3565), .ZN(n3568) );
  NAND2_X1 U4534 ( .A1(n3568), .A2(n3567), .ZN(n3601) );
  OAI211_X1 U4535 ( .C1(n3568), .C2(n3567), .A(n3601), .B(n6668), .ZN(n3569)
         );
  INV_X1 U4536 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U4537 ( .A1(n6295), .A2(n6294), .ZN(n3573) );
  NAND2_X1 U4538 ( .A1(n3571), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3572)
         );
  NAND2_X1 U4539 ( .A1(n3573), .A2(n3572), .ZN(n4942) );
  INV_X1 U4540 ( .A(n3590), .ZN(n3588) );
  NAND2_X1 U4541 ( .A1(n3676), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4542 ( .A1(n4019), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4543 ( .A1(n4133), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4544 ( .A1(n4132), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4545 ( .A1(n4135), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4546 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3584)
         );
  AOI22_X1 U4547 ( .A1(n3111), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4548 ( .A1(n3115), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3581) );
  INV_X1 U4549 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U4550 ( .A1(n3093), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4551 ( .A1(n4094), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4552 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3583)
         );
  NAND2_X1 U4553 ( .A1(n3683), .A2(n3602), .ZN(n3585) );
  INV_X1 U4554 ( .A(n3589), .ZN(n3587) );
  NAND2_X1 U4555 ( .A1(n3588), .A2(n3587), .ZN(n3600) );
  NAND2_X1 U4556 ( .A1(n3600), .A2(n3655), .ZN(n3610) );
  NAND2_X1 U4557 ( .A1(n3590), .A2(n3589), .ZN(n3737) );
  INV_X1 U4558 ( .A(n3737), .ZN(n3593) );
  XNOR2_X1 U4559 ( .A(n3601), .B(n3602), .ZN(n3591) );
  NAND2_X1 U4560 ( .A1(n3591), .A2(n6668), .ZN(n3592) );
  INV_X1 U4561 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4946) );
  XNOR2_X1 U4562 ( .A(n3594), .B(n4946), .ZN(n4943) );
  NAND2_X1 U4563 ( .A1(n4942), .A2(n4943), .ZN(n3596) );
  NAND2_X1 U4564 ( .A1(n3594), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3595)
         );
  NAND2_X1 U4565 ( .A1(n3596), .A2(n3595), .ZN(n5043) );
  NAND2_X1 U4566 ( .A1(n3683), .A2(n3612), .ZN(n3597) );
  OAI21_X1 U4567 ( .B1(n3598), .B2(n3419), .A(n3597), .ZN(n3599) );
  INV_X1 U4568 ( .A(n3743), .ZN(n3606) );
  INV_X1 U4569 ( .A(n3601), .ZN(n3603) );
  NAND2_X1 U4570 ( .A1(n3603), .A2(n3602), .ZN(n3611) );
  XNOR2_X1 U4571 ( .A(n3611), .B(n3612), .ZN(n3604) );
  NAND2_X1 U4572 ( .A1(n3604), .A2(n6668), .ZN(n3605) );
  OAI21_X2 U4573 ( .B1(n3606), .B2(n3673), .A(n3605), .ZN(n3607) );
  INV_X1 U4574 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U4575 ( .A1(n3607), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3608)
         );
  INV_X1 U4576 ( .A(n3611), .ZN(n3613) );
  NAND3_X1 U4577 ( .A1(n3613), .A2(n6668), .A3(n3612), .ZN(n3614) );
  NAND2_X1 U4578 ( .A1(n3619), .A2(n3614), .ZN(n3615) );
  XNOR2_X1 U4579 ( .A(n3615), .B(n6974), .ZN(n5067) );
  INV_X1 U4580 ( .A(n5154), .ZN(n3616) );
  INV_X2 U4581 ( .A(n3619), .ZN(n3617) );
  INV_X1 U4582 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U4583 ( .A1(n5892), .A2(n6360), .ZN(n3618) );
  INV_X1 U4584 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6349) );
  AND2_X1 U4585 ( .A1(n5892), .A2(n6349), .ZN(n5201) );
  NAND2_X1 U4586 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5200) );
  INV_X1 U4587 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U4588 ( .A1(n5892), .A2(n5215), .ZN(n5211) );
  NOR2_X1 U4589 ( .A1(n5892), .A2(n5215), .ZN(n5213) );
  NAND2_X1 U4590 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U4591 ( .A1(n5277), .A2(n5276), .ZN(n3621) );
  INV_X1 U4592 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4593 ( .A1(n5892), .A2(n3620), .ZN(n5275) );
  XNOR2_X1 U4594 ( .A(n5892), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5342)
         );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U4596 ( .A1(n5892), .A2(n5352), .ZN(n3622) );
  INV_X1 U4597 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U4598 ( .A1(n5892), .A2(n6860), .ZN(n3624) );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6818) );
  AND2_X1 U4600 ( .A1(n5892), .A2(n6818), .ZN(n5787) );
  NAND2_X1 U4601 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U4602 ( .A1(n5892), .A2(n5987), .ZN(n3626) );
  NAND2_X1 U4603 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4301) );
  INV_X1 U4604 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5887) );
  INV_X1 U4605 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5902) );
  NAND3_X1 U4606 ( .A1(n5887), .A2(n5902), .A3(n5987), .ZN(n3627) );
  NAND2_X1 U4607 ( .A1(n3617), .A2(n3627), .ZN(n3628) );
  AND2_X2 U4608 ( .A1(n4163), .A2(n3628), .ZN(n5771) );
  INV_X1 U4609 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3629) );
  NOR2_X1 U4610 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3630) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6693) );
  INV_X1 U4612 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4276) );
  INV_X1 U4613 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U4614 ( .A1(n3630), .A2(n6693), .A3(n4276), .A4(n4166), .ZN(n3631)
         );
  NAND2_X1 U4615 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U4616 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4313) );
  NOR2_X1 U4617 ( .A1(n5843), .A2(n4313), .ZN(n4337) );
  NAND2_X1 U4618 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5862) );
  INV_X1 U4619 ( .A(n5862), .ZN(n5742) );
  XNOR2_X1 U4620 ( .A(n5892), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5732)
         );
  NAND2_X1 U4621 ( .A1(n5892), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U4622 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5807) );
  INV_X1 U4623 ( .A(n3635), .ZN(n3634) );
  INV_X1 U4624 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5447) );
  AOI21_X1 U4625 ( .B1(n5434), .B2(n3634), .A(n5447), .ZN(n3636) );
  OAI22_X1 U4626 ( .A1(n3636), .A2(n5433), .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5434), .ZN(n4320) );
  NAND2_X1 U4627 ( .A1(n6701), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4628 ( .A1(n5462), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4629 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6799), .ZN(n3650) );
  INV_X1 U4630 ( .A(n3650), .ZN(n3640) );
  INV_X1 U4631 ( .A(n3638), .ZN(n3639) );
  NAND2_X1 U4632 ( .A1(n6526), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4633 ( .A1(n3379), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U4634 ( .A1(n3642), .A2(n3641), .ZN(n3664) );
  INV_X1 U4635 ( .A(n3672), .ZN(n3643) );
  AOI222_X1 U4636 ( .A1(n3645), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n3645), .B2(n6796), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n6796), 
        .ZN(n4179) );
  NAND2_X1 U4637 ( .A1(n3645), .A2(n6796), .ZN(n3646) );
  AOI22_X1 U4638 ( .A1(n3647), .A2(n3676), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6786), .ZN(n3681) );
  INV_X1 U4639 ( .A(n3647), .ZN(n4177) );
  NAND2_X1 U4640 ( .A1(n3683), .A2(n3489), .ZN(n3648) );
  NAND2_X1 U4641 ( .A1(n3648), .A2(n3299), .ZN(n3654) );
  INV_X1 U4642 ( .A(n3654), .ZN(n3660) );
  XNOR2_X1 U4643 ( .A(n3649), .B(n3650), .ZN(n4175) );
  NAND2_X1 U4644 ( .A1(n4175), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3658) );
  OAI21_X1 U4645 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6799), .A(n3650), 
        .ZN(n3652) );
  OAI21_X1 U4646 ( .B1(n3691), .B2(n3652), .A(n4490), .ZN(n3651) );
  NAND2_X1 U4647 ( .A1(n3651), .A2(n3668), .ZN(n3659) );
  NOR2_X1 U4648 ( .A1(n3667), .A2(n3652), .ZN(n3653) );
  OAI211_X1 U4649 ( .C1(n4175), .C2(n3654), .A(n3659), .B(n3653), .ZN(n3657)
         );
  INV_X1 U4650 ( .A(n3684), .ZN(n3656) );
  OAI211_X1 U4651 ( .C1(n3660), .C2(n3658), .A(n3657), .B(n3656), .ZN(n3663)
         );
  INV_X1 U4652 ( .A(n3659), .ZN(n3661) );
  NAND3_X1 U4653 ( .A1(n3661), .A2(n4175), .A3(n3660), .ZN(n3662) );
  NAND2_X1 U4654 ( .A1(n3663), .A2(n3662), .ZN(n3675) );
  INV_X1 U4655 ( .A(n3664), .ZN(n3665) );
  XNOR2_X1 U4656 ( .A(n3666), .B(n3665), .ZN(n4174) );
  INV_X1 U4657 ( .A(n4174), .ZN(n3670) );
  AOI211_X1 U4658 ( .C1(n3675), .C2(n3668), .A(n3670), .B(n3667), .ZN(n3678)
         );
  INV_X1 U4659 ( .A(n3668), .ZN(n3669) );
  AOI21_X1 U4660 ( .B1(n3676), .B2(n3670), .A(n3669), .ZN(n3674) );
  XNOR2_X1 U4661 ( .A(n3672), .B(n3671), .ZN(n4176) );
  OAI22_X1 U4662 ( .A1(n3675), .A2(n3674), .B1(n4176), .B2(n3673), .ZN(n3677)
         );
  OAI22_X1 U4663 ( .A1(n3678), .A2(n3677), .B1(n3676), .B2(n4176), .ZN(n3679)
         );
  AOI222_X1 U4664 ( .A1(n3681), .A2(n3680), .B1(n3681), .B2(n3679), .C1(n3680), 
        .C2(n3679), .ZN(n3682) );
  AOI21_X1 U4665 ( .B1(n3683), .B2(n4179), .A(n3682), .ZN(n3686) );
  NAND2_X1 U4666 ( .A1(n3310), .A2(n4678), .ZN(n3689) );
  AND2_X1 U4667 ( .A1(n5454), .A2(n3342), .ZN(n3690) );
  AND2_X1 U4668 ( .A1(n4194), .A2(n3691), .ZN(n6535) );
  NAND2_X1 U4669 ( .A1(n4320), .A2(n6320), .ZN(n4162) );
  NAND2_X1 U4670 ( .A1(n4461), .A2(n3901), .ZN(n3692) );
  NAND2_X1 U4671 ( .A1(n6455), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4672 ( .A1(n4462), .A2(n3901), .ZN(n3696) );
  AOI22_X1 U4673 ( .A1(n5418), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6455), .ZN(n3694) );
  NOR2_X1 U4674 ( .A1(n3344), .A2(n6455), .ZN(n3709) );
  NAND2_X1 U4675 ( .A1(n3709), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3693) );
  AND2_X1 U4676 ( .A1(n3694), .A2(n3693), .ZN(n3695) );
  NAND2_X1 U4677 ( .A1(n3696), .A2(n3695), .ZN(n4437) );
  AOI21_X1 U4678 ( .B1(n4957), .B2(n3697), .A(n6455), .ZN(n4436) );
  INV_X2 U4679 ( .A(n5416), .ZN(n4344) );
  INV_X1 U4680 ( .A(n3698), .ZN(n6516) );
  AOI22_X1 U4681 ( .A1(n3725), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6455), .ZN(n3700) );
  NAND2_X1 U4682 ( .A1(n3709), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4683 ( .A1(n3700), .A2(n3699), .ZN(n3701) );
  AOI21_X1 U4684 ( .B1(n6516), .B2(n3901), .A(n3701), .ZN(n4434) );
  NAND2_X1 U4685 ( .A1(n4437), .A2(n4438), .ZN(n3707) );
  NAND2_X1 U4686 ( .A1(n3709), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3706) );
  INV_X1 U4687 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4688 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3711) );
  OAI21_X1 U4689 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3711), .ZN(n6311) );
  NAND2_X1 U4690 ( .A1(n4344), .A2(n6311), .ZN(n3702) );
  OAI21_X1 U4691 ( .B1(n3703), .B2(n3824), .A(n3702), .ZN(n3704) );
  AOI21_X1 U4692 ( .B1(n5418), .B2(EAX_REG_2__SCAN_IN), .A(n3704), .ZN(n3705)
         );
  AND2_X1 U4693 ( .A1(n3706), .A2(n3705), .ZN(n4451) );
  NAND2_X1 U4694 ( .A1(n3707), .A2(n4451), .ZN(n3708) );
  INV_X1 U4695 ( .A(n3709), .ZN(n3720) );
  INV_X1 U4696 ( .A(n3711), .ZN(n3713) );
  INV_X1 U4697 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3710) );
  NOR2_X1 U4698 ( .A1(n3711), .A2(n3710), .ZN(n3726) );
  INV_X1 U4699 ( .A(n3726), .ZN(n3712) );
  OAI21_X1 U4700 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3713), .A(n3712), 
        .ZN(n5145) );
  AOI22_X1 U4701 ( .A1(n4344), .A2(n5145), .B1(n5425), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4702 ( .A1(n5418), .A2(EAX_REG_3__SCAN_IN), .ZN(n3714) );
  OAI211_X1 U4703 ( .C1(n3720), .C2(n4635), .A(n3715), .B(n3714), .ZN(n3716)
         );
  NAND2_X1 U4704 ( .A1(n3717), .A2(n3901), .ZN(n3723) );
  XNOR2_X1 U4705 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .B(n3726), .ZN(n6147) );
  INV_X1 U4706 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6944) );
  AOI21_X1 U4707 ( .B1(n6944), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3718) );
  AOI21_X1 U4708 ( .B1(n5418), .B2(EAX_REG_4__SCAN_IN), .A(n3718), .ZN(n3719)
         );
  OAI21_X1 U4709 ( .B1(n3720), .B2(n6796), .A(n3719), .ZN(n3721) );
  OAI21_X1 U4710 ( .B1(n5416), .B2(n6147), .A(n3721), .ZN(n3722) );
  NAND2_X1 U4711 ( .A1(n3723), .A2(n3722), .ZN(n4444) );
  NAND2_X1 U4712 ( .A1(n4443), .A2(n4444), .ZN(n4442) );
  INV_X1 U4713 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U4714 ( .A1(n3727), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3732)
         );
  OAI21_X1 U4715 ( .B1(n3727), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3732), 
        .ZN(n6297) );
  AOI22_X1 U4716 ( .A1(n6297), .A2(n4344), .B1(n5425), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3728) );
  OAI21_X1 U4717 ( .B1(n3928), .B2(n4812), .A(n3728), .ZN(n3729) );
  INV_X1 U4718 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4814) );
  AND2_X1 U4719 ( .A1(n3732), .A2(n6107), .ZN(n3733) );
  OR2_X1 U4720 ( .A1(n3733), .A2(n3739), .ZN(n6099) );
  NOR2_X1 U4721 ( .A1(n3824), .A2(n6107), .ZN(n3734) );
  AOI21_X1 U4722 ( .B1(n6099), .B2(n4344), .A(n3734), .ZN(n3735) );
  OAI21_X1 U4723 ( .B1(n3928), .B2(n4814), .A(n3735), .ZN(n3736) );
  AOI21_X1 U4724 ( .B1(n3737), .B2(n3901), .A(n3736), .ZN(n4783) );
  INV_X1 U4725 ( .A(n4783), .ZN(n3738) );
  INV_X1 U4726 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U4727 ( .A1(n3739), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3740)
         );
  OR2_X1 U4728 ( .A1(n3758), .A2(n3740), .ZN(n6287) );
  AOI22_X1 U4729 ( .A1(n6287), .A2(n4344), .B1(n5425), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3741) );
  OAI21_X1 U4730 ( .B1(n3928), .B2(n5000), .A(n3741), .ZN(n3742) );
  AOI22_X1 U4731 ( .A1(n4132), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4732 ( .A1(n4133), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4733 ( .A1(n3093), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4734 ( .A1(n4094), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3744) );
  NAND4_X1 U4735 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3753)
         );
  AOI22_X1 U4736 ( .A1(n4134), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4737 ( .A1(n5395), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4738 ( .A1(n3115), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4739 ( .A1(n4135), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4740 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  OAI21_X1 U4741 ( .B1(n3753), .B2(n3752), .A(n3901), .ZN(n3757) );
  NAND2_X1 U4742 ( .A1(n5418), .A2(EAX_REG_8__SCAN_IN), .ZN(n3756) );
  XNOR2_X1 U4743 ( .A(n3758), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U4744 ( .A1(n5159), .A2(n4344), .ZN(n3755) );
  NAND2_X1 U4745 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3754)
         );
  NAND4_X1 U4746 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n4936)
         );
  NAND2_X1 U4747 ( .A1(n4935), .A2(n4936), .ZN(n5059) );
  XNOR2_X1 U4748 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3773), .ZN(n6080) );
  AOI22_X1 U4749 ( .A1(n4094), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4750 ( .A1(n3097), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4751 ( .A1(n4132), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4752 ( .A1(n4134), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4753 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3768)
         );
  AOI22_X1 U4754 ( .A1(n4019), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4755 ( .A1(n5404), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4756 ( .A1(n3122), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4757 ( .A1(n4135), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4758 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3767)
         );
  OR2_X1 U4759 ( .A1(n3768), .A2(n3767), .ZN(n3769) );
  AOI22_X1 U4760 ( .A1(n3901), .A2(n3769), .B1(n5425), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4761 ( .A1(n5418), .A2(EAX_REG_9__SCAN_IN), .ZN(n3770) );
  OAI211_X1 U4762 ( .C1(n6080), .C2(n5416), .A(n3771), .B(n3770), .ZN(n5061)
         );
  INV_X1 U4763 ( .A(n5061), .ZN(n3772) );
  XNOR2_X1 U4764 ( .A(n3789), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5205)
         );
  AOI22_X1 U4765 ( .A1(n4132), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4766 ( .A1(n5404), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4767 ( .A1(n3115), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4768 ( .A1(n4094), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4769 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3783)
         );
  AOI22_X1 U4770 ( .A1(n3111), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4771 ( .A1(n3097), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4772 ( .A1(n4019), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4773 ( .A1(n4135), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4774 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3782)
         );
  OAI21_X1 U4775 ( .B1(n3783), .B2(n3782), .A(n3901), .ZN(n3786) );
  NAND2_X1 U4776 ( .A1(n5418), .A2(EAX_REG_10__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4777 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3784)
         );
  NAND3_X1 U4778 ( .A1(n3786), .A2(n3785), .A3(n3784), .ZN(n3787) );
  AOI21_X1 U4779 ( .B1(n5205), .B2(n4344), .A(n3787), .ZN(n5087) );
  NAND2_X1 U4780 ( .A1(n3789), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3804)
         );
  XNOR2_X1 U4781 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3804), .ZN(n6280)
         );
  AOI22_X1 U4782 ( .A1(n5404), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4783 ( .A1(n4132), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4784 ( .A1(n4135), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4785 ( .A1(n4094), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4786 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3799)
         );
  AOI22_X1 U4787 ( .A1(n3097), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4788 ( .A1(n4134), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4789 ( .A1(n3115), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4790 ( .A1(n4019), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4791 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3798)
         );
  OR2_X1 U4792 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  AOI22_X1 U4793 ( .A1(n3901), .A2(n3800), .B1(n5425), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3802) );
  NAND2_X1 U4794 ( .A1(n5418), .A2(EAX_REG_11__SCAN_IN), .ZN(n3801) );
  OAI211_X1 U4795 ( .C1(n6280), .C2(n5416), .A(n3802), .B(n3801), .ZN(n6064)
         );
  XNOR2_X1 U4796 ( .A(n3821), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5280)
         );
  NAND2_X1 U4797 ( .A1(n5280), .A2(n4344), .ZN(n3820) );
  AOI22_X1 U4798 ( .A1(n4094), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4799 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3311), .B1(n4019), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4800 ( .A1(n5404), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4801 ( .A1(n4135), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4802 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3815)
         );
  AOI22_X1 U4803 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n5395), .B1(n3097), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4804 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3574), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4805 ( .A1(n3111), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4806 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3122), .B1(n3113), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3810) );
  NAND4_X1 U4807 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  OAI21_X1 U4808 ( .B1(n3815), .B2(n3814), .A(n3901), .ZN(n3818) );
  NAND2_X1 U4809 ( .A1(n5418), .A2(EAX_REG_12__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4810 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3816)
         );
  AND3_X1 U4811 ( .A1(n3818), .A2(n3817), .A3(n3816), .ZN(n3819) );
  NAND2_X1 U4812 ( .A1(n3820), .A2(n3819), .ZN(n5188) );
  INV_X1 U4813 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3825) );
  OAI21_X1 U4814 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3822), .A(n3892), 
        .ZN(n6060) );
  NAND2_X1 U4815 ( .A1(n6060), .A2(n4344), .ZN(n3823) );
  OAI21_X1 U4816 ( .B1(n3825), .B2(n3824), .A(n3823), .ZN(n3826) );
  AOI21_X1 U4817 ( .B1(n5418), .B2(EAX_REG_13__SCAN_IN), .A(n3826), .ZN(n3829)
         );
  INV_X1 U4818 ( .A(n3829), .ZN(n3827) );
  AOI22_X1 U4819 ( .A1(n3111), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4820 ( .A1(n4094), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4821 ( .A1(n4019), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4822 ( .A1(n4132), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4823 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3840)
         );
  AOI22_X1 U4824 ( .A1(n3097), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4825 ( .A1(n3093), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4826 ( .A1(n3122), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4827 ( .A1(n4135), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4828 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  OR2_X1 U4829 ( .A1(n3840), .A2(n3839), .ZN(n3841) );
  AND2_X1 U4830 ( .A1(n3901), .A2(n3841), .ZN(n5272) );
  NAND2_X1 U4831 ( .A1(n5273), .A2(n5272), .ZN(n5271) );
  NAND2_X1 U4832 ( .A1(n5420), .A2(n5416), .ZN(n3982) );
  NAND2_X1 U4833 ( .A1(n5395), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3844)
         );
  NAND2_X1 U4834 ( .A1(n3115), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3843) );
  AND3_X1 U4835 ( .A1(n3844), .A2(n3843), .A3(n5416), .ZN(n3848) );
  AOI22_X1 U4836 ( .A1(n4094), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4135), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4837 ( .A1(n3111), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4838 ( .A1(n3118), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4839 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3854)
         );
  AOI22_X1 U4840 ( .A1(n5404), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4841 ( .A1(n3097), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4842 ( .A1(n3311), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4843 ( .A1(n5396), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4844 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3853)
         );
  OR2_X1 U4845 ( .A1(n3854), .A2(n3853), .ZN(n3855) );
  NAND2_X1 U4846 ( .A1(n3982), .A2(n3855), .ZN(n3859) );
  AOI22_X1 U4847 ( .A1(n3725), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6455), .ZN(n3858) );
  INV_X1 U4848 ( .A(n3891), .ZN(n3856) );
  NAND2_X1 U4849 ( .A1(n3874), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3911)
         );
  XNOR2_X1 U4850 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n3911), .ZN(n6033)
         );
  AND2_X1 U4851 ( .A1(n6033), .A2(n4344), .ZN(n3857) );
  AOI21_X1 U4852 ( .B1(n3859), .B2(n3858), .A(n3857), .ZN(n5971) );
  AOI22_X1 U4853 ( .A1(n5404), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4854 ( .A1(n4019), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4855 ( .A1(n3097), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4856 ( .A1(n3095), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4857 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3869)
         );
  AOI22_X1 U4858 ( .A1(n3311), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4859 ( .A1(n4094), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4135), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4860 ( .A1(n4134), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4861 ( .A1(n3120), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3864) );
  NAND4_X1 U4862 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3868)
         );
  OR2_X1 U4863 ( .A1(n3869), .A2(n3868), .ZN(n3873) );
  INV_X1 U4864 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3871) );
  XOR2_X1 U4865 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3874), .Z(n5594) );
  INV_X1 U4866 ( .A(n5594), .ZN(n5783) );
  AOI22_X1 U4867 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n4344), 
        .B2(n5783), .ZN(n3870) );
  OAI21_X1 U4868 ( .B1(n3928), .B2(n3871), .A(n3870), .ZN(n3872) );
  AOI21_X1 U4869 ( .B1(n4146), .B2(n3873), .A(n3872), .ZN(n5592) );
  OR2_X1 U4870 ( .A1(n3891), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3876)
         );
  INV_X1 U4871 ( .A(n3874), .ZN(n3875) );
  NAND2_X1 U4872 ( .A1(n3876), .A2(n3875), .ZN(n5792) );
  AOI22_X1 U4873 ( .A1(n3097), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4874 ( .A1(n3115), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4875 ( .A1(n3095), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4876 ( .A1(n4135), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4877 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3886)
         );
  AOI22_X1 U4878 ( .A1(n3111), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4879 ( .A1(n4132), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4880 ( .A1(n5395), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4881 ( .A1(n4094), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4882 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3885)
         );
  OAI21_X1 U4883 ( .B1(n3886), .B2(n3885), .A(n3901), .ZN(n3889) );
  NAND2_X1 U4884 ( .A1(n5418), .A2(EAX_REG_15__SCAN_IN), .ZN(n3888) );
  NAND2_X1 U4885 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3887)
         );
  NAND3_X1 U4886 ( .A1(n3889), .A2(n3888), .A3(n3887), .ZN(n3890) );
  AOI21_X1 U4887 ( .B1(n5792), .B2(n4344), .A(n3890), .ZN(n5607) );
  NOR2_X1 U4888 ( .A1(n5592), .A2(n5607), .ZN(n5590) );
  AND2_X1 U4889 ( .A1(n5971), .A2(n5590), .ZN(n3909) );
  AOI21_X1 U4890 ( .B1(n6814), .B2(n3892), .A(n3891), .ZN(n6045) );
  OR2_X1 U4891 ( .A1(n6045), .A2(n5416), .ZN(n3908) );
  AOI22_X1 U4892 ( .A1(n4019), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4893 ( .A1(n5404), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4894 ( .A1(n3122), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4895 ( .A1(n4135), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4896 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3903)
         );
  AOI22_X1 U4897 ( .A1(n4094), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4898 ( .A1(n4133), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4899 ( .A1(n4132), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4900 ( .A1(n4134), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4901 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3902)
         );
  OAI21_X1 U4902 ( .B1(n3903), .B2(n3902), .A(n3901), .ZN(n3906) );
  NAND2_X1 U4903 ( .A1(n3725), .A2(EAX_REG_14__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U4904 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3904)
         );
  AND3_X1 U4905 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(n3907) );
  NAND2_X1 U4906 ( .A1(n3908), .A2(n3907), .ZN(n5665) );
  AND2_X1 U4907 ( .A1(n3909), .A2(n5665), .ZN(n3910) );
  INV_X1 U4908 ( .A(n3948), .ZN(n3914) );
  OR2_X1 U4909 ( .A1(n3912), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3913)
         );
  NAND2_X1 U4910 ( .A1(n3914), .A2(n3913), .ZN(n5969) );
  AOI22_X1 U4911 ( .A1(n4094), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4912 ( .A1(n3097), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4913 ( .A1(n5404), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4914 ( .A1(n4135), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4915 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3924)
         );
  AOI22_X1 U4916 ( .A1(n3311), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4917 ( .A1(n5395), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4918 ( .A1(n3111), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4919 ( .A1(n3115), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3919) );
  NAND4_X1 U4920 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3923)
         );
  NOR2_X1 U4921 ( .A1(n3924), .A2(n3923), .ZN(n3925) );
  NOR2_X1 U4922 ( .A1(n5420), .A2(n3925), .ZN(n3930) );
  INV_X1 U4923 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4924 ( .A1(n6455), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3926)
         );
  OAI211_X1 U4925 ( .C1(n3928), .C2(n3927), .A(n5416), .B(n3926), .ZN(n3929)
         );
  OAI22_X1 U4926 ( .A1(n5969), .A2(n5416), .B1(n3930), .B2(n3929), .ZN(n5578)
         );
  INV_X1 U4927 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3931) );
  XNOR2_X1 U4928 ( .A(n3948), .B(n3931), .ZN(n5774) );
  NAND2_X1 U4929 ( .A1(n5774), .A2(n4344), .ZN(n3947) );
  AOI22_X1 U4930 ( .A1(n4094), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3097), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4931 ( .A1(n3115), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4932 ( .A1(n5404), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4933 ( .A1(n4019), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4934 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3943)
         );
  AOI22_X1 U4935 ( .A1(n3122), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4936 ( .A1(n5395), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3937)
         );
  NAND2_X1 U4937 ( .A1(n3111), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3936) );
  AND3_X1 U4938 ( .A1(n3937), .A2(n3936), .A3(n5416), .ZN(n3940) );
  AOI22_X1 U4939 ( .A1(n4135), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4940 ( .A1(n3120), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4941 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3942)
         );
  OAI21_X1 U4942 ( .B1(n3943), .B2(n3942), .A(n3982), .ZN(n3945) );
  AOI22_X1 U4943 ( .A1(n3725), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6455), .ZN(n3944) );
  NAND2_X1 U4944 ( .A1(n3945), .A2(n3944), .ZN(n3946) );
  NAND2_X1 U4945 ( .A1(n3947), .A2(n3946), .ZN(n5563) );
  INV_X1 U4946 ( .A(n3951), .ZN(n3950) );
  INV_X1 U4947 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3949) );
  NAND2_X1 U4948 ( .A1(n3950), .A2(n3949), .ZN(n3952) );
  AND2_X1 U4949 ( .A1(n3952), .A2(n4000), .ZN(n5946) );
  AOI22_X1 U4950 ( .A1(n5404), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4951 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5395), .B1(n4019), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4952 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3095), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4953 ( .A1(n4094), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4954 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3962)
         );
  AOI22_X1 U4955 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3311), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4956 ( .A1(n3097), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4957 ( .A1(n3111), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4958 ( .A1(n4135), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4959 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3961)
         );
  OR2_X1 U4960 ( .A1(n3962), .A2(n3961), .ZN(n3966) );
  INV_X1 U4961 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3964) );
  NAND2_X1 U4962 ( .A1(n6455), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3963)
         );
  OAI211_X1 U4963 ( .C1(n3928), .C2(n3964), .A(n5416), .B(n3963), .ZN(n3965)
         );
  AOI21_X1 U4964 ( .B1(n4146), .B2(n3966), .A(n3965), .ZN(n3967) );
  AOI21_X1 U4965 ( .B1(n5946), .B2(n4344), .A(n3967), .ZN(n5649) );
  AOI21_X1 U4966 ( .B1(n3120), .B2(INSTQUEUE_REG_6__5__SCAN_IN), .A(n4344), 
        .ZN(n3970) );
  NAND2_X1 U4967 ( .A1(n3097), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3969)
         );
  AND2_X1 U4968 ( .A1(n3970), .A2(n3969), .ZN(n3974) );
  AOI22_X1 U4969 ( .A1(n3115), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4970 ( .A1(n5404), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4971 ( .A1(n4019), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4972 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4973 ( .A1(n3311), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4974 ( .A1(n3317), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4135), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4975 ( .A1(n3111), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4976 ( .A1(n4094), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4977 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  OR2_X1 U4978 ( .A1(n3980), .A2(n3979), .ZN(n3981) );
  NAND2_X1 U4979 ( .A1(n3982), .A2(n3981), .ZN(n3985) );
  AOI22_X1 U4980 ( .A1(n3725), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6455), .ZN(n3984) );
  XNOR2_X1 U4981 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4000), .ZN(n5936)
         );
  AND2_X1 U4982 ( .A1(n5936), .A2(n4344), .ZN(n3983) );
  AOI21_X1 U4983 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n5643) );
  AOI22_X1 U4984 ( .A1(n3097), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4985 ( .A1(n3311), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4986 ( .A1(n5404), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4987 ( .A1(n3574), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U4988 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3995)
         );
  AOI22_X1 U4989 ( .A1(n3115), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4990 ( .A1(n4019), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4135), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4991 ( .A1(n3111), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4992 ( .A1(n4094), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U4993 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3994)
         );
  NOR2_X1 U4994 ( .A1(n3995), .A2(n3994), .ZN(n3999) );
  NAND2_X1 U4995 ( .A1(n6455), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3996)
         );
  NAND2_X1 U4996 ( .A1(n5416), .A2(n3996), .ZN(n3997) );
  AOI21_X1 U4997 ( .B1(n5418), .B2(EAX_REG_22__SCAN_IN), .A(n3997), .ZN(n3998)
         );
  OAI21_X1 U4998 ( .B1(n5420), .B2(n3999), .A(n3998), .ZN(n4008) );
  INV_X1 U4999 ( .A(n4050), .ZN(n4006) );
  INV_X1 U5000 ( .A(n4002), .ZN(n4004) );
  INV_X1 U5001 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4003) );
  NAND2_X1 U5002 ( .A1(n4004), .A2(n4003), .ZN(n4005) );
  NAND2_X1 U5003 ( .A1(n4006), .A2(n4005), .ZN(n5921) );
  OR2_X1 U5004 ( .A1(n5921), .A2(n5416), .ZN(n4007) );
  NAND2_X1 U5005 ( .A1(n4008), .A2(n4007), .ZN(n5638) );
  AOI22_X1 U5006 ( .A1(n3097), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U5007 ( .A1(n5397), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U5008 ( .A1(n3095), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5009 ( .A1(n4135), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U5010 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4018)
         );
  AOI22_X1 U5011 ( .A1(n3111), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5012 ( .A1(n4132), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5013 ( .A1(n3115), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5014 ( .A1(n4094), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4013) );
  NAND4_X1 U5015 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4017)
         );
  NOR2_X1 U5016 ( .A1(n4018), .A2(n4017), .ZN(n4038) );
  AOI22_X1 U5017 ( .A1(n4094), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5018 ( .A1(n4135), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5019 ( .A1(n4132), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5020 ( .A1(n5395), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U5021 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4029)
         );
  AOI22_X1 U5022 ( .A1(n3111), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5023 ( .A1(n3115), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5024 ( .A1(n3122), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5025 ( .A1(n4133), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4024) );
  NAND4_X1 U5026 ( .A1(n4027), .A2(n4026), .A3(n4025), .A4(n4024), .ZN(n4028)
         );
  NOR2_X1 U5027 ( .A1(n4029), .A2(n4028), .ZN(n4037) );
  XOR2_X1 U5028 ( .A(n4038), .B(n4037), .Z(n4030) );
  NAND2_X1 U5029 ( .A1(n4030), .A2(n4146), .ZN(n4033) );
  INV_X1 U5030 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5749) );
  OAI21_X1 U5031 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5749), .A(n5416), .ZN(
        n4031) );
  AOI21_X1 U5032 ( .B1(n5418), .B2(EAX_REG_23__SCAN_IN), .A(n4031), .ZN(n4032)
         );
  NAND2_X1 U5033 ( .A1(n4033), .A2(n4032), .ZN(n4035) );
  XNOR2_X1 U5034 ( .A(n4050), .B(n5749), .ZN(n5747) );
  NAND2_X1 U5035 ( .A1(n5747), .A2(n4344), .ZN(n4034) );
  NAND2_X1 U5036 ( .A1(n4035), .A2(n4034), .ZN(n5551) );
  NOR2_X1 U5037 ( .A1(n4038), .A2(n4037), .ZN(n4066) );
  AOI22_X1 U5038 ( .A1(n4019), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5039 ( .A1(n4133), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5040 ( .A1(n4132), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5041 ( .A1(n4135), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U5042 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4048)
         );
  AOI22_X1 U5043 ( .A1(n4134), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5044 ( .A1(n3115), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5045 ( .A1(n3093), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5046 ( .A1(n4094), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4043) );
  NAND4_X1 U5047 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(n4047)
         );
  INV_X1 U5048 ( .A(n4065), .ZN(n4049) );
  XNOR2_X1 U5049 ( .A(n4066), .B(n4049), .ZN(n4054) );
  XNOR2_X1 U5050 ( .A(n4069), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5913)
         );
  NAND2_X1 U5051 ( .A1(n3725), .A2(EAX_REG_24__SCAN_IN), .ZN(n4052) );
  NAND2_X1 U5052 ( .A1(n5425), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4051)
         );
  OAI211_X1 U5053 ( .C1(n5913), .C2(n5416), .A(n4052), .B(n4051), .ZN(n4053)
         );
  AOI21_X1 U5054 ( .B1(n4054), .B2(n4146), .A(n4053), .ZN(n5625) );
  AOI22_X1 U5055 ( .A1(n4134), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5056 ( .A1(n3115), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5057 ( .A1(n3093), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5058 ( .A1(n4094), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U5059 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4064)
         );
  AOI22_X1 U5060 ( .A1(n5397), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5061 ( .A1(n3097), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5062 ( .A1(n3311), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5063 ( .A1(n4135), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5064 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  NOR2_X1 U5065 ( .A1(n4064), .A2(n4063), .ZN(n4074) );
  NAND2_X1 U5066 ( .A1(n4066), .A2(n4065), .ZN(n4073) );
  XOR2_X1 U5067 ( .A(n4074), .B(n4073), .Z(n4067) );
  NAND2_X1 U5068 ( .A1(n4067), .A2(n4146), .ZN(n4072) );
  INV_X1 U5069 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5729) );
  AOI21_X1 U5070 ( .B1(n5729), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4068) );
  AOI21_X1 U5071 ( .B1(n5418), .B2(EAX_REG_25__SCAN_IN), .A(n4068), .ZN(n4071)
         );
  XNOR2_X1 U5072 ( .A(n4088), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5731)
         );
  AOI22_X1 U5073 ( .A1(n4072), .A2(n4071), .B1(n4344), .B2(n5731), .ZN(n5537)
         );
  NAND2_X1 U5074 ( .A1(n5535), .A2(n5537), .ZN(n5526) );
  NOR2_X1 U5075 ( .A1(n4074), .A2(n4073), .ZN(n4093) );
  AOI22_X1 U5076 ( .A1(n4019), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5077 ( .A1(n4133), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5078 ( .A1(n4132), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5079 ( .A1(n4135), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5080 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4084)
         );
  AOI22_X1 U5081 ( .A1(n3111), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5082 ( .A1(n3115), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5083 ( .A1(n3093), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5084 ( .A1(n4094), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U5085 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4083)
         );
  OR2_X1 U5086 ( .A1(n4084), .A2(n4083), .ZN(n4092) );
  XNOR2_X1 U5087 ( .A(n4093), .B(n4092), .ZN(n4085) );
  NOR2_X1 U5088 ( .A1(n4085), .A2(n5420), .ZN(n4091) );
  INV_X1 U5089 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6228) );
  NOR2_X1 U5090 ( .A1(n6941), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4086)
         );
  OAI22_X1 U5091 ( .A1(n3928), .A2(n6228), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4086), .ZN(n4090) );
  INV_X1 U5092 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6863) );
  OAI21_X1 U5093 ( .B1(n4088), .B2(n5729), .A(n6863), .ZN(n4089) );
  NAND2_X1 U5094 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U5095 ( .A1(n4089), .A2(n4108), .ZN(n5725) );
  OAI22_X1 U5096 ( .A1(n4091), .A2(n4090), .B1(n5416), .B2(n5725), .ZN(n5527)
         );
  NOR2_X2 U5097 ( .A1(n5526), .A2(n5527), .ZN(n5509) );
  NAND2_X1 U5098 ( .A1(n4093), .A2(n4092), .ZN(n4114) );
  AOI22_X1 U5099 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3311), .B1(n3317), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5100 ( .A1(n4019), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4135), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5101 ( .A1(n3115), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5102 ( .A1(n4094), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4095) );
  NAND4_X1 U5103 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4104)
         );
  AOI22_X1 U5104 ( .A1(n4134), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5105 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3096), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5106 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3122), .B1(n3395), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5107 ( .A1(n3574), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5108 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4103)
         );
  NOR2_X1 U5109 ( .A1(n4104), .A2(n4103), .ZN(n4115) );
  XOR2_X1 U5110 ( .A(n4114), .B(n4115), .Z(n4105) );
  NAND2_X1 U5111 ( .A1(n4105), .A2(n4146), .ZN(n4111) );
  INV_X1 U5112 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6862) );
  NOR2_X1 U5113 ( .A1(n6862), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4106) );
  AOI211_X1 U5114 ( .C1(n5418), .C2(EAX_REG_27__SCAN_IN), .A(n4344), .B(n4106), 
        .ZN(n4110) );
  NAND2_X1 U5115 ( .A1(n4108), .A2(n6862), .ZN(n4109) );
  AND2_X1 U5116 ( .A1(n4112), .A2(n4109), .ZN(n5716) );
  AOI22_X1 U5117 ( .A1(n4111), .A2(n4110), .B1(n4344), .B2(n5716), .ZN(n5510)
         );
  NAND2_X1 U5118 ( .A1(n4112), .A2(n6688), .ZN(n4113) );
  NAND2_X1 U5119 ( .A1(n4348), .A2(n4113), .ZN(n5705) );
  NOR2_X1 U5120 ( .A1(n4115), .A2(n4114), .ZN(n4131) );
  AOI22_X1 U5121 ( .A1(n5397), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5122 ( .A1(n3097), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5123 ( .A1(n4132), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5124 ( .A1(n4135), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4116) );
  NAND4_X1 U5125 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4125)
         );
  AOI22_X1 U5126 ( .A1(n3111), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5404), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5127 ( .A1(n3115), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5128 ( .A1(n3093), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5129 ( .A1(n4094), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4120) );
  NAND4_X1 U5130 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4124)
         );
  OR2_X1 U5131 ( .A1(n4125), .A2(n4124), .ZN(n4130) );
  XNOR2_X1 U5132 ( .A(n4131), .B(n4130), .ZN(n4128) );
  NOR2_X1 U5133 ( .A1(n6688), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4126) );
  AOI211_X1 U5134 ( .C1(n5418), .C2(EAX_REG_28__SCAN_IN), .A(n4344), .B(n4126), 
        .ZN(n4127) );
  OAI21_X1 U5135 ( .B1(n4128), .B2(n5420), .A(n4127), .ZN(n4129) );
  OAI21_X1 U5136 ( .B1(n5416), .B2(n5705), .A(n4129), .ZN(n5500) );
  NAND2_X1 U5137 ( .A1(n4131), .A2(n4130), .ZN(n5411) );
  AOI22_X1 U5138 ( .A1(n4132), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5397), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5139 ( .A1(n3097), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5140 ( .A1(n4134), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5141 ( .A1(n4135), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4136) );
  NAND4_X1 U5142 ( .A1(n4139), .A2(n4138), .A3(n4137), .A4(n4136), .ZN(n4145)
         );
  AOI22_X1 U5143 ( .A1(n3115), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5144 ( .A1(n3317), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5145 ( .A1(n5404), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5146 ( .A1(n4094), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4140) );
  NAND4_X1 U5147 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4144)
         );
  NOR2_X1 U5148 ( .A1(n4145), .A2(n4144), .ZN(n5412) );
  XOR2_X1 U5149 ( .A(n5411), .B(n5412), .Z(n4147) );
  NAND2_X1 U5150 ( .A1(n4147), .A2(n4146), .ZN(n4150) );
  INV_X1 U5151 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4157) );
  NOR2_X1 U5152 ( .A1(n4157), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4148) );
  AOI211_X1 U5153 ( .C1(n5418), .C2(EAX_REG_29__SCAN_IN), .A(n4344), .B(n4148), 
        .ZN(n4149) );
  XNOR2_X1 U5154 ( .A(n4348), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4371)
         );
  AOI22_X1 U5155 ( .A1(n4150), .A2(n4149), .B1(n4344), .B2(n4371), .ZN(n4152)
         );
  NAND2_X1 U5156 ( .A1(n4345), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6562) );
  NAND2_X1 U5157 ( .A1(n6452), .A2(n4156), .ZN(n6664) );
  NAND2_X1 U5158 ( .A1(n6664), .A2(n6786), .ZN(n4153) );
  NAND2_X1 U5159 ( .A1(n6786), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5160 ( .A1(n6941), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5161 ( .A1(n4155), .A2(n4154), .ZN(n6321) );
  NAND2_X1 U5162 ( .A1(n6375), .A2(REIP_REG_29__SCAN_IN), .ZN(n4335) );
  OAI21_X1 U5163 ( .B1(n6304), .B2(n4157), .A(n4335), .ZN(n4158) );
  AOI21_X1 U5164 ( .B1(n6298), .B2(n4371), .A(n4158), .ZN(n4159) );
  NAND2_X1 U5165 ( .A1(n4162), .A2(n4161), .ZN(U2957) );
  NAND2_X1 U5166 ( .A1(n5772), .A2(n3617), .ZN(n4165) );
  OR2_X1 U5167 ( .A1(n4163), .A2(n3629), .ZN(n4164) );
  NAND2_X1 U5168 ( .A1(n4165), .A2(n4164), .ZN(n5765) );
  XNOR2_X1 U5169 ( .A(n5892), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5766)
         );
  NOR2_X1 U5170 ( .A1(n5892), .A2(n4166), .ZN(n4167) );
  XNOR2_X1 U5171 ( .A(n5892), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5761)
         );
  NOR2_X1 U5172 ( .A1(n5892), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5753)
         );
  NAND2_X1 U5173 ( .A1(n3101), .A2(n5753), .ZN(n5744) );
  OAI21_X1 U5174 ( .B1(n3617), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5759), 
        .ZN(n5755) );
  NAND3_X1 U5175 ( .A1(n5892), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4168) );
  XNOR2_X1 U5176 ( .A(n4169), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5741)
         );
  INV_X1 U5177 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6573) );
  NAND3_X1 U5178 ( .A1(n4170), .A2(n4354), .A3(n6666), .ZN(n4172) );
  NAND3_X1 U5179 ( .A1(n4172), .A2(n4490), .A3(n3344), .ZN(n4173) );
  NAND2_X1 U5180 ( .A1(n4622), .A2(n4173), .ZN(n4183) );
  NAND2_X1 U5181 ( .A1(n3489), .A2(n6671), .ZN(n4181) );
  AND3_X1 U5182 ( .A1(n4176), .A2(n4175), .A3(n4174), .ZN(n4178) );
  OAI21_X1 U5183 ( .B1(n4179), .B2(n4178), .A(n4177), .ZN(n4405) );
  INV_X1 U5184 ( .A(n4405), .ZN(n4180) );
  NOR2_X1 U5185 ( .A1(n4180), .A2(READY_N), .ZN(n4614) );
  NAND2_X1 U5186 ( .A1(n4181), .A2(n4614), .ZN(n4182) );
  MUX2_X1 U5187 ( .A(n4183), .B(n4182), .S(n3346), .Z(n4192) );
  INV_X1 U5188 ( .A(n4622), .ZN(n4185) );
  INV_X1 U5189 ( .A(n5454), .ZN(n6514) );
  NAND2_X1 U5190 ( .A1(n6514), .A2(n3489), .ZN(n4287) );
  INV_X1 U5191 ( .A(n4287), .ZN(n4184) );
  NAND2_X1 U5192 ( .A1(n4185), .A2(n4184), .ZN(n4626) );
  INV_X1 U5193 ( .A(n3368), .ZN(n4186) );
  NAND2_X1 U5194 ( .A1(n4186), .A2(n6668), .ZN(n4187) );
  AND2_X1 U5195 ( .A1(n4188), .A2(n4187), .ZN(n4294) );
  NAND2_X1 U5196 ( .A1(n4194), .A2(n4294), .ZN(n4190) );
  INV_X1 U5197 ( .A(n4189), .ZN(n4404) );
  NAND2_X1 U5198 ( .A1(n4190), .A2(n4404), .ZN(n4286) );
  AND2_X1 U5199 ( .A1(n4194), .A2(n4673), .ZN(n4613) );
  INV_X1 U5200 ( .A(n4613), .ZN(n4604) );
  INV_X1 U5201 ( .A(n6535), .ZN(n4198) );
  INV_X1 U5202 ( .A(n4282), .ZN(n4195) );
  AOI22_X1 U5203 ( .A1(n4195), .A2(n3310), .B1(n4170), .B2(n4382), .ZN(n4197)
         );
  NAND4_X1 U5204 ( .A1(n4604), .A2(n4198), .A3(n4197), .A4(n6003), .ZN(n4199)
         );
  INV_X2 U5205 ( .A(n4382), .ZN(n4430) );
  NAND2_X1 U5206 ( .A1(n4200), .A2(n4490), .ZN(n4219) );
  NAND2_X1 U5207 ( .A1(n4219), .A2(n6836), .ZN(n4202) );
  OAI211_X1 U5208 ( .C1(n4430), .C2(EBX_REG_1__SCAN_IN), .A(n4202), .B(n4226), 
        .ZN(n4205) );
  INV_X1 U5209 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4203) );
  NAND2_X1 U5210 ( .A1(n5652), .A2(n4203), .ZN(n4204) );
  NAND2_X1 U5211 ( .A1(n4205), .A2(n4204), .ZN(n4209) );
  NAND2_X1 U5212 ( .A1(n4219), .A2(EBX_REG_0__SCAN_IN), .ZN(n4207) );
  INV_X1 U5213 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5214 ( .A1(n4226), .A2(n5080), .ZN(n4206) );
  NAND2_X1 U5215 ( .A1(n4207), .A2(n4206), .ZN(n4208) );
  XNOR2_X1 U5216 ( .A(n4209), .B(n4208), .ZN(n4383) );
  NAND2_X1 U5217 ( .A1(n4383), .A2(n4382), .ZN(n4385) );
  INV_X1 U5218 ( .A(n4208), .ZN(n4432) );
  OR2_X1 U5219 ( .A1(n4209), .A2(n4432), .ZN(n4210) );
  NAND2_X1 U5220 ( .A1(n4385), .A2(n4210), .ZN(n4457) );
  INV_X1 U5221 ( .A(n4457), .ZN(n4214) );
  MUX2_X1 U5222 ( .A(n5384), .B(n4219), .S(EBX_REG_2__SCAN_IN), .Z(n4212) );
  NAND2_X1 U5223 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4211)
         );
  AND2_X1 U5224 ( .A1(n4212), .A2(n4211), .ZN(n4456) );
  OR2_X1 U5225 ( .A1(n4332), .A2(EBX_REG_3__SCAN_IN), .ZN(n4217) );
  NAND2_X1 U5226 ( .A1(n5384), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4215)
         );
  OAI211_X1 U5227 ( .C1(n4430), .C2(EBX_REG_3__SCAN_IN), .A(n4219), .B(n4215), 
        .ZN(n4216) );
  NAND2_X1 U5228 ( .A1(n4217), .A2(n4216), .ZN(n4755) );
  NAND2_X1 U5229 ( .A1(n4219), .A2(n4218), .ZN(n4220) );
  OAI211_X1 U5230 ( .C1(n4430), .C2(EBX_REG_4__SCAN_IN), .A(n4220), .B(n4226), 
        .ZN(n4223) );
  INV_X1 U5231 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4221) );
  NAND2_X1 U5232 ( .A1(n5652), .A2(n4221), .ZN(n4222) );
  AND2_X1 U5233 ( .A1(n4223), .A2(n4222), .ZN(n4446) );
  MUX2_X1 U5234 ( .A(n4332), .B(n4226), .S(EBX_REG_5__SCAN_IN), .Z(n4225) );
  OR2_X1 U5235 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4224)
         );
  AND2_X1 U5236 ( .A1(n4225), .A2(n4224), .ZN(n6108) );
  NAND2_X1 U5237 ( .A1(n4219), .A2(n4946), .ZN(n4227) );
  OAI211_X1 U5238 ( .C1(n4430), .C2(EBX_REG_6__SCAN_IN), .A(n4227), .B(n5384), 
        .ZN(n4229) );
  INV_X1 U5239 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U5240 ( .A1(n5652), .A2(n6731), .ZN(n4228) );
  MUX2_X1 U5241 ( .A(n4332), .B(n5384), .S(EBX_REG_7__SCAN_IN), .Z(n4231) );
  OR2_X1 U5242 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4230)
         );
  NAND2_X1 U5243 ( .A1(n4231), .A2(n4230), .ZN(n5048) );
  NAND2_X1 U5244 ( .A1(n4219), .A2(n6974), .ZN(n4232) );
  OAI211_X1 U5245 ( .C1(n4430), .C2(EBX_REG_8__SCAN_IN), .A(n4232), .B(n5384), 
        .ZN(n4235) );
  INV_X1 U5246 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4233) );
  NAND2_X1 U5247 ( .A1(n5652), .A2(n4233), .ZN(n4234) );
  NAND2_X1 U5248 ( .A1(n4235), .A2(n4234), .ZN(n4937) );
  OR2_X1 U5249 ( .A1(n4332), .A2(EBX_REG_9__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U5250 ( .A1(n5384), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4236)
         );
  OAI211_X1 U5251 ( .C1(n4430), .C2(EBX_REG_9__SCAN_IN), .A(n4219), .B(n4236), 
        .ZN(n4237) );
  AND2_X1 U5252 ( .A1(n4238), .A2(n4237), .ZN(n6071) );
  MUX2_X1 U5253 ( .A(n5384), .B(n4219), .S(EBX_REG_10__SCAN_IN), .Z(n4240) );
  NAND2_X1 U5254 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4239) );
  NAND2_X1 U5255 ( .A1(n4240), .A2(n4239), .ZN(n5093) );
  INV_X1 U5256 ( .A(n5093), .ZN(n4241) );
  OR2_X1 U5257 ( .A1(n4332), .A2(EBX_REG_11__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U5258 ( .A1(n5384), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4242) );
  OAI211_X1 U5259 ( .C1(n4430), .C2(EBX_REG_11__SCAN_IN), .A(n4219), .B(n4242), 
        .ZN(n4243) );
  NAND2_X1 U5260 ( .A1(n4244), .A2(n4243), .ZN(n5216) );
  OR2_X1 U5261 ( .A1(n4332), .A2(EBX_REG_13__SCAN_IN), .ZN(n4247) );
  NAND2_X1 U5262 ( .A1(n5384), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4245) );
  OAI211_X1 U5263 ( .C1(n4430), .C2(EBX_REG_13__SCAN_IN), .A(n4219), .B(n4245), 
        .ZN(n4246) );
  AND2_X1 U5264 ( .A1(n4247), .A2(n4246), .ZN(n5354) );
  MUX2_X1 U5265 ( .A(n5384), .B(n4219), .S(EBX_REG_12__SCAN_IN), .Z(n4249) );
  NAND2_X1 U5266 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4248) );
  NAND2_X1 U5267 ( .A1(n4249), .A2(n4248), .ZN(n5355) );
  MUX2_X1 U5268 ( .A(n5384), .B(n4219), .S(EBX_REG_14__SCAN_IN), .Z(n4251) );
  NAND2_X1 U5269 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4250) );
  NAND2_X1 U5270 ( .A1(n4251), .A2(n4250), .ZN(n5668) );
  NAND2_X1 U5271 ( .A1(n5669), .A2(n5668), .ZN(n5671) );
  NAND2_X1 U5272 ( .A1(n5390), .A2(EBX_REG_15__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5273 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U5274 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  XNOR2_X1 U5275 ( .A(n4254), .B(n5652), .ZN(n5610) );
  MUX2_X1 U5276 ( .A(n5384), .B(n4219), .S(EBX_REG_16__SCAN_IN), .Z(n4256) );
  NAND2_X1 U5277 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4255) );
  OR2_X1 U5278 ( .A1(n4332), .A2(EBX_REG_17__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U5279 ( .A1(n5384), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4257) );
  OAI211_X1 U5280 ( .C1(n4430), .C2(EBX_REG_17__SCAN_IN), .A(n4219), .B(n4257), 
        .ZN(n4258) );
  NAND2_X1 U5281 ( .A1(n4259), .A2(n4258), .ZN(n5896) );
  NAND2_X1 U5282 ( .A1(n4219), .A2(n3629), .ZN(n4260) );
  OAI211_X1 U5283 ( .C1(n4430), .C2(EBX_REG_19__SCAN_IN), .A(n4260), .B(n5384), 
        .ZN(n4262) );
  INV_X1 U5284 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U5285 ( .A1(n5652), .A2(n5657), .ZN(n4261) );
  NAND2_X1 U5286 ( .A1(n5390), .A2(EBX_REG_18__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U5287 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4263) );
  NAND2_X1 U5288 ( .A1(n4264), .A2(n4263), .ZN(n5653) );
  XNOR2_X1 U5289 ( .A(n5653), .B(n5652), .ZN(n5582) );
  OR2_X1 U5290 ( .A1(n4430), .A2(EBX_REG_20__SCAN_IN), .ZN(n4266) );
  OR2_X1 U5291 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4265)
         );
  NAND2_X1 U5292 ( .A1(n4265), .A2(n4266), .ZN(n5654) );
  MUX2_X1 U5293 ( .A(n4266), .B(n5654), .S(n5384), .Z(n4267) );
  MUX2_X1 U5294 ( .A(n4332), .B(n5384), .S(EBX_REG_21__SCAN_IN), .Z(n4269) );
  OR2_X1 U5295 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4268)
         );
  AND2_X2 U5296 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  OR2_X1 U5297 ( .A1(n4332), .A2(EBX_REG_23__SCAN_IN), .ZN(n4272) );
  NAND2_X1 U5298 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4270) );
  OAI211_X1 U5299 ( .C1(n4430), .C2(EBX_REG_23__SCAN_IN), .A(n4219), .B(n4270), 
        .ZN(n4271) );
  AND2_X1 U5300 ( .A1(n4272), .A2(n4271), .ZN(n5552) );
  MUX2_X1 U5301 ( .A(n5384), .B(n4219), .S(EBX_REG_22__SCAN_IN), .Z(n4274) );
  NAND2_X1 U5302 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U5303 ( .A1(n4274), .A2(n4273), .ZN(n5639) );
  AND2_X1 U5304 ( .A1(n5552), .A2(n5639), .ZN(n4275) );
  NAND2_X1 U5305 ( .A1(n4219), .A2(n4276), .ZN(n4277) );
  OAI211_X1 U5306 ( .C1(n4430), .C2(EBX_REG_24__SCAN_IN), .A(n4277), .B(n5384), 
        .ZN(n4279) );
  INV_X1 U5307 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U5308 ( .A1(n5652), .A2(n5629), .ZN(n4278) );
  NAND2_X1 U5309 ( .A1(n5555), .A2(n4280), .ZN(n4281) );
  NAND2_X1 U5310 ( .A1(n4170), .A2(n6668), .ZN(n4417) );
  OAI21_X1 U5311 ( .B1(n4282), .B2(n3310), .A(n4417), .ZN(n4283) );
  NAND2_X1 U5312 ( .A1(n6375), .A2(REIP_REG_24__SCAN_IN), .ZN(n5736) );
  INV_X1 U5313 ( .A(n5736), .ZN(n4284) );
  AOI21_X1 U5314 ( .B1(n5916), .B2(n6377), .A(n4284), .ZN(n4318) );
  NAND2_X1 U5315 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6330) );
  NOR2_X1 U5316 ( .A1(n5352), .A2(n6330), .ZN(n5998) );
  NAND2_X1 U5317 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5998), .ZN(n5979) );
  INV_X1 U5318 ( .A(n5979), .ZN(n4300) );
  OR2_X1 U5319 ( .A1(n5077), .A2(n3346), .ZN(n4285) );
  NAND2_X1 U5320 ( .A1(n4286), .A2(n4285), .ZN(n4618) );
  NOR2_X1 U5321 ( .A1(n5057), .A2(n6974), .ZN(n6342) );
  NAND3_X1 U5322 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6342), .ZN(n4288) );
  AOI21_X1 U5323 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4754) );
  NAND2_X1 U5324 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4763) );
  NOR2_X1 U5325 ( .A1(n4754), .A2(n4763), .ZN(n6363) );
  NAND2_X1 U5326 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6363), .ZN(n4945)
         );
  NOR2_X1 U5327 ( .A1(n4946), .A2(n4945), .ZN(n5054) );
  INV_X1 U5328 ( .A(n5054), .ZN(n5046) );
  OR2_X1 U5329 ( .A1(n4288), .A2(n5046), .ZN(n4303) );
  NAND2_X1 U5330 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U5331 ( .A1(n4752), .A2(n4763), .ZN(n6362) );
  NAND3_X1 U5332 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6362), .ZN(n5051) );
  NOR2_X1 U5333 ( .A1(n5051), .A2(n4288), .ZN(n5353) );
  OAI21_X1 U5334 ( .B1(n5390), .B2(n4290), .A(n4289), .ZN(n4293) );
  NAND2_X1 U5335 ( .A1(n3344), .A2(n3346), .ZN(n4292) );
  NAND2_X1 U5336 ( .A1(n3367), .A2(n5652), .ZN(n4291) );
  AND4_X1 U5337 ( .A1(n4294), .A2(n4293), .A3(n4292), .A4(n4291), .ZN(n4295)
         );
  NAND2_X1 U5338 ( .A1(n4296), .A2(n4295), .ZN(n4603) );
  OAI21_X1 U5339 ( .B1(n3362), .B2(n4490), .A(n4632), .ZN(n4297) );
  OR2_X1 U5340 ( .A1(n4603), .A2(n4297), .ZN(n4298) );
  NAND2_X1 U5341 ( .A1(n4299), .A2(n4298), .ZN(n5344) );
  AND2_X1 U5342 ( .A1(n4189), .A2(n3489), .ZN(n6517) );
  NAND2_X1 U5343 ( .A1(n5344), .A2(n5359), .ZN(n5052) );
  NAND2_X1 U5344 ( .A1(n5353), .A2(n6384), .ZN(n5863) );
  NAND2_X1 U5345 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5984) );
  INV_X1 U5346 ( .A(n4301), .ZN(n4308) );
  NAND2_X1 U5347 ( .A1(n5903), .A2(n4308), .ZN(n5875) );
  NOR3_X1 U5348 ( .A1(n5861), .A2(n5843), .A3(n6693), .ZN(n4316) );
  NAND2_X1 U5349 ( .A1(n4302), .A2(n6001), .ZN(n4508) );
  OAI21_X1 U5350 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5344), .A(n4508), 
        .ZN(n5050) );
  AOI21_X1 U5351 ( .B1(n6378), .B2(n4303), .A(n5050), .ZN(n4304) );
  OAI21_X1 U5352 ( .B1(n4305), .B2(n5353), .A(n4304), .ZN(n6328) );
  INV_X1 U5353 ( .A(n6328), .ZN(n4307) );
  NAND2_X1 U5354 ( .A1(n5864), .A2(n5344), .ZN(n5348) );
  OAI21_X1 U5355 ( .B1(n5984), .B2(n5979), .A(n6339), .ZN(n4306) );
  NAND2_X1 U5356 ( .A1(n4307), .A2(n4306), .ZN(n5901) );
  NAND2_X1 U5357 ( .A1(n4308), .A2(n5742), .ZN(n4309) );
  AND2_X1 U5358 ( .A1(n6339), .A2(n4309), .ZN(n4310) );
  AND2_X1 U5359 ( .A1(n6339), .A2(n5843), .ZN(n4311) );
  NOR2_X1 U5360 ( .A1(n5858), .A2(n4311), .ZN(n5840) );
  INV_X1 U5361 ( .A(n6384), .ZN(n4312) );
  NAND2_X1 U5362 ( .A1(n5864), .A2(n4312), .ZN(n4314) );
  NAND2_X1 U5363 ( .A1(n4314), .A2(n4313), .ZN(n4315) );
  OAI21_X1 U5364 ( .B1(n4316), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5836), 
        .ZN(n4317) );
  OAI21_X1 U5365 ( .B1(n5741), .B2(n6370), .A(n4319), .ZN(U2994) );
  NAND2_X1 U5366 ( .A1(n4320), .A2(n6382), .ZN(n4342) );
  INV_X1 U5367 ( .A(n6339), .ZN(n5379) );
  NAND2_X1 U5368 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U5369 ( .A1(n6339), .A2(n4339), .ZN(n4321) );
  OAI21_X1 U5370 ( .B1(n5808), .B2(n5379), .A(n5816), .ZN(n5378) );
  INV_X1 U5371 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5542) );
  MUX2_X1 U5372 ( .A(n5384), .B(n4332), .S(n5542), .Z(n4324) );
  OR2_X1 U5373 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4323)
         );
  NAND2_X1 U5374 ( .A1(n4324), .A2(n4323), .ZN(n5540) );
  MUX2_X1 U5375 ( .A(n4332), .B(n5384), .S(EBX_REG_27__SCAN_IN), .Z(n4326) );
  OR2_X1 U5376 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4325)
         );
  NAND2_X1 U5377 ( .A1(n4326), .A2(n4325), .ZN(n5513) );
  INV_X1 U5378 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U5379 ( .A1(n4219), .A2(n5701), .ZN(n4327) );
  OAI211_X1 U5380 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4430), .A(n4327), .B(n4226), 
        .ZN(n4329) );
  INV_X1 U5381 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U5382 ( .A1(n5652), .A2(n5623), .ZN(n4328) );
  AND2_X1 U5383 ( .A1(n4329), .A2(n4328), .ZN(n5512) );
  MUX2_X1 U5384 ( .A(n5384), .B(n4219), .S(EBX_REG_28__SCAN_IN), .Z(n4331) );
  NAND2_X1 U5385 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4330) );
  NAND2_X1 U5386 ( .A1(n4331), .A2(n4330), .ZN(n5501) );
  NOR2_X1 U5387 ( .A1(n5390), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5383)
         );
  MUX2_X1 U5388 ( .A(EBX_REG_29__SCAN_IN), .B(n5383), .S(n4226), .Z(n4334) );
  NOR2_X1 U5389 ( .A1(n4332), .A2(EBX_REG_29__SCAN_IN), .ZN(n4333) );
  OR2_X1 U5390 ( .A1(n4334), .A2(n4333), .ZN(n5387) );
  XNOR2_X1 U5391 ( .A(n5388), .B(n5387), .ZN(n5620) );
  OAI21_X1 U5392 ( .B1(n5620), .B2(n6352), .A(n4335), .ZN(n4336) );
  AOI21_X1 U5393 ( .B1(n5378), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4336), 
        .ZN(n4340) );
  INV_X1 U5394 ( .A(n4337), .ZN(n4338) );
  NAND2_X1 U5395 ( .A1(n5820), .A2(n5808), .ZN(n5448) );
  NAND2_X1 U5396 ( .A1(n4342), .A2(n4341), .ZN(U2989) );
  NAND2_X1 U5397 ( .A1(n4419), .A2(n4402), .ZN(n4393) );
  NAND2_X1 U5398 ( .A1(n4399), .A2(n6543), .ZN(n4394) );
  AND2_X1 U5399 ( .A1(n4345), .A2(n4344), .ZN(n6556) );
  OR2_X1 U5400 ( .A1(n6333), .A2(n6556), .ZN(n4346) );
  NOR3_X1 U5401 ( .A1(n6786), .A2(n6959), .A3(n6560), .ZN(n6548) );
  INV_X1 U5402 ( .A(n4348), .ZN(n4349) );
  NAND2_X1 U5403 ( .A1(n4349), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5422)
         );
  INV_X1 U5404 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5467) );
  NOR2_X1 U5405 ( .A1(n5429), .A2(n6645), .ZN(n4352) );
  NAND2_X1 U5406 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n4357) );
  NAND2_X1 U5407 ( .A1(n6666), .A2(n6941), .ZN(n6542) );
  INV_X1 U5408 ( .A(n6542), .ZN(n4353) );
  INV_X2 U5409 ( .A(n6137), .ZN(n6118) );
  INV_X1 U5410 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6592) );
  INV_X1 U5411 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6589) );
  INV_X1 U5412 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6586) );
  INV_X1 U5413 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6583) );
  NAND3_X1 U5414 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6134) );
  NOR2_X1 U5415 ( .A1(n6583), .A2(n6134), .ZN(n6117) );
  NAND2_X1 U5416 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6117), .ZN(n6094) );
  NOR2_X1 U5417 ( .A1(n6586), .A2(n6094), .ZN(n6087) );
  NAND2_X1 U5418 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6087), .ZN(n5163) );
  NOR2_X1 U5419 ( .A1(n6589), .A2(n5163), .ZN(n6078) );
  NAND2_X1 U5420 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6078), .ZN(n5091) );
  OR2_X1 U5421 ( .A1(n6592), .A2(n5091), .ZN(n6061) );
  NOR2_X1 U5422 ( .A1(n6718), .A2(n6061), .ZN(n5195) );
  NAND2_X1 U5423 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5195), .ZN(n6050) );
  INV_X1 U5424 ( .A(n6050), .ZN(n4356) );
  NAND2_X1 U5425 ( .A1(REIP_REG_13__SCAN_IN), .A2(n4356), .ZN(n6042) );
  NOR2_X1 U5426 ( .A1(n6597), .A2(n6042), .ZN(n4358) );
  AND2_X2 U5427 ( .A1(n6118), .A2(n4358), .ZN(n5611) );
  NAND2_X1 U5428 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5611), .ZN(n5596) );
  NOR2_X2 U5429 ( .A1(n6601), .A2(n5596), .ZN(n6036) );
  NAND2_X1 U5430 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6036), .ZN(n5566) );
  NAND2_X1 U5431 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5945), .ZN(n5941) );
  NAND3_X1 U5432 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4359) );
  NOR2_X1 U5433 ( .A1(n5941), .A2(n4359), .ZN(n5546) );
  NAND2_X1 U5434 ( .A1(n5546), .A2(REIP_REG_24__SCAN_IN), .ZN(n5543) );
  INV_X1 U5435 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5723) );
  INV_X1 U5436 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6617) );
  OR3_X2 U5437 ( .A1(n5543), .A2(n5723), .A3(n6617), .ZN(n5523) );
  NAND2_X1 U5438 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4365) );
  NOR2_X1 U5439 ( .A1(n5523), .A2(n4365), .ZN(n5481) );
  INV_X1 U5440 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6624) );
  AND2_X1 U5441 ( .A1(n5481), .A2(n6624), .ZN(n5477) );
  INV_X1 U5442 ( .A(n5477), .ZN(n4380) );
  INV_X1 U5443 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6604) );
  INV_X1 U5444 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U5445 ( .A1(n4358), .A2(n6092), .ZN(n5615) );
  NOR4_X1 U5446 ( .A1(n6604), .A2(n6601), .A3(n6599), .A4(n5615), .ZN(n5564)
         );
  NAND4_X1 U5447 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5564), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5922) );
  INV_X1 U5448 ( .A(n5922), .ZN(n4361) );
  INV_X1 U5449 ( .A(n4359), .ZN(n4360) );
  NAND2_X1 U5450 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  NAND2_X1 U5451 ( .A1(n6137), .A2(n6092), .ZN(n5923) );
  INV_X1 U5452 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6756) );
  OR3_X1 U5453 ( .A1(n6756), .A2(n5723), .A3(n6617), .ZN(n4363) );
  AND2_X1 U5454 ( .A1(n5923), .A2(n4363), .ZN(n4364) );
  NOR2_X1 U5455 ( .A1(n5914), .A2(n4364), .ZN(n5534) );
  NAND2_X1 U5456 ( .A1(n6118), .A2(n4365), .ZN(n4366) );
  NAND2_X1 U5457 ( .A1(n5534), .A2(n4366), .ZN(n5507) );
  INV_X1 U5458 ( .A(n5078), .ZN(n4369) );
  NAND2_X1 U5459 ( .A1(EBX_REG_31__SCAN_IN), .A2(n6542), .ZN(n4367) );
  NOR2_X1 U5460 ( .A1(n4430), .A2(n4367), .ZN(n4368) );
  AOI22_X1 U5461 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6126), .B1(n6081), 
        .B2(n4371), .ZN(n4377) );
  OAI21_X1 U5462 ( .B1(n6542), .B2(n6671), .A(n6668), .ZN(n4372) );
  NOR2_X1 U5463 ( .A1(n5078), .A2(n4372), .ZN(n5491) );
  INV_X1 U5464 ( .A(n5491), .ZN(n4375) );
  INV_X1 U5465 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6724) );
  NAND3_X1 U5466 ( .A1(n4373), .A2(n6542), .A3(n6724), .ZN(n4374) );
  NAND2_X1 U5467 ( .A1(n6125), .A2(EBX_REG_29__SCAN_IN), .ZN(n4376) );
  OAI211_X1 U5468 ( .C1(n5620), .C2(n6130), .A(n4377), .B(n4376), .ZN(n4378)
         );
  INV_X1 U5469 ( .A(n4378), .ZN(n4379) );
  NAND4_X1 U5470 ( .A1(n3207), .A2(n4380), .A3(n3206), .A4(n4379), .ZN(U2798)
         );
  INV_X1 U5471 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U5472 ( .A1(n5345), .A2(n5348), .ZN(n4514) );
  INV_X1 U5473 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6836) );
  AOI21_X1 U5474 ( .B1(n4508), .B2(n4514), .A(n6836), .ZN(n4392) );
  NOR3_X1 U5475 ( .A1(n5379), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4381), 
        .ZN(n4391) );
  OR2_X1 U5476 ( .A1(n4383), .A2(n4382), .ZN(n4384) );
  AND2_X1 U5477 ( .A1(n4385), .A2(n4384), .ZN(n5182) );
  NOR2_X1 U5478 ( .A1(n6352), .A2(n5182), .ZN(n4390) );
  OAI21_X1 U5479 ( .B1(n4388), .B2(n4387), .A(n4386), .ZN(n6312) );
  INV_X1 U5480 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5186) );
  OAI22_X1 U5481 ( .A1(n6370), .A2(n6312), .B1(n6001), .B2(n5186), .ZN(n4389)
         );
  OR4_X1 U5482 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(U3017) );
  INV_X1 U5483 ( .A(n4393), .ZN(n4412) );
  AND2_X1 U5484 ( .A1(n6447), .A2(n6645), .ZN(n5095) );
  NOR2_X1 U5485 ( .A1(n4412), .A2(n5095), .ZN(n4396) );
  INV_X1 U5486 ( .A(n4394), .ZN(n4398) );
  NOR2_X1 U5487 ( .A1(n4398), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4395) );
  INV_X1 U5488 ( .A(n5077), .ZN(n6672) );
  OR2_X1 U5489 ( .A1(n6672), .A2(n6668), .ZN(n4400) );
  AOI22_X1 U5490 ( .A1(n4396), .A2(n4395), .B1(n6663), .B2(n4400), .ZN(U3474)
         );
  INV_X1 U5491 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4397) );
  OAI21_X1 U5492 ( .B1(n4398), .B2(n4397), .A(n4396), .ZN(U2788) );
  OAI22_X1 U5493 ( .A1(n4622), .A2(n4673), .B1(n4402), .B2(n4399), .ZN(n6009)
         );
  AOI21_X1 U5494 ( .B1(n4400), .B2(n6671), .A(READY_N), .ZN(n4401) );
  NOR2_X1 U5495 ( .A1(n6009), .A2(n4401), .ZN(n6537) );
  NOR2_X1 U5496 ( .A1(n6537), .A2(n6554), .ZN(n6015) );
  INV_X1 U5497 ( .A(MORE_REG_SCAN_IN), .ZN(n4411) );
  OR2_X1 U5498 ( .A1(n6535), .A2(n4402), .ZN(n4403) );
  NOR2_X1 U5499 ( .A1(n4403), .A2(n4613), .ZN(n4409) );
  OR2_X1 U5500 ( .A1(n4405), .A2(n4404), .ZN(n4408) );
  NAND2_X1 U5501 ( .A1(n4622), .A2(n4406), .ZN(n4407) );
  OAI211_X1 U5502 ( .C1(n4622), .C2(n4409), .A(n4408), .B(n4407), .ZN(n6534)
         );
  NAND2_X1 U5503 ( .A1(n6015), .A2(n6534), .ZN(n4410) );
  OAI21_X1 U5504 ( .B1(n6015), .B2(n4411), .A(n4410), .ZN(U3471) );
  OAI21_X2 U5505 ( .B1(n6668), .B2(n6666), .A(n4412), .ZN(n6263) );
  INV_X1 U5506 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6771) );
  INV_X1 U5507 ( .A(n6278), .ZN(n4415) );
  NOR2_X1 U5508 ( .A1(n4430), .A2(READY_N), .ZN(n4413) );
  INV_X1 U5509 ( .A(DATAI_13_), .ZN(n4414) );
  NOR2_X1 U5510 ( .A1(n6239), .A2(n4414), .ZN(n6235) );
  AOI21_X1 U5511 ( .B1(EAX_REG_13__SCAN_IN), .B2(n4415), .A(n6235), .ZN(n4416)
         );
  OAI21_X1 U5512 ( .B1(n6222), .B2(n6771), .A(n4416), .ZN(U2952) );
  INV_X1 U5513 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U5514 ( .A1(n6681), .A2(UWORD_REG_6__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4420) );
  OAI21_X1 U5515 ( .B1(n6821), .B2(n4779), .A(n4420), .ZN(U2901) );
  AOI22_X1 U5516 ( .A1(n6681), .A2(UWORD_REG_4__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4421) );
  OAI21_X1 U5517 ( .B1(n3964), .B2(n4779), .A(n4421), .ZN(U2903) );
  INV_X1 U5518 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6214) );
  AOI22_X1 U5519 ( .A1(n6681), .A2(UWORD_REG_5__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4422) );
  OAI21_X1 U5520 ( .B1(n6214), .B2(n4779), .A(n4422), .ZN(U2902) );
  AOI22_X1 U5521 ( .A1(n6681), .A2(UWORD_REG_2__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4423) );
  OAI21_X1 U5522 ( .B1(n3927), .B2(n4779), .A(n4423), .ZN(U2905) );
  INV_X1 U5523 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6210) );
  AOI22_X1 U5524 ( .A1(n6681), .A2(UWORD_REG_3__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4424) );
  OAI21_X1 U5525 ( .B1(n6210), .B2(n4779), .A(n4424), .ZN(U2904) );
  AOI22_X1 U5526 ( .A1(n6681), .A2(UWORD_REG_0__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4425) );
  OAI21_X1 U5527 ( .B1(n3871), .B2(n4779), .A(n4425), .ZN(U2907) );
  INV_X1 U5528 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6206) );
  AOI22_X1 U5529 ( .A1(n6681), .A2(UWORD_REG_1__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4426) );
  OAI21_X1 U5530 ( .B1(n6206), .B2(n4779), .A(n4426), .ZN(U2906) );
  INV_X1 U5531 ( .A(n4678), .ZN(n5672) );
  NAND3_X1 U5532 ( .A1(n4427), .A2(n3324), .A3(n5672), .ZN(n4429) );
  OAI22_X1 U5533 ( .A1(n4622), .A2(n4605), .B1(n4430), .B2(n4674), .ZN(n4431)
         );
  INV_X1 U5534 ( .A(n5390), .ZN(n4433) );
  AOI21_X1 U5535 ( .B1(n4433), .B2(n5345), .A(n4432), .ZN(n5079) );
  INV_X1 U5536 ( .A(n5079), .ZN(n4518) );
  INV_X1 U5537 ( .A(n4434), .ZN(n4435) );
  XNOR2_X1 U5538 ( .A(n4436), .B(n4435), .ZN(n6326) );
  OAI222_X1 U5539 ( .A1(n6153), .A2(n4518), .B1(n5080), .B2(n6170), .C1(n6148), 
        .C2(n6326), .ZN(U2859) );
  OR2_X1 U5540 ( .A1(n4438), .A2(n4437), .ZN(n4439) );
  INV_X1 U5541 ( .A(n6313), .ZN(n4786) );
  INV_X1 U5542 ( .A(n5182), .ZN(n4440) );
  AOI22_X1 U5543 ( .A1(n6165), .A2(n4440), .B1(EBX_REG_1__SCAN_IN), .B2(n5663), 
        .ZN(n4441) );
  OAI21_X1 U5544 ( .B1(n6148), .B2(n4786), .A(n4441), .ZN(U2858) );
  OR2_X1 U5545 ( .A1(n3107), .A2(n4444), .ZN(n4445) );
  AND2_X1 U5546 ( .A1(n4442), .A2(n4445), .ZN(n6132) );
  INV_X1 U5547 ( .A(n6132), .ZN(n4787) );
  AND2_X1 U5548 ( .A1(n4758), .A2(n4446), .ZN(n4447) );
  OR2_X1 U5549 ( .A1(n4447), .A2(n6109), .ZN(n6129) );
  INV_X1 U5550 ( .A(n6129), .ZN(n4448) );
  AOI22_X1 U5551 ( .A1(n6165), .A2(n4448), .B1(EBX_REG_4__SCAN_IN), .B2(n5663), 
        .ZN(n4449) );
  OAI21_X1 U5552 ( .B1(n4787), .B2(n6148), .A(n4449), .ZN(U2855) );
  INV_X1 U5553 ( .A(n3707), .ZN(n4454) );
  INV_X1 U5554 ( .A(n4451), .ZN(n4453) );
  OR3_X1 U5555 ( .A1(n4454), .A2(n4453), .A3(n4452), .ZN(n4455) );
  AND2_X1 U5556 ( .A1(n4450), .A2(n4455), .ZN(n6308) );
  INV_X1 U5557 ( .A(n6308), .ZN(n4789) );
  NAND2_X1 U5558 ( .A1(n4457), .A2(n4456), .ZN(n4458) );
  AND2_X1 U5559 ( .A1(n4756), .A2(n4458), .ZN(n6376) );
  AOI22_X1 U5560 ( .A1(n6165), .A2(n6376), .B1(EBX_REG_2__SCAN_IN), .B2(n5663), 
        .ZN(n4459) );
  OAI21_X1 U5561 ( .B1(n6148), .B2(n4789), .A(n4459), .ZN(U2857) );
  NAND2_X1 U5562 ( .A1(n4500), .A2(n4460), .ZN(n5125) );
  AOI21_X1 U5563 ( .B1(n4657), .B2(n5906), .A(n6325), .ZN(n4470) );
  NAND2_X1 U5564 ( .A1(n6447), .A2(n6941), .ZN(n5222) );
  INV_X1 U5565 ( .A(n5222), .ZN(n5005) );
  AND2_X1 U5566 ( .A1(n4464), .A2(n6516), .ZN(n5109) );
  INV_X1 U5567 ( .A(n6398), .ZN(n4565) );
  INV_X1 U5568 ( .A(n4507), .ZN(n4469) );
  AOI21_X1 U5569 ( .B1(n5109), .B2(n4565), .A(n4469), .ZN(n4475) );
  OAI21_X1 U5570 ( .B1(n4470), .B2(n5005), .A(n4475), .ZN(n4472) );
  OAI21_X1 U5571 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6959), .A(n4689), 
        .ZN(n6451) );
  INV_X1 U5572 ( .A(n6451), .ZN(n5111) );
  OAI211_X1 U5573 ( .C1(n6447), .C2(n4473), .A(n4472), .B(n5111), .ZN(n4504)
         );
  INV_X1 U5574 ( .A(DATAI_30_), .ZN(n4474) );
  INV_X1 U5575 ( .A(n6495), .ZN(n5304) );
  AND2_X1 U5576 ( .A1(n5906), .A2(n5115), .ZN(n4571) );
  NAND2_X1 U5577 ( .A1(n6314), .A2(DATAI_22_), .ZN(n6500) );
  INV_X1 U5578 ( .A(n6500), .ZN(n5302) );
  OAI22_X1 U5579 ( .A1(n4475), .A2(n6452), .B1(n4688), .B2(n6455), .ZN(n4501)
         );
  AOI22_X1 U5580 ( .A1(n4663), .A2(n5302), .B1(n6497), .B2(n4501), .ZN(n4476)
         );
  OAI21_X1 U5581 ( .B1(n5304), .B2(n4717), .A(n4476), .ZN(n4477) );
  AOI21_X1 U5582 ( .B1(INSTQUEUE_REG_15__6__SCAN_IN), .B2(n4504), .A(n4477), 
        .ZN(n4478) );
  OAI21_X1 U5583 ( .B1(n4507), .B2(n5125), .A(n4478), .ZN(U3146) );
  NAND2_X1 U5584 ( .A1(n4500), .A2(n3299), .ZN(n5128) );
  INV_X1 U5585 ( .A(DATAI_29_), .ZN(n4479) );
  INV_X1 U5586 ( .A(n6489), .ZN(n5316) );
  NAND2_X1 U5587 ( .A1(n6314), .A2(DATAI_21_), .ZN(n6494) );
  INV_X1 U5588 ( .A(n6494), .ZN(n5314) );
  AOI22_X1 U5589 ( .A1(n4663), .A2(n5314), .B1(n6491), .B2(n4501), .ZN(n4480)
         );
  OAI21_X1 U5590 ( .B1(n5316), .B2(n4717), .A(n4480), .ZN(n4481) );
  AOI21_X1 U5591 ( .B1(INSTQUEUE_REG_15__5__SCAN_IN), .B2(n4504), .A(n4481), 
        .ZN(n4482) );
  OAI21_X1 U5592 ( .B1(n4507), .B2(n5128), .A(n4482), .ZN(U3145) );
  INV_X1 U5593 ( .A(DATAI_27_), .ZN(n4483) );
  INV_X1 U5594 ( .A(n6475), .ZN(n5310) );
  NAND2_X1 U5595 ( .A1(n6314), .A2(DATAI_19_), .ZN(n6480) );
  INV_X1 U5596 ( .A(n6480), .ZN(n5308) );
  AOI22_X1 U5597 ( .A1(n4663), .A2(n5308), .B1(n6477), .B2(n4501), .ZN(n4484)
         );
  OAI21_X1 U5598 ( .B1(n5310), .B2(n4717), .A(n4484), .ZN(n4485) );
  AOI21_X1 U5599 ( .B1(INSTQUEUE_REG_15__3__SCAN_IN), .B2(n4504), .A(n4485), 
        .ZN(n4486) );
  OAI21_X1 U5600 ( .B1(n4507), .B2(n5119), .A(n4486), .ZN(U3143) );
  NAND2_X1 U5601 ( .A1(n4500), .A2(n3346), .ZN(n5137) );
  INV_X1 U5602 ( .A(DATAI_2_), .ZN(n4788) );
  NAND2_X1 U5603 ( .A1(n6471), .A2(n4501), .ZN(n4489) );
  NAND2_X1 U5604 ( .A1(n6314), .A2(DATAI_26_), .ZN(n6442) );
  NAND2_X1 U5605 ( .A1(n6314), .A2(DATAI_18_), .ZN(n6474) );
  OAI22_X1 U5606 ( .A1(n6442), .A2(n4717), .B1(n4552), .B2(n6474), .ZN(n4487)
         );
  AOI21_X1 U5607 ( .B1(INSTQUEUE_REG_15__2__SCAN_IN), .B2(n4504), .A(n4487), 
        .ZN(n4488) );
  OAI211_X1 U5608 ( .C1(n5137), .C2(n4507), .A(n4489), .B(n4488), .ZN(U3142)
         );
  NAND2_X1 U5609 ( .A1(n4500), .A2(n4490), .ZN(n5134) );
  INV_X1 U5610 ( .A(DATAI_0_), .ZN(n4870) );
  NAND2_X1 U5611 ( .A1(n6459), .A2(n4501), .ZN(n4493) );
  NAND2_X1 U5612 ( .A1(n6314), .A2(DATAI_24_), .ZN(n6462) );
  NAND2_X1 U5613 ( .A1(n6314), .A2(DATAI_16_), .ZN(n6407) );
  OAI22_X1 U5614 ( .A1(n6462), .A2(n4717), .B1(n4552), .B2(n6407), .ZN(n4491)
         );
  AOI21_X1 U5615 ( .B1(INSTQUEUE_REG_15__0__SCAN_IN), .B2(n4504), .A(n4491), 
        .ZN(n4492) );
  OAI211_X1 U5616 ( .C1(n5134), .C2(n4507), .A(n4493), .B(n4492), .ZN(U3140)
         );
  NAND2_X1 U5617 ( .A1(n4500), .A2(n3310), .ZN(n5131) );
  NAND2_X1 U5618 ( .A1(n6484), .A2(n4501), .ZN(n4496) );
  NAND2_X1 U5619 ( .A1(n6314), .A2(DATAI_28_), .ZN(n6488) );
  NAND2_X1 U5620 ( .A1(n6314), .A2(DATAI_20_), .ZN(n6417) );
  OAI22_X1 U5621 ( .A1(n6488), .A2(n4717), .B1(n4552), .B2(n6417), .ZN(n4494)
         );
  AOI21_X1 U5622 ( .B1(INSTQUEUE_REG_15__4__SCAN_IN), .B2(n4504), .A(n4494), 
        .ZN(n4495) );
  OAI211_X1 U5623 ( .C1(n5131), .C2(n4507), .A(n4496), .B(n4495), .ZN(U3144)
         );
  NAND2_X1 U5624 ( .A1(n4500), .A2(n3489), .ZN(n5143) );
  INV_X1 U5625 ( .A(DATAI_1_), .ZN(n4785) );
  NAND2_X1 U5626 ( .A1(n6465), .A2(n4501), .ZN(n4499) );
  NAND2_X1 U5627 ( .A1(n6314), .A2(DATAI_25_), .ZN(n6433) );
  NAND2_X1 U5628 ( .A1(n6314), .A2(DATAI_17_), .ZN(n6468) );
  OAI22_X1 U5629 ( .A1(n6433), .A2(n4717), .B1(n4552), .B2(n6468), .ZN(n4497)
         );
  AOI21_X1 U5630 ( .B1(INSTQUEUE_REG_15__1__SCAN_IN), .B2(n4504), .A(n4497), 
        .ZN(n4498) );
  OAI211_X1 U5631 ( .C1(n5143), .C2(n4507), .A(n4499), .B(n4498), .ZN(U3141)
         );
  NAND2_X1 U5632 ( .A1(n4500), .A2(n4678), .ZN(n5122) );
  NAND2_X1 U5633 ( .A1(n6506), .A2(n4501), .ZN(n4506) );
  INV_X1 U5634 ( .A(DATAI_31_), .ZN(n4502) );
  NOR2_X1 U5635 ( .A1(n6325), .A2(n4502), .ZN(n6502) );
  INV_X1 U5636 ( .A(n6502), .ZN(n5298) );
  NAND2_X1 U5637 ( .A1(n6314), .A2(DATAI_23_), .ZN(n6511) );
  OAI22_X1 U5638 ( .A1(n5298), .A2(n4717), .B1(n4552), .B2(n6511), .ZN(n4503)
         );
  AOI21_X1 U5639 ( .B1(INSTQUEUE_REG_15__7__SCAN_IN), .B2(n4504), .A(n4503), 
        .ZN(n4505) );
  OAI211_X1 U5640 ( .C1(n5122), .C2(n4507), .A(n4506), .B(n4505), .ZN(U3147)
         );
  INV_X1 U5641 ( .A(n4508), .ZN(n4509) );
  OAI21_X1 U5642 ( .B1(n4510), .B2(n4509), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4517) );
  INV_X1 U5643 ( .A(n4511), .ZN(n4513) );
  AOI21_X1 U5644 ( .B1(n4513), .B2(n5345), .A(n4512), .ZN(n6319) );
  INV_X1 U5645 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6658) );
  OAI21_X1 U5646 ( .B1(n6001), .B2(n6658), .A(n4514), .ZN(n4515) );
  AOI21_X1 U5647 ( .B1(n6382), .B2(n6319), .A(n4515), .ZN(n4516) );
  OAI211_X1 U5648 ( .C1(n6352), .C2(n4518), .A(n4517), .B(n4516), .ZN(U3018)
         );
  NAND3_X1 U5649 ( .A1(n6532), .A2(n6526), .A3(n6701), .ZN(n4728) );
  NOR2_X1 U5650 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4728), .ZN(n4667)
         );
  INV_X1 U5651 ( .A(n4667), .ZN(n4520) );
  AND2_X1 U5652 ( .A1(n4526), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6391) );
  INV_X1 U5653 ( .A(n4961), .ZN(n4519) );
  NOR2_X1 U5654 ( .A1(n4519), .A2(n4962), .ZN(n5010) );
  OAI21_X1 U5655 ( .B1(n5010), .B2(n6455), .A(n4689), .ZN(n5006) );
  AOI211_X1 U5656 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4520), .A(n6391), .B(
        n5006), .ZN(n4525) );
  NOR2_X1 U5657 ( .A1(n4822), .A2(n5906), .ZN(n4522) );
  NOR3_X1 U5658 ( .A1(n4748), .A2(n4663), .A3(n6452), .ZN(n4523) );
  NAND2_X1 U5659 ( .A1(n4466), .A2(n5907), .ZN(n5107) );
  OR2_X1 U5660 ( .A1(n4464), .A2(n5107), .ZN(n4723) );
  OAI21_X1 U5661 ( .B1(n4523), .B2(n5005), .A(n4723), .ZN(n4524) );
  INV_X1 U5662 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4532) );
  OR2_X1 U5663 ( .A1(n4723), .A2(n6452), .ZN(n4528) );
  NAND2_X1 U5664 ( .A1(n5010), .A2(n6400), .ZN(n4527) );
  NAND2_X1 U5665 ( .A1(n4528), .A2(n4527), .ZN(n4662) );
  AOI22_X1 U5666 ( .A1(n4663), .A2(n6489), .B1(n6491), .B2(n4662), .ZN(n4529)
         );
  OAI21_X1 U5667 ( .B1(n4665), .B2(n6494), .A(n4529), .ZN(n4530) );
  AOI21_X1 U5668 ( .B1(n6490), .B2(n4667), .A(n4530), .ZN(n4531) );
  OAI21_X1 U5669 ( .B1(n4670), .B2(n4532), .A(n4531), .ZN(U3025) );
  INV_X1 U5670 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4536) );
  AOI22_X1 U5671 ( .A1(n4663), .A2(n6495), .B1(n6497), .B2(n4662), .ZN(n4533)
         );
  OAI21_X1 U5672 ( .B1(n4665), .B2(n6500), .A(n4533), .ZN(n4534) );
  AOI21_X1 U5673 ( .B1(n6496), .B2(n4667), .A(n4534), .ZN(n4535) );
  OAI21_X1 U5674 ( .B1(n4670), .B2(n4536), .A(n4535), .ZN(U3026) );
  OAI22_X1 U5675 ( .A1(n4665), .A2(n6407), .B1(n6462), .B2(n4552), .ZN(n4537)
         );
  AOI21_X1 U5676 ( .B1(n6445), .B2(n4667), .A(n4537), .ZN(n4539) );
  NAND2_X1 U5677 ( .A1(n6459), .A2(n4662), .ZN(n4538) );
  OAI211_X1 U5678 ( .C1(n4670), .C2(n4540), .A(n4539), .B(n4538), .ZN(U3020)
         );
  INV_X1 U5679 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4544) );
  OAI22_X1 U5680 ( .A1(n4665), .A2(n6417), .B1(n6488), .B2(n4552), .ZN(n4541)
         );
  AOI21_X1 U5681 ( .B1(n6483), .B2(n4667), .A(n4541), .ZN(n4543) );
  NAND2_X1 U5682 ( .A1(n6484), .A2(n4662), .ZN(n4542) );
  OAI211_X1 U5683 ( .C1(n4670), .C2(n4544), .A(n4543), .B(n4542), .ZN(U3024)
         );
  OAI22_X1 U5684 ( .A1(n4665), .A2(n6474), .B1(n6442), .B2(n4552), .ZN(n4545)
         );
  AOI21_X1 U5685 ( .B1(n6470), .B2(n4667), .A(n4545), .ZN(n4547) );
  NAND2_X1 U5686 ( .A1(n6471), .A2(n4662), .ZN(n4546) );
  OAI211_X1 U5687 ( .C1(n4670), .C2(n4548), .A(n4547), .B(n4546), .ZN(U3022)
         );
  OAI22_X1 U5688 ( .A1(n4665), .A2(n6511), .B1(n5298), .B2(n4552), .ZN(n4549)
         );
  AOI21_X1 U5689 ( .B1(n6504), .B2(n4667), .A(n4549), .ZN(n4551) );
  NAND2_X1 U5690 ( .A1(n6506), .A2(n4662), .ZN(n4550) );
  OAI211_X1 U5691 ( .C1(n4670), .C2(n3419), .A(n4551), .B(n4550), .ZN(U3027)
         );
  OAI22_X1 U5692 ( .A1(n4665), .A2(n6468), .B1(n6433), .B2(n4552), .ZN(n4553)
         );
  AOI21_X1 U5693 ( .B1(n6464), .B2(n4667), .A(n4553), .ZN(n4555) );
  NAND2_X1 U5694 ( .A1(n6465), .A2(n4662), .ZN(n4554) );
  OAI211_X1 U5695 ( .C1(n4670), .C2(n4556), .A(n4555), .B(n4554), .ZN(U3021)
         );
  XNOR2_X1 U5696 ( .A(n4558), .B(n3106), .ZN(n4762) );
  AND2_X1 U5697 ( .A1(n4450), .A2(n4559), .ZN(n4560) );
  OR2_X1 U5698 ( .A1(n4560), .A2(n3107), .ZN(n4686) );
  INV_X1 U5699 ( .A(n4686), .ZN(n6167) );
  AND2_X1 U5700 ( .A1(n6333), .A2(REIP_REG_3__SCAN_IN), .ZN(n4759) );
  AOI21_X1 U5701 ( .B1(n6322), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4759), 
        .ZN(n4561) );
  OAI21_X1 U5702 ( .B1(n5145), .B2(n6318), .A(n4561), .ZN(n4562) );
  AOI21_X1 U5703 ( .B1(n6314), .B2(n6167), .A(n4562), .ZN(n4563) );
  OAI21_X1 U5704 ( .B1(n6284), .B2(n4762), .A(n4563), .ZN(U2983) );
  OR2_X1 U5705 ( .A1(n3698), .A2(n5004), .ZN(n4585) );
  INV_X1 U5706 ( .A(n4585), .ZN(n4564) );
  INV_X1 U5707 ( .A(n4582), .ZN(n6436) );
  AOI21_X1 U5708 ( .B1(n4565), .B2(n4564), .A(n6436), .ZN(n4570) );
  NAND2_X1 U5709 ( .A1(n4583), .A2(n6446), .ZN(n4658) );
  NAND3_X1 U5710 ( .A1(n6447), .A2(n4570), .A3(n4658), .ZN(n4567) );
  OAI211_X1 U5711 ( .C1(n4568), .C2(n6447), .A(n5111), .B(n4567), .ZN(n6438)
         );
  NAND2_X1 U5712 ( .A1(n6447), .A2(n4658), .ZN(n4569) );
  INV_X1 U5713 ( .A(n4568), .ZN(n6395) );
  OAI22_X1 U5714 ( .A1(n4570), .A2(n4569), .B1(n6455), .B2(n6395), .ZN(n6437)
         );
  AOI22_X1 U5715 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6438), .B1(n6497), 
        .B2(n6437), .ZN(n4573) );
  AOI22_X1 U5716 ( .A1(n6396), .A2(n6495), .B1(n6434), .B2(n5302), .ZN(n4572)
         );
  OAI211_X1 U5717 ( .C1(n4582), .C2(n5125), .A(n4573), .B(n4572), .ZN(U3082)
         );
  AOI22_X1 U5718 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6438), .B1(n6506), 
        .B2(n6437), .ZN(n4575) );
  INV_X1 U5719 ( .A(n6511), .ZN(n5296) );
  AOI22_X1 U5720 ( .A1(n6396), .A2(n6502), .B1(n6434), .B2(n5296), .ZN(n4574)
         );
  OAI211_X1 U5721 ( .C1(n4582), .C2(n5122), .A(n4575), .B(n4574), .ZN(U3083)
         );
  AOI22_X1 U5722 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6438), .B1(n6484), 
        .B2(n6437), .ZN(n4577) );
  INV_X1 U5723 ( .A(n6488), .ZN(n6414) );
  INV_X1 U5724 ( .A(n6417), .ZN(n6482) );
  AOI22_X1 U5725 ( .A1(n6396), .A2(n6414), .B1(n6434), .B2(n6482), .ZN(n4576)
         );
  OAI211_X1 U5726 ( .C1(n4582), .C2(n5131), .A(n4577), .B(n4576), .ZN(U3080)
         );
  AOI22_X1 U5727 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6438), .B1(n6491), 
        .B2(n6437), .ZN(n4579) );
  AOI22_X1 U5728 ( .A1(n6396), .A2(n6489), .B1(n6434), .B2(n5314), .ZN(n4578)
         );
  OAI211_X1 U5729 ( .C1(n4582), .C2(n5128), .A(n4579), .B(n4578), .ZN(U3081)
         );
  AOI22_X1 U5730 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6438), .B1(n6477), 
        .B2(n6437), .ZN(n4581) );
  AOI22_X1 U5731 ( .A1(n6396), .A2(n6475), .B1(n6434), .B2(n5308), .ZN(n4580)
         );
  OAI211_X1 U5732 ( .C1(n4582), .C2(n5119), .A(n4581), .B(n4580), .ZN(U3079)
         );
  NAND2_X1 U5733 ( .A1(n4583), .A2(n4656), .ZN(n4591) );
  OAI21_X1 U5734 ( .B1(n4591), .B2(n6941), .A(n6447), .ZN(n5009) );
  INV_X1 U5735 ( .A(n5009), .ZN(n4587) );
  NAND2_X1 U5736 ( .A1(n6701), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4856) );
  OR2_X1 U5737 ( .A1(n4856), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5002)
         );
  NOR2_X1 U5738 ( .A1(n6799), .A2(n5002), .ZN(n4805) );
  INV_X1 U5739 ( .A(n4805), .ZN(n4584) );
  OAI21_X1 U5740 ( .B1(n5003), .B2(n4585), .A(n4584), .ZN(n4589) );
  INV_X1 U5741 ( .A(n5002), .ZN(n4586) );
  AOI21_X1 U5742 ( .B1(n6452), .B2(n5002), .A(n6451), .ZN(n4588) );
  OAI21_X1 U5743 ( .B1(n5009), .B2(n4589), .A(n4588), .ZN(n4804) );
  AOI22_X1 U5744 ( .A1(n6496), .A2(n4805), .B1(n4804), .B2(
        INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4593) );
  INV_X1 U5745 ( .A(n4591), .ZN(n4590) );
  NAND2_X1 U5746 ( .A1(n4590), .A2(n4957), .ZN(n5037) );
  NOR2_X2 U5747 ( .A1(n4591), .A2(n4957), .ZN(n6424) );
  AOI22_X1 U5748 ( .A1(n5031), .A2(n6495), .B1(n6424), .B2(n5302), .ZN(n4592)
         );
  OAI211_X1 U5749 ( .C1(n4808), .C2(n5307), .A(n4593), .B(n4592), .ZN(U3066)
         );
  AOI22_X1 U5750 ( .A1(n6490), .A2(n4805), .B1(n4804), .B2(
        INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5751 ( .A1(n5031), .A2(n6489), .B1(n6424), .B2(n5314), .ZN(n4594)
         );
  OAI211_X1 U5752 ( .C1(n4808), .C2(n5319), .A(n4595), .B(n4594), .ZN(U3065)
         );
  XNOR2_X1 U5753 ( .A(n4597), .B(n3104), .ZN(n4770) );
  NOR2_X1 U5754 ( .A1(n6001), .A2(n6583), .ZN(n4766) );
  AOI21_X1 U5755 ( .B1(n6322), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4766), 
        .ZN(n4598) );
  OAI21_X1 U5756 ( .B1(n6147), .B2(n6318), .A(n4598), .ZN(n4599) );
  AOI21_X1 U5757 ( .B1(n6132), .B2(n6314), .A(n4599), .ZN(n4600) );
  OAI21_X1 U5758 ( .B1(n6284), .B2(n4770), .A(n4600), .ZN(U2982) );
  INV_X1 U5759 ( .A(n4170), .ZN(n4621) );
  NAND4_X1 U5760 ( .A1(n6003), .A2(n3362), .A3(n4621), .A4(n4601), .ZN(n4602)
         );
  NOR2_X1 U5761 ( .A1(n4603), .A2(n4602), .ZN(n6512) );
  OR2_X1 U5762 ( .A1(n4466), .A2(n6512), .ZN(n4612) );
  NAND2_X1 U5763 ( .A1(n4605), .A2(n4604), .ZN(n4641) );
  INV_X1 U5764 ( .A(n4606), .ZN(n5365) );
  NAND2_X1 U5765 ( .A1(n5365), .A2(n3379), .ZN(n4629) );
  NAND2_X1 U5766 ( .A1(n4606), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U5767 ( .A1(n4629), .A2(n4631), .ZN(n4610) );
  XNOR2_X1 U5768 ( .A(n3379), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4607)
         );
  NAND2_X1 U5769 ( .A1(n6517), .A2(n4607), .ZN(n4608) );
  OAI21_X1 U5770 ( .B1(n4610), .B2(n4632), .A(n4608), .ZN(n4609) );
  AOI21_X1 U5771 ( .B1(n4641), .B2(n4610), .A(n4609), .ZN(n4611) );
  AND2_X1 U5772 ( .A1(n4612), .A2(n4611), .ZN(n5366) );
  NAND2_X1 U5773 ( .A1(n4622), .A2(n4613), .ZN(n4617) );
  INV_X1 U5774 ( .A(n4614), .ZN(n4615) );
  INV_X1 U5775 ( .A(n4676), .ZN(n4628) );
  INV_X1 U5776 ( .A(n4618), .ZN(n4627) );
  INV_X1 U5777 ( .A(n6671), .ZN(n4619) );
  NAND2_X1 U5778 ( .A1(n4619), .A2(n6666), .ZN(n4620) );
  AOI21_X1 U5779 ( .B1(n4637), .B2(n4621), .A(n4620), .ZN(n4623) );
  OAI21_X1 U5780 ( .B1(n4624), .B2(n4623), .A(n4622), .ZN(n4625) );
  NAND4_X1 U5781 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n6518)
         );
  MUX2_X1 U5782 ( .A(n3379), .B(n5366), .S(n6518), .Z(n6523) );
  NOR2_X1 U5783 ( .A1(n6523), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4644) );
  INV_X1 U5784 ( .A(n4464), .ZN(n6392) );
  INV_X1 U5785 ( .A(n4629), .ZN(n4630) );
  XNOR2_X1 U5786 ( .A(n4630), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4640)
         );
  AOI21_X1 U5787 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4631), .A(n4133), 
        .ZN(n6641) );
  NOR2_X1 U5788 ( .A1(n4632), .A2(n6641), .ZN(n4639) );
  MUX2_X1 U5789 ( .A(n4635), .B(n4634), .S(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .Z(n4636) );
  NOR3_X1 U5790 ( .A1(n4637), .A2(n4633), .A3(n4636), .ZN(n4638) );
  AOI211_X1 U5791 ( .C1(n4641), .C2(n4640), .A(n4639), .B(n4638), .ZN(n4642)
         );
  OAI21_X1 U5792 ( .B1(n6392), .B2(n6512), .A(n4642), .ZN(n6639) );
  MUX2_X1 U5793 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6639), .S(n6518), 
        .Z(n6533) );
  OR2_X1 U5794 ( .A1(n6645), .A2(FLUSH_REG_SCAN_IN), .ZN(n4646) );
  INV_X1 U5795 ( .A(n4646), .ZN(n4643) );
  AOI22_X1 U5796 ( .A1(n4644), .A2(n6533), .B1(n4634), .B2(n4643), .ZN(n6540)
         );
  OAI21_X1 U5797 ( .B1(n6518), .B2(STATE2_REG_1__SCAN_IN), .A(n4646), .ZN(
        n4650) );
  INV_X1 U5798 ( .A(n5004), .ZN(n4647) );
  OR2_X1 U5799 ( .A1(n3469), .A2(n4647), .ZN(n4648) );
  XNOR2_X1 U5800 ( .A(n4648), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6138)
         );
  NOR2_X1 U5801 ( .A1(n6003), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5802 ( .A1(n4650), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n6138), .B2(n4649), .ZN(n6539) );
  OAI21_X1 U5803 ( .B1(n6540), .B2(n4645), .A(n6539), .ZN(n4653) );
  NOR2_X1 U5804 ( .A1(n6786), .A2(n4652), .ZN(n6561) );
  OAI21_X1 U5805 ( .B1(n4653), .B2(FLUSH_REG_SCAN_IN), .A(n6561), .ZN(n4651)
         );
  NAND2_X1 U5806 ( .A1(n4651), .A2(n4963), .ZN(n6389) );
  NOR2_X1 U5807 ( .A1(n4653), .A2(n4652), .ZN(n6549) );
  AND2_X1 U5808 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6959), .ZN(n5910) );
  OAI22_X1 U5809 ( .A1(n4957), .A2(n6452), .B1(n3698), .B2(n5910), .ZN(n4654)
         );
  OAI21_X1 U5810 ( .B1(n6549), .B2(n4654), .A(n6389), .ZN(n4655) );
  OAI21_X1 U5811 ( .B1(n6389), .B2(n6799), .A(n4655), .ZN(U3465) );
  NAND2_X1 U5812 ( .A1(n4858), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4859) );
  AND2_X1 U5813 ( .A1(n4859), .A2(n6449), .ZN(n4815) );
  AOI21_X1 U5814 ( .B1(n4815), .B2(n4658), .A(n6452), .ZN(n4660) );
  INV_X1 U5815 ( .A(n4822), .ZN(n4824) );
  OAI22_X1 U5816 ( .A1(n4824), .A2(n5222), .B1(n6392), .B2(n5910), .ZN(n4659)
         );
  OAI21_X1 U5817 ( .B1(n4660), .B2(n4659), .A(n6389), .ZN(n4661) );
  OAI21_X1 U5818 ( .B1(n6389), .B2(n6532), .A(n4661), .ZN(U3462) );
  INV_X1 U5819 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4669) );
  AOI22_X1 U5820 ( .A1(n4663), .A2(n6475), .B1(n6477), .B2(n4662), .ZN(n4664)
         );
  OAI21_X1 U5821 ( .B1(n4665), .B2(n6480), .A(n4664), .ZN(n4666) );
  AOI21_X1 U5822 ( .B1(n6476), .B2(n4667), .A(n4666), .ZN(n4668) );
  OAI21_X1 U5823 ( .B1(n4670), .B2(n4669), .A(n4668), .ZN(U3023) );
  AOI22_X1 U5824 ( .A1(n6476), .A2(n4805), .B1(n4804), .B2(
        INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5825 ( .A1(n5031), .A2(n6475), .B1(n6424), .B2(n5308), .ZN(n4671)
         );
  OAI211_X1 U5826 ( .C1(n4808), .C2(n5313), .A(n4672), .B(n4671), .ZN(U3063)
         );
  NOR2_X1 U5827 ( .A1(n4674), .A2(n5076), .ZN(n4675) );
  AND2_X1 U5828 ( .A1(n4679), .A2(n4678), .ZN(n4682) );
  INV_X1 U5829 ( .A(n4682), .ZN(n4680) );
  INV_X1 U5830 ( .A(n6177), .ZN(n4684) );
  INV_X1 U5831 ( .A(n6180), .ZN(n4683) );
  AOI22_X1 U5832 ( .A1(n6183), .A2(DATAI_3_), .B1(EAX_REG_3__SCAN_IN), .B2(
        n6179), .ZN(n4685) );
  OAI21_X1 U5833 ( .B1(n5951), .B2(n4686), .A(n4685), .ZN(U2888) );
  NOR2_X1 U5834 ( .A1(n6398), .A2(n6452), .ZN(n6393) );
  INV_X1 U5835 ( .A(n4962), .ZN(n4687) );
  NOR2_X1 U5836 ( .A1(n4687), .A2(n6532), .ZN(n5289) );
  AOI22_X1 U5837 ( .A1(n6393), .A2(n4464), .B1(n6391), .B2(n5289), .ZN(n4722)
         );
  NOR2_X1 U5838 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4688), .ZN(n4719)
         );
  OAI21_X1 U5839 ( .B1(n4962), .B2(n6455), .A(n4689), .ZN(n6399) );
  NOR3_X1 U5840 ( .A1(n6399), .A2(n6532), .A3(n6400), .ZN(n4693) );
  OAI21_X1 U5841 ( .B1(n4894), .B2(n4690), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4691) );
  NAND3_X1 U5842 ( .A1(n6398), .A2(n6447), .A3(n4691), .ZN(n4692) );
  NAND2_X1 U5843 ( .A1(n4716), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4696)
         );
  OAI22_X1 U5844 ( .A1(n4879), .A2(n5298), .B1(n6511), .B2(n4717), .ZN(n4694)
         );
  AOI21_X1 U5845 ( .B1(n6504), .B2(n4719), .A(n4694), .ZN(n4695) );
  OAI211_X1 U5846 ( .C1(n4722), .C2(n5301), .A(n4696), .B(n4695), .ZN(U3139)
         );
  INV_X1 U5847 ( .A(n4719), .ZN(n4712) );
  NAND2_X1 U5848 ( .A1(n4716), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4699)
         );
  OAI22_X1 U5849 ( .A1(n4717), .A2(n6494), .B1(n4722), .B2(n5319), .ZN(n4697)
         );
  AOI21_X1 U5850 ( .B1(n6489), .B2(n4894), .A(n4697), .ZN(n4698) );
  OAI211_X1 U5851 ( .C1(n4712), .C2(n5128), .A(n4699), .B(n4698), .ZN(U3137)
         );
  NAND2_X1 U5852 ( .A1(n4716), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4702)
         );
  OAI22_X1 U5853 ( .A1(n4879), .A2(n6442), .B1(n6474), .B2(n4717), .ZN(n4700)
         );
  AOI21_X1 U5854 ( .B1(n6470), .B2(n4719), .A(n4700), .ZN(n4701) );
  OAI211_X1 U5855 ( .C1(n4722), .C2(n5323), .A(n4702), .B(n4701), .ZN(U3134)
         );
  NAND2_X1 U5856 ( .A1(n4716), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4705)
         );
  OAI22_X1 U5857 ( .A1(n4879), .A2(n6433), .B1(n6468), .B2(n4717), .ZN(n4703)
         );
  AOI21_X1 U5858 ( .B1(n6464), .B2(n4719), .A(n4703), .ZN(n4704) );
  OAI211_X1 U5859 ( .C1(n4722), .C2(n5331), .A(n4705), .B(n4704), .ZN(U3133)
         );
  NAND2_X1 U5860 ( .A1(n4716), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4708)
         );
  OAI22_X1 U5861 ( .A1(n4717), .A2(n6500), .B1(n4722), .B2(n5307), .ZN(n4706)
         );
  AOI21_X1 U5862 ( .B1(n6495), .B2(n4894), .A(n4706), .ZN(n4707) );
  OAI211_X1 U5863 ( .C1(n4712), .C2(n5125), .A(n4708), .B(n4707), .ZN(U3138)
         );
  NAND2_X1 U5864 ( .A1(n4716), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4711)
         );
  OAI22_X1 U5865 ( .A1(n4717), .A2(n6480), .B1(n4722), .B2(n5313), .ZN(n4709)
         );
  AOI21_X1 U5866 ( .B1(n6475), .B2(n4894), .A(n4709), .ZN(n4710) );
  OAI211_X1 U5867 ( .C1(n4712), .C2(n5119), .A(n4711), .B(n4710), .ZN(U3135)
         );
  NAND2_X1 U5868 ( .A1(n4716), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4715)
         );
  OAI22_X1 U5869 ( .A1(n4879), .A2(n6462), .B1(n6407), .B2(n4717), .ZN(n4713)
         );
  AOI21_X1 U5870 ( .B1(n6445), .B2(n4719), .A(n4713), .ZN(n4714) );
  OAI211_X1 U5871 ( .C1(n4722), .C2(n5339), .A(n4715), .B(n4714), .ZN(U3132)
         );
  NAND2_X1 U5872 ( .A1(n4716), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4721)
         );
  OAI22_X1 U5873 ( .A1(n4879), .A2(n6488), .B1(n6417), .B2(n4717), .ZN(n4718)
         );
  AOI21_X1 U5874 ( .B1(n6483), .B2(n4719), .A(n4718), .ZN(n4720) );
  OAI211_X1 U5875 ( .C1(n4722), .C2(n5327), .A(n4721), .B(n4720), .ZN(U3136)
         );
  NOR2_X1 U5876 ( .A1(n6799), .A2(n4728), .ZN(n4724) );
  INV_X1 U5877 ( .A(n4723), .ZN(n4725) );
  AOI21_X1 U5878 ( .B1(n4725), .B2(n6516), .A(n4724), .ZN(n4729) );
  AOI21_X1 U5879 ( .B1(n4731), .B2(STATEBS16_REG_SCAN_IN), .A(n6452), .ZN(
        n4727) );
  AOI22_X1 U5880 ( .A1(n4729), .A2(n4727), .B1(n6452), .B2(n4728), .ZN(n4726)
         );
  NAND2_X1 U5881 ( .A1(n5111), .A2(n4726), .ZN(n4747) );
  INV_X1 U5882 ( .A(n4727), .ZN(n4730) );
  OAI22_X1 U5883 ( .A1(n4730), .A2(n4729), .B1(n6455), .B2(n4728), .ZN(n4746)
         );
  AOI22_X1 U5884 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4747), .B1(n6471), 
        .B2(n4746), .ZN(n4733) );
  INV_X1 U5885 ( .A(n6442), .ZN(n6469) );
  INV_X1 U5886 ( .A(n6474), .ZN(n6435) );
  AOI22_X1 U5887 ( .A1(n4748), .A2(n6469), .B1(n4931), .B2(n6435), .ZN(n4732)
         );
  OAI211_X1 U5888 ( .C1(n4751), .C2(n5137), .A(n4733), .B(n4732), .ZN(U3030)
         );
  AOI22_X1 U5889 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4747), .B1(n6459), 
        .B2(n4746), .ZN(n4735) );
  INV_X1 U5890 ( .A(n6462), .ZN(n6404) );
  INV_X1 U5891 ( .A(n6407), .ZN(n6444) );
  AOI22_X1 U5892 ( .A1(n6404), .A2(n4748), .B1(n4931), .B2(n6444), .ZN(n4734)
         );
  OAI211_X1 U5893 ( .C1(n4751), .C2(n5134), .A(n4735), .B(n4734), .ZN(U3028)
         );
  AOI22_X1 U5894 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4747), .B1(n6484), 
        .B2(n4746), .ZN(n4737) );
  AOI22_X1 U5895 ( .A1(n4748), .A2(n6414), .B1(n4931), .B2(n6482), .ZN(n4736)
         );
  OAI211_X1 U5896 ( .C1(n4751), .C2(n5131), .A(n4737), .B(n4736), .ZN(U3032)
         );
  AOI22_X1 U5897 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4747), .B1(n6506), 
        .B2(n4746), .ZN(n4739) );
  AOI22_X1 U5898 ( .A1(n4748), .A2(n6502), .B1(n4931), .B2(n5296), .ZN(n4738)
         );
  OAI211_X1 U5899 ( .C1(n4751), .C2(n5122), .A(n4739), .B(n4738), .ZN(U3035)
         );
  AOI22_X1 U5900 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4747), .B1(n6477), 
        .B2(n4746), .ZN(n4741) );
  AOI22_X1 U5901 ( .A1(n4748), .A2(n6475), .B1(n4931), .B2(n5308), .ZN(n4740)
         );
  OAI211_X1 U5902 ( .C1(n4751), .C2(n5119), .A(n4741), .B(n4740), .ZN(U3031)
         );
  AOI22_X1 U5903 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4747), .B1(n6491), 
        .B2(n4746), .ZN(n4743) );
  AOI22_X1 U5904 ( .A1(n4748), .A2(n6489), .B1(n4931), .B2(n5314), .ZN(n4742)
         );
  OAI211_X1 U5905 ( .C1(n4751), .C2(n5128), .A(n4743), .B(n4742), .ZN(U3033)
         );
  AOI22_X1 U5906 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4747), .B1(n6465), 
        .B2(n4746), .ZN(n4745) );
  INV_X1 U5907 ( .A(n6433), .ZN(n6463) );
  INV_X1 U5908 ( .A(n6468), .ZN(n6430) );
  AOI22_X1 U5909 ( .A1(n4748), .A2(n6463), .B1(n4931), .B2(n6430), .ZN(n4744)
         );
  OAI211_X1 U5910 ( .C1(n4751), .C2(n5143), .A(n4745), .B(n4744), .ZN(U3029)
         );
  AOI22_X1 U5911 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4747), .B1(n6497), 
        .B2(n4746), .ZN(n4750) );
  AOI22_X1 U5912 ( .A1(n4748), .A2(n6495), .B1(n4931), .B2(n5302), .ZN(n4749)
         );
  OAI211_X1 U5913 ( .C1(n4751), .C2(n5125), .A(n4750), .B(n4749), .ZN(U3034)
         );
  AOI21_X1 U5914 ( .B1(n5052), .B2(n4752), .A(n5050), .ZN(n6380) );
  NAND2_X1 U5915 ( .A1(n6378), .A2(n4754), .ZN(n6386) );
  NAND2_X1 U5916 ( .A1(n6380), .A2(n6386), .ZN(n4767) );
  INV_X1 U5917 ( .A(n4752), .ZN(n4753) );
  AOI21_X1 U5918 ( .B1(n4753), .B2(n6384), .A(n6378), .ZN(n5045) );
  NOR2_X1 U5919 ( .A1(n4754), .A2(n5045), .ZN(n4764) );
  AOI22_X1 U5920 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4767), .B1(n4764), 
        .B2(n6694), .ZN(n4761) );
  NAND2_X1 U5921 ( .A1(n4756), .A2(n4755), .ZN(n4757) );
  AND2_X1 U5922 ( .A1(n4758), .A2(n4757), .ZN(n6164) );
  AOI21_X1 U5923 ( .B1(n6377), .B2(n6164), .A(n4759), .ZN(n4760) );
  OAI211_X1 U5924 ( .C1(n6370), .C2(n4762), .A(n4761), .B(n4760), .ZN(U3015)
         );
  OAI211_X1 U5925 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4764), .B(n4763), .ZN(n4769) );
  NOR2_X1 U5926 ( .A1(n6352), .A2(n6129), .ZN(n4765) );
  AOI211_X1 U5927 ( .C1(n4767), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4766), 
        .B(n4765), .ZN(n4768) );
  OAI211_X1 U5928 ( .C1(n6370), .C2(n4770), .A(n4769), .B(n4768), .ZN(U3014)
         );
  INV_X1 U5929 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U5930 ( .A1(n6665), .A2(UWORD_REG_14__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4771) );
  OAI21_X1 U5931 ( .B1(n6958), .B2(n4779), .A(n4771), .ZN(U2893) );
  INV_X1 U5932 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6225) );
  AOI22_X1 U5933 ( .A1(n6665), .A2(UWORD_REG_9__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4772) );
  OAI21_X1 U5934 ( .B1(n6225), .B2(n4779), .A(n4772), .ZN(U2898) );
  INV_X1 U5935 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6956) );
  AOI22_X1 U5936 ( .A1(n6665), .A2(UWORD_REG_8__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4773) );
  OAI21_X1 U5937 ( .B1(n6956), .B2(n4779), .A(n4773), .ZN(U2899) );
  INV_X1 U5938 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6219) );
  AOI22_X1 U5939 ( .A1(n6665), .A2(UWORD_REG_7__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4774) );
  OAI21_X1 U5940 ( .B1(n6219), .B2(n4779), .A(n4774), .ZN(U2900) );
  AOI22_X1 U5941 ( .A1(n6665), .A2(UWORD_REG_10__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4775) );
  OAI21_X1 U5942 ( .B1(n6228), .B2(n4779), .A(n4775), .ZN(U2897) );
  INV_X1 U5943 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6237) );
  AOI22_X1 U5944 ( .A1(n6665), .A2(UWORD_REG_13__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4776) );
  OAI21_X1 U5945 ( .B1(n6237), .B2(n4779), .A(n4776), .ZN(U2894) );
  INV_X1 U5946 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6234) );
  AOI22_X1 U5947 ( .A1(n6665), .A2(UWORD_REG_12__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4777) );
  OAI21_X1 U5948 ( .B1(n6234), .B2(n4779), .A(n4777), .ZN(U2895) );
  INV_X1 U5949 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6231) );
  AOI22_X1 U5950 ( .A1(n6665), .A2(UWORD_REG_11__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4778) );
  OAI21_X1 U5951 ( .B1(n6231), .B2(n4779), .A(n4778), .ZN(U2896) );
  INV_X1 U5952 ( .A(n4781), .ZN(n4782) );
  AOI21_X1 U5953 ( .B1(n4783), .B2(n4780), .A(n4782), .ZN(n4953) );
  INV_X1 U5954 ( .A(n4953), .ZN(n6101) );
  XNOR2_X1 U5955 ( .A(n6110), .B(n3208), .ZN(n6098) );
  AOI22_X1 U5956 ( .A1(n6165), .A2(n6098), .B1(EBX_REG_6__SCAN_IN), .B2(n5663), 
        .ZN(n4784) );
  OAI21_X1 U5957 ( .B1(n6101), .B2(n6148), .A(n4784), .ZN(U2853) );
  INV_X1 U5958 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6768) );
  OAI222_X1 U5959 ( .A1(n4786), .A2(n5951), .B1(n5001), .B2(n4785), .C1(n6186), 
        .C2(n6768), .ZN(U2890) );
  INV_X1 U5960 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6253) );
  OAI222_X1 U5961 ( .A1(n4787), .A2(n5951), .B1(n5001), .B2(n6962), .C1(n6253), 
        .C2(n6186), .ZN(U2887) );
  INV_X1 U5962 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6247) );
  OAI222_X1 U5963 ( .A1(n4789), .A2(n5951), .B1(n5001), .B2(n4788), .C1(n6186), 
        .C2(n6247), .ZN(U2889) );
  INV_X1 U5964 ( .A(n6424), .ZN(n4802) );
  OAI22_X1 U5965 ( .A1(n4802), .A2(n6511), .B1(n5298), .B2(n5037), .ZN(n4790)
         );
  AOI21_X1 U5966 ( .B1(INSTQUEUE_REG_5__7__SCAN_IN), .B2(n4804), .A(n4790), 
        .ZN(n4792) );
  NAND2_X1 U5967 ( .A1(n6504), .A2(n4805), .ZN(n4791) );
  OAI211_X1 U5968 ( .C1(n5301), .C2(n4808), .A(n4792), .B(n4791), .ZN(U3067)
         );
  OAI22_X1 U5969 ( .A1(n4802), .A2(n6417), .B1(n6488), .B2(n5037), .ZN(n4793)
         );
  AOI21_X1 U5970 ( .B1(INSTQUEUE_REG_5__4__SCAN_IN), .B2(n4804), .A(n4793), 
        .ZN(n4795) );
  NAND2_X1 U5971 ( .A1(n6483), .A2(n4805), .ZN(n4794) );
  OAI211_X1 U5972 ( .C1(n5327), .C2(n4808), .A(n4795), .B(n4794), .ZN(U3064)
         );
  OAI22_X1 U5973 ( .A1(n4802), .A2(n6407), .B1(n6462), .B2(n5037), .ZN(n4796)
         );
  AOI21_X1 U5974 ( .B1(INSTQUEUE_REG_5__0__SCAN_IN), .B2(n4804), .A(n4796), 
        .ZN(n4798) );
  NAND2_X1 U5975 ( .A1(n6445), .A2(n4805), .ZN(n4797) );
  OAI211_X1 U5976 ( .C1(n5339), .C2(n4808), .A(n4798), .B(n4797), .ZN(U3060)
         );
  OAI22_X1 U5977 ( .A1(n4802), .A2(n6474), .B1(n6442), .B2(n5037), .ZN(n4799)
         );
  AOI21_X1 U5978 ( .B1(INSTQUEUE_REG_5__2__SCAN_IN), .B2(n4804), .A(n4799), 
        .ZN(n4801) );
  NAND2_X1 U5979 ( .A1(n6470), .A2(n4805), .ZN(n4800) );
  OAI211_X1 U5980 ( .C1(n5323), .C2(n4808), .A(n4801), .B(n4800), .ZN(U3062)
         );
  OAI22_X1 U5981 ( .A1(n4802), .A2(n6468), .B1(n6433), .B2(n5037), .ZN(n4803)
         );
  AOI21_X1 U5982 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(n4804), .A(n4803), 
        .ZN(n4807) );
  NAND2_X1 U5983 ( .A1(n6464), .A2(n4805), .ZN(n4806) );
  OAI211_X1 U5984 ( .C1(n5331), .C2(n4808), .A(n4807), .B(n4806), .ZN(U3061)
         );
  INV_X1 U5985 ( .A(n4809), .ZN(n4810) );
  NAND2_X1 U5986 ( .A1(n4442), .A2(n4810), .ZN(n4811) );
  INV_X1 U5987 ( .A(n6300), .ZN(n4813) );
  INV_X1 U5988 ( .A(DATAI_5_), .ZN(n6212) );
  OAI222_X1 U5989 ( .A1(n4813), .A2(n5951), .B1(n6212), .B2(n5001), .C1(n4812), 
        .C2(n6186), .ZN(U2886) );
  INV_X1 U5990 ( .A(DATAI_6_), .ZN(n6215) );
  OAI222_X1 U5991 ( .A1(n6101), .A2(n5951), .B1(n6215), .B2(n5001), .C1(n4814), 
        .C2(n6186), .ZN(U2885) );
  NAND3_X1 U5992 ( .A1(n4815), .A2(n6446), .A3(n4823), .ZN(n4816) );
  NAND2_X1 U5993 ( .A1(n4816), .A2(n6447), .ZN(n4828) );
  INV_X1 U5994 ( .A(n4828), .ZN(n4820) );
  NAND2_X1 U5995 ( .A1(n4466), .A2(n4468), .ZN(n5287) );
  OR2_X1 U5996 ( .A1(n4464), .A2(n5287), .ZN(n4901) );
  OR2_X1 U5997 ( .A1(n4901), .A2(n3698), .ZN(n4818) );
  INV_X1 U5998 ( .A(n6443), .ZN(n4817) );
  NAND2_X1 U5999 ( .A1(n4817), .A2(n6532), .ZN(n4850) );
  NAND2_X1 U6000 ( .A1(n4818), .A2(n4850), .ZN(n4827) );
  NAND3_X1 U6001 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6532), .A3(n6526), .ZN(n4899) );
  INV_X1 U6002 ( .A(n4899), .ZN(n4819) );
  INV_X1 U6003 ( .A(n4850), .ZN(n4838) );
  INV_X1 U6004 ( .A(n4821), .ZN(n5285) );
  NOR3_X1 U6005 ( .A1(n4822), .A2(n3110), .A3(n5285), .ZN(n4900) );
  NAND4_X1 U6006 ( .A1(n4824), .A2(n5115), .A3(n4823), .A4(n5906), .ZN(n5036)
         );
  OAI22_X1 U6007 ( .A1(n4929), .A2(n6462), .B1(n6407), .B2(n5036), .ZN(n4825)
         );
  AOI21_X1 U6008 ( .B1(n6445), .B2(n4838), .A(n4825), .ZN(n4830) );
  AOI21_X1 U6009 ( .B1(n6452), .B2(n4899), .A(n6451), .ZN(n4826) );
  NAND2_X1 U6010 ( .A1(n4853), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4829) );
  OAI211_X1 U6011 ( .C1(n5339), .C2(n4855), .A(n4830), .B(n4829), .ZN(U3044)
         );
  OAI22_X1 U6012 ( .A1(n4929), .A2(n5316), .B1(n6494), .B2(n5036), .ZN(n4831)
         );
  AOI21_X1 U6013 ( .B1(n6490), .B2(n4838), .A(n4831), .ZN(n4833) );
  NAND2_X1 U6014 ( .A1(n4853), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4832) );
  OAI211_X1 U6015 ( .C1(n4855), .C2(n5319), .A(n4833), .B(n4832), .ZN(U3049)
         );
  OAI22_X1 U6016 ( .A1(n4929), .A2(n5304), .B1(n6500), .B2(n5036), .ZN(n4834)
         );
  AOI21_X1 U6017 ( .B1(n6496), .B2(n4838), .A(n4834), .ZN(n4836) );
  NAND2_X1 U6018 ( .A1(n4853), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4835) );
  OAI211_X1 U6019 ( .C1(n4855), .C2(n5307), .A(n4836), .B(n4835), .ZN(U3050)
         );
  OAI22_X1 U6020 ( .A1(n4929), .A2(n5310), .B1(n6480), .B2(n5036), .ZN(n4837)
         );
  AOI21_X1 U6021 ( .B1(n6476), .B2(n4838), .A(n4837), .ZN(n4840) );
  NAND2_X1 U6022 ( .A1(n4853), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4839) );
  OAI211_X1 U6023 ( .C1(n4855), .C2(n5313), .A(n4840), .B(n4839), .ZN(U3047)
         );
  OAI22_X1 U6024 ( .A1(n4929), .A2(n6433), .B1(n6468), .B2(n5036), .ZN(n4842)
         );
  NOR2_X1 U6025 ( .A1(n5143), .A2(n4850), .ZN(n4841) );
  AOI211_X1 U6026 ( .C1(n4853), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4842), 
        .B(n4841), .ZN(n4843) );
  OAI21_X1 U6027 ( .B1(n5331), .B2(n4855), .A(n4843), .ZN(U3045) );
  OAI22_X1 U6028 ( .A1(n4929), .A2(n5298), .B1(n6511), .B2(n5036), .ZN(n4845)
         );
  NOR2_X1 U6029 ( .A1(n5122), .A2(n4850), .ZN(n4844) );
  AOI211_X1 U6030 ( .C1(n4853), .C2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4845), 
        .B(n4844), .ZN(n4846) );
  OAI21_X1 U6031 ( .B1(n5301), .B2(n4855), .A(n4846), .ZN(U3051) );
  OAI22_X1 U6032 ( .A1(n4929), .A2(n6442), .B1(n6474), .B2(n5036), .ZN(n4848)
         );
  NOR2_X1 U6033 ( .A1(n5137), .A2(n4850), .ZN(n4847) );
  AOI211_X1 U6034 ( .C1(n4853), .C2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4848), 
        .B(n4847), .ZN(n4849) );
  OAI21_X1 U6035 ( .B1(n5323), .B2(n4855), .A(n4849), .ZN(U3046) );
  OAI22_X1 U6036 ( .A1(n4929), .A2(n6488), .B1(n6417), .B2(n5036), .ZN(n4852)
         );
  NOR2_X1 U6037 ( .A1(n5131), .A2(n4850), .ZN(n4851) );
  AOI211_X1 U6038 ( .C1(n4853), .C2(INSTQUEUE_REG_3__4__SCAN_IN), .A(n4852), 
        .B(n4851), .ZN(n4854) );
  OAI21_X1 U6039 ( .B1(n5327), .B2(n4855), .A(n4854), .ZN(U3048) );
  INV_X1 U6040 ( .A(n5003), .ZN(n4960) );
  NOR2_X1 U6041 ( .A1(n6532), .A2(n4856), .ZN(n4956) );
  AND2_X1 U6042 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4956), .ZN(n4883)
         );
  AOI21_X1 U6043 ( .B1(n5109), .B2(n4960), .A(n4883), .ZN(n4860) );
  NAND2_X1 U6044 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4857) );
  OAI22_X1 U6045 ( .A1(n4860), .A2(n6452), .B1(n4857), .B2(n4856), .ZN(n4891)
         );
  NAND2_X1 U6046 ( .A1(n4858), .A2(n4957), .ZN(n4991) );
  INV_X1 U6047 ( .A(n4991), .ZN(n4877) );
  NAND2_X1 U6048 ( .A1(n4860), .A2(n4859), .ZN(n4863) );
  INV_X1 U6049 ( .A(n4956), .ZN(n4861) );
  NAND2_X1 U6050 ( .A1(n6452), .A2(n4861), .ZN(n4862) );
  OAI211_X1 U6051 ( .C1(n6452), .C2(n4863), .A(n5111), .B(n4862), .ZN(n4890)
         );
  AOI22_X1 U6052 ( .A1(n4877), .A2(n6414), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4890), .ZN(n4864) );
  OAI21_X1 U6053 ( .B1(n6417), .B2(n4879), .A(n4864), .ZN(n4865) );
  AOI21_X1 U6054 ( .B1(n6483), .B2(n4883), .A(n4865), .ZN(n4866) );
  OAI21_X1 U6055 ( .B1(n5327), .B2(n4882), .A(n4866), .ZN(U3128) );
  AOI22_X1 U6056 ( .A1(n4877), .A2(n6404), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4890), .ZN(n4867) );
  OAI21_X1 U6057 ( .B1(n6407), .B2(n4879), .A(n4867), .ZN(n4868) );
  AOI21_X1 U6058 ( .B1(n6445), .B2(n4883), .A(n4868), .ZN(n4869) );
  OAI21_X1 U6059 ( .B1(n5339), .B2(n4882), .A(n4869), .ZN(U3124) );
  INV_X1 U6060 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6723) );
  OAI222_X1 U6061 ( .A1(n5951), .A2(n6326), .B1(n6186), .B2(n6723), .C1(n4870), 
        .C2(n5001), .ZN(U2891) );
  AOI22_X1 U6062 ( .A1(n4877), .A2(n6502), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4890), .ZN(n4871) );
  OAI21_X1 U6063 ( .B1(n6511), .B2(n4879), .A(n4871), .ZN(n4872) );
  AOI21_X1 U6064 ( .B1(n6504), .B2(n4883), .A(n4872), .ZN(n4873) );
  OAI21_X1 U6065 ( .B1(n5301), .B2(n4882), .A(n4873), .ZN(U3131) );
  AOI22_X1 U6066 ( .A1(n4877), .A2(n6469), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4890), .ZN(n4874) );
  OAI21_X1 U6067 ( .B1(n6474), .B2(n4879), .A(n4874), .ZN(n4875) );
  AOI21_X1 U6068 ( .B1(n6470), .B2(n4883), .A(n4875), .ZN(n4876) );
  OAI21_X1 U6069 ( .B1(n5323), .B2(n4882), .A(n4876), .ZN(U3126) );
  AOI22_X1 U6070 ( .A1(n4877), .A2(n6463), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4890), .ZN(n4878) );
  OAI21_X1 U6071 ( .B1(n6468), .B2(n4879), .A(n4878), .ZN(n4880) );
  AOI21_X1 U6072 ( .B1(n6464), .B2(n4883), .A(n4880), .ZN(n4881) );
  OAI21_X1 U6073 ( .B1(n5331), .B2(n4882), .A(n4881), .ZN(U3125) );
  INV_X1 U6074 ( .A(n4883), .ZN(n4896) );
  AOI22_X1 U6075 ( .A1(n4891), .A2(n6497), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4890), .ZN(n4884) );
  OAI21_X1 U6076 ( .B1(n4991), .B2(n5304), .A(n4884), .ZN(n4885) );
  AOI21_X1 U6077 ( .B1(n5302), .B2(n4894), .A(n4885), .ZN(n4886) );
  OAI21_X1 U6078 ( .B1(n5125), .B2(n4896), .A(n4886), .ZN(U3130) );
  AOI22_X1 U6079 ( .A1(n4891), .A2(n6477), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4890), .ZN(n4887) );
  OAI21_X1 U6080 ( .B1(n4991), .B2(n5310), .A(n4887), .ZN(n4888) );
  AOI21_X1 U6081 ( .B1(n5308), .B2(n4894), .A(n4888), .ZN(n4889) );
  OAI21_X1 U6082 ( .B1(n5119), .B2(n4896), .A(n4889), .ZN(U3127) );
  AOI22_X1 U6083 ( .A1(n4891), .A2(n6491), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4890), .ZN(n4892) );
  OAI21_X1 U6084 ( .B1(n4991), .B2(n5316), .A(n4892), .ZN(n4893) );
  AOI21_X1 U6085 ( .B1(n5314), .B2(n4894), .A(n4893), .ZN(n4895) );
  OAI21_X1 U6086 ( .B1(n5128), .B2(n4896), .A(n4895), .ZN(U3129) );
  OR2_X1 U6087 ( .A1(n4901), .A2(n6452), .ZN(n4898) );
  AND2_X1 U6088 ( .A1(n4962), .A2(n6532), .ZN(n6390) );
  NAND2_X1 U6089 ( .A1(n6400), .A2(n6390), .ZN(n4897) );
  NOR2_X1 U6090 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4899), .ZN(n4924)
         );
  OAI21_X1 U6091 ( .B1(n4931), .B2(n4900), .A(n5222), .ZN(n4902) );
  AOI21_X1 U6092 ( .B1(n4902), .B2(n4901), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4903) );
  NOR2_X1 U6093 ( .A1(n6391), .A2(n6399), .ZN(n5295) );
  NAND2_X1 U6094 ( .A1(n4927), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4906) );
  INV_X1 U6095 ( .A(n4931), .ZN(n4922) );
  OAI22_X1 U6096 ( .A1(n4922), .A2(n6488), .B1(n4929), .B2(n6417), .ZN(n4904)
         );
  AOI21_X1 U6097 ( .B1(n6483), .B2(n4924), .A(n4904), .ZN(n4905) );
  OAI211_X1 U6098 ( .C1(n4928), .C2(n5327), .A(n4906), .B(n4905), .ZN(U3040)
         );
  NAND2_X1 U6099 ( .A1(n4927), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4909) );
  OAI22_X1 U6100 ( .A1(n4922), .A2(n6462), .B1(n6407), .B2(n4929), .ZN(n4907)
         );
  AOI21_X1 U6101 ( .B1(n6445), .B2(n4924), .A(n4907), .ZN(n4908) );
  OAI211_X1 U6102 ( .C1(n4928), .C2(n5339), .A(n4909), .B(n4908), .ZN(U3036)
         );
  INV_X1 U6103 ( .A(n4924), .ZN(n4934) );
  NAND2_X1 U6104 ( .A1(n4927), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4912) );
  OAI22_X1 U6105 ( .A1(n4929), .A2(n6494), .B1(n4928), .B2(n5319), .ZN(n4910)
         );
  AOI21_X1 U6106 ( .B1(n4931), .B2(n6489), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6107 ( .C1(n4934), .C2(n5128), .A(n4912), .B(n4911), .ZN(U3041)
         );
  NAND2_X1 U6108 ( .A1(n4927), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4915) );
  OAI22_X1 U6109 ( .A1(n4929), .A2(n6480), .B1(n4928), .B2(n5313), .ZN(n4913)
         );
  AOI21_X1 U6110 ( .B1(n4931), .B2(n6475), .A(n4913), .ZN(n4914) );
  OAI211_X1 U6111 ( .C1(n4934), .C2(n5119), .A(n4915), .B(n4914), .ZN(U3039)
         );
  NAND2_X1 U6112 ( .A1(n4927), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4918) );
  OAI22_X1 U6113 ( .A1(n4922), .A2(n6442), .B1(n4929), .B2(n6474), .ZN(n4916)
         );
  AOI21_X1 U6114 ( .B1(n6470), .B2(n4924), .A(n4916), .ZN(n4917) );
  OAI211_X1 U6115 ( .C1(n4928), .C2(n5323), .A(n4918), .B(n4917), .ZN(U3038)
         );
  NAND2_X1 U6116 ( .A1(n4927), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4921) );
  OAI22_X1 U6117 ( .A1(n4922), .A2(n6433), .B1(n4929), .B2(n6468), .ZN(n4919)
         );
  AOI21_X1 U6118 ( .B1(n6464), .B2(n4924), .A(n4919), .ZN(n4920) );
  OAI211_X1 U6119 ( .C1(n4928), .C2(n5331), .A(n4921), .B(n4920), .ZN(U3037)
         );
  NAND2_X1 U6120 ( .A1(n4927), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4926) );
  OAI22_X1 U6121 ( .A1(n4922), .A2(n5298), .B1(n4929), .B2(n6511), .ZN(n4923)
         );
  AOI21_X1 U6122 ( .B1(n6504), .B2(n4924), .A(n4923), .ZN(n4925) );
  OAI211_X1 U6123 ( .C1(n4928), .C2(n5301), .A(n4926), .B(n4925), .ZN(U3043)
         );
  NAND2_X1 U6124 ( .A1(n4927), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4933) );
  OAI22_X1 U6125 ( .A1(n4929), .A2(n6500), .B1(n4928), .B2(n5307), .ZN(n4930)
         );
  AOI21_X1 U6126 ( .B1(n4931), .B2(n6495), .A(n4930), .ZN(n4932) );
  OAI211_X1 U6127 ( .C1(n4934), .C2(n5125), .A(n4933), .B(n4932), .ZN(U3042)
         );
  XNOR2_X1 U6128 ( .A(n4999), .B(n4936), .ZN(n5167) );
  NOR2_X1 U6129 ( .A1(n5047), .A2(n4937), .ZN(n4938) );
  OR2_X1 U6130 ( .A1(n6072), .A2(n4938), .ZN(n5160) );
  INV_X1 U6131 ( .A(n5160), .ZN(n4939) );
  AOI22_X1 U6132 ( .A1(n6165), .A2(n4939), .B1(EBX_REG_8__SCAN_IN), .B2(n5663), 
        .ZN(n4940) );
  OAI21_X1 U6133 ( .B1(n5167), .B2(n6148), .A(n4940), .ZN(U2851) );
  AOI22_X1 U6134 ( .A1(n6183), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6179), .ZN(n4941) );
  OAI21_X1 U6135 ( .B1(n5167), .B2(n5951), .A(n4941), .ZN(U2883) );
  XNOR2_X1 U6136 ( .A(n4943), .B(n4942), .ZN(n4955) );
  NOR2_X1 U6137 ( .A1(n6001), .A2(n6586), .ZN(n4950) );
  INV_X1 U6139 ( .A(n6380), .ZN(n4944) );
  AOI21_X1 U6140 ( .B1(n6339), .B2(n4945), .A(n4944), .ZN(n6365) );
  OAI33_X1 U6141 ( .A1(1'b0), .A2(n6365), .A3(n4946), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4945), .B3(n5045), .ZN(n4948) );
  AOI211_X1 U6142 ( .C1(n6377), .C2(n6098), .A(n4950), .B(n4948), .ZN(n4949)
         );
  OAI21_X1 U6143 ( .B1(n6370), .B2(n4955), .A(n4949), .ZN(U3012) );
  AOI21_X1 U6144 ( .B1(n6322), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4950), 
        .ZN(n4951) );
  OAI21_X1 U6145 ( .B1(n6099), .B2(n6318), .A(n4951), .ZN(n4952) );
  AOI21_X1 U6146 ( .B1(n4953), .B2(n6314), .A(n4952), .ZN(n4954) );
  OAI21_X1 U6147 ( .B1(n6284), .B2(n4955), .A(n4954), .ZN(U2980) );
  AND2_X1 U6148 ( .A1(n6799), .A2(n4956), .ZN(n4993) );
  INV_X1 U6149 ( .A(n4993), .ZN(n4980) );
  INV_X1 U6150 ( .A(n5116), .ZN(n4958) );
  AOI21_X1 U6151 ( .B1(n6510), .B2(n4991), .A(n6941), .ZN(n4959) );
  AOI211_X1 U6152 ( .C1(n4960), .C2(n5004), .A(n6452), .B(n4959), .ZN(n4966)
         );
  INV_X1 U6153 ( .A(n6400), .ZN(n4964) );
  OR2_X1 U6154 ( .A1(n4962), .A2(n4961), .ZN(n4967) );
  AOI21_X1 U6155 ( .B1(n4967), .B2(STATE2_REG_2__SCAN_IN), .A(n4963), .ZN(
        n5225) );
  OAI211_X1 U6156 ( .C1(n6959), .C2(n4993), .A(n4964), .B(n5225), .ZN(n4965)
         );
  NAND2_X1 U6157 ( .A1(n4990), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4970)
         );
  NOR2_X1 U6158 ( .A1(n5003), .A2(n6452), .ZN(n5011) );
  INV_X1 U6159 ( .A(n4967), .ZN(n5231) );
  AOI22_X1 U6160 ( .A1(n5011), .A2(n4464), .B1(n5231), .B2(n6391), .ZN(n4996)
         );
  OAI22_X1 U6161 ( .A1(n4991), .A2(n6500), .B1(n4996), .B2(n5307), .ZN(n4968)
         );
  AOI21_X1 U6162 ( .B1(n6481), .B2(n6495), .A(n4968), .ZN(n4969) );
  OAI211_X1 U6163 ( .C1(n4980), .C2(n5125), .A(n4970), .B(n4969), .ZN(U3122)
         );
  NAND2_X1 U6164 ( .A1(n4990), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4973)
         );
  OAI22_X1 U6165 ( .A1(n4991), .A2(n6494), .B1(n4996), .B2(n5319), .ZN(n4971)
         );
  AOI21_X1 U6166 ( .B1(n6481), .B2(n6489), .A(n4971), .ZN(n4972) );
  OAI211_X1 U6167 ( .C1(n4980), .C2(n5128), .A(n4973), .B(n4972), .ZN(U3121)
         );
  NAND2_X1 U6168 ( .A1(n4990), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4976)
         );
  OAI22_X1 U6169 ( .A1(n6510), .A2(n6488), .B1(n6417), .B2(n4991), .ZN(n4974)
         );
  AOI21_X1 U6170 ( .B1(n6483), .B2(n4993), .A(n4974), .ZN(n4975) );
  OAI211_X1 U6171 ( .C1(n4996), .C2(n5327), .A(n4976), .B(n4975), .ZN(U3120)
         );
  NAND2_X1 U6172 ( .A1(n4990), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4979)
         );
  OAI22_X1 U6173 ( .A1(n4991), .A2(n6480), .B1(n4996), .B2(n5313), .ZN(n4977)
         );
  AOI21_X1 U6174 ( .B1(n6481), .B2(n6475), .A(n4977), .ZN(n4978) );
  OAI211_X1 U6175 ( .C1(n4980), .C2(n5119), .A(n4979), .B(n4978), .ZN(U3119)
         );
  NAND2_X1 U6176 ( .A1(n4990), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4983)
         );
  OAI22_X1 U6177 ( .A1(n6510), .A2(n6442), .B1(n6474), .B2(n4991), .ZN(n4981)
         );
  AOI21_X1 U6178 ( .B1(n6470), .B2(n4993), .A(n4981), .ZN(n4982) );
  OAI211_X1 U6179 ( .C1(n4996), .C2(n5323), .A(n4983), .B(n4982), .ZN(U3118)
         );
  NAND2_X1 U6180 ( .A1(n4990), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4986)
         );
  OAI22_X1 U6181 ( .A1(n6510), .A2(n6433), .B1(n6468), .B2(n4991), .ZN(n4984)
         );
  AOI21_X1 U6182 ( .B1(n6464), .B2(n4993), .A(n4984), .ZN(n4985) );
  OAI211_X1 U6183 ( .C1(n4996), .C2(n5331), .A(n4986), .B(n4985), .ZN(U3117)
         );
  NAND2_X1 U6184 ( .A1(n4990), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4989)
         );
  OAI22_X1 U6185 ( .A1(n6510), .A2(n6462), .B1(n6407), .B2(n4991), .ZN(n4987)
         );
  AOI21_X1 U6186 ( .B1(n6445), .B2(n4993), .A(n4987), .ZN(n4988) );
  OAI211_X1 U6187 ( .C1(n4996), .C2(n5339), .A(n4989), .B(n4988), .ZN(U3116)
         );
  NAND2_X1 U6188 ( .A1(n4990), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4995)
         );
  OAI22_X1 U6189 ( .A1(n6510), .A2(n5298), .B1(n6511), .B2(n4991), .ZN(n4992)
         );
  AOI21_X1 U6190 ( .B1(n6504), .B2(n4993), .A(n4992), .ZN(n4994) );
  OAI211_X1 U6191 ( .C1(n4996), .C2(n5301), .A(n4995), .B(n4994), .ZN(U3123)
         );
  AND2_X1 U6192 ( .A1(n4781), .A2(n4997), .ZN(n4998) );
  NOR2_X1 U6193 ( .A1(n4999), .A2(n4998), .ZN(n6289) );
  INV_X1 U6194 ( .A(n6289), .ZN(n5064) );
  INV_X1 U6195 ( .A(DATAI_7_), .ZN(n6217) );
  OAI222_X1 U6196 ( .A1(n5064), .A2(n5951), .B1(n6217), .B2(n5001), .C1(n5000), 
        .C2(n6186), .ZN(U2884) );
  NOR2_X1 U6197 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5002), .ZN(n5039)
         );
  INV_X1 U6198 ( .A(n5039), .ZN(n5034) );
  OAI22_X1 U6199 ( .A1(n5036), .A2(n5005), .B1(n5004), .B2(n5003), .ZN(n5008)
         );
  AOI211_X1 U6200 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5034), .A(n6400), .B(
        n5006), .ZN(n5007) );
  NAND2_X1 U6201 ( .A1(n5035), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U6202 ( .A1(n5011), .A2(n6392), .B1(n6391), .B2(n5010), .ZN(n5042)
         );
  OAI22_X1 U6203 ( .A1(n5036), .A2(n5310), .B1(n5042), .B2(n5313), .ZN(n5012)
         );
  AOI21_X1 U6204 ( .B1(n5308), .B2(n5031), .A(n5012), .ZN(n5013) );
  OAI211_X1 U6205 ( .C1(n5034), .C2(n5119), .A(n5014), .B(n5013), .ZN(U3055)
         );
  NAND2_X1 U6206 ( .A1(n5035), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5017) );
  OAI22_X1 U6207 ( .A1(n5036), .A2(n5304), .B1(n5042), .B2(n5307), .ZN(n5015)
         );
  AOI21_X1 U6208 ( .B1(n5302), .B2(n5031), .A(n5015), .ZN(n5016) );
  OAI211_X1 U6209 ( .C1(n5034), .C2(n5125), .A(n5017), .B(n5016), .ZN(U3058)
         );
  NAND2_X1 U6210 ( .A1(n5035), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5020) );
  OAI22_X1 U6211 ( .A1(n5037), .A2(n6407), .B1(n5036), .B2(n6462), .ZN(n5018)
         );
  AOI21_X1 U6212 ( .B1(n6445), .B2(n5039), .A(n5018), .ZN(n5019) );
  OAI211_X1 U6213 ( .C1(n5042), .C2(n5339), .A(n5020), .B(n5019), .ZN(U3052)
         );
  NAND2_X1 U6214 ( .A1(n5035), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5023) );
  OAI22_X1 U6215 ( .A1(n5037), .A2(n6468), .B1(n5036), .B2(n6433), .ZN(n5021)
         );
  AOI21_X1 U6216 ( .B1(n6464), .B2(n5039), .A(n5021), .ZN(n5022) );
  OAI211_X1 U6217 ( .C1(n5042), .C2(n5331), .A(n5023), .B(n5022), .ZN(U3053)
         );
  NAND2_X1 U6218 ( .A1(n5035), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5026) );
  OAI22_X1 U6219 ( .A1(n5037), .A2(n6511), .B1(n5036), .B2(n5298), .ZN(n5024)
         );
  AOI21_X1 U6220 ( .B1(n6504), .B2(n5039), .A(n5024), .ZN(n5025) );
  OAI211_X1 U6221 ( .C1(n5042), .C2(n5301), .A(n5026), .B(n5025), .ZN(U3059)
         );
  NAND2_X1 U6222 ( .A1(n5035), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5029) );
  OAI22_X1 U6223 ( .A1(n5037), .A2(n6417), .B1(n5036), .B2(n6488), .ZN(n5027)
         );
  AOI21_X1 U6224 ( .B1(n6483), .B2(n5039), .A(n5027), .ZN(n5028) );
  OAI211_X1 U6225 ( .C1(n5042), .C2(n5327), .A(n5029), .B(n5028), .ZN(U3056)
         );
  NAND2_X1 U6226 ( .A1(n5035), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5033) );
  OAI22_X1 U6227 ( .A1(n5036), .A2(n5316), .B1(n5042), .B2(n5319), .ZN(n5030)
         );
  AOI21_X1 U6228 ( .B1(n5314), .B2(n5031), .A(n5030), .ZN(n5032) );
  OAI211_X1 U6229 ( .C1(n5034), .C2(n5128), .A(n5033), .B(n5032), .ZN(U3057)
         );
  NAND2_X1 U6230 ( .A1(n5035), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5041) );
  OAI22_X1 U6231 ( .A1(n5037), .A2(n6474), .B1(n5036), .B2(n6442), .ZN(n5038)
         );
  AOI21_X1 U6232 ( .B1(n6470), .B2(n5039), .A(n5038), .ZN(n5040) );
  OAI211_X1 U6233 ( .C1(n5042), .C2(n5323), .A(n5041), .B(n5040), .ZN(U3054)
         );
  XNOR2_X1 U6234 ( .A(n5043), .B(n5044), .ZN(n6286) );
  NOR2_X1 U6235 ( .A1(n5046), .A2(n5045), .ZN(n6341) );
  AOI21_X1 U6236 ( .B1(n5049), .B2(n5048), .A(n5047), .ZN(n6086) );
  INV_X1 U6237 ( .A(n6086), .ZN(n5065) );
  AOI21_X1 U6238 ( .B1(n5052), .B2(n5051), .A(n5050), .ZN(n5053) );
  OAI21_X1 U6239 ( .B1(n5054), .B2(n5864), .A(n5053), .ZN(n6338) );
  NAND2_X1 U6240 ( .A1(n6338), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5055)
         );
  NAND2_X1 U6241 ( .A1(n6375), .A2(REIP_REG_7__SCAN_IN), .ZN(n6291) );
  OAI211_X1 U6242 ( .C1(n6352), .C2(n5065), .A(n5055), .B(n6291), .ZN(n5056)
         );
  AOI21_X1 U6243 ( .B1(n6341), .B2(n5057), .A(n5056), .ZN(n5058) );
  OAI21_X1 U6244 ( .B1(n6370), .B2(n6286), .A(n5058), .ZN(U3011) );
  INV_X1 U6245 ( .A(n5059), .ZN(n5062) );
  INV_X1 U6246 ( .A(n5060), .ZN(n5088) );
  OAI21_X1 U6247 ( .B1(n5062), .B2(n5061), .A(n5088), .ZN(n6079) );
  AOI22_X1 U6248 ( .A1(n6183), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6179), .ZN(n5063) );
  OAI21_X1 U6249 ( .B1(n6079), .B2(n5951), .A(n5063), .ZN(U2882) );
  INV_X1 U6250 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6774) );
  OAI222_X1 U6251 ( .A1(n5065), .A2(n6153), .B1(n6170), .B2(n6774), .C1(n5064), 
        .C2(n6148), .ZN(U2852) );
  XNOR2_X1 U6252 ( .A(n5066), .B(n5067), .ZN(n5075) );
  INV_X1 U6253 ( .A(n5167), .ZN(n5070) );
  AOI22_X1 U6254 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6375), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5068) );
  OAI21_X1 U6255 ( .B1(n5159), .B2(n6318), .A(n5068), .ZN(n5069) );
  AOI21_X1 U6256 ( .B1(n5070), .B2(n6314), .A(n5069), .ZN(n5071) );
  OAI21_X1 U6257 ( .B1(n5075), .B2(n6284), .A(n5071), .ZN(U2978) );
  INV_X1 U6258 ( .A(n6342), .ZN(n6340) );
  OAI211_X1 U6259 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6341), .B(n6340), .ZN(n5074) );
  OAI22_X1 U6260 ( .A1(n6352), .A2(n5160), .B1(n6589), .B2(n6001), .ZN(n5072)
         );
  AOI21_X1 U6261 ( .B1(n6338), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5072), 
        .ZN(n5073) );
  OAI211_X1 U6262 ( .C1(n6370), .C2(n5075), .A(n5074), .B(n5073), .ZN(U3010)
         );
  OAI21_X1 U6263 ( .B1(n5078), .B2(n5076), .A(n6100), .ZN(n6133) );
  INV_X1 U6264 ( .A(n6133), .ZN(n5085) );
  NOR2_X1 U6265 ( .A1(n5078), .A2(n5077), .ZN(n6139) );
  AOI22_X1 U6266 ( .A1(n6112), .A2(n5079), .B1(n6139), .B2(n6516), .ZN(n5084)
         );
  NAND2_X1 U6267 ( .A1(n6106), .A2(n6146), .ZN(n5082) );
  INV_X1 U6268 ( .A(n5923), .ZN(n5565) );
  OAI22_X1 U6269 ( .A1(n5565), .A2(n6658), .B1(n6123), .B2(n5080), .ZN(n5081)
         );
  AOI21_X1 U6270 ( .B1(n5082), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5081), 
        .ZN(n5083) );
  OAI211_X1 U6271 ( .C1(n5085), .C2(n6326), .A(n5084), .B(n5083), .ZN(U2827)
         );
  AND2_X1 U6272 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  NOR2_X1 U6273 ( .A1(n5086), .A2(n5089), .ZN(n5207) );
  INV_X1 U6274 ( .A(n5207), .ZN(n5104) );
  AOI22_X1 U6275 ( .A1(n6183), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6179), .ZN(n5090) );
  OAI21_X1 U6276 ( .B1(n5104), .B2(n5951), .A(n5090), .ZN(U2881) );
  NOR3_X1 U6277 ( .A1(n6137), .A2(REIP_REG_10__SCAN_IN), .A3(n5091), .ZN(n5099) );
  INV_X1 U6278 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5103) );
  INV_X1 U6279 ( .A(n5092), .ZN(n5094) );
  OAI21_X1 U6280 ( .B1(n5094), .B2(n5093), .A(n5217), .ZN(n6345) );
  OAI22_X1 U6281 ( .A1(n6123), .A2(n5103), .B1(n6130), .B2(n6345), .ZN(n5096)
         );
  AOI211_X1 U6282 ( .C1(n6126), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5096), 
        .B(n6113), .ZN(n5097) );
  OAI21_X1 U6283 ( .B1(n6146), .B2(n5205), .A(n5097), .ZN(n5098) );
  NOR2_X1 U6284 ( .A1(n5099), .A2(n5098), .ZN(n5102) );
  INV_X1 U6285 ( .A(n6078), .ZN(n5100) );
  NAND2_X1 U6286 ( .A1(n6118), .A2(n5100), .ZN(n5162) );
  NAND2_X1 U6287 ( .A1(n5162), .A2(n6092), .ZN(n6074) );
  NOR2_X1 U6288 ( .A1(n6137), .A2(REIP_REG_9__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U6289 ( .B1(n6074), .B2(n6077), .A(REIP_REG_10__SCAN_IN), .ZN(n5101) );
  OAI211_X1 U6290 ( .C1(n5104), .C2(n6100), .A(n5102), .B(n5101), .ZN(U2817)
         );
  OAI222_X1 U6291 ( .A1(n5104), .A2(n6148), .B1(n6170), .B2(n5103), .C1(n6345), 
        .C2(n6153), .ZN(U2849) );
  NAND3_X1 U6292 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6526), .A3(n6701), .ZN(n5224) );
  NOR2_X1 U6293 ( .A1(n6799), .A2(n5224), .ZN(n5108) );
  OR2_X1 U6294 ( .A1(n5906), .A2(n6941), .ZN(n5105) );
  OR2_X1 U6295 ( .A1(n6449), .A2(n5105), .ZN(n5106) );
  AND2_X1 U6296 ( .A1(n5106), .A2(n6447), .ZN(n5112) );
  INV_X1 U6297 ( .A(n5107), .ZN(n5221) );
  AOI21_X1 U6298 ( .B1(n5109), .B2(n5221), .A(n5108), .ZN(n5114) );
  AOI22_X1 U6299 ( .A1(n5112), .A2(n5114), .B1(n6452), .B2(n5224), .ZN(n5110)
         );
  NAND2_X1 U6300 ( .A1(n5111), .A2(n5110), .ZN(n5139) );
  INV_X1 U6301 ( .A(n5112), .ZN(n5113) );
  OAI22_X1 U6302 ( .A1(n5114), .A2(n5113), .B1(n6455), .B2(n5224), .ZN(n5138)
         );
  AOI22_X1 U6303 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5139), .B1(n6477), 
        .B2(n5138), .ZN(n5118) );
  NOR3_X2 U6304 ( .A1(n6449), .A2(n5115), .A3(n5906), .ZN(n5229) );
  AOI22_X1 U6305 ( .A1(n6475), .A2(n5229), .B1(n5290), .B2(n5308), .ZN(n5117)
         );
  OAI211_X1 U6306 ( .C1(n5119), .C2(n5142), .A(n5118), .B(n5117), .ZN(U3095)
         );
  AOI22_X1 U6307 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5139), .B1(n6506), 
        .B2(n5138), .ZN(n5121) );
  AOI22_X1 U6308 ( .A1(n6502), .A2(n5229), .B1(n5290), .B2(n5296), .ZN(n5120)
         );
  OAI211_X1 U6309 ( .C1(n5122), .C2(n5142), .A(n5121), .B(n5120), .ZN(U3099)
         );
  AOI22_X1 U6310 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5139), .B1(n6497), 
        .B2(n5138), .ZN(n5124) );
  AOI22_X1 U6311 ( .A1(n6495), .A2(n5229), .B1(n5290), .B2(n5302), .ZN(n5123)
         );
  OAI211_X1 U6312 ( .C1(n5125), .C2(n5142), .A(n5124), .B(n5123), .ZN(U3098)
         );
  AOI22_X1 U6313 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5139), .B1(n6491), 
        .B2(n5138), .ZN(n5127) );
  AOI22_X1 U6314 ( .A1(n6489), .A2(n5229), .B1(n5290), .B2(n5314), .ZN(n5126)
         );
  OAI211_X1 U6315 ( .C1(n5128), .C2(n5142), .A(n5127), .B(n5126), .ZN(U3097)
         );
  AOI22_X1 U6316 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5139), .B1(n6484), 
        .B2(n5138), .ZN(n5130) );
  AOI22_X1 U6317 ( .A1(n6414), .A2(n5229), .B1(n5290), .B2(n6482), .ZN(n5129)
         );
  OAI211_X1 U6318 ( .C1(n5131), .C2(n5142), .A(n5130), .B(n5129), .ZN(U3096)
         );
  AOI22_X1 U6319 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5139), .B1(n6459), 
        .B2(n5138), .ZN(n5133) );
  AOI22_X1 U6320 ( .A1(n6404), .A2(n5229), .B1(n5290), .B2(n6444), .ZN(n5132)
         );
  OAI211_X1 U6321 ( .C1(n5134), .C2(n5142), .A(n5133), .B(n5132), .ZN(U3092)
         );
  AOI22_X1 U6322 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5139), .B1(n6471), 
        .B2(n5138), .ZN(n5136) );
  AOI22_X1 U6323 ( .A1(n6469), .A2(n5229), .B1(n5290), .B2(n6435), .ZN(n5135)
         );
  OAI211_X1 U6324 ( .C1(n5137), .C2(n5142), .A(n5136), .B(n5135), .ZN(U3094)
         );
  AOI22_X1 U6325 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5139), .B1(n6465), 
        .B2(n5138), .ZN(n5141) );
  AOI22_X1 U6326 ( .A1(n6463), .A2(n5229), .B1(n5290), .B2(n6430), .ZN(n5140)
         );
  OAI211_X1 U6327 ( .C1(n5143), .C2(n5142), .A(n5141), .B(n5140), .ZN(U3093)
         );
  INV_X1 U6328 ( .A(n6092), .ZN(n5178) );
  OAI21_X1 U6329 ( .B1(n5178), .B2(n5186), .A(n5923), .ZN(n5144) );
  NAND2_X1 U6330 ( .A1(n5144), .A2(REIP_REG_2__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6331 ( .A1(n6118), .A2(n6134), .ZN(n5153) );
  AOI22_X1 U6332 ( .A1(n6112), .A2(n6164), .B1(n6139), .B2(n4464), .ZN(n5150)
         );
  INV_X1 U6333 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6334 ( .A1(n6092), .A2(n5153), .ZN(n6124) );
  AOI22_X1 U6335 ( .A1(n6081), .A2(n5146), .B1(REIP_REG_3__SCAN_IN), .B2(n6124), .ZN(n5149) );
  NAND2_X1 U6336 ( .A1(n6133), .A2(n6167), .ZN(n5148) );
  NAND2_X1 U6337 ( .A1(n6126), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5147)
         );
  NAND4_X1 U6338 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n5151)
         );
  AOI21_X1 U6339 ( .B1(EBX_REG_3__SCAN_IN), .B2(n6125), .A(n5151), .ZN(n5152)
         );
  OAI21_X1 U6340 ( .B1(n5176), .B2(n5153), .A(n5152), .ZN(U2824) );
  XNOR2_X1 U6341 ( .A(n5892), .B(n6360), .ZN(n5155) );
  XNOR2_X1 U6342 ( .A(n5154), .B(n5155), .ZN(n6354) );
  NAND2_X1 U6343 ( .A1(n6354), .A2(n6320), .ZN(n5158) );
  NAND2_X1 U6344 ( .A1(n6375), .A2(REIP_REG_9__SCAN_IN), .ZN(n6350) );
  OAI21_X1 U6345 ( .B1(n6304), .B2(n6075), .A(n6350), .ZN(n5156) );
  AOI21_X1 U6346 ( .B1(n6298), .B2(n6080), .A(n5156), .ZN(n5157) );
  OAI211_X1 U6347 ( .C1(n6325), .C2(n6079), .A(n5158), .B(n5157), .ZN(U2977)
         );
  OAI22_X1 U6348 ( .A1(n6130), .A2(n5160), .B1(n6146), .B2(n5159), .ZN(n5165)
         );
  AOI22_X1 U6349 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6126), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6074), .ZN(n5161) );
  OAI211_X1 U6350 ( .C1(n5163), .C2(n5162), .A(n5161), .B(n6128), .ZN(n5164)
         );
  AOI211_X1 U6351 ( .C1(EBX_REG_8__SCAN_IN), .C2(n6125), .A(n5165), .B(n5164), 
        .ZN(n5166) );
  OAI21_X1 U6352 ( .B1(n5167), .B2(n6100), .A(n5166), .ZN(U2819) );
  INV_X1 U6353 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6739) );
  OAI21_X1 U6354 ( .B1(n6137), .B2(n5186), .A(n6739), .ZN(n5175) );
  NAND2_X1 U6355 ( .A1(n6125), .A2(EBX_REG_2__SCAN_IN), .ZN(n5173) );
  AOI22_X1 U6356 ( .A1(n6112), .A2(n6376), .B1(n6133), .B2(n6308), .ZN(n5172)
         );
  INV_X1 U6357 ( .A(n6311), .ZN(n5168) );
  AOI22_X1 U6358 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6126), .B1(n6081), 
        .B2(n5168), .ZN(n5171) );
  INV_X1 U6359 ( .A(n4466), .ZN(n5169) );
  NAND2_X1 U6360 ( .A1(n6139), .A2(n5169), .ZN(n5170) );
  NAND4_X1 U6361 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n5174)
         );
  AOI21_X1 U6362 ( .B1(n5176), .B2(n5175), .A(n5174), .ZN(n5177) );
  INV_X1 U6363 ( .A(n5177), .ZN(U2825) );
  INV_X1 U6364 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6365 ( .A1(n6133), .A2(n6313), .ZN(n5180) );
  AOI22_X1 U6366 ( .A1(n6081), .A2(n5181), .B1(n5178), .B2(REIP_REG_1__SCAN_IN), .ZN(n5179) );
  OAI211_X1 U6367 ( .C1(n5181), .C2(n6106), .A(n5180), .B(n5179), .ZN(n5185)
         );
  INV_X1 U6368 ( .A(n6139), .ZN(n5183) );
  OAI22_X1 U6369 ( .A1(n5183), .A2(n5907), .B1(n5182), .B2(n6130), .ZN(n5184)
         );
  AOI211_X1 U6370 ( .C1(n6118), .C2(n5186), .A(n5185), .B(n5184), .ZN(n5187)
         );
  OAI21_X1 U6371 ( .B1(n6123), .B2(n4203), .A(n5187), .ZN(U2826) );
  XOR2_X1 U6372 ( .A(n5188), .B(n6065), .Z(n5282) );
  AOI22_X1 U6373 ( .A1(n6183), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6179), .ZN(n5189) );
  OAI21_X1 U6374 ( .B1(n5198), .B2(n5951), .A(n5189), .ZN(U2879) );
  XOR2_X1 U6375 ( .A(n5355), .B(n5356), .Z(n6331) );
  AOI22_X1 U6376 ( .A1(n6165), .A2(n6331), .B1(EBX_REG_12__SCAN_IN), .B2(n5663), .ZN(n5190) );
  OAI21_X1 U6377 ( .B1(n5198), .B2(n6148), .A(n5190), .ZN(U2847) );
  INV_X1 U6378 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5192) );
  OAI21_X1 U6379 ( .B1(n6137), .B2(n5195), .A(n6092), .ZN(n6063) );
  AOI22_X1 U6380 ( .A1(n6112), .A2(n6331), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6063), .ZN(n5191) );
  OAI211_X1 U6381 ( .C1(n6106), .C2(n5192), .A(n5191), .B(n6128), .ZN(n5194)
         );
  NOR2_X1 U6382 ( .A1(n6146), .A2(n5280), .ZN(n5193) );
  AOI211_X1 U6383 ( .C1(EBX_REG_12__SCAN_IN), .C2(n6125), .A(n5194), .B(n5193), 
        .ZN(n5197) );
  NOR2_X1 U6384 ( .A1(n6137), .A2(REIP_REG_12__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U6385 ( .A1(n6057), .A2(n5195), .ZN(n5196) );
  OAI211_X1 U6386 ( .C1(n5198), .C2(n6100), .A(n5197), .B(n5196), .ZN(U2815)
         );
  INV_X1 U6387 ( .A(n5200), .ZN(n5202) );
  NOR2_X1 U6388 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  XNOR2_X1 U6389 ( .A(n3105), .B(n5203), .ZN(n6347) );
  INV_X1 U6390 ( .A(n6347), .ZN(n5209) );
  AOI22_X1 U6391 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6375), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5204) );
  OAI21_X1 U6392 ( .B1(n5205), .B2(n6318), .A(n5204), .ZN(n5206) );
  AOI21_X1 U6393 ( .B1(n5207), .B2(n6314), .A(n5206), .ZN(n5208) );
  OAI21_X1 U6394 ( .B1(n5209), .B2(n6284), .A(n5208), .ZN(U2976) );
  INV_X1 U6395 ( .A(n5211), .ZN(n5212) );
  NOR2_X1 U6396 ( .A1(n5213), .A2(n5212), .ZN(n5214) );
  XNOR2_X1 U6397 ( .A(n5210), .B(n5214), .ZN(n6285) );
  AOI22_X1 U6398 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6328), .B1(n6327), .B2(n5215), .ZN(n5220) );
  AND2_X1 U6399 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NOR2_X1 U6400 ( .A1(n5356), .A2(n5218), .ZN(n6158) );
  AOI22_X1 U6401 ( .A1(n6377), .A2(n6158), .B1(n6375), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5219) );
  OAI211_X1 U6402 ( .C1(n6285), .C2(n6370), .A(n5220), .B(n5219), .ZN(U3007)
         );
  NAND2_X1 U6403 ( .A1(n5221), .A2(n4464), .ZN(n5230) );
  NAND2_X1 U6404 ( .A1(n5262), .A2(n6447), .ZN(n5223) );
  OAI21_X1 U6405 ( .B1(n5229), .B2(n5223), .A(n5222), .ZN(n5228) );
  NOR2_X1 U6406 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5224), .ZN(n5265)
         );
  INV_X1 U6407 ( .A(n6391), .ZN(n5226) );
  OAI211_X1 U6408 ( .C1(n6959), .C2(n5265), .A(n5226), .B(n5225), .ZN(n5227)
         );
  INV_X1 U6409 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5237) );
  INV_X1 U6410 ( .A(n5229), .ZN(n5263) );
  OR2_X1 U6411 ( .A1(n5230), .A2(n6452), .ZN(n5233) );
  NAND2_X1 U6412 ( .A1(n6400), .A2(n5231), .ZN(n5232) );
  NAND2_X1 U6413 ( .A1(n5233), .A2(n5232), .ZN(n5266) );
  AOI22_X1 U6414 ( .A1(n6434), .A2(n6495), .B1(n6497), .B2(n5266), .ZN(n5234)
         );
  OAI21_X1 U6415 ( .B1(n5263), .B2(n6500), .A(n5234), .ZN(n5235) );
  AOI21_X1 U6416 ( .B1(n6496), .B2(n5265), .A(n5235), .ZN(n5236) );
  OAI21_X1 U6417 ( .B1(n5270), .B2(n5237), .A(n5236), .ZN(U3090) );
  INV_X1 U6418 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5241) );
  AOI22_X1 U6419 ( .A1(n6434), .A2(n6489), .B1(n6491), .B2(n5266), .ZN(n5238)
         );
  OAI21_X1 U6420 ( .B1(n5263), .B2(n6494), .A(n5238), .ZN(n5239) );
  AOI21_X1 U6421 ( .B1(n6490), .B2(n5265), .A(n5239), .ZN(n5240) );
  OAI21_X1 U6422 ( .B1(n5270), .B2(n5241), .A(n5240), .ZN(U3089) );
  INV_X1 U6423 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5245) );
  AOI22_X1 U6424 ( .A1(n6434), .A2(n6475), .B1(n6477), .B2(n5266), .ZN(n5242)
         );
  OAI21_X1 U6425 ( .B1(n5263), .B2(n6480), .A(n5242), .ZN(n5243) );
  AOI21_X1 U6426 ( .B1(n6476), .B2(n5265), .A(n5243), .ZN(n5244) );
  OAI21_X1 U6427 ( .B1(n5270), .B2(n5245), .A(n5244), .ZN(U3087) );
  INV_X1 U6428 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5249) );
  OAI22_X1 U6429 ( .A1(n5263), .A2(n6474), .B1(n6442), .B2(n5262), .ZN(n5246)
         );
  AOI21_X1 U6430 ( .B1(n6470), .B2(n5265), .A(n5246), .ZN(n5248) );
  NAND2_X1 U6431 ( .A1(n6471), .A2(n5266), .ZN(n5247) );
  OAI211_X1 U6432 ( .C1(n5270), .C2(n5249), .A(n5248), .B(n5247), .ZN(U3086)
         );
  INV_X1 U6433 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5253) );
  OAI22_X1 U6434 ( .A1(n5263), .A2(n6417), .B1(n6488), .B2(n5262), .ZN(n5250)
         );
  AOI21_X1 U6435 ( .B1(n6483), .B2(n5265), .A(n5250), .ZN(n5252) );
  NAND2_X1 U6436 ( .A1(n6484), .A2(n5266), .ZN(n5251) );
  OAI211_X1 U6437 ( .C1(n5270), .C2(n5253), .A(n5252), .B(n5251), .ZN(U3088)
         );
  INV_X1 U6438 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5257) );
  OAI22_X1 U6439 ( .A1(n5263), .A2(n6468), .B1(n6433), .B2(n5262), .ZN(n5254)
         );
  AOI21_X1 U6440 ( .B1(n6464), .B2(n5265), .A(n5254), .ZN(n5256) );
  NAND2_X1 U6441 ( .A1(n6465), .A2(n5266), .ZN(n5255) );
  OAI211_X1 U6442 ( .C1(n5270), .C2(n5257), .A(n5256), .B(n5255), .ZN(U3085)
         );
  INV_X1 U6443 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5261) );
  OAI22_X1 U6444 ( .A1(n5263), .A2(n6407), .B1(n6462), .B2(n5262), .ZN(n5258)
         );
  AOI21_X1 U6445 ( .B1(n6445), .B2(n5265), .A(n5258), .ZN(n5260) );
  NAND2_X1 U6446 ( .A1(n6459), .A2(n5266), .ZN(n5259) );
  OAI211_X1 U6447 ( .C1(n5270), .C2(n5261), .A(n5260), .B(n5259), .ZN(U3084)
         );
  INV_X1 U6448 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5269) );
  OAI22_X1 U6449 ( .A1(n5263), .A2(n6511), .B1(n5298), .B2(n5262), .ZN(n5264)
         );
  AOI21_X1 U6450 ( .B1(n6504), .B2(n5265), .A(n5264), .ZN(n5268) );
  NAND2_X1 U6451 ( .A1(n6506), .A2(n5266), .ZN(n5267) );
  OAI211_X1 U6452 ( .C1(n5270), .C2(n5269), .A(n5268), .B(n5267), .ZN(U3091)
         );
  OAI21_X1 U6453 ( .B1(n5273), .B2(n5272), .A(n5271), .ZN(n6154) );
  AOI22_X1 U6454 ( .A1(n6183), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6179), .ZN(n5274) );
  OAI21_X1 U6455 ( .B1(n6154), .B2(n5951), .A(n5274), .ZN(U2878) );
  NAND2_X1 U6456 ( .A1(n5276), .A2(n5275), .ZN(n5278) );
  XOR2_X1 U6457 ( .A(n5278), .B(n5277), .Z(n6332) );
  INV_X1 U6458 ( .A(n6332), .ZN(n5284) );
  AOI22_X1 U6459 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6375), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5279) );
  OAI21_X1 U6460 ( .B1(n5280), .B2(n6318), .A(n5279), .ZN(n5281) );
  AOI21_X1 U6461 ( .B1(n5282), .B2(n6314), .A(n5281), .ZN(n5283) );
  OAI21_X1 U6462 ( .B1(n5284), .B2(n6284), .A(n5283), .ZN(U2974) );
  OR2_X1 U6463 ( .A1(n6501), .A2(n5290), .ZN(n5286) );
  AOI21_X1 U6464 ( .B1(n5286), .B2(STATEBS16_REG_SCAN_IN), .A(n6452), .ZN(
        n5293) );
  INV_X1 U6465 ( .A(n5287), .ZN(n5288) );
  NAND3_X1 U6466 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6526), .ZN(n6456) );
  NOR2_X1 U6467 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6456), .ZN(n5336)
         );
  INV_X1 U6468 ( .A(n6450), .ZN(n5292) );
  INV_X1 U6469 ( .A(n5336), .ZN(n5291) );
  AOI22_X1 U6470 ( .A1(n5293), .A2(n5292), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5291), .ZN(n5294) );
  OAI211_X1 U6471 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6455), .A(n5295), .B(n5294), .ZN(n5332) );
  AOI22_X1 U6472 ( .A1(n6501), .A2(n5296), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5332), .ZN(n5297) );
  OAI21_X1 U6473 ( .B1(n5334), .B2(n5298), .A(n5297), .ZN(n5299) );
  AOI21_X1 U6474 ( .B1(n6504), .B2(n5336), .A(n5299), .ZN(n5300) );
  OAI21_X1 U6475 ( .B1(n5301), .B2(n5338), .A(n5300), .ZN(U3107) );
  AOI22_X1 U6476 ( .A1(n6501), .A2(n5302), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5332), .ZN(n5303) );
  OAI21_X1 U6477 ( .B1(n5334), .B2(n5304), .A(n5303), .ZN(n5305) );
  AOI21_X1 U6478 ( .B1(n6496), .B2(n5336), .A(n5305), .ZN(n5306) );
  OAI21_X1 U6479 ( .B1(n5338), .B2(n5307), .A(n5306), .ZN(U3106) );
  AOI22_X1 U6480 ( .A1(n6501), .A2(n5308), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5332), .ZN(n5309) );
  OAI21_X1 U6481 ( .B1(n5334), .B2(n5310), .A(n5309), .ZN(n5311) );
  AOI21_X1 U6482 ( .B1(n6476), .B2(n5336), .A(n5311), .ZN(n5312) );
  OAI21_X1 U6483 ( .B1(n5338), .B2(n5313), .A(n5312), .ZN(U3103) );
  AOI22_X1 U6484 ( .A1(n6501), .A2(n5314), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5332), .ZN(n5315) );
  OAI21_X1 U6485 ( .B1(n5334), .B2(n5316), .A(n5315), .ZN(n5317) );
  AOI21_X1 U6486 ( .B1(n6490), .B2(n5336), .A(n5317), .ZN(n5318) );
  OAI21_X1 U6487 ( .B1(n5338), .B2(n5319), .A(n5318), .ZN(U3105) );
  AOI22_X1 U6488 ( .A1(n6501), .A2(n6435), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5332), .ZN(n5320) );
  OAI21_X1 U6489 ( .B1(n5334), .B2(n6442), .A(n5320), .ZN(n5321) );
  AOI21_X1 U6490 ( .B1(n6470), .B2(n5336), .A(n5321), .ZN(n5322) );
  OAI21_X1 U6491 ( .B1(n5323), .B2(n5338), .A(n5322), .ZN(U3102) );
  AOI22_X1 U6492 ( .A1(n6501), .A2(n6482), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5332), .ZN(n5324) );
  OAI21_X1 U6493 ( .B1(n5334), .B2(n6488), .A(n5324), .ZN(n5325) );
  AOI21_X1 U6494 ( .B1(n6483), .B2(n5336), .A(n5325), .ZN(n5326) );
  OAI21_X1 U6495 ( .B1(n5327), .B2(n5338), .A(n5326), .ZN(U3104) );
  AOI22_X1 U6496 ( .A1(n6501), .A2(n6430), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5332), .ZN(n5328) );
  OAI21_X1 U6497 ( .B1(n5334), .B2(n6433), .A(n5328), .ZN(n5329) );
  AOI21_X1 U6498 ( .B1(n6464), .B2(n5336), .A(n5329), .ZN(n5330) );
  OAI21_X1 U6499 ( .B1(n5331), .B2(n5338), .A(n5330), .ZN(U3101) );
  AOI22_X1 U6500 ( .A1(n6501), .A2(n6444), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5332), .ZN(n5333) );
  OAI21_X1 U6501 ( .B1(n5334), .B2(n6462), .A(n5333), .ZN(n5335) );
  AOI21_X1 U6502 ( .B1(n6445), .B2(n5336), .A(n5335), .ZN(n5337) );
  OAI21_X1 U6503 ( .B1(n5339), .B2(n5338), .A(n5337), .ZN(U3100) );
  OAI21_X1 U6504 ( .B1(n5340), .B2(n5342), .A(n5341), .ZN(n5976) );
  INV_X1 U6505 ( .A(n5976), .ZN(n5364) );
  INV_X1 U6506 ( .A(n5353), .ZN(n5343) );
  OR3_X1 U6507 ( .A1(n5345), .A2(n5344), .A3(n5343), .ZN(n5346) );
  AOI211_X1 U6508 ( .C1(n5347), .C2(n5346), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n6330), .ZN(n5350) );
  AOI211_X1 U6509 ( .C1(n5348), .C2(n6330), .A(n5350), .B(n6328), .ZN(n5349)
         );
  OAI21_X1 U6510 ( .B1(n5998), .B2(n5359), .A(n5349), .ZN(n5997) );
  OAI21_X1 U6511 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5350), .A(n5997), 
        .ZN(n5363) );
  INV_X1 U6512 ( .A(n6330), .ZN(n5351) );
  NAND3_X1 U6513 ( .A1(n5353), .A2(n5352), .A3(n5351), .ZN(n5360) );
  AOI21_X1 U6514 ( .B1(n5356), .B2(n5355), .A(n5354), .ZN(n5357) );
  OR2_X1 U6515 ( .A1(n5669), .A2(n5357), .ZN(n6152) );
  OR2_X1 U6516 ( .A1(n6352), .A2(n6152), .ZN(n5358) );
  NAND2_X1 U6517 ( .A1(n6375), .A2(REIP_REG_13__SCAN_IN), .ZN(n5977) );
  OAI211_X1 U6518 ( .C1(n5360), .C2(n5359), .A(n5358), .B(n5977), .ZN(n5361)
         );
  INV_X1 U6519 ( .A(n5361), .ZN(n5362) );
  OAI211_X1 U6520 ( .C1(n5364), .C2(n6370), .A(n5363), .B(n5362), .ZN(U3005)
         );
  AOI22_X1 U6521 ( .A1(n6518), .A2(n6543), .B1(FLUSH_REG_SCAN_IN), .B2(n6561), 
        .ZN(n6002) );
  NAND2_X1 U6522 ( .A1(n6002), .A2(n6637), .ZN(n6649) );
  INV_X1 U6523 ( .A(n6649), .ZN(n6643) );
  AOI21_X1 U6524 ( .B1(n5365), .B2(n5460), .A(n6643), .ZN(n5371) );
  INV_X1 U6525 ( .A(n5366), .ZN(n5369) );
  INV_X1 U6526 ( .A(n6651), .ZN(n6004) );
  INV_X1 U6527 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5380) );
  AOI22_X1 U6528 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5380), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6836), .ZN(n5458) );
  NAND2_X1 U6529 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5453) );
  NAND3_X1 U6530 ( .A1(n4606), .A2(n3379), .A3(n5460), .ZN(n5367) );
  OAI21_X1 U6531 ( .B1(n5458), .B2(n5453), .A(n5367), .ZN(n5368) );
  AOI21_X1 U6532 ( .B1(n5369), .B2(n6004), .A(n5368), .ZN(n5370) );
  OAI22_X1 U6533 ( .A1(n5371), .A2(n3379), .B1(n5370), .B2(n6643), .ZN(U3459)
         );
  NAND2_X1 U6534 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5376) );
  INV_X1 U6535 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5373) );
  NAND4_X1 U6536 ( .A1(n5718), .A2(n5807), .A3(n5373), .A4(n5447), .ZN(n5374)
         );
  OR2_X1 U6537 ( .A1(n5372), .A2(n5374), .ZN(n5375) );
  XNOR2_X1 U6538 ( .A(n5377), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5432)
         );
  AOI21_X1 U6539 ( .B1(n5447), .B2(n6339), .A(n5378), .ZN(n5438) );
  OAI21_X1 U6540 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5379), .A(n5438), 
        .ZN(n5394) );
  NAND3_X1 U6541 ( .A1(n5380), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5381) );
  NOR2_X1 U6542 ( .A1(n5448), .A2(n5381), .ZN(n5393) );
  NOR2_X1 U6543 ( .A1(n4430), .A2(EBX_REG_29__SCAN_IN), .ZN(n5382) );
  OR3_X2 U6544 ( .A1(n5388), .A2(n5383), .A3(n5382), .ZN(n5442) );
  NAND2_X1 U6545 ( .A1(n5442), .A2(n5384), .ZN(n5439) );
  NAND2_X1 U6546 ( .A1(n5390), .A2(EBX_REG_30__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6547 ( .A1(n4430), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6548 ( .A1(n5386), .A2(n5385), .ZN(n5441) );
  OR3_X1 U6549 ( .A1(n5388), .A2(n5441), .A3(n5387), .ZN(n5389) );
  NAND2_X1 U6550 ( .A1(n5439), .A2(n5389), .ZN(n5392) );
  AOI22_X1 U6551 ( .A1(n5390), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4430), .ZN(n5391) );
  NAND2_X1 U6552 ( .A1(n6375), .A2(REIP_REG_31__SCAN_IN), .ZN(n5428) );
  AOI22_X1 U6553 ( .A1(n3096), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5395), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5402) );
  AOI22_X1 U6554 ( .A1(n5397), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5396), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5401) );
  AOI22_X1 U6555 ( .A1(n3111), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5400) );
  AOI22_X1 U6556 ( .A1(n3113), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5398), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5399) );
  NAND4_X1 U6557 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n5410)
         );
  AOI22_X1 U6558 ( .A1(n3115), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3095), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5408) );
  AOI22_X1 U6559 ( .A1(n4094), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4135), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5407) );
  AOI22_X1 U6560 ( .A1(n3311), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3574), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5406) );
  AOI22_X1 U6561 ( .A1(n5404), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3093), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5405) );
  NAND4_X1 U6562 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n5409)
         );
  NOR2_X1 U6563 ( .A1(n5410), .A2(n5409), .ZN(n5414) );
  NOR2_X1 U6564 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  XOR2_X1 U6565 ( .A(n5414), .B(n5413), .Z(n5421) );
  NAND2_X1 U6566 ( .A1(n6455), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5415)
         );
  NAND2_X1 U6567 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  AOI21_X1 U6568 ( .B1(n5418), .B2(EAX_REG_30__SCAN_IN), .A(n5417), .ZN(n5419)
         );
  OAI21_X1 U6569 ( .B1(n5421), .B2(n5420), .A(n5419), .ZN(n5424) );
  XNOR2_X1 U6570 ( .A(n5422), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5478)
         );
  NAND2_X1 U6571 ( .A1(n5478), .A2(n4344), .ZN(n5423) );
  NAND2_X1 U6572 ( .A1(n5424), .A2(n5423), .ZN(n5464) );
  AOI22_X1 U6573 ( .A1(n3725), .A2(EAX_REG_31__SCAN_IN), .B1(n5425), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6574 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5427)
         );
  OAI211_X1 U6575 ( .C1(n6318), .C2(n5429), .A(n5428), .B(n5427), .ZN(n5430)
         );
  AOI21_X1 U6576 ( .B1(n5673), .B2(n6314), .A(n5430), .ZN(n5431) );
  OAI21_X1 U6577 ( .B1(n5432), .B2(n6284), .A(n5431), .ZN(U2955) );
  INV_X1 U6578 ( .A(n5433), .ZN(n5436) );
  NAND2_X1 U6579 ( .A1(n5434), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6580 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  XNOR2_X1 U6581 ( .A(n5437), .B(n5373), .ZN(n5475) );
  INV_X1 U6582 ( .A(n5438), .ZN(n5451) );
  INV_X1 U6583 ( .A(n5442), .ZN(n5440) );
  OAI211_X1 U6584 ( .C1(n5440), .C2(n5388), .A(n5439), .B(n5441), .ZN(n5446)
         );
  INV_X1 U6585 ( .A(n5388), .ZN(n5444) );
  INV_X1 U6586 ( .A(n5441), .ZN(n5443) );
  OAI211_X1 U6587 ( .C1(n5444), .C2(n5384), .A(n5443), .B(n5442), .ZN(n5445)
         );
  NAND2_X1 U6588 ( .A1(n5446), .A2(n5445), .ZN(n5488) );
  NAND2_X1 U6589 ( .A1(n6375), .A2(REIP_REG_30__SCAN_IN), .ZN(n5466) );
  OAI21_X1 U6590 ( .B1(n5488), .B2(n6352), .A(n5466), .ZN(n5450) );
  NOR3_X1 U6591 ( .A1(n5448), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5447), 
        .ZN(n5449) );
  AOI211_X1 U6592 ( .C1(n5451), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5450), .B(n5449), .ZN(n5452) );
  OAI21_X1 U6593 ( .B1(n5475), .B2(n6370), .A(n5452), .ZN(U2988) );
  OAI21_X1 U6594 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6640), .A(n6649), 
        .ZN(n6647) );
  INV_X1 U6595 ( .A(n6647), .ZN(n5463) );
  INV_X1 U6596 ( .A(n5453), .ZN(n5457) );
  NOR3_X1 U6597 ( .A1(n5454), .A2(n4645), .A3(n4606), .ZN(n5455) );
  AOI21_X1 U6598 ( .B1(n6517), .B2(n5462), .A(n5455), .ZN(n5456) );
  OAI21_X1 U6599 ( .B1(n5907), .B2(n6512), .A(n5456), .ZN(n6519) );
  AOI222_X1 U6600 ( .A1(n5460), .A2(n5459), .B1(n5458), .B2(n5457), .C1(n6519), 
        .C2(n6004), .ZN(n5461) );
  OAI22_X1 U6601 ( .A1(n5463), .A2(n5462), .B1(n6643), .B2(n5461), .ZN(U3460)
         );
  XNOR2_X2 U6602 ( .A(n5465), .B(n5464), .ZN(n5476) );
  INV_X1 U6603 ( .A(n5478), .ZN(n5470) );
  OAI21_X1 U6604 ( .B1(n6304), .B2(n5467), .A(n5466), .ZN(n5468) );
  INV_X1 U6605 ( .A(n5468), .ZN(n5469) );
  INV_X1 U6606 ( .A(n5471), .ZN(n5472) );
  INV_X1 U6607 ( .A(n5473), .ZN(n5474) );
  OAI21_X1 U6608 ( .B1(n5475), .B2(n6284), .A(n5474), .ZN(U2956) );
  NOR2_X1 U6609 ( .A1(n5477), .A2(n5507), .ZN(n5490) );
  INV_X1 U6610 ( .A(n5490), .ZN(n5484) );
  AOI22_X1 U6611 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6126), .B1(n6081), 
        .B2(n5478), .ZN(n5480) );
  NAND2_X1 U6612 ( .A1(n6125), .A2(EBX_REG_30__SCAN_IN), .ZN(n5479) );
  OAI211_X1 U6613 ( .C1(n5488), .C2(n6130), .A(n5480), .B(n5479), .ZN(n5483)
         );
  INV_X1 U6614 ( .A(n5481), .ZN(n5493) );
  NOR3_X1 U6615 ( .A1(n5493), .A2(REIP_REG_30__SCAN_IN), .A3(n6624), .ZN(n5482) );
  AOI211_X1 U6616 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5484), .A(n5483), .B(n5482), .ZN(n5485) );
  OAI21_X1 U6617 ( .B1(n5476), .B2(n6100), .A(n5485), .ZN(U2797) );
  AOI22_X1 U6618 ( .A1(n6177), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6179), .ZN(n5487) );
  NAND2_X1 U6619 ( .A1(n6180), .A2(DATAI_14_), .ZN(n5486) );
  OAI211_X1 U6620 ( .C1(n5476), .C2(n5951), .A(n5487), .B(n5486), .ZN(U2861)
         );
  INV_X1 U6621 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5489) );
  OAI222_X1 U6622 ( .A1(n6148), .A2(n5476), .B1(n5489), .B2(n6170), .C1(n5488), 
        .C2(n6153), .ZN(U2829) );
  INV_X1 U6623 ( .A(n5673), .ZN(n5498) );
  OAI21_X1 U6624 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6137), .A(n5490), .ZN(n5496) );
  AOI22_X1 U6625 ( .A1(n5491), .A2(EBX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n6126), .ZN(n5492) );
  OAI21_X1 U6626 ( .B1(n5618), .B2(n6130), .A(n5492), .ZN(n5495) );
  INV_X1 U6627 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6968) );
  NOR4_X1 U6628 ( .A1(n5493), .A2(REIP_REG_31__SCAN_IN), .A3(n6968), .A4(n6624), .ZN(n5494) );
  OAI21_X1 U6629 ( .B1(n5498), .B2(n6100), .A(n5497), .ZN(U2796) );
  INV_X1 U6630 ( .A(n5707), .ZN(n5680) );
  OR2_X1 U6631 ( .A1(n5516), .A2(n5501), .ZN(n5502) );
  NAND2_X1 U6632 ( .A1(n5388), .A2(n5502), .ZN(n5803) );
  OAI22_X1 U6633 ( .A1(n6688), .A2(n6106), .B1(n6146), .B2(n5705), .ZN(n5503)
         );
  AOI21_X1 U6634 ( .B1(EBX_REG_28__SCAN_IN), .B2(n6125), .A(n5503), .ZN(n5504)
         );
  OAI21_X1 U6635 ( .B1(n5803), .B2(n6130), .A(n5504), .ZN(n5506) );
  INV_X1 U6636 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6621) );
  NOR3_X1 U6637 ( .A1(n5523), .A2(REIP_REG_28__SCAN_IN), .A3(n6621), .ZN(n5505) );
  AOI211_X1 U6638 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5507), .A(n5506), .B(n5505), .ZN(n5508) );
  OAI21_X1 U6639 ( .B1(n5680), .B2(n6100), .A(n5508), .ZN(U2799) );
  INV_X1 U6640 ( .A(n5713), .ZN(n5511) );
  NAND2_X1 U6641 ( .A1(n5511), .A2(n6091), .ZN(n5522) );
  INV_X1 U6642 ( .A(n5512), .ZN(n5528) );
  INV_X1 U6643 ( .A(n5513), .ZN(n5514) );
  AOI21_X1 U6644 ( .B1(n5538), .B2(n5528), .A(n5514), .ZN(n5515) );
  OR2_X1 U6645 ( .A1(n5516), .A2(n5515), .ZN(n5815) );
  AOI22_X1 U6646 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6126), .B1(n6081), 
        .B2(n5716), .ZN(n5518) );
  NAND2_X1 U6647 ( .A1(n6125), .A2(EBX_REG_27__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U6648 ( .C1(n5815), .C2(n6130), .A(n5518), .B(n5517), .ZN(n5520)
         );
  NOR2_X1 U6649 ( .A1(n5534), .A2(n6621), .ZN(n5519) );
  NOR2_X1 U6650 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  OAI211_X1 U6651 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5523), .A(n5522), .B(n5521), .ZN(U2800) );
  INV_X1 U6652 ( .A(n5543), .ZN(n5524) );
  AOI21_X1 U6653 ( .B1(n5524), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5533) );
  AOI21_X1 U6654 ( .B1(n5527), .B2(n5526), .A(n5525), .ZN(n5727) );
  NAND2_X1 U6655 ( .A1(n5727), .A2(n6091), .ZN(n5532) );
  OAI22_X1 U6656 ( .A1(n6863), .A2(n6106), .B1(n6146), .B2(n5725), .ZN(n5530)
         );
  XNOR2_X1 U6657 ( .A(n5538), .B(n5528), .ZN(n5823) );
  NOR2_X1 U6658 ( .A1(n5823), .A2(n6130), .ZN(n5529) );
  AOI211_X1 U6659 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6125), .A(n5530), .B(n5529), 
        .ZN(n5531) );
  OAI211_X1 U6660 ( .C1(n5534), .C2(n5533), .A(n5532), .B(n5531), .ZN(U2801)
         );
  XNOR2_X1 U6661 ( .A(n5536), .B(n5537), .ZN(n5735) );
  AOI21_X1 U6662 ( .B1(n5540), .B2(n5539), .A(n5538), .ZN(n5832) );
  AOI22_X1 U6663 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6126), .B1(n6081), 
        .B2(n5731), .ZN(n5541) );
  OAI21_X1 U6664 ( .B1(n6123), .B2(n5542), .A(n5541), .ZN(n5545) );
  NOR2_X1 U6665 ( .A1(n5543), .A2(REIP_REG_25__SCAN_IN), .ZN(n5544) );
  AOI211_X1 U6666 ( .C1(n5832), .C2(n6112), .A(n5545), .B(n5544), .ZN(n5549)
         );
  NAND2_X1 U6667 ( .A1(n5546), .A2(n6756), .ZN(n5917) );
  INV_X1 U6668 ( .A(n5917), .ZN(n5547) );
  OAI21_X1 U6669 ( .B1(n5547), .B2(n5914), .A(REIP_REG_25__SCAN_IN), .ZN(n5548) );
  OAI211_X1 U6670 ( .C1(n5735), .C2(n6100), .A(n5549), .B(n5548), .ZN(U2802)
         );
  INV_X1 U6671 ( .A(n5550), .ZN(n5635) );
  XOR2_X1 U6672 ( .A(n5551), .B(n5635), .Z(n5751) );
  NAND2_X1 U6673 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5927) );
  INV_X1 U6674 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6614) );
  OAI21_X1 U6675 ( .B1(n5927), .B2(n5941), .A(n6614), .ZN(n5560) );
  NAND2_X1 U6676 ( .A1(n5647), .A2(n5639), .ZN(n5554) );
  INV_X1 U6677 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U6678 ( .A1(n5554), .A2(n5553), .ZN(n5556) );
  NAND2_X1 U6679 ( .A1(n5556), .A2(n5555), .ZN(n5842) );
  INV_X1 U6680 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5632) );
  OAI22_X1 U6681 ( .A1(n6123), .A2(n5632), .B1(n5749), .B2(n6106), .ZN(n5557)
         );
  AOI21_X1 U6682 ( .B1(n6081), .B2(n5747), .A(n5557), .ZN(n5558) );
  OAI21_X1 U6683 ( .B1(n5842), .B2(n6130), .A(n5558), .ZN(n5559) );
  AOI21_X1 U6684 ( .B1(n5560), .B2(n5914), .A(n5559), .ZN(n5561) );
  OAI21_X1 U6685 ( .B1(n5690), .B2(n6100), .A(n5561), .ZN(U2804) );
  AOI21_X1 U6686 ( .B1(n5563), .B2(n3123), .A(n5650), .ZN(n5778) );
  INV_X1 U6687 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6606) );
  NOR3_X1 U6688 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6606), .A3(n5566), .ZN(n5576) );
  NOR2_X1 U6689 ( .A1(n5565), .A2(n5564), .ZN(n6035) );
  NOR2_X1 U6690 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5566), .ZN(n5584) );
  OAI21_X1 U6691 ( .B1(n6035), .B2(n5584), .A(REIP_REG_19__SCAN_IN), .ZN(n5574) );
  AOI22_X1 U6692 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6125), .B1(n5774), .B2(n6081), .ZN(n5573) );
  INV_X1 U6693 ( .A(n5582), .ZN(n5567) );
  NAND2_X1 U6694 ( .A1(n5898), .A2(n5567), .ZN(n5568) );
  NAND2_X1 U6695 ( .A1(n5568), .A2(n3137), .ZN(n5569) );
  NAND2_X1 U6696 ( .A1(n3126), .A2(n5569), .ZN(n5874) );
  NAND2_X1 U6697 ( .A1(n6126), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5570)
         );
  OAI211_X1 U6698 ( .C1(n5874), .C2(n6130), .A(n5570), .B(n6128), .ZN(n5571)
         );
  INV_X1 U6699 ( .A(n5571), .ZN(n5572) );
  NAND3_X1 U6700 ( .A1(n5574), .A2(n5573), .A3(n5572), .ZN(n5575) );
  AOI211_X1 U6701 ( .C1(n5778), .C2(n6091), .A(n5576), .B(n5575), .ZN(n5577)
         );
  INV_X1 U6702 ( .A(n5577), .ZN(U2808) );
  NAND2_X1 U6703 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  NAND2_X1 U6704 ( .A1(n6171), .A2(n6091), .ZN(n5588) );
  INV_X1 U6705 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6802) );
  INV_X1 U6706 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6865) );
  OAI22_X1 U6707 ( .A1(n6123), .A2(n6802), .B1(n6865), .B2(n6106), .ZN(n5581)
         );
  AOI211_X1 U6708 ( .C1(n6035), .C2(REIP_REG_18__SCAN_IN), .A(n6113), .B(n5581), .ZN(n5587) );
  XNOR2_X1 U6709 ( .A(n5898), .B(n5582), .ZN(n5890) );
  INV_X1 U6710 ( .A(n5969), .ZN(n5583) );
  AOI22_X1 U6711 ( .A1(n5890), .A2(n6112), .B1(n5583), .B2(n6081), .ZN(n5586)
         );
  INV_X1 U6712 ( .A(n5584), .ZN(n5585) );
  NAND4_X1 U6713 ( .A1(n5588), .A2(n5587), .A3(n5586), .A4(n5585), .ZN(U2809)
         );
  AOI22_X1 U6714 ( .A1(n5611), .A2(n6599), .B1(n5923), .B2(n5615), .ZN(n5604)
         );
  AND2_X1 U6715 ( .A1(n5589), .A2(n5665), .ZN(n5591) );
  NAND2_X1 U6716 ( .A1(n5589), .A2(n5665), .ZN(n5666) );
  OR2_X1 U6717 ( .A1(n5666), .A2(n5607), .ZN(n5605) );
  AND2_X1 U6718 ( .A1(n5605), .A2(n5592), .ZN(n5593) );
  NAND2_X1 U6719 ( .A1(n6178), .A2(n6091), .ZN(n5603) );
  AOI22_X1 U6720 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6126), .B1(n5594), 
        .B2(n6081), .ZN(n5595) );
  OAI211_X1 U6721 ( .C1(REIP_REG_16__SCAN_IN), .C2(n5596), .A(n5595), .B(n6128), .ZN(n5601) );
  NAND2_X1 U6722 ( .A1(n5608), .A2(n5597), .ZN(n5598) );
  NAND2_X1 U6723 ( .A1(n5897), .A2(n5598), .ZN(n5980) );
  NAND2_X1 U6724 ( .A1(n6125), .A2(EBX_REG_16__SCAN_IN), .ZN(n5599) );
  OAI21_X1 U6725 ( .B1(n5980), .B2(n6130), .A(n5599), .ZN(n5600) );
  NOR2_X1 U6726 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  OAI211_X1 U6727 ( .C1(n5604), .C2(n6601), .A(n5603), .B(n5602), .ZN(U2811)
         );
  INV_X1 U6728 ( .A(n5605), .ZN(n5606) );
  AOI21_X1 U6729 ( .B1(n5607), .B2(n5666), .A(n5606), .ZN(n5794) );
  INV_X1 U6730 ( .A(n5794), .ZN(n5695) );
  INV_X1 U6731 ( .A(n5608), .ZN(n5609) );
  AOI21_X1 U6732 ( .B1(n5610), .B2(n5671), .A(n5609), .ZN(n5990) );
  AOI22_X1 U6733 ( .A1(n6112), .A2(n5990), .B1(n5611), .B2(n6599), .ZN(n5612)
         );
  OAI211_X1 U6734 ( .C1(n6106), .C2(n6849), .A(n5612), .B(n6128), .ZN(n5614)
         );
  NOR2_X1 U6735 ( .A1(n6146), .A2(n5792), .ZN(n5613) );
  AOI211_X1 U6736 ( .C1(EBX_REG_15__SCAN_IN), .C2(n6125), .A(n5614), .B(n5613), 
        .ZN(n5617) );
  AND2_X1 U6737 ( .A1(n5923), .A2(n5615), .ZN(n6044) );
  NAND2_X1 U6738 ( .A1(n6044), .A2(REIP_REG_15__SCAN_IN), .ZN(n5616) );
  OAI211_X1 U6739 ( .C1(n5695), .C2(n6100), .A(n5617), .B(n5616), .ZN(U2812)
         );
  OAI22_X1 U6740 ( .A1(n5618), .A2(n6153), .B1(n6170), .B2(n6724), .ZN(U2828)
         );
  INV_X1 U6741 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5621) );
  OAI222_X1 U6742 ( .A1(n6148), .A2(n5619), .B1(n5621), .B2(n6170), .C1(n5620), 
        .C2(n6153), .ZN(U2830) );
  INV_X1 U6743 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6734) );
  OAI222_X1 U6744 ( .A1(n6148), .A2(n5680), .B1(n6734), .B2(n6170), .C1(n5803), 
        .C2(n6153), .ZN(U2831) );
  INV_X1 U6745 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5622) );
  INV_X1 U6746 ( .A(n5727), .ZN(n5685) );
  OAI222_X1 U6747 ( .A1(n5685), .A2(n6148), .B1(n5623), .B2(n6170), .C1(n6153), 
        .C2(n5823), .ZN(U2833) );
  AOI22_X1 U6748 ( .A1(n5832), .A2(n6165), .B1(EBX_REG_25__SCAN_IN), .B2(n5663), .ZN(n5624) );
  OAI21_X1 U6749 ( .B1(n5735), .B2(n6148), .A(n5624), .ZN(U2834) );
  INV_X1 U6750 ( .A(n5536), .ZN(n5628) );
  NAND2_X1 U6751 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  NAND2_X1 U6752 ( .A1(n5628), .A2(n5627), .ZN(n5915) );
  NOR2_X1 U6753 ( .A1(n6170), .A2(n5629), .ZN(n5630) );
  AOI21_X1 U6754 ( .B1(n5916), .B2(n6165), .A(n5630), .ZN(n5631) );
  OAI21_X1 U6755 ( .B1(n5915), .B2(n6148), .A(n5631), .ZN(U2835) );
  OAI22_X1 U6756 ( .A1(n5842), .A2(n6153), .B1(n5632), .B2(n6170), .ZN(n5633)
         );
  INV_X1 U6757 ( .A(n5633), .ZN(n5634) );
  OAI21_X1 U6758 ( .B1(n5690), .B2(n6148), .A(n5634), .ZN(U2836) );
  INV_X1 U6759 ( .A(n5635), .ZN(n5636) );
  AOI21_X1 U6760 ( .B1(n5638), .B2(n5637), .A(n5636), .ZN(n5955) );
  INV_X1 U6761 ( .A(n5955), .ZN(n5641) );
  INV_X1 U6762 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5640) );
  XNOR2_X1 U6763 ( .A(n5647), .B(n5639), .ZN(n5925) );
  OAI222_X1 U6764 ( .A1(n6148), .A2(n5641), .B1(n5640), .B2(n6170), .C1(n6153), 
        .C2(n5925), .ZN(U2837) );
  XNOR2_X1 U6765 ( .A(n5642), .B(n5643), .ZN(n5958) );
  INV_X1 U6766 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5648) );
  NOR2_X1 U6767 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  OR2_X1 U6768 ( .A1(n5647), .A2(n5646), .ZN(n5937) );
  OAI222_X1 U6769 ( .A1(n5958), .A2(n6148), .B1(n5648), .B2(n6170), .C1(n6153), 
        .C2(n5937), .ZN(U2838) );
  NOR2_X1 U6770 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  MUX2_X1 U6771 ( .A(n5653), .B(n5652), .S(n3135), .Z(n5655) );
  XNOR2_X1 U6772 ( .A(n5655), .B(n5654), .ZN(n5943) );
  AOI22_X1 U6773 ( .A1(n5943), .A2(n6165), .B1(EBX_REG_20__SCAN_IN), .B2(n5663), .ZN(n5656) );
  OAI21_X1 U6774 ( .B1(n5942), .B2(n6148), .A(n5656), .ZN(U2839) );
  INV_X1 U6775 ( .A(n5778), .ZN(n5693) );
  OAI22_X1 U6776 ( .A1(n5874), .A2(n6153), .B1(n5657), .B2(n6170), .ZN(n5658)
         );
  INV_X1 U6777 ( .A(n5658), .ZN(n5659) );
  OAI21_X1 U6778 ( .B1(n5693), .B2(n6148), .A(n5659), .ZN(U2840) );
  INV_X1 U6779 ( .A(n6171), .ZN(n5661) );
  INV_X1 U6780 ( .A(n5890), .ZN(n5660) );
  OAI222_X1 U6781 ( .A1(n6148), .A2(n5661), .B1(n6170), .B2(n6802), .C1(n6153), 
        .C2(n5660), .ZN(U2841) );
  INV_X1 U6782 ( .A(n6178), .ZN(n5662) );
  INV_X1 U6783 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6703) );
  OAI222_X1 U6784 ( .A1(n5662), .A2(n6148), .B1(n6170), .B2(n6703), .C1(n5980), 
        .C2(n6153), .ZN(U2843) );
  AOI22_X1 U6785 ( .A1(n5990), .A2(n6165), .B1(EBX_REG_15__SCAN_IN), .B2(n5663), .ZN(n5664) );
  OAI21_X1 U6786 ( .B1(n5695), .B2(n6148), .A(n5664), .ZN(U2844) );
  OR2_X1 U6787 ( .A1(n5589), .A2(n5665), .ZN(n5667) );
  INV_X1 U6788 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6940) );
  OR2_X1 U6789 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND2_X1 U6790 ( .A1(n5671), .A2(n5670), .ZN(n6040) );
  OAI222_X1 U6791 ( .A1(n5697), .A2(n6148), .B1(n6170), .B2(n6940), .C1(n6040), 
        .C2(n6153), .ZN(U2845) );
  NAND3_X1 U6792 ( .A1(n5673), .A2(n5672), .A3(n6186), .ZN(n5675) );
  AOI22_X1 U6793 ( .A1(n6177), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6179), .ZN(n5674) );
  NAND2_X1 U6794 ( .A1(n5675), .A2(n5674), .ZN(U2860) );
  AOI22_X1 U6795 ( .A1(n6177), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6179), .ZN(n5677) );
  NAND2_X1 U6796 ( .A1(n6180), .A2(DATAI_13_), .ZN(n5676) );
  OAI211_X1 U6797 ( .C1(n5619), .C2(n5951), .A(n5677), .B(n5676), .ZN(U2862)
         );
  AOI22_X1 U6798 ( .A1(n6177), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6179), .ZN(n5679) );
  NAND2_X1 U6799 ( .A1(n6180), .A2(DATAI_12_), .ZN(n5678) );
  OAI211_X1 U6800 ( .C1(n5680), .C2(n5951), .A(n5679), .B(n5678), .ZN(U2863)
         );
  AOI22_X1 U6801 ( .A1(n6177), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6179), .ZN(n5682) );
  NAND2_X1 U6802 ( .A1(n6180), .A2(DATAI_11_), .ZN(n5681) );
  OAI211_X1 U6803 ( .C1(n5713), .C2(n5951), .A(n5682), .B(n5681), .ZN(U2864)
         );
  AOI22_X1 U6804 ( .A1(n6177), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6179), .ZN(n5684) );
  NAND2_X1 U6805 ( .A1(n6180), .A2(DATAI_10_), .ZN(n5683) );
  OAI211_X1 U6806 ( .C1(n5685), .C2(n5951), .A(n5684), .B(n5683), .ZN(U2865)
         );
  AOI22_X1 U6807 ( .A1(n6177), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6179), .ZN(n5687) );
  NAND2_X1 U6808 ( .A1(n6180), .A2(DATAI_9_), .ZN(n5686) );
  OAI211_X1 U6809 ( .C1(n5735), .C2(n5951), .A(n5687), .B(n5686), .ZN(U2866)
         );
  AOI22_X1 U6810 ( .A1(n6177), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6179), .ZN(n5689) );
  NAND2_X1 U6811 ( .A1(n6180), .A2(DATAI_7_), .ZN(n5688) );
  OAI211_X1 U6812 ( .C1(n5690), .C2(n5951), .A(n5689), .B(n5688), .ZN(U2868)
         );
  AOI22_X1 U6813 ( .A1(n6177), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6179), .ZN(n5692) );
  NAND2_X1 U6814 ( .A1(n6180), .A2(DATAI_3_), .ZN(n5691) );
  OAI211_X1 U6815 ( .C1(n5693), .C2(n5951), .A(n5692), .B(n5691), .ZN(U2872)
         );
  AOI22_X1 U6816 ( .A1(n6183), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6179), .ZN(n5694) );
  OAI21_X1 U6817 ( .B1(n5695), .B2(n5951), .A(n5694), .ZN(U2876) );
  AOI22_X1 U6818 ( .A1(n6183), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6179), .ZN(n5696) );
  OAI21_X1 U6819 ( .B1(n5697), .B2(n5951), .A(n5696), .ZN(U2877) );
  INV_X1 U6820 ( .A(n5698), .ZN(n5722) );
  NAND3_X1 U6821 ( .A1(n5722), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5892), .ZN(n5702) );
  AND2_X1 U6822 ( .A1(n5718), .A2(n3632), .ZN(n5700) );
  NAND2_X1 U6823 ( .A1(n5699), .A2(n5700), .ZN(n5710) );
  AOI22_X1 U6824 ( .A1(n5702), .A2(n5710), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5701), .ZN(n5703) );
  XNOR2_X1 U6825 ( .A(n5703), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5813)
         );
  INV_X1 U6826 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6989) );
  NOR2_X1 U6827 ( .A1(n6001), .A2(n6989), .ZN(n5805) );
  AOI21_X1 U6828 ( .B1(n6322), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5805), 
        .ZN(n5704) );
  OAI21_X1 U6829 ( .B1(n5705), .B2(n6318), .A(n5704), .ZN(n5706) );
  AOI21_X1 U6830 ( .B1(n5707), .B2(n6314), .A(n5706), .ZN(n5708) );
  OAI21_X1 U6831 ( .B1(n6284), .B2(n5813), .A(n5708), .ZN(U2958) );
  INV_X1 U6832 ( .A(n5709), .ZN(n5711) );
  NAND2_X1 U6833 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  XNOR2_X1 U6834 ( .A(n5712), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5822)
         );
  NAND2_X1 U6835 ( .A1(n6375), .A2(REIP_REG_27__SCAN_IN), .ZN(n5814) );
  OAI21_X1 U6836 ( .B1(n6304), .B2(n6862), .A(n5814), .ZN(n5715) );
  NOR2_X1 U6837 ( .A1(n5713), .A2(n6325), .ZN(n5714) );
  INV_X1 U6838 ( .A(n5718), .ZN(n5720) );
  NAND2_X1 U6839 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  XNOR2_X1 U6840 ( .A(n5722), .B(n5721), .ZN(n5830) );
  NOR2_X1 U6841 ( .A1(n6001), .A2(n5723), .ZN(n5825) );
  AOI21_X1 U6842 ( .B1(n6322), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5825), 
        .ZN(n5724) );
  OAI21_X1 U6843 ( .B1(n5725), .B2(n6318), .A(n5724), .ZN(n5726) );
  AOI21_X1 U6844 ( .B1(n5727), .B2(n6314), .A(n5726), .ZN(n5728) );
  OAI21_X1 U6845 ( .B1(n5830), .B2(n6284), .A(n5728), .ZN(U2960) );
  NAND2_X1 U6846 ( .A1(n6375), .A2(REIP_REG_25__SCAN_IN), .ZN(n5833) );
  OAI21_X1 U6847 ( .B1(n6304), .B2(n5729), .A(n5833), .ZN(n5730) );
  AOI21_X1 U6848 ( .B1(n6298), .B2(n5731), .A(n5730), .ZN(n5734) );
  OAI21_X1 U6849 ( .B1(n5699), .B2(n5732), .A(n5372), .ZN(n5831) );
  NAND2_X1 U6850 ( .A1(n5831), .A2(n6320), .ZN(n5733) );
  OAI211_X1 U6851 ( .C1(n5735), .C2(n6325), .A(n5734), .B(n5733), .ZN(U2961)
         );
  INV_X1 U6852 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5737) );
  OAI21_X1 U6853 ( .B1(n6304), .B2(n5737), .A(n5736), .ZN(n5739) );
  NOR2_X1 U6854 ( .A1(n5915), .A2(n6325), .ZN(n5738) );
  AOI211_X1 U6855 ( .C1(n6298), .C2(n5913), .A(n5739), .B(n5738), .ZN(n5740)
         );
  OAI21_X1 U6856 ( .B1(n5741), .B2(n6284), .A(n5740), .ZN(U2962) );
  INV_X1 U6857 ( .A(n5843), .ZN(n5743) );
  NAND3_X1 U6858 ( .A1(n5892), .A2(n5743), .A3(n5742), .ZN(n5745) );
  OAI21_X1 U6859 ( .B1(n4163), .B2(n5745), .A(n5744), .ZN(n5746) );
  XNOR2_X1 U6860 ( .A(n5746), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5848)
         );
  NAND2_X1 U6861 ( .A1(n6298), .A2(n5747), .ZN(n5748) );
  NAND2_X1 U6862 ( .A1(n6375), .A2(REIP_REG_23__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U6863 ( .C1(n6304), .C2(n5749), .A(n5748), .B(n5841), .ZN(n5750)
         );
  AOI21_X1 U6864 ( .B1(n5751), .B2(n6314), .A(n5750), .ZN(n5752) );
  OAI21_X1 U6865 ( .B1(n5848), .B2(n6284), .A(n5752), .ZN(U2963) );
  AOI21_X1 U6866 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5892), .A(n5753), 
        .ZN(n5754) );
  XNOR2_X1 U6867 ( .A(n5755), .B(n5754), .ZN(n5854) );
  NAND2_X1 U6868 ( .A1(n6375), .A2(REIP_REG_22__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U6869 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5756)
         );
  OAI211_X1 U6870 ( .C1(n6318), .C2(n5921), .A(n5849), .B(n5756), .ZN(n5757)
         );
  AOI21_X1 U6871 ( .B1(n5955), .B2(n6314), .A(n5757), .ZN(n5758) );
  OAI21_X1 U6872 ( .B1(n5854), .B2(n6284), .A(n5758), .ZN(U2964) );
  OAI21_X1 U6873 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5855) );
  NAND2_X1 U6874 ( .A1(n5855), .A2(n6320), .ZN(n5764) );
  INV_X1 U6875 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U6876 ( .A1(n6375), .A2(REIP_REG_21__SCAN_IN), .ZN(n5856) );
  OAI21_X1 U6877 ( .B1(n6304), .B2(n5934), .A(n5856), .ZN(n5762) );
  AOI21_X1 U6878 ( .B1(n6298), .B2(n5936), .A(n5762), .ZN(n5763) );
  OAI211_X1 U6879 ( .C1(n6325), .C2(n5958), .A(n5764), .B(n5763), .ZN(U2965)
         );
  XOR2_X1 U6880 ( .A(n5766), .B(n5765), .Z(n5871) );
  NAND2_X1 U6881 ( .A1(n5871), .A2(n6320), .ZN(n5770) );
  AND2_X1 U6882 ( .A1(n6375), .A2(REIP_REG_20__SCAN_IN), .ZN(n5866) );
  INV_X1 U6883 ( .A(n5946), .ZN(n5767) );
  NOR2_X1 U6884 ( .A1(n6318), .A2(n5767), .ZN(n5768) );
  AOI211_X1 U6885 ( .C1(n6322), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5866), 
        .B(n5768), .ZN(n5769) );
  OAI211_X1 U6886 ( .C1(n6325), .C2(n5942), .A(n5770), .B(n5769), .ZN(U2966)
         );
  OAI21_X1 U6887 ( .B1(n5771), .B2(n3629), .A(n5772), .ZN(n5773) );
  XNOR2_X1 U6888 ( .A(n5773), .B(n5892), .ZN(n5880) );
  INV_X1 U6889 ( .A(n5774), .ZN(n5776) );
  NAND2_X1 U6890 ( .A1(n6375), .A2(REIP_REG_19__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U6891 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5775)
         );
  OAI211_X1 U6892 ( .C1(n6318), .C2(n5776), .A(n5873), .B(n5775), .ZN(n5777)
         );
  AOI21_X1 U6893 ( .B1(n5778), .B2(n6314), .A(n5777), .ZN(n5779) );
  OAI21_X1 U6894 ( .B1(n5880), .B2(n6284), .A(n5779), .ZN(U2967) );
  XNOR2_X1 U6895 ( .A(n5892), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5781)
         );
  XNOR2_X1 U6896 ( .A(n5780), .B(n5781), .ZN(n5981) );
  AOI22_X1 U6897 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6375), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5782) );
  OAI21_X1 U6898 ( .B1(n5783), .B2(n6318), .A(n5782), .ZN(n5784) );
  AOI21_X1 U6899 ( .B1(n6178), .B2(n6314), .A(n5784), .ZN(n5785) );
  OAI21_X1 U6900 ( .B1(n5981), .B2(n6284), .A(n5785), .ZN(U2970) );
  INV_X1 U6901 ( .A(n5786), .ZN(n5788) );
  NOR2_X1 U6902 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  XNOR2_X1 U6903 ( .A(n5790), .B(n5789), .ZN(n5991) );
  INV_X1 U6904 ( .A(n5991), .ZN(n5796) );
  AOI22_X1 U6905 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6375), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U6906 ( .B1(n5792), .B2(n6318), .A(n5791), .ZN(n5793) );
  AOI21_X1 U6907 ( .B1(n5794), .B2(n6314), .A(n5793), .ZN(n5795) );
  OAI21_X1 U6908 ( .B1(n6284), .B2(n5796), .A(n5795), .ZN(U2971) );
  XNOR2_X1 U6909 ( .A(n5892), .B(n6860), .ZN(n5798) );
  XNOR2_X1 U6910 ( .A(n5797), .B(n5798), .ZN(n5995) );
  INV_X1 U6911 ( .A(n6045), .ZN(n5800) );
  AOI22_X1 U6912 ( .A1(n6322), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6375), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5799) );
  OAI21_X1 U6913 ( .B1(n6318), .B2(n5800), .A(n5799), .ZN(n5801) );
  AOI21_X1 U6914 ( .B1(n6046), .B2(n6314), .A(n5801), .ZN(n5802) );
  OAI21_X1 U6915 ( .B1(n5995), .B2(n6284), .A(n5802), .ZN(U2972) );
  INV_X1 U6916 ( .A(n5816), .ZN(n5806) );
  NOR2_X1 U6917 ( .A1(n5803), .A2(n6352), .ZN(n5804) );
  AOI211_X1 U6918 ( .C1(n5806), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5805), .B(n5804), .ZN(n5812) );
  INV_X1 U6919 ( .A(n5807), .ZN(n5810) );
  INV_X1 U6920 ( .A(n5808), .ZN(n5809) );
  NAND3_X1 U6921 ( .A1(n5820), .A2(n5810), .A3(n5809), .ZN(n5811) );
  OAI211_X1 U6922 ( .C1(n5813), .C2(n6370), .A(n5812), .B(n5811), .ZN(U2990)
         );
  INV_X1 U6923 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5819) );
  OAI21_X1 U6924 ( .B1(n5815), .B2(n6352), .A(n5814), .ZN(n5818) );
  NOR2_X1 U6925 ( .A1(n5816), .A2(n5819), .ZN(n5817) );
  AOI211_X1 U6926 ( .C1(n5820), .C2(n5819), .A(n5818), .B(n5817), .ZN(n5821)
         );
  OAI21_X1 U6927 ( .B1(n5822), .B2(n6370), .A(n5821), .ZN(U2991) );
  NOR2_X1 U6928 ( .A1(n5823), .A2(n6352), .ZN(n5824) );
  AOI211_X1 U6929 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5836), .A(n5825), .B(n5824), .ZN(n5829) );
  INV_X1 U6930 ( .A(n5839), .ZN(n5827) );
  XNOR2_X1 U6931 ( .A(n3632), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5826)
         );
  NAND2_X1 U6932 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  OAI211_X1 U6933 ( .C1(n5830), .C2(n6370), .A(n5829), .B(n5828), .ZN(U2992)
         );
  NAND2_X1 U6934 ( .A1(n5831), .A2(n6382), .ZN(n5838) );
  INV_X1 U6935 ( .A(n5832), .ZN(n5834) );
  OAI21_X1 U6936 ( .B1(n5834), .B2(n6352), .A(n5833), .ZN(n5835) );
  AOI21_X1 U6937 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5836), .A(n5835), 
        .ZN(n5837) );
  OAI211_X1 U6938 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5839), .A(n5838), .B(n5837), .ZN(U2993) );
  INV_X1 U6939 ( .A(n5840), .ZN(n5846) );
  OAI21_X1 U6940 ( .B1(n5842), .B2(n6352), .A(n5841), .ZN(n5845) );
  NOR3_X1 U6941 ( .A1(n5861), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5843), 
        .ZN(n5844) );
  AOI211_X1 U6942 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5846), .A(n5845), .B(n5844), .ZN(n5847) );
  OAI21_X1 U6943 ( .B1(n5848), .B2(n6370), .A(n5847), .ZN(U2995) );
  OAI21_X1 U6944 ( .B1(n5925), .B2(n6352), .A(n5849), .ZN(n5852) );
  XNOR2_X1 U6945 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .B(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5850) );
  NOR2_X1 U6946 ( .A1(n5861), .A2(n5850), .ZN(n5851) );
  AOI211_X1 U6947 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5858), .A(n5852), .B(n5851), .ZN(n5853) );
  OAI21_X1 U6948 ( .B1(n5854), .B2(n6370), .A(n5853), .ZN(U2996) );
  NAND2_X1 U6949 ( .A1(n5855), .A2(n6382), .ZN(n5860) );
  OAI21_X1 U6950 ( .B1(n5937), .B2(n6352), .A(n5856), .ZN(n5857) );
  AOI21_X1 U6951 ( .B1(n5858), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5857), 
        .ZN(n5859) );
  OAI211_X1 U6952 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5861), .A(n5860), .B(n5859), .ZN(U2997) );
  OAI21_X1 U6953 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5862), .ZN(n5869) );
  NAND2_X1 U6954 ( .A1(n5864), .A2(n5863), .ZN(n6329) );
  AOI21_X1 U6955 ( .B1(n5902), .B2(n6329), .A(n5901), .ZN(n5886) );
  NAND2_X1 U6956 ( .A1(n6339), .A2(n5887), .ZN(n5865) );
  NAND2_X1 U6957 ( .A1(n5886), .A2(n5865), .ZN(n5878) );
  NAND2_X1 U6958 ( .A1(n5878), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5868) );
  AOI21_X1 U6959 ( .B1(n5943), .B2(n6377), .A(n5866), .ZN(n5867) );
  OAI211_X1 U6960 ( .C1(n5875), .C2(n5869), .A(n5868), .B(n5867), .ZN(n5870)
         );
  AOI21_X1 U6961 ( .B1(n5871), .B2(n6382), .A(n5870), .ZN(n5872) );
  INV_X1 U6962 ( .A(n5872), .ZN(U2998) );
  OAI21_X1 U6963 ( .B1(n5874), .B2(n6352), .A(n5873), .ZN(n5877) );
  NOR2_X1 U6964 ( .A1(n5875), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5876)
         );
  AOI211_X1 U6965 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5878), .A(n5877), .B(n5876), .ZN(n5879) );
  OAI21_X1 U6966 ( .B1(n5880), .B2(n6370), .A(n5879), .ZN(U2999) );
  NOR3_X1 U6967 ( .A1(n5780), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5883) );
  NOR2_X1 U6968 ( .A1(n5881), .A2(n5902), .ZN(n5882) );
  MUX2_X1 U6969 ( .A(n5883), .B(n5882), .S(n5892), .Z(n5884) );
  XNOR2_X1 U6970 ( .A(n5884), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5965)
         );
  NAND2_X1 U6971 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5903), .ZN(n5888) );
  NAND2_X1 U6972 ( .A1(n6333), .A2(REIP_REG_18__SCAN_IN), .ZN(n5885) );
  OAI221_X1 U6973 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5888), .C1(
        n5887), .C2(n5886), .A(n5885), .ZN(n5889) );
  AOI21_X1 U6974 ( .B1(n6377), .B2(n5890), .A(n5889), .ZN(n5891) );
  OAI21_X1 U6975 ( .B1(n5965), .B2(n6370), .A(n5891), .ZN(U3000) );
  NAND2_X1 U6976 ( .A1(n3617), .A2(n5987), .ZN(n5894) );
  NAND3_X1 U6977 ( .A1(n5780), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5892), .ZN(n5893) );
  OAI21_X1 U6978 ( .B1(n5780), .B2(n5894), .A(n5893), .ZN(n5895) );
  XNOR2_X1 U6979 ( .A(n5895), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5974)
         );
  AND2_X1 U6980 ( .A1(n5897), .A2(n5896), .ZN(n5899) );
  OR2_X1 U6981 ( .A1(n5899), .A2(n5898), .ZN(n6034) );
  OAI22_X1 U6982 ( .A1(n6034), .A2(n6352), .B1(n6001), .B2(n6604), .ZN(n5900)
         );
  AOI21_X1 U6983 ( .B1(n5901), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5900), 
        .ZN(n5905) );
  NAND2_X1 U6984 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  OAI211_X1 U6985 ( .C1(n5974), .C2(n6370), .A(n5905), .B(n5904), .ZN(U3001)
         );
  OAI21_X1 U6986 ( .B1(n5906), .B2(STATEBS16_REG_SCAN_IN), .A(n6447), .ZN(
        n5908) );
  OAI22_X1 U6987 ( .A1(n5908), .A2(n6446), .B1(n5907), .B2(n5910), .ZN(n5909)
         );
  MUX2_X1 U6988 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5909), .S(n6389), 
        .Z(U3464) );
  XNOR2_X1 U6989 ( .A(n3110), .B(n6446), .ZN(n5911) );
  OAI22_X1 U6990 ( .A1(n5911), .A2(n6452), .B1(n4466), .B2(n5910), .ZN(n5912)
         );
  MUX2_X1 U6991 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5912), .S(n6389), 
        .Z(U3463) );
  AND2_X1 U6992 ( .A1(n6680), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6993 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6125), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6126), .ZN(n5920) );
  AOI22_X1 U6994 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5914), .B1(n5913), .B2(
        n6081), .ZN(n5919) );
  INV_X1 U6995 ( .A(n5915), .ZN(n5952) );
  AOI22_X1 U6996 ( .A1(n5952), .A2(n6091), .B1(n5916), .B2(n6112), .ZN(n5918)
         );
  NAND4_X1 U6997 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(U2803)
         );
  AOI22_X1 U6998 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6125), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6126), .ZN(n5932) );
  INV_X1 U6999 ( .A(n5921), .ZN(n5924) );
  AND2_X1 U7000 ( .A1(n5923), .A2(n5922), .ZN(n5944) );
  AOI22_X1 U7001 ( .A1(n5924), .A2(n6081), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5944), .ZN(n5931) );
  INV_X1 U7002 ( .A(n5925), .ZN(n5926) );
  AOI22_X1 U7003 ( .A1(n5955), .A2(n6091), .B1(n6112), .B2(n5926), .ZN(n5930)
         );
  INV_X1 U7004 ( .A(n5941), .ZN(n5928) );
  OAI211_X1 U7005 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5928), .B(n5927), .ZN(n5929) );
  NAND4_X1 U7006 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(U2805)
         );
  AOI22_X1 U7007 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6125), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5944), .ZN(n5933) );
  OAI21_X1 U7008 ( .B1(n5934), .B2(n6106), .A(n5933), .ZN(n5935) );
  AOI21_X1 U7009 ( .B1(n5936), .B2(n6081), .A(n5935), .ZN(n5940) );
  OAI22_X1 U7010 ( .A1(n5958), .A2(n6100), .B1(n6130), .B2(n5937), .ZN(n5938)
         );
  INV_X1 U7011 ( .A(n5938), .ZN(n5939) );
  OAI211_X1 U7012 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5941), .A(n5940), .B(n5939), .ZN(U2806) );
  AOI22_X1 U7013 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6125), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6126), .ZN(n5950) );
  INV_X1 U7014 ( .A(n5942), .ZN(n5962) );
  AOI22_X1 U7015 ( .A1(n5962), .A2(n6091), .B1(n6112), .B2(n5943), .ZN(n5949)
         );
  OAI21_X1 U7016 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5945), .A(n5944), .ZN(n5948) );
  NAND2_X1 U7017 ( .A1(n5946), .A2(n6081), .ZN(n5947) );
  NAND4_X1 U7018 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(U2807)
         );
  AOI22_X1 U7019 ( .A1(n5952), .A2(n6184), .B1(n6177), .B2(DATAI_24_), .ZN(
        n5954) );
  AOI22_X1 U7020 ( .A1(n6180), .A2(DATAI_8_), .B1(n6179), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7021 ( .A1(n5954), .A2(n5953), .ZN(U2867) );
  AOI22_X1 U7022 ( .A1(n5955), .A2(n6184), .B1(n6177), .B2(DATAI_22_), .ZN(
        n5957) );
  AOI22_X1 U7023 ( .A1(n6180), .A2(DATAI_6_), .B1(n6179), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7024 ( .A1(n5957), .A2(n5956), .ZN(U2869) );
  INV_X1 U7025 ( .A(n5958), .ZN(n5959) );
  AOI22_X1 U7026 ( .A1(n5959), .A2(n6184), .B1(n6177), .B2(DATAI_21_), .ZN(
        n5961) );
  AOI22_X1 U7027 ( .A1(n6180), .A2(DATAI_5_), .B1(n6179), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7028 ( .A1(n5961), .A2(n5960), .ZN(U2870) );
  AOI22_X1 U7029 ( .A1(n5962), .A2(n6184), .B1(n6177), .B2(DATAI_20_), .ZN(
        n5964) );
  AOI22_X1 U7030 ( .A1(n6180), .A2(DATAI_4_), .B1(n6179), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7031 ( .A1(n5964), .A2(n5963), .ZN(U2871) );
  AOI22_X1 U7032 ( .A1(n6333), .A2(REIP_REG_18__SCAN_IN), .B1(n6322), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5968) );
  INV_X1 U7033 ( .A(n5965), .ZN(n5966) );
  AOI22_X1 U7034 ( .A1(n5966), .A2(n6320), .B1(n6314), .B2(n6171), .ZN(n5967)
         );
  OAI211_X1 U7035 ( .C1(n6318), .C2(n5969), .A(n5968), .B(n5967), .ZN(U2968)
         );
  AOI22_X1 U7036 ( .A1(n6333), .A2(REIP_REG_17__SCAN_IN), .B1(n6322), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5973) );
  XOR2_X1 U7037 ( .A(n5971), .B(n5970), .Z(n6174) );
  AOI22_X1 U7038 ( .A1(n6174), .A2(n6314), .B1(n6298), .B2(n6033), .ZN(n5972)
         );
  OAI211_X1 U7039 ( .C1(n5974), .C2(n6284), .A(n5973), .B(n5972), .ZN(U2969)
         );
  OAI22_X1 U7040 ( .A1(n6154), .A2(n6325), .B1(n6060), .B2(n6318), .ZN(n5975)
         );
  AOI21_X1 U7041 ( .B1(n6320), .B2(n5976), .A(n5975), .ZN(n5978) );
  OAI211_X1 U7042 ( .C1(n3825), .C2(n6304), .A(n5978), .B(n5977), .ZN(U2973)
         );
  AOI21_X1 U7043 ( .B1(n6339), .B2(n5979), .A(n6328), .ZN(n5988) );
  AOI21_X1 U7044 ( .B1(n6818), .B2(n5987), .A(n5994), .ZN(n5985) );
  NOR2_X1 U7045 ( .A1(n6001), .A2(n6601), .ZN(n5983) );
  OAI22_X1 U7046 ( .A1(n5981), .A2(n6370), .B1(n6352), .B2(n5980), .ZN(n5982)
         );
  AOI211_X1 U7047 ( .C1(n5985), .C2(n5984), .A(n5983), .B(n5982), .ZN(n5986)
         );
  OAI21_X1 U7048 ( .B1(n5988), .B2(n5987), .A(n5986), .ZN(U3002) );
  INV_X1 U7049 ( .A(n5988), .ZN(n5989) );
  AOI22_X1 U7050 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5989), .B1(n6333), .B2(REIP_REG_15__SCAN_IN), .ZN(n5993) );
  AOI22_X1 U7051 ( .A1(n5991), .A2(n6382), .B1(n6377), .B2(n5990), .ZN(n5992)
         );
  OAI211_X1 U7052 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5994), .A(n5993), .B(n5992), .ZN(U3003) );
  OAI22_X1 U7053 ( .A1(n5995), .A2(n6370), .B1(n6352), .B2(n6040), .ZN(n5996)
         );
  AOI21_X1 U7054 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5997), .A(n5996), 
        .ZN(n6000) );
  NAND3_X1 U7055 ( .A1(n5998), .A2(n6860), .A3(n6327), .ZN(n5999) );
  OAI211_X1 U7056 ( .C1(n6597), .C2(n6001), .A(n6000), .B(n5999), .ZN(U3004)
         );
  INV_X1 U7057 ( .A(n6002), .ZN(n6006) );
  INV_X1 U7058 ( .A(n6003), .ZN(n6005) );
  NAND4_X1 U7059 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6138), .ZN(n6007)
         );
  OAI21_X1 U7060 ( .B1(n6649), .B2(n6796), .A(n6007), .ZN(U3455) );
  AOI21_X1 U7061 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6564), .A(n6573), .ZN(n6012) );
  INV_X1 U7062 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6008) );
  INV_X1 U7063 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6569) );
  NOR2_X2 U7064 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6569), .ZN(n6679) );
  AOI21_X1 U7065 ( .B1(n6012), .B2(n6008), .A(n6679), .ZN(U2789) );
  OAI21_X1 U7066 ( .B1(n6009), .B2(n6554), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6010) );
  OAI21_X1 U7067 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6555), .A(n6010), .ZN(
        U2790) );
  INV_X2 U7068 ( .A(n6679), .ZN(n6662) );
  NOR2_X1 U7069 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6013) );
  OAI21_X1 U7070 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6013), .A(n6662), .ZN(n6011)
         );
  OAI21_X1 U7071 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6662), .A(n6011), .ZN(
        U2791) );
  OAI21_X1 U7072 ( .B1(n6013), .B2(BS16_N), .A(n6635), .ZN(n6633) );
  OAI21_X1 U7073 ( .B1(n6635), .B2(n6941), .A(n6633), .ZN(U2792) );
  INV_X1 U7074 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7075 ( .B1(n6015), .B2(n6014), .A(n6284), .ZN(U2793) );
  NOR4_X1 U7076 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6019) );
  NOR4_X1 U7077 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6018) );
  NOR4_X1 U7078 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6017) );
  NOR4_X1 U7079 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6016) );
  NAND4_X1 U7080 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n6025)
         );
  NOR4_X1 U7081 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6023) );
  AOI211_X1 U7082 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_17__SCAN_IN), .B(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6022) );
  NOR4_X1 U7083 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n6021) );
  NOR4_X1 U7084 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n6020) );
  NAND4_X1 U7085 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n6024)
         );
  NOR2_X1 U7086 ( .A1(n6025), .A2(n6024), .ZN(n6656) );
  INV_X1 U7087 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6027) );
  NOR3_X1 U7088 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7089 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6028), .A(n6656), .ZN(n6026)
         );
  OAI21_X1 U7090 ( .B1(n6656), .B2(n6027), .A(n6026), .ZN(U2794) );
  INV_X1 U7091 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6634) );
  AOI21_X1 U7092 ( .B1(n5186), .B2(n6634), .A(n6028), .ZN(n6030) );
  INV_X1 U7093 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6029) );
  INV_X1 U7094 ( .A(n6656), .ZN(n6659) );
  AOI22_X1 U7095 ( .A1(n6656), .A2(n6030), .B1(n6029), .B2(n6659), .ZN(U2795)
         );
  INV_X1 U7096 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6151) );
  OAI22_X1 U7097 ( .A1(n6123), .A2(n6151), .B1(n6031), .B2(n6106), .ZN(n6032)
         );
  AOI211_X1 U7098 ( .C1(n6081), .C2(n6033), .A(n6113), .B(n6032), .ZN(n6039)
         );
  INV_X1 U7099 ( .A(n6034), .ZN(n6149) );
  AOI22_X1 U7100 ( .A1(n6174), .A2(n6091), .B1(n6112), .B2(n6149), .ZN(n6038)
         );
  OAI21_X1 U7101 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6036), .A(n6035), .ZN(n6037) );
  NAND3_X1 U7102 ( .A1(n6039), .A2(n6038), .A3(n6037), .ZN(U2810) );
  INV_X1 U7103 ( .A(n6040), .ZN(n6041) );
  AOI22_X1 U7104 ( .A1(n6125), .A2(EBX_REG_14__SCAN_IN), .B1(n6112), .B2(n6041), .ZN(n6049) );
  OAI21_X1 U7105 ( .B1(n6137), .B2(n6042), .A(n6597), .ZN(n6043) );
  AOI22_X1 U7106 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6126), .B1(n6044), 
        .B2(n6043), .ZN(n6048) );
  AOI22_X1 U7107 ( .A1(n6046), .A2(n6091), .B1(n6081), .B2(n6045), .ZN(n6047)
         );
  NAND4_X1 U7108 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6128), .ZN(U2813)
         );
  NOR2_X1 U7109 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6050), .ZN(n6053) );
  NAND2_X1 U7110 ( .A1(n6126), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6051)
         );
  OAI211_X1 U7111 ( .C1(n6130), .C2(n6152), .A(n6128), .B(n6051), .ZN(n6052)
         );
  AOI21_X1 U7112 ( .B1(n6118), .B2(n6053), .A(n6052), .ZN(n6055) );
  NAND2_X1 U7113 ( .A1(n6125), .A2(EBX_REG_13__SCAN_IN), .ZN(n6054) );
  OAI211_X1 U7114 ( .C1(n6154), .C2(n6100), .A(n6055), .B(n6054), .ZN(n6056)
         );
  INV_X1 U7115 ( .A(n6056), .ZN(n6059) );
  OAI21_X1 U7116 ( .B1(n6063), .B2(n6057), .A(REIP_REG_13__SCAN_IN), .ZN(n6058) );
  OAI211_X1 U7117 ( .C1(n6146), .C2(n6060), .A(n6059), .B(n6058), .ZN(U2814)
         );
  OAI21_X1 U7118 ( .B1(n6137), .B2(n6061), .A(n6718), .ZN(n6062) );
  AOI22_X1 U7119 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6125), .B1(n6063), .B2(n6062), .ZN(n6070) );
  AOI22_X1 U7120 ( .A1(n6112), .A2(n6158), .B1(PHYADDRPOINTER_REG_11__SCAN_IN), 
        .B2(n6126), .ZN(n6069) );
  INV_X1 U7121 ( .A(n6064), .ZN(n6067) );
  INV_X1 U7122 ( .A(n5086), .ZN(n6066) );
  AOI21_X1 U7123 ( .B1(n6067), .B2(n6066), .A(n6065), .ZN(n6281) );
  AOI22_X1 U7124 ( .A1(n6281), .A2(n6091), .B1(n6081), .B2(n6280), .ZN(n6068)
         );
  NAND4_X1 U7125 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6128), .ZN(U2816)
         );
  OR2_X1 U7126 ( .A1(n6072), .A2(n6071), .ZN(n6073) );
  NAND2_X1 U7127 ( .A1(n5092), .A2(n6073), .ZN(n6351) );
  INV_X1 U7128 ( .A(n6351), .ZN(n6160) );
  AOI22_X1 U7129 ( .A1(n6074), .A2(REIP_REG_9__SCAN_IN), .B1(n6112), .B2(n6160), .ZN(n6084) );
  INV_X1 U7130 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6990) );
  OAI22_X1 U7131 ( .A1(n6123), .A2(n6990), .B1(n6075), .B2(n6106), .ZN(n6076)
         );
  AOI211_X1 U7132 ( .C1(n6078), .C2(n6077), .A(n6113), .B(n6076), .ZN(n6083)
         );
  INV_X1 U7133 ( .A(n6079), .ZN(n6161) );
  AOI22_X1 U7134 ( .A1(n6161), .A2(n6091), .B1(n6081), .B2(n6080), .ZN(n6082)
         );
  NAND3_X1 U7135 ( .A1(n6084), .A2(n6083), .A3(n6082), .ZN(U2818) );
  INV_X1 U7136 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6293) );
  OAI21_X1 U7137 ( .B1(n6106), .B2(n6293), .A(n6128), .ZN(n6085) );
  AOI21_X1 U7138 ( .B1(n6112), .B2(n6086), .A(n6085), .ZN(n6089) );
  INV_X1 U7139 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6831) );
  NAND3_X1 U7140 ( .A1(n6118), .A2(n6831), .A3(n6087), .ZN(n6088) );
  OAI211_X1 U7141 ( .C1(n6123), .C2(n6774), .A(n6089), .B(n6088), .ZN(n6090)
         );
  AOI21_X1 U7142 ( .B1(n6091), .B2(n6289), .A(n6090), .ZN(n6096) );
  INV_X1 U7143 ( .A(n6094), .ZN(n6093) );
  OAI21_X1 U7144 ( .B1(n6137), .B2(n6093), .A(n6092), .ZN(n6119) );
  NOR3_X1 U7145 ( .A1(n6137), .A2(REIP_REG_6__SCAN_IN), .A3(n6094), .ZN(n6097)
         );
  OAI21_X1 U7146 ( .B1(n6119), .B2(n6097), .A(REIP_REG_7__SCAN_IN), .ZN(n6095)
         );
  OAI211_X1 U7147 ( .C1(n6146), .C2(n6287), .A(n6096), .B(n6095), .ZN(U2820)
         );
  AOI211_X1 U7148 ( .C1(n6112), .C2(n6098), .A(n6113), .B(n6097), .ZN(n6105)
         );
  NOR2_X1 U7149 ( .A1(n6123), .A2(n6731), .ZN(n6103) );
  OAI22_X1 U7150 ( .A1(n6101), .A2(n6100), .B1(n6099), .B2(n6146), .ZN(n6102)
         );
  AOI211_X1 U7151 ( .C1(n6119), .C2(REIP_REG_6__SCAN_IN), .A(n6103), .B(n6102), 
        .ZN(n6104) );
  OAI211_X1 U7152 ( .C1(n6107), .C2(n6106), .A(n6105), .B(n6104), .ZN(U2821)
         );
  INV_X1 U7153 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6691) );
  OR2_X1 U7154 ( .A1(n6109), .A2(n6108), .ZN(n6111) );
  AND2_X1 U7155 ( .A1(n6111), .A2(n6110), .ZN(n6367) );
  NAND2_X1 U7156 ( .A1(n6112), .A2(n6367), .ZN(n6115) );
  AOI21_X1 U7157 ( .B1(n6126), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6113), 
        .ZN(n6114) );
  OAI211_X1 U7158 ( .C1(n6146), .C2(n6297), .A(n6115), .B(n6114), .ZN(n6116)
         );
  AOI21_X1 U7159 ( .B1(n6300), .B2(n6133), .A(n6116), .ZN(n6122) );
  AND2_X1 U7160 ( .A1(n6118), .A2(n6117), .ZN(n6120) );
  OAI21_X1 U7161 ( .B1(n6120), .B2(REIP_REG_5__SCAN_IN), .A(n6119), .ZN(n6121)
         );
  OAI211_X1 U7162 ( .C1(n6123), .C2(n6691), .A(n6122), .B(n6121), .ZN(U2822)
         );
  AOI22_X1 U7163 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6125), .B1(
        REIP_REG_4__SCAN_IN), .B2(n6124), .ZN(n6145) );
  NAND2_X1 U7164 ( .A1(n6126), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6127)
         );
  OAI211_X1 U7165 ( .C1(n6130), .C2(n6129), .A(n6128), .B(n6127), .ZN(n6131)
         );
  INV_X1 U7166 ( .A(n6131), .ZN(n6143) );
  NAND2_X1 U7167 ( .A1(n6133), .A2(n6132), .ZN(n6142) );
  INV_X1 U7168 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7169 ( .A1(n6583), .A2(n6135), .ZN(n6136) );
  OR2_X1 U7170 ( .A1(n6137), .A2(n6136), .ZN(n6141) );
  NAND2_X1 U7171 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  OAI211_X1 U7172 ( .C1(n6147), .C2(n6146), .A(n6145), .B(n6144), .ZN(U2823)
         );
  AOI22_X1 U7173 ( .A1(n6174), .A2(n6166), .B1(n6165), .B2(n6149), .ZN(n6150)
         );
  OAI21_X1 U7174 ( .B1(n6170), .B2(n6151), .A(n6150), .ZN(U2842) );
  INV_X1 U7175 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6157) );
  OAI22_X1 U7176 ( .A1(n6154), .A2(n6148), .B1(n6153), .B2(n6152), .ZN(n6155)
         );
  INV_X1 U7177 ( .A(n6155), .ZN(n6156) );
  OAI21_X1 U7178 ( .B1(n6170), .B2(n6157), .A(n6156), .ZN(U2846) );
  INV_X1 U7179 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7180 ( .A1(n6281), .A2(n6166), .B1(n6165), .B2(n6158), .ZN(n6159)
         );
  OAI21_X1 U7181 ( .B1(n6170), .B2(n6721), .A(n6159), .ZN(U2848) );
  AOI22_X1 U7182 ( .A1(n6161), .A2(n6166), .B1(n6165), .B2(n6160), .ZN(n6162)
         );
  OAI21_X1 U7183 ( .B1(n6170), .B2(n6990), .A(n6162), .ZN(U2850) );
  AOI22_X1 U7184 ( .A1(n6300), .A2(n6166), .B1(n6165), .B2(n6367), .ZN(n6163)
         );
  OAI21_X1 U7185 ( .B1(n6170), .B2(n6691), .A(n6163), .ZN(U2854) );
  INV_X1 U7186 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6169) );
  AOI22_X1 U7187 ( .A1(n6167), .A2(n6166), .B1(n6165), .B2(n6164), .ZN(n6168)
         );
  OAI21_X1 U7188 ( .B1(n6170), .B2(n6169), .A(n6168), .ZN(U2856) );
  AOI22_X1 U7189 ( .A1(n6171), .A2(n6184), .B1(n6177), .B2(DATAI_18_), .ZN(
        n6173) );
  AOI22_X1 U7190 ( .A1(n6180), .A2(DATAI_2_), .B1(n6179), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7191 ( .A1(n6173), .A2(n6172), .ZN(U2873) );
  AOI22_X1 U7192 ( .A1(n6174), .A2(n6184), .B1(n6177), .B2(DATAI_17_), .ZN(
        n6176) );
  AOI22_X1 U7193 ( .A1(n6180), .A2(DATAI_1_), .B1(n6179), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7194 ( .A1(n6176), .A2(n6175), .ZN(U2874) );
  AOI22_X1 U7195 ( .A1(n6178), .A2(n6184), .B1(n6177), .B2(DATAI_16_), .ZN(
        n6182) );
  AOI22_X1 U7196 ( .A1(n6180), .A2(DATAI_0_), .B1(n6179), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7197 ( .A1(n6182), .A2(n6181), .ZN(U2875) );
  INV_X1 U7198 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U7199 ( .A1(n6281), .A2(n6184), .B1(DATAI_11_), .B2(n6183), .ZN(
        n6185) );
  OAI21_X1 U7200 ( .B1(n6765), .B2(n6186), .A(n6185), .ZN(U2880) );
  INV_X1 U7201 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6279) );
  AOI22_X1 U7202 ( .A1(n6681), .A2(LWORD_REG_15__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6187) );
  OAI21_X1 U7203 ( .B1(n6279), .B2(n6203), .A(n6187), .ZN(U2908) );
  INV_X1 U7204 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6749) );
  AOI22_X1 U7205 ( .A1(n6681), .A2(LWORD_REG_14__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6188) );
  OAI21_X1 U7206 ( .B1(n6749), .B2(n6203), .A(n6188), .ZN(U2909) );
  INV_X1 U7207 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6273) );
  AOI22_X1 U7208 ( .A1(n6681), .A2(LWORD_REG_12__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6189) );
  OAI21_X1 U7209 ( .B1(n6273), .B2(n6203), .A(n6189), .ZN(U2911) );
  AOI22_X1 U7210 ( .A1(n6681), .A2(LWORD_REG_11__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6190) );
  OAI21_X1 U7211 ( .B1(n6765), .B2(n6203), .A(n6190), .ZN(U2912) );
  INV_X1 U7212 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6972) );
  AOI22_X1 U7213 ( .A1(n6681), .A2(LWORD_REG_10__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6191) );
  OAI21_X1 U7214 ( .B1(n6972), .B2(n6203), .A(n6191), .ZN(U2913) );
  INV_X1 U7215 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7216 ( .A1(n6681), .A2(LWORD_REG_9__SCAN_IN), .B1(n6192), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6193) );
  OAI21_X1 U7217 ( .B1(n6265), .B2(n6203), .A(n6193), .ZN(U2914) );
  INV_X1 U7218 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U7219 ( .A1(n6681), .A2(LWORD_REG_8__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6194) );
  OAI21_X1 U7220 ( .B1(n6866), .B2(n6203), .A(n6194), .ZN(U2915) );
  AOI22_X1 U7221 ( .A1(n6681), .A2(LWORD_REG_7__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6195) );
  OAI21_X1 U7222 ( .B1(n5000), .B2(n6203), .A(n6195), .ZN(U2916) );
  AOI22_X1 U7223 ( .A1(n6681), .A2(LWORD_REG_6__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6196) );
  OAI21_X1 U7224 ( .B1(n4814), .B2(n6203), .A(n6196), .ZN(U2917) );
  AOI22_X1 U7225 ( .A1(n6681), .A2(LWORD_REG_5__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6197) );
  OAI21_X1 U7226 ( .B1(n4812), .B2(n6203), .A(n6197), .ZN(U2918) );
  AOI22_X1 U7227 ( .A1(n6681), .A2(LWORD_REG_4__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6198) );
  OAI21_X1 U7228 ( .B1(n6253), .B2(n6203), .A(n6198), .ZN(U2919) );
  INV_X1 U7229 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6250) );
  AOI22_X1 U7230 ( .A1(n6681), .A2(LWORD_REG_3__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6199) );
  OAI21_X1 U7231 ( .B1(n6250), .B2(n6203), .A(n6199), .ZN(U2920) );
  AOI22_X1 U7232 ( .A1(n6681), .A2(LWORD_REG_2__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6200) );
  OAI21_X1 U7233 ( .B1(n6247), .B2(n6203), .A(n6200), .ZN(U2921) );
  AOI22_X1 U7234 ( .A1(n6681), .A2(LWORD_REG_1__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6201) );
  OAI21_X1 U7235 ( .B1(n6768), .B2(n6203), .A(n6201), .ZN(U2922) );
  AOI22_X1 U7236 ( .A1(n6681), .A2(LWORD_REG_0__SCAN_IN), .B1(n6680), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7237 ( .B1(n6723), .B2(n6203), .A(n6202), .ZN(U2923) );
  INV_X1 U7238 ( .A(n6239), .ZN(n6276) );
  AND2_X1 U7239 ( .A1(n6276), .A2(DATAI_0_), .ZN(n6241) );
  AOI21_X1 U7240 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6271), .A(n6241), .ZN(n6204) );
  OAI21_X1 U7241 ( .B1(n3871), .B2(n6278), .A(n6204), .ZN(U2924) );
  AND2_X1 U7242 ( .A1(n6276), .A2(DATAI_1_), .ZN(n6243) );
  AOI21_X1 U7243 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6271), .A(n6243), .ZN(n6205) );
  OAI21_X1 U7244 ( .B1(n6206), .B2(n6278), .A(n6205), .ZN(U2925) );
  AND2_X1 U7245 ( .A1(n6276), .A2(DATAI_2_), .ZN(n6245) );
  AOI21_X1 U7246 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6271), .A(n6245), .ZN(n6207) );
  OAI21_X1 U7247 ( .B1(n3927), .B2(n6278), .A(n6207), .ZN(U2926) );
  INV_X1 U7248 ( .A(DATAI_3_), .ZN(n6208) );
  NOR2_X1 U7249 ( .A1(n6239), .A2(n6208), .ZN(n6248) );
  AOI21_X1 U7250 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6271), .A(n6248), .ZN(n6209) );
  OAI21_X1 U7251 ( .B1(n6210), .B2(n6278), .A(n6209), .ZN(U2927) );
  AND2_X1 U7252 ( .A1(n6276), .A2(DATAI_4_), .ZN(n6251) );
  AOI21_X1 U7253 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6271), .A(n6251), .ZN(n6211) );
  OAI21_X1 U7254 ( .B1(n3964), .B2(n6278), .A(n6211), .ZN(U2928) );
  NOR2_X1 U7255 ( .A1(n6239), .A2(n6212), .ZN(n6254) );
  AOI21_X1 U7256 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6271), .A(n6254), .ZN(n6213) );
  OAI21_X1 U7257 ( .B1(n6214), .B2(n6278), .A(n6213), .ZN(U2929) );
  NOR2_X1 U7258 ( .A1(n6239), .A2(n6215), .ZN(n6256) );
  AOI21_X1 U7259 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6271), .A(n6256), .ZN(n6216) );
  OAI21_X1 U7260 ( .B1(n6821), .B2(n6278), .A(n6216), .ZN(U2930) );
  NOR2_X1 U7261 ( .A1(n6239), .A2(n6217), .ZN(n6258) );
  AOI21_X1 U7262 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6271), .A(n6258), .ZN(n6218) );
  OAI21_X1 U7263 ( .B1(n6219), .B2(n6278), .A(n6218), .ZN(U2931) );
  INV_X1 U7264 ( .A(DATAI_8_), .ZN(n6220) );
  NOR2_X1 U7265 ( .A1(n6239), .A2(n6220), .ZN(n6260) );
  AOI21_X1 U7266 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6271), .A(n6260), .ZN(n6221) );
  OAI21_X1 U7267 ( .B1(n6956), .B2(n6278), .A(n6221), .ZN(U2932) );
  INV_X1 U7268 ( .A(DATAI_9_), .ZN(n6223) );
  NOR2_X1 U7269 ( .A1(n6239), .A2(n6223), .ZN(n6262) );
  AOI21_X1 U7270 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6263), .A(n6262), .ZN(n6224) );
  OAI21_X1 U7271 ( .B1(n6225), .B2(n6278), .A(n6224), .ZN(U2933) );
  INV_X1 U7272 ( .A(DATAI_10_), .ZN(n6226) );
  NOR2_X1 U7273 ( .A1(n6239), .A2(n6226), .ZN(n6266) );
  AOI21_X1 U7274 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6263), .A(n6266), .ZN(
        n6227) );
  OAI21_X1 U7275 ( .B1(n6228), .B2(n6278), .A(n6227), .ZN(U2934) );
  INV_X1 U7276 ( .A(DATAI_11_), .ZN(n6229) );
  NOR2_X1 U7277 ( .A1(n6239), .A2(n6229), .ZN(n6268) );
  AOI21_X1 U7278 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6263), .A(n6268), .ZN(
        n6230) );
  OAI21_X1 U7279 ( .B1(n6231), .B2(n6278), .A(n6230), .ZN(U2935) );
  INV_X1 U7280 ( .A(DATAI_12_), .ZN(n6232) );
  NOR2_X1 U7281 ( .A1(n6239), .A2(n6232), .ZN(n6270) );
  AOI21_X1 U7282 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6263), .A(n6270), .ZN(
        n6233) );
  OAI21_X1 U7283 ( .B1(n6234), .B2(n6278), .A(n6233), .ZN(U2936) );
  AOI21_X1 U7284 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6263), .A(n6235), .ZN(
        n6236) );
  OAI21_X1 U7285 ( .B1(n6237), .B2(n6278), .A(n6236), .ZN(U2937) );
  INV_X1 U7286 ( .A(DATAI_14_), .ZN(n6238) );
  NOR2_X1 U7287 ( .A1(n6239), .A2(n6238), .ZN(n6274) );
  AOI21_X1 U7288 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6263), .A(n6274), .ZN(
        n6240) );
  OAI21_X1 U7289 ( .B1(n6958), .B2(n6278), .A(n6240), .ZN(U2938) );
  AOI21_X1 U7290 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6263), .A(n6241), .ZN(n6242) );
  OAI21_X1 U7291 ( .B1(n6723), .B2(n6278), .A(n6242), .ZN(U2939) );
  AOI21_X1 U7292 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6263), .A(n6243), .ZN(n6244) );
  OAI21_X1 U7293 ( .B1(n6768), .B2(n6278), .A(n6244), .ZN(U2940) );
  AOI21_X1 U7294 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6263), .A(n6245), .ZN(n6246) );
  OAI21_X1 U7295 ( .B1(n6247), .B2(n6278), .A(n6246), .ZN(U2941) );
  AOI21_X1 U7296 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6263), .A(n6248), .ZN(n6249) );
  OAI21_X1 U7297 ( .B1(n6250), .B2(n6278), .A(n6249), .ZN(U2942) );
  AOI21_X1 U7298 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6271), .A(n6251), .ZN(n6252) );
  OAI21_X1 U7299 ( .B1(n6253), .B2(n6278), .A(n6252), .ZN(U2943) );
  AOI21_X1 U7300 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6263), .A(n6254), .ZN(n6255) );
  OAI21_X1 U7301 ( .B1(n4812), .B2(n6278), .A(n6255), .ZN(U2944) );
  AOI21_X1 U7302 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6263), .A(n6256), .ZN(n6257) );
  OAI21_X1 U7303 ( .B1(n4814), .B2(n6278), .A(n6257), .ZN(U2945) );
  AOI21_X1 U7304 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6263), .A(n6258), .ZN(n6259) );
  OAI21_X1 U7305 ( .B1(n5000), .B2(n6278), .A(n6259), .ZN(U2946) );
  AOI21_X1 U7306 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6263), .A(n6260), .ZN(n6261) );
  OAI21_X1 U7307 ( .B1(n6866), .B2(n6278), .A(n6261), .ZN(U2947) );
  AOI21_X1 U7308 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6263), .A(n6262), .ZN(n6264) );
  OAI21_X1 U7309 ( .B1(n6265), .B2(n6278), .A(n6264), .ZN(U2948) );
  AOI21_X1 U7310 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6263), .A(n6266), .ZN(
        n6267) );
  OAI21_X1 U7311 ( .B1(n6972), .B2(n6278), .A(n6267), .ZN(U2949) );
  AOI21_X1 U7312 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6271), .A(n6268), .ZN(
        n6269) );
  OAI21_X1 U7313 ( .B1(n6765), .B2(n6278), .A(n6269), .ZN(U2950) );
  AOI21_X1 U7314 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6271), .A(n6270), .ZN(
        n6272) );
  OAI21_X1 U7315 ( .B1(n6273), .B2(n6278), .A(n6272), .ZN(U2951) );
  AOI21_X1 U7316 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6263), .A(n6274), .ZN(
        n6275) );
  OAI21_X1 U7317 ( .B1(n6749), .B2(n6278), .A(n6275), .ZN(U2953) );
  AOI22_X1 U7318 ( .A1(n6263), .A2(LWORD_REG_15__SCAN_IN), .B1(n6276), .B2(
        DATAI_15_), .ZN(n6277) );
  OAI21_X1 U7319 ( .B1(n6279), .B2(n6278), .A(n6277), .ZN(U2954) );
  AOI22_X1 U7320 ( .A1(n6333), .A2(REIP_REG_11__SCAN_IN), .B1(n6322), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6283) );
  AOI22_X1 U7321 ( .A1(n6281), .A2(n6314), .B1(n6298), .B2(n6280), .ZN(n6282)
         );
  OAI211_X1 U7322 ( .C1(n6285), .C2(n6284), .A(n6283), .B(n6282), .ZN(U2975)
         );
  INV_X1 U7323 ( .A(n6286), .ZN(n6290) );
  INV_X1 U7324 ( .A(n6287), .ZN(n6288) );
  AOI222_X1 U7325 ( .A1(n6290), .A2(n6320), .B1(n6289), .B2(n6314), .C1(n6288), 
        .C2(n6298), .ZN(n6292) );
  OAI211_X1 U7326 ( .C1(n6293), .C2(n6304), .A(n6292), .B(n6291), .ZN(U2979)
         );
  INV_X1 U7327 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U7328 ( .A(n6294), .B(n6296), .ZN(n6371) );
  INV_X1 U7329 ( .A(n6371), .ZN(n6301) );
  INV_X1 U7330 ( .A(n6297), .ZN(n6299) );
  AOI222_X1 U7331 ( .A1(n6301), .A2(n6320), .B1(n6300), .B2(n6314), .C1(n6299), 
        .C2(n6298), .ZN(n6303) );
  AND2_X1 U7332 ( .A1(n6333), .A2(REIP_REG_5__SCAN_IN), .ZN(n6366) );
  INV_X1 U7333 ( .A(n6366), .ZN(n6302) );
  OAI211_X1 U7334 ( .C1(n6738), .C2(n6304), .A(n6303), .B(n6302), .ZN(U2981)
         );
  AOI22_X1 U7335 ( .A1(n6333), .A2(REIP_REG_2__SCAN_IN), .B1(n6322), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6310) );
  XNOR2_X1 U7336 ( .A(n6305), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6307)
         );
  XNOR2_X1 U7337 ( .A(n6307), .B(n6306), .ZN(n6381) );
  AOI22_X1 U7338 ( .A1(n6381), .A2(n6320), .B1(n6308), .B2(n6314), .ZN(n6309)
         );
  OAI211_X1 U7339 ( .C1(n6318), .C2(n6311), .A(n6310), .B(n6309), .ZN(U2984)
         );
  AOI22_X1 U7340 ( .A1(n6333), .A2(REIP_REG_1__SCAN_IN), .B1(n6322), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6317) );
  INV_X1 U7341 ( .A(n6312), .ZN(n6315) );
  AOI22_X1 U7342 ( .A1(n6320), .A2(n6315), .B1(n6314), .B2(n6313), .ZN(n6316)
         );
  OAI211_X1 U7343 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6318), .A(n6317), 
        .B(n6316), .ZN(U2985) );
  AOI22_X1 U7344 ( .A1(n6320), .A2(n6319), .B1(n6375), .B2(REIP_REG_0__SCAN_IN), .ZN(n6324) );
  OAI21_X1 U7345 ( .B1(n6322), .B2(n6321), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6323) );
  OAI211_X1 U7346 ( .C1(n6326), .C2(n6325), .A(n6324), .B(n6323), .ZN(U2986)
         );
  AOI21_X1 U7347 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6327), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6337) );
  AOI21_X1 U7348 ( .B1(n6330), .B2(n6329), .A(n6328), .ZN(n6336) );
  AOI22_X1 U7349 ( .A1(n6332), .A2(n6382), .B1(n6377), .B2(n6331), .ZN(n6335)
         );
  NAND2_X1 U7350 ( .A1(n6333), .A2(REIP_REG_12__SCAN_IN), .ZN(n6334) );
  OAI211_X1 U7351 ( .C1(n6337), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3006)
         );
  AOI21_X1 U7352 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6361) );
  NAND2_X1 U7353 ( .A1(n6342), .A2(n6341), .ZN(n6357) );
  AOI221_X1 U7354 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6360), .C2(n6349), .A(n6357), 
        .ZN(n6343) );
  AOI21_X1 U7355 ( .B1(n6375), .B2(REIP_REG_10__SCAN_IN), .A(n6343), .ZN(n6344) );
  OAI21_X1 U7356 ( .B1(n6352), .B2(n6345), .A(n6344), .ZN(n6346) );
  AOI21_X1 U7357 ( .B1(n6347), .B2(n6382), .A(n6346), .ZN(n6348) );
  OAI21_X1 U7358 ( .B1(n6361), .B2(n6349), .A(n6348), .ZN(U3008) );
  OAI21_X1 U7359 ( .B1(n6352), .B2(n6351), .A(n6350), .ZN(n6353) );
  INV_X1 U7360 ( .A(n6353), .ZN(n6356) );
  NAND2_X1 U7361 ( .A1(n6354), .A2(n6382), .ZN(n6355) );
  OAI211_X1 U7362 ( .C1(n6357), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6356), 
        .B(n6355), .ZN(n6358) );
  INV_X1 U7363 ( .A(n6358), .ZN(n6359) );
  OAI21_X1 U7364 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(U3009) );
  NAND2_X1 U7365 ( .A1(n6362), .A2(n6384), .ZN(n6374) );
  AOI21_X1 U7366 ( .B1(n6378), .B2(n6363), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6364) );
  OR2_X1 U7367 ( .A1(n6365), .A2(n6364), .ZN(n6369) );
  AOI21_X1 U7368 ( .B1(n6377), .B2(n6367), .A(n6366), .ZN(n6368) );
  OAI211_X1 U7369 ( .C1(n6371), .C2(n6370), .A(n6369), .B(n6368), .ZN(n6372)
         );
  INV_X1 U7370 ( .A(n6372), .ZN(n6373) );
  OAI21_X1 U7371 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6374), .A(n6373), 
        .ZN(U3013) );
  AOI22_X1 U7372 ( .A1(n6377), .A2(n6376), .B1(n6375), .B2(REIP_REG_2__SCAN_IN), .ZN(n6388) );
  NAND3_X1 U7373 ( .A1(n6378), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U7374 ( .A1(n6380), .A2(n6379), .ZN(n6383) );
  AOI22_X1 U7375 ( .A1(n6383), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6382), 
        .B2(n6381), .ZN(n6387) );
  INV_X1 U7376 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6685) );
  NAND3_X1 U7377 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6384), .A3(n6685), 
        .ZN(n6385) );
  NAND4_X1 U7378 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(U3016)
         );
  NOR2_X1 U7379 ( .A1(n6530), .A2(n6389), .ZN(U3019) );
  AOI22_X1 U7380 ( .A1(n6393), .A2(n6392), .B1(n6391), .B2(n6390), .ZN(n6394)
         );
  INV_X1 U7381 ( .A(n6394), .ZN(n6423) );
  NOR2_X1 U7382 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6395), .ZN(n6422)
         );
  AOI22_X1 U7383 ( .A1(n6459), .A2(n6423), .B1(n6445), .B2(n6422), .ZN(n6406)
         );
  OAI21_X1 U7384 ( .B1(n6424), .B2(n6396), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6397) );
  NAND3_X1 U7385 ( .A1(n6398), .A2(n6447), .A3(n6397), .ZN(n6403) );
  INV_X1 U7386 ( .A(n6422), .ZN(n6401) );
  AOI211_X1 U7387 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6401), .A(n6400), .B(
        n6399), .ZN(n6402) );
  NAND3_X1 U7388 ( .A1(n6532), .A2(n6403), .A3(n6402), .ZN(n6425) );
  AOI22_X1 U7389 ( .A1(n6425), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6404), 
        .B2(n6424), .ZN(n6405) );
  OAI211_X1 U7390 ( .C1(n6407), .C2(n6441), .A(n6406), .B(n6405), .ZN(U3068)
         );
  AOI22_X1 U7391 ( .A1(n6465), .A2(n6423), .B1(n6464), .B2(n6422), .ZN(n6409)
         );
  AOI22_X1 U7392 ( .A1(n6425), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6463), 
        .B2(n6424), .ZN(n6408) );
  OAI211_X1 U7393 ( .C1(n6468), .C2(n6441), .A(n6409), .B(n6408), .ZN(U3069)
         );
  AOI22_X1 U7394 ( .A1(n6471), .A2(n6423), .B1(n6470), .B2(n6422), .ZN(n6411)
         );
  AOI22_X1 U7395 ( .A1(n6425), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6469), 
        .B2(n6424), .ZN(n6410) );
  OAI211_X1 U7396 ( .C1(n6474), .C2(n6441), .A(n6411), .B(n6410), .ZN(U3070)
         );
  AOI22_X1 U7397 ( .A1(n6476), .A2(n6422), .B1(n6477), .B2(n6423), .ZN(n6413)
         );
  AOI22_X1 U7398 ( .A1(n6425), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6475), 
        .B2(n6424), .ZN(n6412) );
  OAI211_X1 U7399 ( .C1(n6480), .C2(n6441), .A(n6413), .B(n6412), .ZN(U3071)
         );
  AOI22_X1 U7400 ( .A1(n6484), .A2(n6423), .B1(n6483), .B2(n6422), .ZN(n6416)
         );
  AOI22_X1 U7401 ( .A1(n6425), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6414), 
        .B2(n6424), .ZN(n6415) );
  OAI211_X1 U7402 ( .C1(n6417), .C2(n6441), .A(n6416), .B(n6415), .ZN(U3072)
         );
  AOI22_X1 U7403 ( .A1(n6490), .A2(n6422), .B1(n6491), .B2(n6423), .ZN(n6419)
         );
  AOI22_X1 U7404 ( .A1(n6425), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6489), 
        .B2(n6424), .ZN(n6418) );
  OAI211_X1 U7405 ( .C1(n6494), .C2(n6441), .A(n6419), .B(n6418), .ZN(U3073)
         );
  AOI22_X1 U7406 ( .A1(n6496), .A2(n6422), .B1(n6497), .B2(n6423), .ZN(n6421)
         );
  AOI22_X1 U7407 ( .A1(n6425), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6495), 
        .B2(n6424), .ZN(n6420) );
  OAI211_X1 U7408 ( .C1(n6500), .C2(n6441), .A(n6421), .B(n6420), .ZN(U3074)
         );
  AOI22_X1 U7409 ( .A1(n6506), .A2(n6423), .B1(n6504), .B2(n6422), .ZN(n6427)
         );
  AOI22_X1 U7410 ( .A1(n6425), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6502), 
        .B2(n6424), .ZN(n6426) );
  OAI211_X1 U7411 ( .C1(n6511), .C2(n6441), .A(n6427), .B(n6426), .ZN(U3075)
         );
  AOI22_X1 U7412 ( .A1(n6445), .A2(n6436), .B1(n6444), .B2(n6434), .ZN(n6429)
         );
  AOI22_X1 U7413 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6438), .B1(n6459), 
        .B2(n6437), .ZN(n6428) );
  OAI211_X1 U7414 ( .C1(n6462), .C2(n6441), .A(n6429), .B(n6428), .ZN(U3076)
         );
  AOI22_X1 U7415 ( .A1(n6464), .A2(n6436), .B1(n6430), .B2(n6434), .ZN(n6432)
         );
  AOI22_X1 U7416 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6438), .B1(n6465), 
        .B2(n6437), .ZN(n6431) );
  OAI211_X1 U7417 ( .C1(n6433), .C2(n6441), .A(n6432), .B(n6431), .ZN(U3077)
         );
  AOI22_X1 U7418 ( .A1(n6470), .A2(n6436), .B1(n6435), .B2(n6434), .ZN(n6440)
         );
  AOI22_X1 U7419 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6438), .B1(n6471), 
        .B2(n6437), .ZN(n6439) );
  OAI211_X1 U7420 ( .C1(n6442), .C2(n6441), .A(n6440), .B(n6439), .ZN(U3078)
         );
  NOR2_X1 U7421 ( .A1(n6443), .A2(n6532), .ZN(n6503) );
  AOI22_X1 U7422 ( .A1(n6445), .A2(n6503), .B1(n6444), .B2(n6481), .ZN(n6461)
         );
  INV_X1 U7423 ( .A(n6446), .ZN(n6448) );
  OAI21_X1 U7424 ( .B1(n6449), .B2(n6448), .A(n6447), .ZN(n6458) );
  AOI21_X1 U7425 ( .B1(n6450), .B2(n6516), .A(n6503), .ZN(n6457) );
  INV_X1 U7426 ( .A(n6457), .ZN(n6454) );
  AOI21_X1 U7427 ( .B1(n6452), .B2(n6456), .A(n6451), .ZN(n6453) );
  OAI21_X1 U7428 ( .B1(n6458), .B2(n6454), .A(n6453), .ZN(n6507) );
  OAI22_X1 U7429 ( .A1(n6458), .A2(n6457), .B1(n6456), .B2(n6455), .ZN(n6505)
         );
  AOI22_X1 U7430 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6507), .B1(n6459), 
        .B2(n6505), .ZN(n6460) );
  OAI211_X1 U7431 ( .C1(n6462), .C2(n6487), .A(n6461), .B(n6460), .ZN(U3108)
         );
  AOI22_X1 U7432 ( .A1(n6464), .A2(n6503), .B1(n6463), .B2(n6501), .ZN(n6467)
         );
  AOI22_X1 U7433 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6507), .B1(n6465), 
        .B2(n6505), .ZN(n6466) );
  OAI211_X1 U7434 ( .C1(n6468), .C2(n6510), .A(n6467), .B(n6466), .ZN(U3109)
         );
  AOI22_X1 U7435 ( .A1(n6470), .A2(n6503), .B1(n6469), .B2(n6501), .ZN(n6473)
         );
  AOI22_X1 U7436 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6507), .B1(n6471), 
        .B2(n6505), .ZN(n6472) );
  OAI211_X1 U7437 ( .C1(n6474), .C2(n6510), .A(n6473), .B(n6472), .ZN(U3110)
         );
  AOI22_X1 U7438 ( .A1(n6476), .A2(n6503), .B1(n6475), .B2(n6501), .ZN(n6479)
         );
  AOI22_X1 U7439 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6507), .B1(n6477), 
        .B2(n6505), .ZN(n6478) );
  OAI211_X1 U7440 ( .C1(n6480), .C2(n6510), .A(n6479), .B(n6478), .ZN(U3111)
         );
  AOI22_X1 U7441 ( .A1(n6483), .A2(n6503), .B1(n6482), .B2(n6481), .ZN(n6486)
         );
  AOI22_X1 U7442 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6507), .B1(n6484), 
        .B2(n6505), .ZN(n6485) );
  OAI211_X1 U7443 ( .C1(n6488), .C2(n6487), .A(n6486), .B(n6485), .ZN(U3112)
         );
  AOI22_X1 U7444 ( .A1(n6490), .A2(n6503), .B1(n6489), .B2(n6501), .ZN(n6493)
         );
  AOI22_X1 U7445 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6507), .B1(n6491), 
        .B2(n6505), .ZN(n6492) );
  OAI211_X1 U7446 ( .C1(n6494), .C2(n6510), .A(n6493), .B(n6492), .ZN(U3113)
         );
  AOI22_X1 U7447 ( .A1(n6496), .A2(n6503), .B1(n6495), .B2(n6501), .ZN(n6499)
         );
  AOI22_X1 U7448 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6507), .B1(n6497), 
        .B2(n6505), .ZN(n6498) );
  OAI211_X1 U7449 ( .C1(n6500), .C2(n6510), .A(n6499), .B(n6498), .ZN(U3114)
         );
  AOI22_X1 U7450 ( .A1(n6504), .A2(n6503), .B1(n6502), .B2(n6501), .ZN(n6509)
         );
  AOI22_X1 U7451 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6507), .B1(n6506), 
        .B2(n6505), .ZN(n6508) );
  OAI211_X1 U7452 ( .C1(n6511), .C2(n6510), .A(n6509), .B(n6508), .ZN(U3115)
         );
  INV_X1 U7453 ( .A(n6533), .ZN(n6529) );
  INV_X1 U7454 ( .A(n6512), .ZN(n6515) );
  AOI22_X1 U7455 ( .A1(n6516), .A2(n6515), .B1(n6514), .B2(n6513), .ZN(n6646)
         );
  NAND2_X1 U7456 ( .A1(n6517), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6652) );
  NAND3_X1 U7457 ( .A1(n6646), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6652), .ZN(n6520) );
  OAI211_X1 U7458 ( .C1(n6701), .C2(n6520), .A(n6519), .B(n6518), .ZN(n6522)
         );
  NAND2_X1 U7459 ( .A1(n6701), .A2(n6520), .ZN(n6521) );
  NAND2_X1 U7460 ( .A1(n6522), .A2(n6521), .ZN(n6527) );
  INV_X1 U7461 ( .A(n6527), .ZN(n6524) );
  OAI21_X1 U7462 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6524), .A(n6523), 
        .ZN(n6525) );
  OAI21_X1 U7463 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(n6528) );
  OAI21_X1 U7464 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6529), .A(n6528), 
        .ZN(n6531) );
  OAI211_X1 U7465 ( .C1(n6533), .C2(n6532), .A(n6531), .B(n6530), .ZN(n6541)
         );
  OR2_X1 U7466 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6536) );
  AOI211_X1 U7467 ( .C1(n6537), .C2(n6536), .A(n6535), .B(n6534), .ZN(n6538)
         );
  AND4_X1 U7468 ( .A1(n6541), .A2(n6540), .A3(n6539), .A4(n6538), .ZN(n6552)
         );
  NOR2_X1 U7469 ( .A1(n6671), .A2(n6542), .ZN(n6546) );
  AOI22_X1 U7470 ( .A1(n6552), .A2(n6543), .B1(READY_N), .B2(n6681), .ZN(n6544) );
  AOI21_X1 U7471 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6547) );
  INV_X1 U7472 ( .A(n6547), .ZN(n6638) );
  OAI21_X1 U7473 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6666), .A(n6638), .ZN(
        n6553) );
  AOI221_X1 U7474 ( .B1(n6549), .B2(STATE2_REG_0__SCAN_IN), .C1(n6553), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6548), .ZN(n6551) );
  OAI211_X1 U7475 ( .C1(n6560), .C2(n6640), .A(n6786), .B(n6638), .ZN(n6550)
         );
  OAI211_X1 U7476 ( .C1(n6552), .C2(n6554), .A(n6551), .B(n6550), .ZN(U3148)
         );
  OAI211_X1 U7477 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6553), .ZN(n6559) );
  OAI21_X1 U7478 ( .B1(READY_N), .B2(n6555), .A(n6554), .ZN(n6557) );
  AOI21_X1 U7479 ( .B1(n6557), .B2(n6638), .A(n6556), .ZN(n6558) );
  NAND2_X1 U7480 ( .A1(n6559), .A2(n6558), .ZN(U3149) );
  INV_X1 U7481 ( .A(n6560), .ZN(n6675) );
  INV_X1 U7482 ( .A(n6561), .ZN(n6636) );
  OAI221_X1 U7483 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6666), .A(n6636), .ZN(n6563) );
  OAI21_X1 U7484 ( .B1(n6675), .B2(n6563), .A(n6562), .ZN(U3150) );
  INV_X1 U7485 ( .A(n6635), .ZN(n6631) );
  AND2_X1 U7486 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6631), .ZN(U3151) );
  AND2_X1 U7487 ( .A1(n6631), .A2(DATAWIDTH_REG_30__SCAN_IN), .ZN(U3152) );
  AND2_X1 U7488 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6631), .ZN(U3153) );
  AND2_X1 U7489 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6631), .ZN(U3154) );
  AND2_X1 U7490 ( .A1(n6631), .A2(DATAWIDTH_REG_27__SCAN_IN), .ZN(U3155) );
  AND2_X1 U7491 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6631), .ZN(U3156) );
  AND2_X1 U7492 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6631), .ZN(U3157) );
  AND2_X1 U7493 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6631), .ZN(U3158) );
  AND2_X1 U7494 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6631), .ZN(U3159) );
  AND2_X1 U7495 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6631), .ZN(U3160) );
  AND2_X1 U7496 ( .A1(n6631), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7497 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6631), .ZN(U3162) );
  AND2_X1 U7498 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6631), .ZN(U3163) );
  AND2_X1 U7499 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6631), .ZN(U3164) );
  AND2_X1 U7500 ( .A1(n6631), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  AND2_X1 U7501 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6631), .ZN(U3166) );
  AND2_X1 U7502 ( .A1(n6631), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7503 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6631), .ZN(U3168) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6631), .ZN(U3169) );
  AND2_X1 U7505 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6631), .ZN(U3170) );
  AND2_X1 U7506 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6631), .ZN(U3171) );
  AND2_X1 U7507 ( .A1(n6631), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6631), .ZN(U3173) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6631), .ZN(U3174) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6631), .ZN(U3175) );
  AND2_X1 U7511 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6631), .ZN(U3176) );
  AND2_X1 U7512 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6631), .ZN(U3177) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6631), .ZN(U3178) );
  AND2_X1 U7514 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6631), .ZN(U3179) );
  AND2_X1 U7515 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6631), .ZN(U3180) );
  NOR2_X1 U7516 ( .A1(n6569), .A2(n6564), .ZN(n6570) );
  AOI22_X1 U7517 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6578) );
  AND2_X1 U7518 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6567) );
  INV_X1 U7519 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6677) );
  INV_X1 U7520 ( .A(NA_N), .ZN(n6571) );
  AOI221_X1 U7521 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6571), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6575) );
  AOI221_X1 U7522 ( .B1(n6567), .B2(n6662), .C1(n6677), .C2(n6662), .A(n6575), 
        .ZN(n6565) );
  OAI21_X1 U7523 ( .B1(n6570), .B2(n6578), .A(n6565), .ZN(U3181) );
  NOR2_X1 U7524 ( .A1(n6573), .A2(n6677), .ZN(n6572) );
  NAND2_X1 U7525 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6566) );
  OAI21_X1 U7526 ( .B1(n6572), .B2(n6567), .A(n6566), .ZN(n6568) );
  OAI211_X1 U7527 ( .C1(n6569), .C2(n6666), .A(n6671), .B(n6568), .ZN(U3182)
         );
  AOI21_X1 U7528 ( .B1(n6572), .B2(n6571), .A(n6570), .ZN(n6577) );
  AOI221_X1 U7529 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6666), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6574) );
  AOI221_X1 U7530 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6574), .C2(HOLD), .A(n6573), .ZN(n6576) );
  OAI22_X1 U7531 ( .A1(n6578), .A2(n6577), .B1(n6576), .B2(n6575), .ZN(U3183)
         );
  NOR2_X2 U7532 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6662), .ZN(n6607) );
  AOI22_X1 U7533 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6662), .ZN(n6579) );
  OAI21_X1 U7534 ( .B1(n5186), .B2(n6625), .A(n6579), .ZN(U3184) );
  AOI22_X1 U7535 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6662), .ZN(n6580) );
  OAI21_X1 U7536 ( .B1(n6739), .B2(n6625), .A(n6580), .ZN(U3185) );
  INV_X1 U7537 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7538 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6662), .ZN(n6581) );
  OAI21_X1 U7539 ( .B1(n6750), .B2(n6625), .A(n6581), .ZN(U3186) );
  INV_X1 U7540 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6829) );
  INV_X1 U7541 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6582) );
  INV_X1 U7542 ( .A(n6607), .ZN(n6628) );
  OAI222_X1 U7543 ( .A1(n6625), .A2(n6583), .B1(n6829), .B2(n6679), .C1(n6582), 
        .C2(n6628), .ZN(U3187) );
  INV_X1 U7544 ( .A(n6625), .ZN(n6626) );
  AOI222_X1 U7545 ( .A1(n6626), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6662), .C1(REIP_REG_6__SCAN_IN), .C2(
        n6607), .ZN(n6584) );
  INV_X1 U7546 ( .A(n6584), .ZN(U3188) );
  AOI22_X1 U7547 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6662), .ZN(n6585) );
  OAI21_X1 U7548 ( .B1(n6586), .B2(n6625), .A(n6585), .ZN(U3189) );
  AOI22_X1 U7549 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6662), .ZN(n6587) );
  OAI21_X1 U7550 ( .B1(n6831), .B2(n6625), .A(n6587), .ZN(U3190) );
  AOI22_X1 U7551 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6662), .ZN(n6588) );
  OAI21_X1 U7552 ( .B1(n6589), .B2(n6625), .A(n6588), .ZN(U3191) );
  AOI222_X1 U7553 ( .A1(n6626), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6662), .C1(REIP_REG_10__SCAN_IN), .C2(
        n6607), .ZN(n6590) );
  INV_X1 U7554 ( .A(n6590), .ZN(U3192) );
  AOI22_X1 U7555 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6662), .ZN(n6591) );
  OAI21_X1 U7556 ( .B1(n6592), .B2(n6625), .A(n6591), .ZN(U3193) );
  INV_X1 U7557 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6593) );
  INV_X1 U7558 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6595) );
  OAI222_X1 U7559 ( .A1(n6625), .A2(n6718), .B1(n6593), .B2(n6679), .C1(n6595), 
        .C2(n6628), .ZN(U3194) );
  AOI22_X1 U7560 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6662), .ZN(n6594) );
  OAI21_X1 U7561 ( .B1(n6595), .B2(n6625), .A(n6594), .ZN(U3195) );
  AOI22_X1 U7562 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6662), .ZN(n6596) );
  OAI21_X1 U7563 ( .B1(n6597), .B2(n6628), .A(n6596), .ZN(U3196) );
  AOI22_X1 U7564 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6662), .ZN(n6598) );
  OAI21_X1 U7565 ( .B1(n6599), .B2(n6628), .A(n6598), .ZN(U3197) );
  AOI22_X1 U7566 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6662), .ZN(n6600) );
  OAI21_X1 U7567 ( .B1(n6601), .B2(n6628), .A(n6600), .ZN(U3198) );
  AOI22_X1 U7568 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6662), .ZN(n6602) );
  OAI21_X1 U7569 ( .B1(n6604), .B2(n6628), .A(n6602), .ZN(U3199) );
  AOI22_X1 U7570 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6662), .ZN(n6603) );
  OAI21_X1 U7571 ( .B1(n6604), .B2(n6625), .A(n6603), .ZN(U3200) );
  AOI22_X1 U7572 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6662), .ZN(n6605) );
  OAI21_X1 U7573 ( .B1(n6606), .B2(n6625), .A(n6605), .ZN(U3201) );
  INV_X1 U7574 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6609) );
  AOI22_X1 U7575 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6607), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6662), .ZN(n6608) );
  OAI21_X1 U7576 ( .B1(n6609), .B2(n6625), .A(n6608), .ZN(U3202) );
  INV_X1 U7577 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6611) );
  AOI22_X1 U7578 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6662), .ZN(n6610) );
  OAI21_X1 U7579 ( .B1(n6611), .B2(n6628), .A(n6610), .ZN(U3203) );
  INV_X1 U7580 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7581 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6662), .ZN(n6612) );
  OAI21_X1 U7582 ( .B1(n6945), .B2(n6628), .A(n6612), .ZN(U3204) );
  AOI22_X1 U7583 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6662), .ZN(n6613) );
  OAI21_X1 U7584 ( .B1(n6614), .B2(n6628), .A(n6613), .ZN(U3205) );
  AOI22_X1 U7585 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6662), .ZN(n6615) );
  OAI21_X1 U7586 ( .B1(n6756), .B2(n6628), .A(n6615), .ZN(U3206) );
  AOI22_X1 U7587 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6662), .ZN(n6616) );
  OAI21_X1 U7588 ( .B1(n6617), .B2(n6628), .A(n6616), .ZN(U3207) );
  AOI22_X1 U7589 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6662), .ZN(n6618) );
  OAI21_X1 U7590 ( .B1(n5723), .B2(n6628), .A(n6618), .ZN(U3208) );
  INV_X1 U7591 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6619) );
  OAI222_X1 U7592 ( .A1(n6625), .A2(n5723), .B1(n6619), .B2(n6679), .C1(n6621), 
        .C2(n6628), .ZN(U3209) );
  INV_X1 U7593 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6620) );
  OAI222_X1 U7594 ( .A1(n6625), .A2(n6621), .B1(n6620), .B2(n6679), .C1(n6989), 
        .C2(n6628), .ZN(U3210) );
  INV_X1 U7595 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6622) );
  OAI222_X1 U7596 ( .A1(n6625), .A2(n6989), .B1(n6622), .B2(n6679), .C1(n6624), 
        .C2(n6628), .ZN(U3211) );
  INV_X1 U7597 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6623) );
  OAI222_X1 U7598 ( .A1(n6625), .A2(n6624), .B1(n6623), .B2(n6679), .C1(n6968), 
        .C2(n6628), .ZN(U3212) );
  INV_X1 U7599 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U7600 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6626), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6662), .ZN(n6627) );
  OAI21_X1 U7601 ( .B1(n6629), .B2(n6628), .A(n6627), .ZN(U3213) );
  MUX2_X1 U7602 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6679), .Z(U3445) );
  MUX2_X1 U7603 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6679), .Z(U3446) );
  MUX2_X1 U7604 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6679), .Z(U3447) );
  MUX2_X1 U7605 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6679), .Z(U3448) );
  INV_X1 U7606 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6632) );
  INV_X1 U7607 ( .A(n6633), .ZN(n6630) );
  AOI21_X1 U7608 ( .B1(n6632), .B2(n6631), .A(n6630), .ZN(U3451) );
  OAI21_X1 U7609 ( .B1(n6635), .B2(n6634), .A(n6633), .ZN(U3452) );
  OAI211_X1 U7610 ( .C1(n6959), .C2(n6638), .A(n6637), .B(n6636), .ZN(U3453)
         );
  INV_X1 U7611 ( .A(n6639), .ZN(n6642) );
  OAI22_X1 U7612 ( .A1(n6642), .A2(n6651), .B1(n6641), .B2(n6640), .ZN(n6644)
         );
  MUX2_X1 U7613 ( .A(n6644), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6643), 
        .Z(U3456) );
  OAI22_X1 U7614 ( .A1(n6646), .A2(n6651), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6645), .ZN(n6648) );
  OAI22_X1 U7615 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6649), .B1(n6648), .B2(n6647), .ZN(n6650) );
  OAI21_X1 U7616 ( .B1(n6652), .B2(n6651), .A(n6650), .ZN(U3461) );
  AOI21_X1 U7617 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6653) );
  AOI22_X1 U7618 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6653), .B2(n5186), .ZN(n6655) );
  INV_X1 U7619 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7620 ( .A1(n6656), .A2(n6655), .B1(n6654), .B2(n6659), .ZN(U3468)
         );
  INV_X1 U7621 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U7622 ( .A1(n6659), .A2(REIP_REG_1__SCAN_IN), .ZN(n6657) );
  AOI22_X1 U7623 ( .A1(n6660), .A2(n6659), .B1(n6658), .B2(n6657), .ZN(U3469)
         );
  NAND2_X1 U7624 ( .A1(n6662), .A2(W_R_N_REG_SCAN_IN), .ZN(n6661) );
  OAI21_X1 U7625 ( .B1(n6662), .B2(READREQUEST_REG_SCAN_IN), .A(n6661), .ZN(
        U3470) );
  AOI211_X1 U7626 ( .C1(n6666), .C2(n6665), .A(n6664), .B(n6663), .ZN(n6667)
         );
  INV_X1 U7627 ( .A(n6667), .ZN(n6678) );
  OAI21_X1 U7628 ( .B1(n6671), .B2(n6941), .A(n6668), .ZN(n6669) );
  NAND3_X1 U7629 ( .A1(n6669), .A2(STATE2_REG_2__SCAN_IN), .A3(n6666), .ZN(
        n6670) );
  AOI21_X1 U7630 ( .B1(n6672), .B2(n6671), .A(n6670), .ZN(n6673) );
  NOR2_X1 U7631 ( .A1(n6673), .A2(n6786), .ZN(n6674) );
  OAI21_X1 U7632 ( .B1(n6675), .B2(n6674), .A(n6678), .ZN(n6676) );
  OAI21_X1 U7633 ( .B1(n6678), .B2(n6677), .A(n6676), .ZN(U3472) );
  MUX2_X1 U7634 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6679), .Z(U3473) );
  AOI222_X1 U7635 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6682), .B1(n6681), .B2(
        LWORD_REG_13__SCAN_IN), .C1(n6680), .C2(DATAO_REG_13__SCAN_IN), .ZN(
        n7009) );
  INV_X1 U7636 ( .A(keyinput50), .ZN(n6684) );
  AOI22_X1 U7637 ( .A1(n6685), .A2(keyinput97), .B1(DATAO_REG_14__SCAN_IN), 
        .B2(n6684), .ZN(n6683) );
  OAI221_X1 U7638 ( .B1(n6685), .B2(keyinput97), .C1(n6684), .C2(
        DATAO_REG_14__SCAN_IN), .A(n6683), .ZN(n6698) );
  INV_X1 U7639 ( .A(keyinput114), .ZN(n6687) );
  AOI22_X1 U7640 ( .A1(n6688), .A2(keyinput4), .B1(ADDRESS_REG_27__SCAN_IN), 
        .B2(n6687), .ZN(n6686) );
  OAI221_X1 U7641 ( .B1(n6688), .B2(keyinput4), .C1(n6687), .C2(
        ADDRESS_REG_27__SCAN_IN), .A(n6686), .ZN(n6697) );
  INV_X1 U7642 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6690) );
  AOI22_X1 U7643 ( .A1(n6691), .A2(keyinput23), .B1(n6690), .B2(keyinput9), 
        .ZN(n6689) );
  OAI221_X1 U7644 ( .B1(n6691), .B2(keyinput23), .C1(n6690), .C2(keyinput9), 
        .A(n6689), .ZN(n6696) );
  AOI22_X1 U7645 ( .A1(n6694), .A2(keyinput79), .B1(n6693), .B2(keyinput53), 
        .ZN(n6692) );
  OAI221_X1 U7646 ( .B1(n6694), .B2(keyinput79), .C1(n6693), .C2(keyinput53), 
        .A(n6692), .ZN(n6695) );
  NOR4_X1 U7647 ( .A1(n6698), .A2(n6697), .A3(n6696), .A4(n6695), .ZN(n6747)
         );
  INV_X1 U7648 ( .A(keyinput82), .ZN(n6700) );
  AOI22_X1 U7649 ( .A1(n6701), .A2(keyinput20), .B1(DATAWIDTH_REG_27__SCAN_IN), 
        .B2(n6700), .ZN(n6699) );
  OAI221_X1 U7650 ( .B1(n6701), .B2(keyinput20), .C1(n6700), .C2(
        DATAWIDTH_REG_27__SCAN_IN), .A(n6699), .ZN(n6713) );
  AOI22_X1 U7651 ( .A1(n6704), .A2(keyinput33), .B1(keyinput122), .B2(n6703), 
        .ZN(n6702) );
  OAI221_X1 U7652 ( .B1(n6704), .B2(keyinput33), .C1(n6703), .C2(keyinput122), 
        .A(n6702), .ZN(n6712) );
  INV_X1 U7653 ( .A(keyinput105), .ZN(n6706) );
  AOI22_X1 U7654 ( .A1(n3949), .A2(keyinput104), .B1(DATAO_REG_15__SCAN_IN), 
        .B2(n6706), .ZN(n6705) );
  OAI221_X1 U7655 ( .B1(n3949), .B2(keyinput104), .C1(n6706), .C2(
        DATAO_REG_15__SCAN_IN), .A(n6705), .ZN(n6711) );
  INV_X1 U7656 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6709) );
  INV_X1 U7657 ( .A(keyinput96), .ZN(n6708) );
  AOI22_X1 U7658 ( .A1(n6709), .A2(keyinput48), .B1(ADDRESS_REG_4__SCAN_IN), 
        .B2(n6708), .ZN(n6707) );
  OAI221_X1 U7659 ( .B1(n6709), .B2(keyinput48), .C1(n6708), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6707), .ZN(n6710) );
  NOR4_X1 U7660 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6746)
         );
  INV_X1 U7661 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U7662 ( .A1(n5241), .A2(keyinput120), .B1(n6715), .B2(keyinput108), 
        .ZN(n6714) );
  OAI221_X1 U7663 ( .B1(n5241), .B2(keyinput120), .C1(n6715), .C2(keyinput108), 
        .A(n6714), .ZN(n6728) );
  INV_X1 U7664 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6717) );
  AOI22_X1 U7665 ( .A1(n6718), .A2(keyinput58), .B1(n6717), .B2(keyinput43), 
        .ZN(n6716) );
  OAI221_X1 U7666 ( .B1(n6718), .B2(keyinput58), .C1(n6717), .C2(keyinput43), 
        .A(n6716), .ZN(n6727) );
  INV_X1 U7667 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6720) );
  AOI22_X1 U7668 ( .A1(n6721), .A2(keyinput101), .B1(n6720), .B2(keyinput1), 
        .ZN(n6719) );
  OAI221_X1 U7669 ( .B1(n6721), .B2(keyinput101), .C1(n6720), .C2(keyinput1), 
        .A(n6719), .ZN(n6726) );
  AOI22_X1 U7670 ( .A1(n6724), .A2(keyinput91), .B1(n6723), .B2(keyinput37), 
        .ZN(n6722) );
  OAI221_X1 U7671 ( .B1(n6724), .B2(keyinput91), .C1(n6723), .C2(keyinput37), 
        .A(n6722), .ZN(n6725) );
  NOR4_X1 U7672 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(n6745)
         );
  INV_X1 U7673 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6730) );
  AOI22_X1 U7674 ( .A1(n6731), .A2(keyinput38), .B1(n6730), .B2(keyinput93), 
        .ZN(n6729) );
  OAI221_X1 U7675 ( .B1(n6731), .B2(keyinput38), .C1(n6730), .C2(keyinput93), 
        .A(n6729), .ZN(n6743) );
  INV_X1 U7676 ( .A(keyinput60), .ZN(n6733) );
  AOI22_X1 U7677 ( .A1(n6734), .A2(keyinput74), .B1(ADDRESS_REG_2__SCAN_IN), 
        .B2(n6733), .ZN(n6732) );
  OAI221_X1 U7678 ( .B1(n6734), .B2(keyinput74), .C1(n6733), .C2(
        ADDRESS_REG_2__SCAN_IN), .A(n6732), .ZN(n6742) );
  INV_X1 U7679 ( .A(keyinput34), .ZN(n6736) );
  AOI22_X1 U7680 ( .A1(n6226), .A2(keyinput99), .B1(ADDRESS_REG_28__SCAN_IN), 
        .B2(n6736), .ZN(n6735) );
  OAI221_X1 U7681 ( .B1(n6226), .B2(keyinput99), .C1(n6736), .C2(
        ADDRESS_REG_28__SCAN_IN), .A(n6735), .ZN(n6741) );
  AOI22_X1 U7682 ( .A1(n6739), .A2(keyinput63), .B1(n6738), .B2(keyinput78), 
        .ZN(n6737) );
  OAI221_X1 U7683 ( .B1(n6739), .B2(keyinput63), .C1(n6738), .C2(keyinput78), 
        .A(n6737), .ZN(n6740) );
  NOR4_X1 U7684 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6744)
         );
  NAND4_X1 U7685 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n7007)
         );
  AOI22_X1 U7686 ( .A1(n6750), .A2(keyinput52), .B1(n6749), .B2(keyinput109), 
        .ZN(n6748) );
  OAI221_X1 U7687 ( .B1(n6750), .B2(keyinput52), .C1(n6749), .C2(keyinput109), 
        .A(n6748), .ZN(n6763) );
  INV_X1 U7688 ( .A(keyinput24), .ZN(n6753) );
  INV_X1 U7689 ( .A(keyinput12), .ZN(n6752) );
  AOI22_X1 U7690 ( .A1(n6753), .A2(ADDRESS_REG_8__SCAN_IN), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(n6752), .ZN(n6751) );
  OAI221_X1 U7691 ( .B1(n6753), .B2(ADDRESS_REG_8__SCAN_IN), .C1(n6752), .C2(
        DATAWIDTH_REG_17__SCAN_IN), .A(n6751), .ZN(n6762) );
  INV_X1 U7692 ( .A(keyinput90), .ZN(n6755) );
  AOI22_X1 U7693 ( .A1(n6756), .A2(keyinput51), .B1(DATAWIDTH_REG_15__SCAN_IN), 
        .B2(n6755), .ZN(n6754) );
  OAI221_X1 U7694 ( .B1(n6756), .B2(keyinput51), .C1(n6755), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6754), .ZN(n6761) );
  INV_X1 U7695 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6759) );
  INV_X1 U7696 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6758) );
  AOI22_X1 U7697 ( .A1(n6759), .A2(keyinput65), .B1(n6758), .B2(keyinput31), 
        .ZN(n6757) );
  OAI221_X1 U7698 ( .B1(n6759), .B2(keyinput65), .C1(n6758), .C2(keyinput31), 
        .A(n6757), .ZN(n6760) );
  NOR4_X1 U7699 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6812)
         );
  INV_X1 U7700 ( .A(keyinput98), .ZN(n6900) );
  AOI22_X1 U7701 ( .A1(n6765), .A2(keyinput40), .B1(DATAO_REG_4__SCAN_IN), 
        .B2(n6900), .ZN(n6764) );
  OAI221_X1 U7702 ( .B1(n6765), .B2(keyinput40), .C1(n6900), .C2(
        DATAO_REG_4__SCAN_IN), .A(n6764), .ZN(n6778) );
  INV_X1 U7703 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7704 ( .A1(n6768), .A2(keyinput55), .B1(n6767), .B2(keyinput123), 
        .ZN(n6766) );
  OAI221_X1 U7705 ( .B1(n6768), .B2(keyinput55), .C1(n6767), .C2(keyinput123), 
        .A(n6766), .ZN(n6777) );
  INV_X1 U7706 ( .A(keyinput86), .ZN(n6770) );
  AOI22_X1 U7707 ( .A1(n6771), .A2(keyinput17), .B1(LWORD_REG_1__SCAN_IN), 
        .B2(n6770), .ZN(n6769) );
  OAI221_X1 U7708 ( .B1(n6771), .B2(keyinput17), .C1(n6770), .C2(
        LWORD_REG_1__SCAN_IN), .A(n6769), .ZN(n6776) );
  INV_X1 U7709 ( .A(keyinput28), .ZN(n6773) );
  AOI22_X1 U7710 ( .A1(n6774), .A2(keyinput80), .B1(UWORD_REG_12__SCAN_IN), 
        .B2(n6773), .ZN(n6772) );
  OAI221_X1 U7711 ( .B1(n6774), .B2(keyinput80), .C1(n6773), .C2(
        UWORD_REG_12__SCAN_IN), .A(n6772), .ZN(n6775) );
  NOR4_X1 U7712 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6811)
         );
  INV_X1 U7713 ( .A(keyinput2), .ZN(n6780) );
  AOI22_X1 U7714 ( .A1(n5261), .A2(keyinput25), .B1(LWORD_REG_4__SCAN_IN), 
        .B2(n6780), .ZN(n6779) );
  OAI221_X1 U7715 ( .B1(n5261), .B2(keyinput25), .C1(n6780), .C2(
        LWORD_REG_4__SCAN_IN), .A(n6779), .ZN(n6793) );
  INV_X1 U7716 ( .A(DATAI_19_), .ZN(n6783) );
  INV_X1 U7717 ( .A(keyinput19), .ZN(n6782) );
  AOI22_X1 U7718 ( .A1(n6783), .A2(keyinput94), .B1(ADS_N_REG_SCAN_IN), .B2(
        n6782), .ZN(n6781) );
  OAI221_X1 U7719 ( .B1(n6783), .B2(keyinput94), .C1(n6782), .C2(
        ADS_N_REG_SCAN_IN), .A(n6781), .ZN(n6792) );
  INV_X1 U7720 ( .A(keyinput68), .ZN(n6785) );
  AOI22_X1 U7721 ( .A1(n6786), .A2(keyinput115), .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n6785), .ZN(n6784) );
  OAI221_X1 U7722 ( .B1(n6786), .B2(keyinput115), .C1(n6785), .C2(
        BYTEENABLE_REG_0__SCAN_IN), .A(n6784), .ZN(n6791) );
  INV_X1 U7723 ( .A(DATAI_16_), .ZN(n6789) );
  INV_X1 U7724 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7725 ( .A1(n6789), .A2(keyinput92), .B1(n6788), .B2(keyinput56), 
        .ZN(n6787) );
  OAI221_X1 U7726 ( .B1(n6789), .B2(keyinput92), .C1(n6788), .C2(keyinput56), 
        .A(n6787), .ZN(n6790) );
  NOR4_X1 U7727 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6810)
         );
  INV_X1 U7728 ( .A(keyinput61), .ZN(n6795) );
  AOI22_X1 U7729 ( .A1(n6796), .A2(keyinput112), .B1(LWORD_REG_8__SCAN_IN), 
        .B2(n6795), .ZN(n6794) );
  OAI221_X1 U7730 ( .B1(n6796), .B2(keyinput112), .C1(n6795), .C2(
        LWORD_REG_8__SCAN_IN), .A(n6794), .ZN(n6808) );
  INV_X1 U7731 ( .A(keyinput125), .ZN(n6798) );
  AOI22_X1 U7732 ( .A1(n6799), .A2(keyinput66), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n6798), .ZN(n6797) );
  OAI221_X1 U7733 ( .B1(n6799), .B2(keyinput66), .C1(n6798), .C2(
        DATAO_REG_31__SCAN_IN), .A(n6797), .ZN(n6807) );
  INV_X1 U7734 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6801) );
  AOI22_X1 U7735 ( .A1(n6802), .A2(keyinput32), .B1(n6801), .B2(keyinput76), 
        .ZN(n6800) );
  OAI221_X1 U7736 ( .B1(n6802), .B2(keyinput32), .C1(n6801), .C2(keyinput76), 
        .A(n6800), .ZN(n6806) );
  XNOR2_X1 U7737 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .B(keyinput88), .ZN(n6804)
         );
  XNOR2_X1 U7738 ( .A(keyinput89), .B(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6803)
         );
  NAND2_X1 U7739 ( .A1(n6804), .A2(n6803), .ZN(n6805) );
  NOR4_X1 U7740 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6809)
         );
  NAND4_X1 U7741 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n7006)
         );
  INV_X1 U7742 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7743 ( .A1(n6815), .A2(keyinput49), .B1(keyinput107), .B2(n6814), 
        .ZN(n6813) );
  OAI221_X1 U7744 ( .B1(n6815), .B2(keyinput49), .C1(n6814), .C2(keyinput107), 
        .A(n6813), .ZN(n6827) );
  INV_X1 U7745 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6817) );
  AOI22_X1 U7746 ( .A1(n6818), .A2(keyinput42), .B1(n6817), .B2(keyinput85), 
        .ZN(n6816) );
  OAI221_X1 U7747 ( .B1(n6818), .B2(keyinput42), .C1(n6817), .C2(keyinput85), 
        .A(n6816), .ZN(n6826) );
  INV_X1 U7748 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U7749 ( .A1(n6821), .A2(keyinput54), .B1(n6820), .B2(keyinput126), 
        .ZN(n6819) );
  OAI221_X1 U7750 ( .B1(n6821), .B2(keyinput54), .C1(n6820), .C2(keyinput126), 
        .A(n6819), .ZN(n6825) );
  INV_X1 U7751 ( .A(keyinput18), .ZN(n6823) );
  AOI22_X1 U7752 ( .A1(n6217), .A2(keyinput75), .B1(BYTEENABLE_REG_3__SCAN_IN), 
        .B2(n6823), .ZN(n6822) );
  OAI221_X1 U7753 ( .B1(n6217), .B2(keyinput75), .C1(n6823), .C2(
        BYTEENABLE_REG_3__SCAN_IN), .A(n6822), .ZN(n6824) );
  NOR4_X1 U7754 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n6874)
         );
  NAND2_X1 U7755 ( .A1(n4350), .A2(keyinput73), .ZN(n6828) );
  OAI221_X1 U7756 ( .B1(n6829), .B2(keyinput127), .C1(n4350), .C2(keyinput73), 
        .A(n6828), .ZN(n6840) );
  INV_X1 U7757 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6832) );
  AOI22_X1 U7758 ( .A1(n6832), .A2(keyinput41), .B1(keyinput11), .B2(n6831), 
        .ZN(n6830) );
  OAI221_X1 U7759 ( .B1(n6832), .B2(keyinput41), .C1(n6831), .C2(keyinput11), 
        .A(n6830), .ZN(n6839) );
  INV_X1 U7760 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7761 ( .A1(n4003), .A2(keyinput29), .B1(n6834), .B2(keyinput119), 
        .ZN(n6833) );
  OAI221_X1 U7762 ( .B1(n4003), .B2(keyinput29), .C1(n6834), .C2(keyinput119), 
        .A(n6833), .ZN(n6838) );
  AOI22_X1 U7763 ( .A1(n6836), .A2(keyinput16), .B1(keyinput81), .B2(n6238), 
        .ZN(n6835) );
  OAI221_X1 U7764 ( .B1(n6836), .B2(keyinput16), .C1(n6238), .C2(keyinput81), 
        .A(n6835), .ZN(n6837) );
  NOR4_X1 U7765 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6873)
         );
  INV_X1 U7766 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6843) );
  INV_X1 U7767 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6842) );
  AOI22_X1 U7768 ( .A1(n6843), .A2(keyinput71), .B1(keyinput103), .B2(n6842), 
        .ZN(n6841) );
  OAI221_X1 U7769 ( .B1(n6843), .B2(keyinput71), .C1(n6842), .C2(keyinput103), 
        .A(n6841), .ZN(n6856) );
  INV_X1 U7770 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6846) );
  INV_X1 U7771 ( .A(DATAI_15_), .ZN(n6845) );
  AOI22_X1 U7772 ( .A1(n6846), .A2(keyinput30), .B1(keyinput77), .B2(n6845), 
        .ZN(n6844) );
  OAI221_X1 U7773 ( .B1(n6846), .B2(keyinput30), .C1(n6845), .C2(keyinput77), 
        .A(n6844), .ZN(n6855) );
  INV_X1 U7774 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6848) );
  INV_X1 U7775 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6852) );
  INV_X1 U7776 ( .A(keyinput62), .ZN(n6851) );
  AOI22_X1 U7777 ( .A1(n6852), .A2(keyinput69), .B1(ADDRESS_REG_25__SCAN_IN), 
        .B2(n6851), .ZN(n6850) );
  OAI221_X1 U7778 ( .B1(n6852), .B2(keyinput69), .C1(n6851), .C2(
        ADDRESS_REG_25__SCAN_IN), .A(n6850), .ZN(n6853) );
  NOR4_X1 U7779 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6872)
         );
  INV_X1 U7780 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6858) );
  AOI22_X1 U7781 ( .A1(n5186), .A2(keyinput39), .B1(n6858), .B2(keyinput83), 
        .ZN(n6857) );
  OAI221_X1 U7782 ( .B1(n5186), .B2(keyinput39), .C1(n6858), .C2(keyinput83), 
        .A(n6857), .ZN(n6870) );
  AOI22_X1 U7783 ( .A1(n5542), .A2(keyinput121), .B1(keyinput113), .B2(n6860), 
        .ZN(n6859) );
  OAI221_X1 U7784 ( .B1(n5542), .B2(keyinput121), .C1(n6860), .C2(keyinput113), 
        .A(n6859), .ZN(n6869) );
  AOI22_X1 U7785 ( .A1(n6863), .A2(keyinput22), .B1(n6862), .B2(keyinput124), 
        .ZN(n6861) );
  OAI221_X1 U7786 ( .B1(n6863), .B2(keyinput22), .C1(n6862), .C2(keyinput124), 
        .A(n6861), .ZN(n6868) );
  AOI22_X1 U7787 ( .A1(n6866), .A2(keyinput102), .B1(n6865), .B2(keyinput72), 
        .ZN(n6864) );
  OAI221_X1 U7788 ( .B1(n6866), .B2(keyinput102), .C1(n6865), .C2(keyinput72), 
        .A(n6864), .ZN(n6867) );
  NOR4_X1 U7789 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n6871)
         );
  NAND4_X1 U7790 ( .A1(n6874), .A2(n6873), .A3(n6872), .A4(n6871), .ZN(n7005)
         );
  INV_X1 U7791 ( .A(keyinput58), .ZN(n6875) );
  NOR4_X1 U7792 ( .A1(keyinput108), .A2(keyinput1), .A3(keyinput91), .A4(n6875), .ZN(n6876) );
  NAND3_X1 U7793 ( .A1(keyinput43), .A2(keyinput101), .A3(n6876), .ZN(n6888)
         );
  NAND4_X1 U7794 ( .A1(keyinput60), .A2(keyinput34), .A3(keyinput99), .A4(
        keyinput63), .ZN(n6877) );
  NOR3_X1 U7795 ( .A1(keyinput93), .A2(keyinput74), .A3(n6877), .ZN(n6886) );
  NAND4_X1 U7796 ( .A1(keyinput50), .A2(keyinput114), .A3(keyinput9), .A4(
        keyinput79), .ZN(n6883) );
  NOR2_X1 U7797 ( .A1(keyinput68), .A2(keyinput23), .ZN(n6878) );
  NAND3_X1 U7798 ( .A1(keyinput97), .A2(keyinput4), .A3(n6878), .ZN(n6882) );
  INV_X1 U7799 ( .A(keyinput122), .ZN(n6879) );
  NAND4_X1 U7800 ( .A1(keyinput105), .A2(keyinput104), .A3(keyinput48), .A4(
        n6879), .ZN(n6881) );
  NAND4_X1 U7801 ( .A1(keyinput53), .A2(keyinput20), .A3(keyinput82), .A4(
        keyinput33), .ZN(n6880) );
  NOR4_X1 U7802 ( .A1(n6883), .A2(n6882), .A3(n6881), .A4(n6880), .ZN(n6885)
         );
  INV_X1 U7803 ( .A(keyinput38), .ZN(n6884) );
  NAND4_X1 U7804 ( .A1(keyinput37), .A2(n6886), .A3(n6885), .A4(n6884), .ZN(
        n6887) );
  NOR4_X1 U7805 ( .A1(keyinput96), .A2(keyinput120), .A3(n6888), .A4(n6887), 
        .ZN(n6935) );
  NAND4_X1 U7806 ( .A1(keyinput113), .A2(keyinput39), .A3(keyinput83), .A4(
        keyinput102), .ZN(n6933) );
  NOR3_X1 U7807 ( .A1(keyinput126), .A2(keyinput22), .A3(keyinput121), .ZN(
        n6889) );
  NAND2_X1 U7808 ( .A1(keyinput72), .A2(n6889), .ZN(n6932) );
  NAND4_X1 U7809 ( .A1(keyinput107), .A2(keyinput75), .A3(keyinput18), .A4(
        keyinput54), .ZN(n6890) );
  NOR3_X1 U7810 ( .A1(keyinput85), .A2(keyinput49), .A3(n6890), .ZN(n6899) );
  INV_X1 U7811 ( .A(keyinput11), .ZN(n6891) );
  NOR4_X1 U7812 ( .A1(keyinput41), .A2(keyinput73), .A3(keyinput16), .A4(n6891), .ZN(n6892) );
  NAND4_X1 U7813 ( .A1(keyinput46), .A2(keyinput81), .A3(keyinput29), .A4(
        n6892), .ZN(n6897) );
  NAND2_X1 U7814 ( .A1(keyinput69), .A2(keyinput103), .ZN(n6893) );
  NOR3_X1 U7815 ( .A1(keyinput62), .A2(keyinput110), .A3(n6893), .ZN(n6895) );
  INV_X1 U7816 ( .A(keyinput124), .ZN(n6894) );
  NAND3_X1 U7817 ( .A1(keyinput30), .A2(n6895), .A3(n6894), .ZN(n6896) );
  NOR4_X1 U7818 ( .A1(keyinput71), .A2(keyinput77), .A3(n6897), .A4(n6896), 
        .ZN(n6898) );
  NAND4_X1 U7819 ( .A1(keyinput119), .A2(keyinput42), .A3(n6899), .A4(n6898), 
        .ZN(n6931) );
  NOR4_X1 U7820 ( .A1(keyinput80), .A2(keyinput28), .A3(keyinput17), .A4(n6900), .ZN(n6929) );
  NAND3_X1 U7821 ( .A1(keyinput40), .A2(keyinput123), .A3(keyinput13), .ZN(
        n6901) );
  NOR2_X1 U7822 ( .A1(keyinput55), .A2(n6901), .ZN(n6928) );
  NOR4_X1 U7823 ( .A1(keyinput109), .A2(keyinput65), .A3(keyinput31), .A4(
        keyinput51), .ZN(n6902) );
  NAND3_X1 U7824 ( .A1(keyinput86), .A2(keyinput24), .A3(n6902), .ZN(n6911) );
  INV_X1 U7825 ( .A(keyinput112), .ZN(n6903) );
  NOR4_X1 U7826 ( .A1(keyinput125), .A2(keyinput61), .A3(keyinput89), .A4(
        n6903), .ZN(n6909) );
  NAND3_X1 U7827 ( .A1(keyinput66), .A2(keyinput76), .A3(keyinput32), .ZN(
        n6904) );
  NOR2_X1 U7828 ( .A1(keyinput90), .A2(n6904), .ZN(n6908) );
  NAND3_X1 U7829 ( .A1(keyinput56), .A2(keyinput19), .A3(keyinput2), .ZN(n6905) );
  NOR2_X1 U7830 ( .A1(keyinput115), .A2(n6905), .ZN(n6907) );
  NOR4_X1 U7831 ( .A1(keyinput88), .A2(keyinput94), .A3(keyinput25), .A4(
        keyinput92), .ZN(n6906) );
  NAND4_X1 U7832 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n6910)
         );
  NOR4_X1 U7833 ( .A1(keyinput12), .A2(keyinput52), .A3(n6911), .A4(n6910), 
        .ZN(n6927) );
  NAND2_X1 U7834 ( .A1(keyinput14), .A2(keyinput0), .ZN(n6912) );
  NOR3_X1 U7835 ( .A1(keyinput5), .A2(keyinput59), .A3(n6912), .ZN(n6913) );
  NAND3_X1 U7836 ( .A1(keyinput87), .A2(keyinput106), .A3(n6913), .ZN(n6925)
         );
  NAND4_X1 U7837 ( .A1(keyinput36), .A2(keyinput67), .A3(keyinput6), .A4(
        keyinput15), .ZN(n6914) );
  NOR3_X1 U7838 ( .A1(keyinput78), .A2(keyinput44), .A3(n6914), .ZN(n6923) );
  INV_X1 U7839 ( .A(keyinput118), .ZN(n6915) );
  NAND4_X1 U7840 ( .A1(keyinput7), .A2(keyinput116), .A3(keyinput111), .A4(
        n6915), .ZN(n6921) );
  OR4_X1 U7841 ( .A1(keyinput95), .A2(keyinput57), .A3(keyinput70), .A4(
        keyinput8), .ZN(n6920) );
  INV_X1 U7842 ( .A(keyinput45), .ZN(n6916) );
  NAND4_X1 U7843 ( .A1(keyinput117), .A2(keyinput64), .A3(keyinput21), .A4(
        n6916), .ZN(n6919) );
  NOR2_X1 U7844 ( .A1(keyinput84), .A2(keyinput35), .ZN(n6917) );
  NAND3_X1 U7845 ( .A1(keyinput47), .A2(keyinput100), .A3(n6917), .ZN(n6918)
         );
  NOR4_X1 U7846 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6922)
         );
  NAND4_X1 U7847 ( .A1(keyinput26), .A2(keyinput27), .A3(n6923), .A4(n6922), 
        .ZN(n6924) );
  NOR4_X1 U7848 ( .A1(keyinput10), .A2(keyinput3), .A3(n6925), .A4(n6924), 
        .ZN(n6926) );
  NAND4_X1 U7849 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6930)
         );
  NOR4_X1 U7850 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n6934)
         );
  AOI21_X1 U7851 ( .B1(n6935), .B2(n6934), .A(keyinput127), .ZN(n7003) );
  INV_X1 U7852 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6938) );
  INV_X1 U7853 ( .A(keyinput67), .ZN(n6937) );
  AOI22_X1 U7854 ( .A1(n6938), .A2(keyinput6), .B1(UWORD_REG_10__SCAN_IN), 
        .B2(n6937), .ZN(n6936) );
  OAI221_X1 U7855 ( .B1(n6938), .B2(keyinput6), .C1(n6937), .C2(
        UWORD_REG_10__SCAN_IN), .A(n6936), .ZN(n6951) );
  AOI22_X1 U7856 ( .A1(n6941), .A2(keyinput15), .B1(n6940), .B2(keyinput95), 
        .ZN(n6939) );
  OAI221_X1 U7857 ( .B1(n6941), .B2(keyinput15), .C1(n6940), .C2(keyinput95), 
        .A(n6939), .ZN(n6950) );
  INV_X1 U7858 ( .A(keyinput36), .ZN(n6943) );
  AOI22_X1 U7859 ( .A1(n6944), .A2(keyinput27), .B1(UWORD_REG_9__SCAN_IN), 
        .B2(n6943), .ZN(n6942) );
  OAI221_X1 U7860 ( .B1(n6944), .B2(keyinput27), .C1(n6943), .C2(
        UWORD_REG_9__SCAN_IN), .A(n6942), .ZN(n6949) );
  XOR2_X1 U7861 ( .A(n6945), .B(keyinput26), .Z(n6947) );
  XNOR2_X1 U7862 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .B(keyinput44), .ZN(n6946) );
  NAND2_X1 U7863 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  NOR4_X1 U7864 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n7002)
         );
  INV_X1 U7865 ( .A(keyinput106), .ZN(n6953) );
  OAI22_X1 U7866 ( .A1(n6223), .A2(keyinput10), .B1(n6953), .B2(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6952) );
  AOI221_X1 U7867 ( .B1(n6223), .B2(keyinput10), .C1(DATAWIDTH_REG_30__SCAN_IN), .C2(n6953), .A(n6952), .ZN(n6966) );
  INV_X1 U7868 ( .A(keyinput3), .ZN(n6955) );
  OAI22_X1 U7869 ( .A1(n6956), .A2(keyinput0), .B1(n6955), .B2(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6954) );
  AOI221_X1 U7870 ( .B1(n6956), .B2(keyinput0), .C1(DATAWIDTH_REG_10__SCAN_IN), 
        .C2(n6955), .A(n6954), .ZN(n6965) );
  OAI22_X1 U7871 ( .A1(n6959), .A2(keyinput5), .B1(n6958), .B2(keyinput14), 
        .ZN(n6957) );
  AOI221_X1 U7872 ( .B1(n6959), .B2(keyinput5), .C1(keyinput14), .C2(n6958), 
        .A(n6957), .ZN(n6964) );
  INV_X1 U7873 ( .A(keyinput46), .ZN(n6961) );
  OAI22_X1 U7874 ( .A1(n6962), .A2(keyinput59), .B1(n6961), .B2(NA_N), .ZN(
        n6960) );
  AOI221_X1 U7875 ( .B1(n6962), .B2(keyinput59), .C1(NA_N), .C2(n6961), .A(
        n6960), .ZN(n6963) );
  NAND4_X1 U7876 ( .A1(n6966), .A2(n6965), .A3(n6964), .A4(n6963), .ZN(n6987)
         );
  OAI22_X1 U7877 ( .A1(n6969), .A2(keyinput35), .B1(n6968), .B2(keyinput84), 
        .ZN(n6967) );
  AOI221_X1 U7878 ( .B1(n6969), .B2(keyinput35), .C1(keyinput84), .C2(n6968), 
        .A(n6967), .ZN(n6978) );
  INV_X1 U7879 ( .A(keyinput117), .ZN(n6971) );
  OAI22_X1 U7880 ( .A1(n6972), .A2(keyinput45), .B1(n6971), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n6970) );
  AOI221_X1 U7881 ( .B1(n6972), .B2(keyinput45), .C1(ADDRESS_REG_26__SCAN_IN), 
        .C2(n6971), .A(n6970), .ZN(n6977) );
  INV_X1 U7882 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6975) );
  OAI22_X1 U7883 ( .A1(n6975), .A2(keyinput21), .B1(n6974), .B2(keyinput87), 
        .ZN(n6973) );
  AOI221_X1 U7884 ( .B1(n6975), .B2(keyinput21), .C1(keyinput87), .C2(n6974), 
        .A(n6973), .ZN(n6976) );
  NAND3_X1 U7885 ( .A1(n6978), .A2(n6977), .A3(n6976), .ZN(n6986) );
  INV_X1 U7886 ( .A(keyinput116), .ZN(n6980) );
  INV_X1 U7887 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6979) );
  XNOR2_X1 U7888 ( .A(n6980), .B(n6979), .ZN(n6984) );
  XNOR2_X1 U7889 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput100), .ZN(n6983) );
  XNOR2_X1 U7890 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput64), .ZN(n6982)
         );
  XNOR2_X1 U7891 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput118), .ZN(
        n6981) );
  NAND4_X1 U7892 ( .A1(n6984), .A2(n6983), .A3(n6982), .A4(n6981), .ZN(n6985)
         );
  NOR3_X1 U7893 ( .A1(n6987), .A2(n6986), .A3(n6985), .ZN(n7000) );
  OAI22_X1 U7894 ( .A1(n6990), .A2(keyinput111), .B1(n6989), .B2(keyinput47), 
        .ZN(n6988) );
  AOI221_X1 U7895 ( .B1(n6990), .B2(keyinput111), .C1(keyinput47), .C2(n6989), 
        .A(n6988), .ZN(n6999) );
  INV_X1 U7896 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6993) );
  INV_X1 U7897 ( .A(keyinput8), .ZN(n6992) );
  OAI22_X1 U7898 ( .A1(n6993), .A2(keyinput7), .B1(n6992), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6991) );
  AOI221_X1 U7899 ( .B1(n6993), .B2(keyinput7), .C1(DATAO_REG_9__SCAN_IN), 
        .C2(n6992), .A(n6991), .ZN(n6998) );
  INV_X1 U7900 ( .A(keyinput57), .ZN(n6996) );
  INV_X1 U7901 ( .A(keyinput70), .ZN(n6995) );
  OAI22_X1 U7902 ( .A1(n6996), .A2(DATAO_REG_1__SCAN_IN), .B1(n6995), .B2(
        ADDRESS_REG_10__SCAN_IN), .ZN(n6994) );
  AOI221_X1 U7903 ( .B1(n6996), .B2(DATAO_REG_1__SCAN_IN), .C1(
        ADDRESS_REG_10__SCAN_IN), .C2(n6995), .A(n6994), .ZN(n6997) );
  AND4_X1 U7904 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), .ZN(n7001)
         );
  OAI211_X1 U7905 ( .C1(ADDRESS_REG_3__SCAN_IN), .C2(n7003), .A(n7002), .B(
        n7001), .ZN(n7004) );
  NOR4_X1 U7906 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n7008)
         );
  XNOR2_X1 U7907 ( .A(n7009), .B(n7008), .ZN(U2910) );
  NAND4_X1 U3642 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3340)
         );
  CLKBUF_X3 U3541 ( .A(n3445), .Z(n3113) );
  CLKBUF_X1 U3546 ( .A(n3490), .Z(n6668) );
  CLKBUF_X1 U3568 ( .A(n6665), .Z(n6681) );
  CLKBUF_X3 U3934 ( .A(n3340), .Z(n4490) );
  CLKBUF_X1 U3935 ( .A(n6192), .Z(n6680) );
endmodule

