

module b20_C_SARLock_k_64_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4287, n4288, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187;

  INV_X1 U4794 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n6609) );
  NAND2_X1 U4795 ( .A1(n9300), .A2(n8859), .ZN(n9295) );
  NAND2_X1 U4796 ( .A1(n5900), .A2(n5899), .ZN(n8508) );
  NAND2_X1 U4797 ( .A1(n4985), .A2(n4984), .ZN(n5091) );
  INV_X1 U4798 ( .A(n5155), .ZN(n5358) );
  CLKBUF_X1 U4799 ( .A(n5693), .Z(n5890) );
  INV_X1 U4800 ( .A(n5636), .ZN(n6501) );
  OR2_X1 U4801 ( .A1(n5774), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5787) );
  INV_X1 U4802 ( .A(n6609), .ZN(n4287) );
  INV_X1 U4803 ( .A(n4287), .ZN(n4288) );
  INV_X1 U4804 ( .A(n4287), .ZN(P1_U3086) );
  NOR2_X1 U4805 ( .A1(n8395), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U4806 ( .A1(n6126), .A2(n4290), .ZN(n6106) );
  AND2_X1 U4807 ( .A1(n8231), .A2(n8232), .ZN(n4734) );
  INV_X1 U4808 ( .A(n8772), .ZN(n5357) );
  OR2_X1 U4809 ( .A1(n5881), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5894) );
  BUF_X1 U4810 ( .A(n5658), .Z(n5858) );
  INV_X1 U4812 ( .A(n7328), .ZN(n7126) );
  CLKBUF_X2 U4814 ( .A(n5663), .Z(n6500) );
  XNOR2_X1 U4815 ( .A(n4499), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6795) );
  AND2_X1 U4816 ( .A1(n8747), .A2(n4359), .ZN(n6575) );
  NAND2_X1 U4817 ( .A1(n4421), .A2(n4323), .ZN(n8747) );
  NAND2_X1 U4818 ( .A1(n5278), .A2(n5277), .ZN(n7947) );
  XNOR2_X1 U4819 ( .A(n4912), .B(SI_1_), .ZN(n5138) );
  NAND2_X4 U4820 ( .A1(n6316), .A2(n6084), .ZN(n6126) );
  NAND2_X2 U4821 ( .A1(n6002), .A2(n6003), .ZN(n5694) );
  AOI21_X2 U4822 ( .B1(n9295), .B2(n9294), .A(n5523), .ZN(n9272) );
  NOR2_X2 U4823 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6760) );
  AOI21_X2 U4824 ( .B1(n8063), .B2(n8062), .A(n7997), .ZN(n8116) );
  NAND2_X2 U4825 ( .A1(n8146), .A2(n7995), .ZN(n8063) );
  OAI21_X2 U4826 ( .B1(n8766), .B2(n9039), .A(n5321), .ZN(n7891) );
  NAND2_X1 U4827 ( .A1(n6316), .A2(n6087), .ZN(n4290) );
  INV_X4 U4828 ( .A(n6108), .ZN(n6311) );
  OAI21_X2 U4829 ( .B1(n5091), .B2(n4989), .A(n4988), .ZN(n5353) );
  INV_X1 U4830 ( .A(n7213), .ZN(n6904) );
  OAI211_X2 U4831 ( .C1(n8772), .C2(n6684), .A(n5157), .B(n5156), .ZN(n7213)
         );
  XNOR2_X2 U4832 ( .A(n5607), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8607) );
  AND2_X4 U4833 ( .A1(n4715), .A2(n4714), .ZN(n4923) );
  NOR2_X2 U4834 ( .A1(n6465), .A2(n4386), .ZN(n6487) );
  INV_X1 U4835 ( .A(n4421), .ZN(n8744) );
  XNOR2_X1 U4836 ( .A(n6217), .B(n6215), .ZN(n8622) );
  OR2_X1 U4837 ( .A1(n10064), .A2(n8203), .ZN(n4743) );
  XNOR2_X1 U4838 ( .A(n6183), .B(n6181), .ZN(n7803) );
  NOR2_X1 U4840 ( .A1(n9960), .A2(n7866), .ZN(n9959) );
  NAND2_X1 U4841 ( .A1(n5233), .A2(n5232), .ZN(n7511) );
  INV_X2 U4842 ( .A(n6125), .ZN(n6219) );
  INV_X1 U4843 ( .A(n9025), .ZN(n4486) );
  INV_X1 U4844 ( .A(n8201), .ZN(n7974) );
  INV_X4 U4845 ( .A(n6161), .ZN(n4291) );
  INV_X1 U4846 ( .A(n9053), .ZN(n4562) );
  CLKBUF_X2 U4847 ( .A(n5634), .Z(n6483) );
  NAND2_X1 U4848 ( .A1(n5694), .A2(n6610), .ZN(n5693) );
  AND2_X1 U4849 ( .A1(n9183), .A2(n9905), .ZN(n4573) );
  OAI211_X1 U4850 ( .C1(n9187), .C2(n4488), .A(n4693), .B(n4692), .ZN(n9183)
         );
  NAND2_X1 U4851 ( .A1(n9187), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U4852 ( .A1(n5478), .A2(n5477), .ZN(n9187) );
  OR2_X1 U4853 ( .A1(n6575), .A2(n6317), .ZN(n6341) );
  OAI21_X1 U4854 ( .B1(n6009), .B2(n8440), .A(n6008), .ZN(n8287) );
  OAI21_X1 U4855 ( .B1(n4533), .B2(n4532), .A(n4335), .ZN(n4531) );
  NAND2_X1 U4856 ( .A1(n9185), .A2(n4574), .ZN(n5533) );
  NAND2_X1 U4857 ( .A1(n4708), .A2(n4300), .ZN(n9203) );
  AND2_X1 U4858 ( .A1(n9181), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U4859 ( .A1(n9010), .A2(n4308), .ZN(n4692) );
  NAND2_X1 U4860 ( .A1(n4838), .A2(n4837), .ZN(n8641) );
  NOR2_X1 U4861 ( .A1(n9010), .A2(n4308), .ZN(n4694) );
  NOR2_X1 U4862 ( .A1(n9743), .A2(n4756), .ZN(n4755) );
  OR2_X1 U4863 ( .A1(n6463), .A2(n8023), .ZN(n6588) );
  NAND2_X1 U4864 ( .A1(n5487), .A2(n5486), .ZN(n9178) );
  AOI21_X1 U4865 ( .B1(n4526), .B2(n6441), .A(n8340), .ZN(n6447) );
  NAND2_X1 U4866 ( .A1(n9400), .A2(n9474), .ZN(n4575) );
  OAI21_X1 U4867 ( .B1(n6184), .B2(n4823), .A(n6192), .ZN(n4821) );
  AND2_X1 U4868 ( .A1(n9299), .A2(n8855), .ZN(n9316) );
  NOR2_X1 U4869 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  OR2_X2 U4870 ( .A1(n8676), .A2(n7895), .ZN(n9372) );
  OR2_X1 U4871 ( .A1(n8394), .A2(n8404), .ZN(n6431) );
  NAND2_X1 U4872 ( .A1(n7459), .A2(n7458), .ZN(n7463) );
  NOR2_X1 U4873 ( .A1(n9959), .A2(n8235), .ZN(n9977) );
  AND2_X1 U4874 ( .A1(n6140), .A2(n4431), .ZN(n4430) );
  AND2_X1 U4875 ( .A1(n4729), .A2(n4725), .ZN(n8234) );
  OAI21_X1 U4876 ( .B1(n4859), .B2(n4858), .A(n4342), .ZN(n4857) );
  MUX2_X1 U4877 ( .A(n6349), .B(n6348), .S(n6605), .Z(n6378) );
  NAND2_X1 U4878 ( .A1(n5293), .A2(n5292), .ZN(n8716) );
  NAND2_X1 U4879 ( .A1(n5264), .A2(n5263), .ZN(n7877) );
  NAND2_X1 U4880 ( .A1(n5251), .A2(n5250), .ZN(n7557) );
  NAND2_X1 U4881 ( .A1(n5288), .A2(n4962), .ZN(n4965) );
  INV_X2 U4882 ( .A(n6946), .ZN(n8474) );
  NAND2_X1 U4883 ( .A1(n5229), .A2(n4896), .ZN(n4948) );
  AND2_X1 U4884 ( .A1(n6367), .A2(n6387), .ZN(n7480) );
  NAND2_X1 U4885 ( .A1(n4506), .A2(n4758), .ZN(n5112) );
  XNOR2_X1 U4886 ( .A(n4689), .B(n5212), .ZN(n6640) );
  INV_X2 U4887 ( .A(n6648), .ZN(n6715) );
  INV_X1 U4888 ( .A(n4419), .ZN(n4418) );
  OAI21_X1 U4889 ( .B1(n6821), .B2(n6820), .A(n6818), .ZN(n4419) );
  NAND4_X1 U4890 ( .A1(n5640), .A2(n5639), .A3(n5638), .A4(n5637), .ZN(n6978)
         );
  AND4_X1 U4891 ( .A1(n5176), .A2(n5175), .A3(n5174), .A4(n5173), .ZN(n7331)
         );
  INV_X1 U4892 ( .A(n7013), .ZN(n4292) );
  CLKBUF_X1 U4893 ( .A(n5624), .Z(n5995) );
  NAND2_X1 U4894 ( .A1(n6010), .A2(n7701), .ZN(n6819) );
  NAND4_X2 U4895 ( .A1(n5136), .A2(n5135), .A3(n5134), .A4(n5133), .ZN(n9053)
         );
  XNOR2_X1 U4896 ( .A(n4410), .B(n5599), .ZN(n6010) );
  INV_X2 U4897 ( .A(n5693), .ZN(n5674) );
  INV_X2 U4898 ( .A(n5182), .ZN(n8878) );
  NAND2_X1 U4899 ( .A1(n4411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4410) );
  INV_X2 U4900 ( .A(n6004), .ZN(n8227) );
  XNOR2_X1 U4901 ( .A(n6043), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U4902 ( .A1(n5141), .A2(n6610), .ZN(n5182) );
  NAND2_X1 U4903 ( .A1(n5560), .A2(n5501), .ZN(n7839) );
  NAND2_X1 U4904 ( .A1(n8604), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5605) );
  XNOR2_X1 U4905 ( .A(n5506), .B(n5505), .ZN(n7779) );
  NOR2_X1 U4906 ( .A1(n5541), .A2(n5534), .ZN(n5559) );
  NAND2_X1 U4907 ( .A1(n5504), .A2(n4313), .ZN(n9018) );
  OR2_X1 U4908 ( .A1(n6034), .A2(n5606), .ZN(n6042) );
  XNOR2_X1 U4909 ( .A(n5057), .B(n5056), .ZN(n9566) );
  NOR3_X1 U4910 ( .A1(n5809), .A2(n4396), .A3(P2_IR_REG_16__SCAN_IN), .ZN(
        n4395) );
  NAND2_X1 U4911 ( .A1(n5093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5339) );
  NAND2_X2 U4912 ( .A1(n5058), .A2(P2_U3151), .ZN(n8618) );
  NAND2_X1 U4913 ( .A1(n5075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5055) );
  OR2_X1 U4914 ( .A1(n5769), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5809) );
  AND2_X1 U4915 ( .A1(n5324), .A2(n5092), .ZN(n5498) );
  CLKBUF_X3 U4916 ( .A(n4923), .Z(n8770) );
  AND2_X1 U4917 ( .A1(n5052), .A2(n5046), .ZN(n4576) );
  NAND2_X1 U4918 ( .A1(n4907), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U4919 ( .A1(n4905), .A2(n7772), .ZN(n4715) );
  NOR2_X1 U4920 ( .A1(n4392), .A2(n4389), .ZN(n5766) );
  AND4_X1 U4921 ( .A1(n5598), .A2(n5865), .A3(n5849), .A4(n5864), .ZN(n4898)
         );
  NOR2_X1 U4922 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4393) );
  NOR2_X1 U4923 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4391) );
  NOR2_X1 U4924 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4390) );
  INV_X1 U4925 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5495) );
  NOR2_X1 U4926 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4579) );
  INV_X1 U4927 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5494) );
  INV_X1 U4928 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5496) );
  INV_X4 U4929 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4930 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5561) );
  NOR2_X1 U4931 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5598) );
  INV_X1 U4932 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5092) );
  INV_X1 U4933 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5865) );
  INV_X1 U4934 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5847) );
  NOR2_X2 U4935 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5177) );
  INV_X1 U4936 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5848) );
  INV_X1 U4937 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5849) );
  INV_X1 U4938 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7354) );
  AOI21_X2 U4939 ( .B1(n8126), .B2(n8122), .A(n8124), .ZN(n8049) );
  XNOR2_X2 U4940 ( .A(n8027), .B(n8298), .ZN(n8020) );
  NAND2_X4 U4941 ( .A1(n5983), .A2(n5982), .ZN(n8298) );
  XNOR2_X1 U4942 ( .A(n5229), .B(n4896), .ZN(n6704) );
  OAI21_X2 U4943 ( .B1(n5112), .B2(n5111), .A(n4941), .ZN(n5229) );
  OR2_X4 U4944 ( .A1(n7980), .A2(n8607), .ZN(n5646) );
  AND2_X4 U4945 ( .A1(n9559), .A2(n5079), .ZN(n5146) );
  NOR3_X4 U4946 ( .A1(n9372), .A2(n9321), .A3(n4450), .ZN(n9320) );
  NAND2_X1 U4947 ( .A1(n4353), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U4948 ( .A1(n4515), .A2(n8437), .ZN(n4514) );
  INV_X1 U4949 ( .A(n4517), .ZN(n4515) );
  INV_X1 U4950 ( .A(n4779), .ZN(n4778) );
  OAI21_X1 U4951 ( .B1(n4975), .B2(n4780), .A(n4974), .ZN(n4779) );
  NAND2_X1 U4952 ( .A1(n5302), .A2(n4971), .ZN(n4780) );
  INV_X1 U4953 ( .A(n7518), .ZN(n4862) );
  NAND2_X1 U4954 ( .A1(n8012), .A2(n8159), .ZN(n8164) );
  AND2_X1 U4956 ( .A1(n5974), .A2(n5973), .ZN(n8295) );
  INV_X1 U4957 ( .A(n8185), .ZN(n8310) );
  MUX2_X1 U4958 ( .A(n6380), .B(n6379), .S(n6593), .Z(n6384) );
  OR2_X1 U4959 ( .A1(n6374), .A2(n4534), .ZN(n6380) );
  NAND2_X1 U4960 ( .A1(n4480), .A2(n8834), .ZN(n4479) );
  AND2_X1 U4961 ( .A1(n4514), .A2(n4511), .ZN(n4510) );
  AND2_X1 U4962 ( .A1(n4512), .A2(n4355), .ZN(n4511) );
  NAND2_X1 U4963 ( .A1(n4516), .A2(n4509), .ZN(n6429) );
  AND2_X1 U4964 ( .A1(n4514), .A2(n4512), .ZN(n4509) );
  AOI211_X1 U4965 ( .C1(n6461), .C2(n6460), .A(n6459), .B(n6458), .ZN(n6465)
         );
  OAI211_X1 U4966 ( .C1(n6455), .C2(n8323), .A(n6454), .B(n6453), .ZN(n6460)
         );
  INV_X1 U4967 ( .A(SI_16_), .ZN(n4976) );
  INV_X1 U4968 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n4966) );
  INV_X1 U4969 ( .A(SI_11_), .ZN(n4955) );
  AOI21_X1 U4970 ( .B1(n4876), .B2(n4873), .A(n4368), .ZN(n4872) );
  OR2_X1 U4971 ( .A1(n4305), .A2(n4874), .ZN(n4873) );
  INV_X1 U4972 ( .A(n5658), .ZN(n5624) );
  NOR2_X1 U4973 ( .A1(n10043), .A2(n4744), .ZN(n8247) );
  NOR2_X1 U4974 ( .A1(n10033), .A2(n4745), .ZN(n4744) );
  INV_X1 U4975 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n4745) );
  NOR3_X1 U4976 ( .A1(n6539), .A2(n4640), .A3(n4644), .ZN(n4637) );
  AOI21_X1 U4977 ( .B1(n4644), .B2(n4642), .A(n4319), .ZN(n4641) );
  INV_X1 U4978 ( .A(n6451), .ZN(n4642) );
  OR2_X1 U4979 ( .A1(n8553), .A2(n8185), .ZN(n5974) );
  INV_X1 U4980 ( .A(n8567), .ZN(n5935) );
  OR2_X1 U4981 ( .A1(n5935), .A2(n8342), .ZN(n6513) );
  AND2_X1 U4982 ( .A1(n8571), .A2(n8188), .ZN(n6442) );
  OR2_X1 U4983 ( .A1(n5910), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5916) );
  OR2_X1 U4984 ( .A1(n8074), .A2(n8378), .ZN(n6436) );
  OR2_X1 U4985 ( .A1(n8168), .A2(n8430), .ZN(n6417) );
  NOR2_X1 U4986 ( .A1(n10081), .A2(n7482), .ZN(n4631) );
  NAND2_X1 U4987 ( .A1(n4630), .A2(n7477), .ZN(n4629) );
  AND2_X1 U4988 ( .A1(n5684), .A2(n4632), .ZN(n4630) );
  NAND2_X1 U4989 ( .A1(n10081), .A2(n7482), .ZN(n4632) );
  NAND2_X1 U4990 ( .A1(n7678), .A2(n4322), .ZN(n4590) );
  OAI21_X1 U4991 ( .B1(n4598), .B2(n4596), .A(n6516), .ZN(n4595) );
  INV_X1 U4992 ( .A(n7782), .ZN(n7246) );
  NOR2_X1 U4993 ( .A1(n4329), .A2(n4881), .ZN(n4880) );
  INV_X1 U4994 ( .A(n5769), .ZN(n4675) );
  INV_X1 U4995 ( .A(n4677), .ZN(n4676) );
  INV_X1 U4996 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6038) );
  AOI21_X1 U4997 ( .B1(n4832), .B2(n4835), .A(n4315), .ZN(n4443) );
  INV_X1 U4998 ( .A(n4812), .ZN(n4809) );
  AOI21_X1 U4999 ( .B1(n4815), .B2(n4814), .A(n4813), .ZN(n4812) );
  INV_X1 U5000 ( .A(n8691), .ZN(n4813) );
  INV_X1 U5001 ( .A(n4817), .ZN(n4814) );
  OAI21_X1 U5002 ( .B1(n6141), .B2(n4831), .A(n4428), .ZN(n6166) );
  INV_X1 U5003 ( .A(n4429), .ZN(n4428) );
  OAI21_X1 U5004 ( .B1(n4430), .B2(n4831), .A(n7543), .ZN(n4429) );
  NOR2_X1 U5005 ( .A1(n6260), .A2(n4839), .ZN(n4836) );
  AND2_X1 U5006 ( .A1(n6085), .A2(n6083), .ZN(n6084) );
  OR2_X1 U5007 ( .A1(n5453), .A2(n6577), .ZN(n5470) );
  OR2_X1 U5008 ( .A1(n9347), .A2(n9379), .ZN(n4451) );
  INV_X1 U5009 ( .A(n4552), .ZN(n4551) );
  NAND2_X1 U5010 ( .A1(n9286), .A2(n9449), .ZN(n4707) );
  OR2_X1 U5011 ( .A1(n8676), .A2(n8763), .ZN(n8831) );
  NAND2_X1 U5012 ( .A1(n6473), .A2(n6472), .ZN(n6494) );
  OR2_X1 U5013 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  OR2_X1 U5014 ( .A1(n6469), .A2(n6468), .ZN(n6473) );
  AOI21_X1 U5015 ( .B1(n4805), .B2(n4802), .A(n4801), .ZN(n4800) );
  INV_X1 U5016 ( .A(n4805), .ZN(n4803) );
  INV_X1 U5017 ( .A(n4999), .ZN(n4801) );
  AOI21_X1 U5018 ( .B1(n4771), .B2(n4775), .A(n4770), .ZN(n4769) );
  NOR2_X1 U5019 ( .A1(n4975), .A2(n4782), .ZN(n4781) );
  INV_X1 U5020 ( .A(n4971), .ZN(n4782) );
  INV_X1 U5021 ( .A(n4786), .ZN(n4785) );
  OAI21_X1 U5022 ( .B1(n4789), .B2(n4296), .A(n4959), .ZN(n4786) );
  NOR2_X1 U5023 ( .A1(n8003), .A2(n8002), .ZN(n4413) );
  NAND2_X1 U5024 ( .A1(n8005), .A2(n8342), .ZN(n8079) );
  AND2_X1 U5025 ( .A1(n8160), .A2(n8010), .ZN(n8080) );
  INV_X1 U5026 ( .A(n7148), .ZN(n4851) );
  NAND2_X1 U5027 ( .A1(n8008), .A2(n8329), .ZN(n8160) );
  AND4_X1 U5028 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n7661)
         );
  OR2_X1 U5029 ( .A1(n5634), .A2(n6748), .ZN(n5647) );
  INV_X1 U5030 ( .A(n5636), .ZN(n5657) );
  XNOR2_X1 U5031 ( .A(n8247), .B(n10051), .ZN(n10064) );
  OR2_X1 U5032 ( .A1(n8077), .A2(n8329), .ZN(n6452) );
  INV_X1 U5033 ( .A(n8186), .ZN(n8329) );
  AOI21_X1 U5034 ( .B1(n4614), .B2(n4294), .A(n4352), .ZN(n4613) );
  OR2_X1 U5035 ( .A1(n8089), .A2(n8441), .ZN(n6420) );
  OR2_X1 U5036 ( .A1(n8461), .A2(n8443), .ZN(n6412) );
  INV_X1 U5037 ( .A(n8460), .ZN(n8440) );
  NAND2_X1 U5038 ( .A1(n6015), .A2(n7967), .ZN(n6975) );
  NAND2_X1 U5039 ( .A1(n8036), .A2(n6599), .ZN(n6600) );
  AND2_X1 U5040 ( .A1(n7843), .A2(n7782), .ZN(n10095) );
  NAND2_X1 U5041 ( .A1(n5766), .A2(n5767), .ZN(n5769) );
  NOR2_X1 U5042 ( .A1(n8884), .A2(n9016), .ZN(n4766) );
  AOI21_X1 U5043 ( .B1(n8883), .B2(n9170), .A(n4490), .ZN(n8884) );
  NAND2_X1 U5044 ( .A1(n9160), .A2(n4491), .ZN(n4490) );
  INV_X1 U5045 ( .A(n4492), .ZN(n4491) );
  AND2_X1 U5046 ( .A1(n9160), .A2(n9163), .ZN(n9016) );
  NAND2_X1 U5047 ( .A1(n9238), .A2(n4452), .ZN(n9169) );
  NOR2_X1 U5048 ( .A1(n9178), .A2(n4453), .ZN(n4452) );
  INV_X1 U5049 ( .A(n4454), .ZN(n4453) );
  NAND2_X1 U5050 ( .A1(n5060), .A2(n5059), .ZN(n9208) );
  AND2_X1 U5051 ( .A1(n5442), .A2(n5441), .ZN(n9263) );
  OR2_X1 U5052 ( .A1(n9241), .A2(n5488), .ZN(n5442) );
  OAI21_X1 U5053 ( .B1(n4701), .B2(n4698), .A(n4695), .ZN(n9251) );
  NAND2_X1 U5054 ( .A1(n4699), .A2(n4895), .ZN(n4698) );
  INV_X1 U5055 ( .A(n4696), .ZN(n4695) );
  INV_X1 U5056 ( .A(n4703), .ZN(n4699) );
  OR2_X1 U5057 ( .A1(n7557), .A2(n9044), .ZN(n5259) );
  NAND2_X1 U5058 ( .A1(n8776), .A2(n8983), .ZN(n4554) );
  AND2_X1 U5059 ( .A1(n8676), .A2(n9368), .ZN(n5336) );
  OAI21_X1 U5060 ( .B1(n9551), .B2(P1_D_REG_0__SCAN_IN), .A(n9553), .ZN(n7132)
         );
  NAND2_X1 U5061 ( .A1(n5525), .A2(n8885), .ZN(n9482) );
  AND2_X1 U5062 ( .A1(n5015), .A2(n5014), .ZN(n5406) );
  NAND2_X1 U5063 ( .A1(n4768), .A2(n4771), .ZN(n5338) );
  OR2_X1 U5064 ( .A1(n5303), .A2(n4775), .ZN(n4768) );
  OR2_X1 U5065 ( .A1(n8018), .A2(n8310), .ZN(n8019) );
  INV_X1 U5066 ( .A(n8559), .ZN(n8167) );
  NAND2_X1 U5067 ( .A1(n6598), .A2(n8460), .ZN(n4669) );
  AOI21_X1 U5068 ( .B1(n4620), .B2(n4618), .A(n4350), .ZN(n6589) );
  AND2_X1 U5069 ( .A1(n4316), .A2(n6585), .ZN(n4618) );
  NAND2_X1 U5070 ( .A1(n4471), .A2(n4470), .ZN(n8787) );
  NAND2_X1 U5071 ( .A1(n8916), .A2(n4486), .ZN(n4471) );
  NAND2_X1 U5072 ( .A1(n4472), .A2(n9025), .ZN(n4470) );
  NOR2_X1 U5073 ( .A1(n6384), .A2(n4523), .ZN(n4522) );
  AND2_X1 U5074 ( .A1(n6394), .A2(n6381), .ZN(n4523) );
  OR2_X1 U5075 ( .A1(n6383), .A2(n6593), .ZN(n4521) );
  NAND2_X1 U5076 ( .A1(n4482), .A2(n4481), .ZN(n4480) );
  NAND2_X1 U5077 ( .A1(n8822), .A2(n4486), .ZN(n4481) );
  NAND2_X1 U5078 ( .A1(n8821), .A2(n9025), .ZN(n4482) );
  NAND2_X1 U5079 ( .A1(n4508), .A2(n4507), .ZN(n6423) );
  NOR2_X1 U5080 ( .A1(n4530), .A2(n6605), .ZN(n4529) );
  NAND2_X1 U5081 ( .A1(n6437), .A2(n4326), .ZN(n4527) );
  INV_X1 U5082 ( .A(n4460), .ZN(n4459) );
  AOI21_X1 U5083 ( .B1(n8844), .B2(n9025), .A(n4461), .ZN(n4460) );
  AND2_X1 U5084 ( .A1(n8843), .A2(n4486), .ZN(n4461) );
  INV_X1 U5085 ( .A(n7968), .ZN(n4658) );
  NAND2_X1 U5086 ( .A1(n8948), .A2(n8894), .ZN(n8867) );
  AND2_X1 U5087 ( .A1(n6462), .A2(n6464), .ZN(n4386) );
  NAND2_X1 U5088 ( .A1(n10100), .A2(n8196), .ZN(n4535) );
  NOR2_X1 U5089 ( .A1(n4631), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U5090 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4634) );
  NAND2_X1 U5091 ( .A1(n4597), .A2(n4602), .ZN(n4596) );
  INV_X1 U5092 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5616) );
  OR2_X1 U5093 ( .A1(n9170), .A2(n8957), .ZN(n8977) );
  NAND2_X1 U5094 ( .A1(n8876), .A2(n8877), .ZN(n4493) );
  NOR2_X1 U5095 ( .A1(n4332), .A2(n4383), .ZN(n4382) );
  INV_X1 U5096 ( .A(n4469), .ZN(n4383) );
  NAND2_X1 U5097 ( .A1(n4493), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U5098 ( .A1(n4493), .A2(n9025), .ZN(n4489) );
  OR2_X1 U5099 ( .A1(n7779), .A2(n9014), .ZN(n6083) );
  OR2_X1 U5100 ( .A1(n9230), .A2(n9244), .ZN(n8948) );
  NAND2_X1 U5101 ( .A1(n5484), .A2(n5483), .ZN(n6471) );
  NAND2_X1 U5102 ( .A1(n4928), .A2(n4927), .ZN(n4505) );
  INV_X1 U5103 ( .A(n7789), .ZN(n4858) );
  NAND2_X1 U5104 ( .A1(n4405), .A2(n4407), .ZN(n4403) );
  INV_X1 U5105 ( .A(n7236), .ZN(n8004) );
  NAND2_X1 U5106 ( .A1(n5588), .A2(n5587), .ZN(n5856) );
  INV_X1 U5107 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5587) );
  INV_X1 U5108 ( .A(n5841), .ZN(n5588) );
  INV_X1 U5109 ( .A(n9944), .ZN(n4733) );
  NAND2_X1 U5110 ( .A1(n9934), .A2(n8259), .ZN(n8260) );
  NAND2_X1 U5111 ( .A1(n9975), .A2(n8240), .ZN(n8242) );
  NAND2_X1 U5112 ( .A1(n4741), .A2(n4740), .ZN(n4384) );
  NAND2_X1 U5113 ( .A1(n8253), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4740) );
  INV_X1 U5114 ( .A(n10010), .ZN(n4741) );
  NAND2_X1 U5115 ( .A1(n10002), .A2(n4494), .ZN(n8268) );
  OR2_X1 U5116 ( .A1(n10001), .A2(n9680), .ZN(n4494) );
  NAND2_X1 U5117 ( .A1(n8167), .A2(n8299), .ZN(n4619) );
  AOI21_X1 U5118 ( .B1(n4610), .B2(n4608), .A(n8363), .ZN(n4607) );
  INV_X1 U5119 ( .A(n4614), .ZN(n4608) );
  INV_X1 U5120 ( .A(n4610), .ZN(n4609) );
  NOR2_X1 U5121 ( .A1(n4294), .A2(n5887), .ZN(n4615) );
  AND2_X1 U5122 ( .A1(n4611), .A2(n4613), .ZN(n4610) );
  OR2_X1 U5123 ( .A1(n8508), .A2(n8387), .ZN(n6430) );
  OR2_X1 U5124 ( .A1(n8145), .A2(n8386), .ZN(n6515) );
  NOR2_X1 U5125 ( .A1(n4585), .A2(n4582), .ZN(n4581) );
  INV_X1 U5126 ( .A(n4589), .ZN(n4582) );
  INV_X1 U5127 ( .A(n4654), .ZN(n4653) );
  OAI21_X1 U5128 ( .B1(n6023), .B2(n4655), .A(n6416), .ZN(n4654) );
  INV_X1 U5129 ( .A(n6412), .ZN(n4655) );
  NAND2_X1 U5130 ( .A1(n4587), .A2(n4312), .ZN(n4586) );
  NAND2_X1 U5131 ( .A1(n4603), .A2(n7983), .ZN(n4602) );
  NOR2_X1 U5132 ( .A1(n5797), .A2(n4601), .ZN(n4600) );
  INV_X1 U5133 ( .A(n5765), .ZN(n4601) );
  AND2_X1 U5134 ( .A1(n6401), .A2(n6020), .ZN(n7846) );
  OR2_X1 U5135 ( .A1(n6483), .A2(n5685), .ZN(n5692) );
  NAND2_X1 U5136 ( .A1(n7430), .A2(n7974), .ZN(n6390) );
  INV_X1 U5137 ( .A(n6975), .ZN(n6352) );
  OR2_X1 U5138 ( .A1(n6622), .A2(n6065), .ZN(n6830) );
  NOR2_X1 U5139 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4849) );
  NAND2_X1 U5140 ( .A1(n4424), .A2(n4423), .ZN(n6183) );
  AOI21_X1 U5141 ( .B1(n4422), .B2(n7650), .A(n4331), .ZN(n4423) );
  NOR2_X1 U5142 ( .A1(n8681), .A2(n4842), .ZN(n4841) );
  INV_X1 U5143 ( .A(n6234), .ZN(n4842) );
  OAI22_X1 U5144 ( .A1(n8830), .A2(n6125), .B1(n8673), .B2(n6161), .ZN(n6226)
         );
  OAI21_X1 U5145 ( .B1(n9170), .B2(n4486), .A(n9038), .ZN(n4492) );
  OR2_X1 U5146 ( .A1(n9280), .A2(n9291), .ZN(n8861) );
  NOR2_X1 U5147 ( .A1(n4542), .A2(n4538), .ZN(n4537) );
  INV_X1 U5148 ( .A(n4546), .ZN(n4538) );
  INV_X1 U5149 ( .A(n9316), .ZN(n4542) );
  NAND2_X1 U5150 ( .A1(n4541), .A2(n9316), .ZN(n4540) );
  INV_X1 U5151 ( .A(n4543), .ZN(n4541) );
  OR2_X1 U5152 ( .A1(n5329), .A2(n8671), .ZN(n5343) );
  NAND2_X1 U5153 ( .A1(n4683), .A2(n4685), .ZN(n4682) );
  OR2_X1 U5154 ( .A1(n7708), .A2(n8714), .ZN(n8835) );
  AND2_X1 U5155 ( .A1(n4566), .A2(n8929), .ZN(n4565) );
  INV_X1 U5156 ( .A(n9000), .ZN(n4566) );
  OR2_X1 U5157 ( .A1(n5280), .A2(n5279), .ZN(n5295) );
  OR2_X1 U5158 ( .A1(n5253), .A2(n5252), .ZN(n5266) );
  OR2_X1 U5159 ( .A1(n7511), .A2(n7547), .ZN(n8810) );
  NAND2_X1 U5160 ( .A1(n7392), .A2(n7394), .ZN(n5227) );
  OR2_X1 U5161 ( .A1(n7192), .A2(n8987), .ZN(n7384) );
  OR2_X1 U5162 ( .A1(n7562), .A2(n7619), .ZN(n8794) );
  OAI21_X1 U5163 ( .B1(n4551), .B2(n8983), .A(n8914), .ZN(n4549) );
  NAND2_X1 U5164 ( .A1(n8886), .A2(n8887), .ZN(n6085) );
  XNOR2_X1 U5165 ( .A(n8909), .B(n4562), .ZN(n8981) );
  AND2_X1 U5166 ( .A1(n4561), .A2(n6810), .ZN(n6955) );
  AND2_X1 U5167 ( .A1(n8887), .A2(n9018), .ZN(n6086) );
  OR2_X1 U5168 ( .A1(n9208), .A2(n9228), .ZN(n8965) );
  OR2_X1 U5169 ( .A1(n9246), .A2(n9263), .ZN(n8894) );
  NAND2_X1 U5170 ( .A1(n5160), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U5171 ( .A1(n5053), .A2(n4847), .ZN(n4846) );
  INV_X1 U5172 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4847) );
  INV_X1 U5173 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5174 ( .A1(n4793), .A2(n4791), .ZN(n5419) );
  AOI21_X1 U5175 ( .B1(n4795), .B2(n4797), .A(n4792), .ZN(n4791) );
  INV_X1 U5176 ( .A(n5015), .ZN(n4792) );
  AND2_X1 U5177 ( .A1(n5498), .A2(n4432), .ZN(n5539) );
  AND2_X1 U5178 ( .A1(n5497), .A2(n4433), .ZN(n4432) );
  NOR2_X1 U5179 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4433) );
  AOI21_X1 U5180 ( .B1(n4774), .B2(n4773), .A(n4772), .ZN(n4771) );
  INV_X1 U5181 ( .A(n4980), .ZN(n4772) );
  INV_X1 U5182 ( .A(n4781), .ZN(n4773) );
  NAND2_X1 U5183 ( .A1(n4968), .A2(n4967), .ZN(n4971) );
  AOI21_X1 U5184 ( .B1(n4785), .B2(n4299), .A(n4349), .ZN(n4784) );
  INV_X1 U5185 ( .A(n4952), .ZN(n4787) );
  NOR2_X1 U5186 ( .A1(n4953), .A2(n4790), .ZN(n4789) );
  INV_X1 U5187 ( .A(n4947), .ZN(n4790) );
  AOI21_X1 U5188 ( .B1(n4759), .B2(n4761), .A(n4345), .ZN(n4758) );
  NAND2_X1 U5189 ( .A1(n5200), .A2(n4759), .ZN(n4506) );
  AND2_X1 U5190 ( .A1(n5199), .A2(n4934), .ZN(n4687) );
  XNOR2_X1 U5191 ( .A(n4915), .B(SI_2_), .ZN(n5153) );
  NAND2_X1 U5192 ( .A1(n8105), .A2(n4413), .ZN(n4853) );
  INV_X1 U5193 ( .A(n8106), .ZN(n4854) );
  AOI21_X1 U5194 ( .B1(n7464), .B2(n4861), .A(n4347), .ZN(n4859) );
  INV_X1 U5195 ( .A(n7463), .ZN(n7461) );
  NAND2_X1 U5196 ( .A1(n4865), .A2(n4863), .ZN(n8146) );
  AOI21_X1 U5197 ( .B1(n4866), .B2(n4869), .A(n4864), .ZN(n4863) );
  NAND2_X1 U5198 ( .A1(n4404), .A2(n4320), .ZN(n4865) );
  INV_X1 U5199 ( .A(n8147), .ZN(n4864) );
  OR2_X1 U5200 ( .A1(n5634), .A2(n5625), .ZN(n5626) );
  NAND2_X1 U5201 ( .A1(n6067), .A2(n7959), .ZN(n6836) );
  AND2_X1 U5202 ( .A1(n8616), .A2(n6623), .ZN(n6067) );
  NAND2_X1 U5203 ( .A1(n6758), .A2(n6759), .ZN(n6922) );
  OR2_X1 U5204 ( .A1(n6927), .A2(n7375), .ZN(n7076) );
  OAI211_X1 U5205 ( .C1(n8233), .C2(n4734), .A(n4732), .B(n4733), .ZN(n4736)
         );
  OR2_X1 U5206 ( .A1(n4734), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U5207 ( .A1(n8233), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4731) );
  XNOR2_X1 U5208 ( .A(n8260), .B(n9950), .ZN(n9952) );
  NAND2_X1 U5209 ( .A1(n9952), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9951) );
  OR2_X1 U5210 ( .A1(n9977), .A2(n9978), .ZN(n9975) );
  OR2_X1 U5211 ( .A1(n9992), .A2(n8243), .ZN(n4737) );
  XNOR2_X1 U5212 ( .A(n8242), .B(n8266), .ZN(n9992) );
  NOR2_X1 U5213 ( .A1(n5809), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U5214 ( .A1(n10003), .A2(n10004), .ZN(n10002) );
  XNOR2_X1 U5215 ( .A(n8268), .B(n10018), .ZN(n10020) );
  XNOR2_X1 U5216 ( .A(n4384), .B(n8269), .ZN(n10027) );
  NOR2_X1 U5217 ( .A1(n10027), .A2(n5840), .ZN(n10026) );
  AND2_X1 U5218 ( .A1(n4743), .A2(n4742), .ZN(n9745) );
  NAND2_X1 U5219 ( .A1(n8248), .A2(n8272), .ZN(n4742) );
  NOR2_X1 U5220 ( .A1(n9745), .A2(n9744), .ZN(n9743) );
  OAI21_X1 U5221 ( .B1(n8279), .B2(n9739), .A(n4377), .ZN(n4753) );
  NAND2_X1 U5222 ( .A1(n4638), .A2(n4636), .ZN(n6592) );
  NOR2_X1 U5223 ( .A1(n4637), .A2(n4340), .ZN(n4636) );
  NOR2_X1 U5224 ( .A1(n6539), .A2(n4640), .ZN(n4639) );
  AND2_X1 U5225 ( .A1(n6588), .A2(n6587), .ZN(n6590) );
  NAND2_X1 U5226 ( .A1(n8298), .A2(n8455), .ZN(n8301) );
  OR2_X1 U5227 ( .A1(n6450), .A2(n4319), .ZN(n8311) );
  NOR2_X1 U5228 ( .A1(n5935), .A2(n8187), .ZN(n5936) );
  OR2_X1 U5229 ( .A1(n6442), .A2(n6440), .ZN(n8340) );
  AOI21_X1 U5230 ( .B1(n8355), .B2(n5995), .A(n5612), .ZN(n8367) );
  AOI21_X1 U5231 ( .B1(n8368), .B2(n5995), .A(n5913), .ZN(n8378) );
  NAND2_X1 U5232 ( .A1(n8401), .A2(n4614), .ZN(n4612) );
  AND2_X1 U5233 ( .A1(n4612), .A2(n4610), .ZN(n8374) );
  AND2_X1 U5234 ( .A1(n6515), .A2(n6514), .ZN(n8402) );
  NOR2_X1 U5235 ( .A1(n8411), .A2(n4661), .ZN(n4660) );
  INV_X1 U5236 ( .A(n6420), .ZN(n4661) );
  NAND2_X1 U5237 ( .A1(n4588), .A2(n4586), .ZN(n8426) );
  NAND2_X1 U5238 ( .A1(n5833), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U5239 ( .A1(n5584), .A2(n5583), .ZN(n5814) );
  INV_X1 U5240 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5583) );
  INV_X1 U5241 ( .A(n5802), .ZN(n5584) );
  AND2_X1 U5242 ( .A1(n4361), .A2(n5796), .ZN(n4598) );
  INV_X1 U5243 ( .A(n4602), .ZN(n4593) );
  NAND2_X1 U5244 ( .A1(n5582), .A2(n7316), .ZN(n5774) );
  INV_X1 U5245 ( .A(n5757), .ZN(n5582) );
  AND2_X1 U5246 ( .A1(n6371), .A2(n6372), .ZN(n4649) );
  NAND2_X1 U5247 ( .A1(n4648), .A2(n4647), .ZN(n7682) );
  AND2_X1 U5248 ( .A1(n7683), .A2(n6375), .ZN(n4647) );
  AOI21_X1 U5249 ( .B1(n7373), .B2(n6392), .A(n4665), .ZN(n4663) );
  INV_X1 U5250 ( .A(n6393), .ZN(n4665) );
  OR2_X1 U5251 ( .A1(n8200), .A2(n10081), .ZN(n7406) );
  INV_X1 U5252 ( .A(n4631), .ZN(n4626) );
  INV_X1 U5253 ( .A(n8457), .ZN(n8444) );
  AND2_X1 U5254 ( .A1(n6567), .A2(n6012), .ZN(n7721) );
  INV_X1 U5255 ( .A(n8455), .ZN(n8442) );
  AND2_X1 U5256 ( .A1(n6052), .A2(n6605), .ZN(n6940) );
  AOI21_X1 U5257 ( .B1(n6047), .B2(n6628), .A(n6046), .ZN(n6943) );
  NAND2_X1 U5258 ( .A1(n6344), .A2(n6343), .ZN(n6463) );
  NAND2_X1 U5259 ( .A1(n5939), .A2(n5938), .ZN(n8077) );
  NAND2_X1 U5260 ( .A1(n5855), .A2(n5854), .ZN(n8089) );
  NAND2_X1 U5261 ( .A1(n5839), .A2(n5838), .ZN(n8168) );
  NAND2_X1 U5262 ( .A1(n6074), .A2(n5994), .ZN(n8460) );
  AND2_X1 U5263 ( .A1(n4880), .A2(n4674), .ZN(n4673) );
  INV_X1 U5264 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4674) );
  XNOR2_X1 U5265 ( .A(n6069), .B(n4883), .ZN(n6743) );
  INV_X1 U5266 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5986) );
  INV_X1 U5267 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5989) );
  INV_X1 U5268 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5888) );
  INV_X1 U5269 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5597) );
  INV_X1 U5270 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5767) );
  OR2_X1 U5271 ( .A1(n5724), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5751) );
  OR2_X1 U5272 ( .A1(n5714), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U5273 ( .A1(n5559), .A2(n5558), .ZN(n6316) );
  NAND2_X1 U5274 ( .A1(n8622), .A2(n8623), .ZN(n8621) );
  AOI21_X1 U5275 ( .B1(n4443), .B2(n4440), .A(n4344), .ZN(n4439) );
  INV_X1 U5276 ( .A(n4832), .ZN(n4440) );
  INV_X1 U5277 ( .A(n7872), .ZN(n4823) );
  NOR2_X1 U5278 ( .A1(n4823), .A2(n4824), .ZN(n4822) );
  INV_X1 U5279 ( .A(n7804), .ZN(n4824) );
  INV_X2 U5280 ( .A(n6126), .ZN(n6295) );
  OR2_X1 U5281 ( .A1(n5410), .A2(n9682), .ZN(n5423) );
  OR2_X1 U5282 ( .A1(n5423), .A2(n5422), .ZN(n5436) );
  NAND2_X1 U5283 ( .A1(n4815), .A2(n4818), .ZN(n4810) );
  NAND2_X1 U5284 ( .A1(n4809), .A2(n4818), .ZN(n4808) );
  INV_X1 U5285 ( .A(n8690), .ZN(n4818) );
  OR2_X1 U5286 ( .A1(n7021), .A2(n4826), .ZN(n4825) );
  INV_X1 U5287 ( .A(n6124), .ZN(n4826) );
  OR2_X1 U5288 ( .A1(n5373), .A2(n8704), .ZN(n5386) );
  NAND2_X1 U5289 ( .A1(n6141), .A2(n4430), .ZN(n7293) );
  INV_X1 U5290 ( .A(n7839), .ZN(n8886) );
  AND2_X1 U5291 ( .A1(n5470), .A2(n5074), .ZN(n9209) );
  OAI21_X1 U5292 ( .B1(n9259), .B2(n4569), .A(n4568), .ZN(n9221) );
  NAND2_X1 U5293 ( .A1(n8901), .A2(n9250), .ZN(n4569) );
  NAND2_X1 U5294 ( .A1(n4570), .A2(n8901), .ZN(n4568) );
  OR2_X1 U5295 ( .A1(n9321), .A2(n9336), .ZN(n9299) );
  AND2_X1 U5296 ( .A1(n9366), .A2(n8841), .ZN(n9345) );
  NAND2_X1 U5297 ( .A1(n7627), .A2(n5520), .ZN(n4567) );
  NAND2_X1 U5298 ( .A1(n4567), .A2(n4565), .ZN(n7815) );
  OR2_X1 U5299 ( .A1(n7947), .A2(n9042), .ZN(n5286) );
  INV_X1 U5300 ( .A(n5286), .ZN(n4685) );
  INV_X1 U5301 ( .A(n4684), .ZN(n4683) );
  OAI21_X1 U5302 ( .B1(n7602), .B2(n4685), .A(n8998), .ZN(n4684) );
  NAND2_X1 U5303 ( .A1(n7603), .A2(n7602), .ZN(n7601) );
  NAND2_X1 U5304 ( .A1(n7487), .A2(n8996), .ZN(n7486) );
  NOR3_X1 U5305 ( .A1(n7557), .A2(n7506), .A3(n7511), .ZN(n7493) );
  OR2_X1 U5306 ( .A1(n7511), .A2(n9045), .ZN(n5241) );
  OR2_X1 U5307 ( .A1(n5219), .A2(n5120), .ZN(n5235) );
  AND4_X1 U5308 ( .A1(n5211), .A2(n5210), .A3(n5209), .A4(n5208), .ZN(n7442)
         );
  NAND2_X1 U5309 ( .A1(n7276), .A2(n5198), .ZN(n7195) );
  NOR2_X1 U5310 ( .A1(n5513), .A2(n4553), .ZN(n4552) );
  NAND2_X1 U5311 ( .A1(n5512), .A2(n5511), .ZN(n8776) );
  AND4_X1 U5312 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n6907)
         );
  INV_X1 U5313 ( .A(n8981), .ZN(n6884) );
  NAND2_X1 U5314 ( .A1(n8909), .A2(n4444), .ZN(n6901) );
  OR2_X1 U5315 ( .A1(n6958), .A2(n9014), .ZN(n9371) );
  AND2_X1 U5316 ( .A1(n5080), .A2(n9563), .ZN(n5220) );
  NAND2_X1 U5317 ( .A1(n5160), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5133) );
  AOI21_X1 U5318 ( .B1(n4295), .B2(n5444), .A(n4339), .ZN(n4709) );
  NAND2_X1 U5319 ( .A1(n9234), .A2(n4295), .ZN(n4708) );
  AND2_X1 U5320 ( .A1(n5435), .A2(n5434), .ZN(n9420) );
  AND2_X1 U5321 ( .A1(n5409), .A2(n5408), .ZN(n9435) );
  OR2_X1 U5322 ( .A1(n4702), .A2(n4705), .ZN(n4700) );
  AND2_X1 U5323 ( .A1(n5405), .A2(n4706), .ZN(n4705) );
  INV_X1 U5324 ( .A(n4707), .ZN(n4702) );
  NAND2_X1 U5325 ( .A1(n4707), .A2(n5393), .ZN(n4703) );
  AND2_X1 U5326 ( .A1(n8775), .A2(n8774), .ZN(n9294) );
  NAND2_X1 U5327 ( .A1(n9452), .A2(n8728), .ZN(n4706) );
  NOR2_X1 U5328 ( .A1(n9338), .A2(n9476), .ZN(n5366) );
  AND2_X1 U5329 ( .A1(n8848), .A2(n8846), .ZN(n9344) );
  NAND2_X1 U5330 ( .A1(n4720), .A2(n4723), .ZN(n4719) );
  INV_X1 U5331 ( .A(n9004), .ZN(n4720) );
  NAND2_X1 U5332 ( .A1(n4721), .A2(n4723), .ZN(n4718) );
  NAND2_X1 U5333 ( .A1(n4722), .A2(n5350), .ZN(n4721) );
  INV_X1 U5334 ( .A(n5336), .ZN(n4722) );
  AND2_X1 U5335 ( .A1(n8841), .A2(n8845), .ZN(n9363) );
  AND2_X1 U5336 ( .A1(n8831), .A2(n9361), .ZN(n9004) );
  NOR2_X1 U5337 ( .A1(n7891), .A2(n9004), .ZN(n7890) );
  AND4_X1 U5338 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n7807)
         );
  AND2_X1 U5339 ( .A1(n9025), .A2(n9018), .ZN(n9895) );
  NAND2_X1 U5340 ( .A1(n5545), .A2(n9569), .ZN(n9551) );
  XNOR2_X1 U5341 ( .A(n6499), .B(n6498), .ZN(n8771) );
  OAI21_X1 U5342 ( .B1(n6494), .B2(n6493), .A(n6492), .ZN(n6499) );
  XNOR2_X1 U5343 ( .A(n5077), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5344 ( .A1(n9555), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U5345 ( .A(n6494), .B(n6493), .ZN(n8879) );
  XNOR2_X1 U5346 ( .A(n5078), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U5347 ( .A1(n4354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U5348 ( .A(n5039), .B(n5038), .ZN(n8612) );
  NAND2_X1 U5349 ( .A1(n5534), .A2(n5053), .ZN(n5543) );
  XNOR2_X1 U5350 ( .A(n5419), .B(n5418), .ZN(n7953) );
  NOR2_X1 U5351 ( .A1(n5394), .A2(n4799), .ZN(n4798) );
  INV_X1 U5352 ( .A(n5003), .ZN(n4799) );
  XNOR2_X1 U5353 ( .A(n5562), .B(n5561), .ZN(n6632) );
  OR2_X1 U5354 ( .A1(n5539), .A2(n9554), .ZN(n5500) );
  INV_X1 U5355 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U5356 ( .A1(n5500), .A2(n5499), .ZN(n5560) );
  NOR2_X1 U5357 ( .A1(n7074), .A2(n7075), .ZN(n4749) );
  OR2_X1 U5358 ( .A1(n6927), .A2(n4750), .ZN(n4747) );
  NAND2_X1 U5359 ( .A1(n4752), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4750) );
  NAND2_X1 U5360 ( .A1(n5824), .A2(n5823), .ZN(n8461) );
  NAND2_X1 U5361 ( .A1(n5976), .A2(n5975), .ZN(n8027) );
  OAI21_X1 U5362 ( .B1(n8116), .B2(n8115), .A(n4871), .ZN(n8070) );
  INV_X1 U5363 ( .A(n4874), .ZN(n4871) );
  AND4_X1 U5364 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n8430)
         );
  AND4_X1 U5365 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n8441)
         );
  NAND2_X1 U5366 ( .A1(n5869), .A2(n5868), .ZN(n8417) );
  NAND2_X1 U5367 ( .A1(n7107), .A2(n7106), .ZN(n4394) );
  NAND2_X1 U5368 ( .A1(n5622), .A2(n5621), .ZN(n8142) );
  NAND2_X1 U5369 ( .A1(n6828), .A2(n8462), .ZN(n8166) );
  NAND2_X1 U5370 ( .A1(n8164), .A2(n8163), .ZN(n4417) );
  INV_X1 U5371 ( .A(n8193), .ZN(n8443) );
  NAND2_X1 U5372 ( .A1(n5972), .A2(n5971), .ZN(n8185) );
  AND3_X1 U5373 ( .A1(n5898), .A2(n5897), .A3(n5896), .ZN(n8404) );
  NAND4_X1 U5374 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n6359)
         );
  OR2_X1 U5375 ( .A1(n5636), .A2(n5644), .ZN(n5650) );
  OR2_X1 U5376 ( .A1(n5658), .A2(n6805), .ZN(n5640) );
  NAND2_X1 U5377 ( .A1(n4757), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4499) );
  INV_X1 U5378 ( .A(n6760), .ZN(n4757) );
  OAI21_X1 U5379 ( .B1(n4754), .B2(n10065), .A(n4502), .ZN(n4501) );
  NOR2_X1 U5380 ( .A1(n4753), .A2(n4503), .ZN(n4502) );
  XNOR2_X1 U5381 ( .A(n4755), .B(n8251), .ZN(n4754) );
  OAI21_X1 U5382 ( .B1(n9931), .B2(n8278), .A(n8277), .ZN(n4503) );
  NAND2_X1 U5383 ( .A1(n5893), .A2(n5892), .ZN(n8394) );
  NAND2_X1 U5384 ( .A1(n6839), .A2(n6827), .ZN(n8462) );
  INV_X1 U5385 ( .A(n8452), .ZN(n8470) );
  NOR2_X1 U5386 ( .A1(n4668), .A2(n10128), .ZN(n4667) );
  INV_X1 U5387 ( .A(n6600), .ZN(n4668) );
  NAND2_X1 U5388 ( .A1(n4669), .A2(n4624), .ZN(n4623) );
  NOR2_X1 U5389 ( .A1(n6597), .A2(n4625), .ZN(n4624) );
  NAND2_X1 U5390 ( .A1(n6600), .A2(n10116), .ZN(n4625) );
  INV_X1 U5391 ( .A(n6463), .ZN(n8033) );
  AND2_X1 U5392 ( .A1(n5952), .A2(n5951), .ZN(n8559) );
  AND2_X1 U5393 ( .A1(n5915), .A2(n5914), .ZN(n8571) );
  INV_X1 U5394 ( .A(n8909), .ZN(n7184) );
  AND4_X1 U5395 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n8626)
         );
  INV_X1 U5396 ( .A(n9432), .ZN(n9278) );
  NAND2_X1 U5397 ( .A1(n5328), .A2(n5327), .ZN(n8676) );
  INV_X1 U5398 ( .A(n9870), .ZN(n7280) );
  INV_X1 U5399 ( .A(n9443), .ZN(n9286) );
  NAND2_X1 U5400 ( .A1(n5096), .A2(n5095), .ZN(n9347) );
  AOI21_X1 U5401 ( .B1(n6324), .B2(n6323), .A(n9865), .ZN(n8754) );
  NOR2_X2 U5402 ( .A1(n6320), .A2(n6327), .ZN(n8746) );
  INV_X1 U5403 ( .A(n4466), .ZN(n4765) );
  NAND2_X1 U5404 ( .A1(n9020), .A2(n9022), .ZN(n4464) );
  INV_X1 U5405 ( .A(n4763), .ZN(n4762) );
  OAI21_X1 U5406 ( .B1(n9023), .B2(n9022), .A(n4341), .ZN(n4763) );
  INV_X1 U5407 ( .A(n7331), .ZN(n9050) );
  AOI22_X1 U5408 ( .A1(n5531), .A2(n9482), .B1(n9161), .B2(n9038), .ZN(n9185)
         );
  NAND2_X1 U5409 ( .A1(n5385), .A2(n5384), .ZN(n9310) );
  NAND2_X1 U5410 ( .A1(n5102), .A2(n5101), .ZN(n8766) );
  INV_X2 U5411 ( .A(n9383), .ZN(n9876) );
  NAND2_X1 U5412 ( .A1(n9908), .A2(n9427), .ZN(n9534) );
  INV_X1 U5413 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U5414 ( .A1(n4311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5057) );
  OAI21_X1 U5415 ( .B1(n4656), .B2(n6354), .A(n6353), .ZN(n6355) );
  OAI21_X1 U5416 ( .B1(n8787), .B2(n8783), .A(n4334), .ZN(n8779) );
  NAND2_X1 U5417 ( .A1(n6373), .A2(n4535), .ZN(n4534) );
  OAI21_X1 U5418 ( .B1(n4522), .B2(n4521), .A(n4520), .ZN(n4519) );
  NAND2_X1 U5419 ( .A1(n4518), .A2(n4513), .ZN(n4512) );
  INV_X1 U5420 ( .A(n6421), .ZN(n4513) );
  AOI21_X1 U5421 ( .B1(n4510), .B2(n4517), .A(n4351), .ZN(n4507) );
  INV_X1 U5422 ( .A(n8776), .ZN(n4472) );
  NAND2_X1 U5423 ( .A1(n4478), .A2(n4477), .ZN(n4476) );
  NOR2_X1 U5424 ( .A1(n8825), .A2(n9025), .ZN(n4477) );
  NAND2_X1 U5425 ( .A1(n4479), .A2(n8826), .ZN(n4478) );
  NAND2_X1 U5426 ( .A1(n4474), .A2(n9025), .ZN(n4473) );
  NAND2_X1 U5427 ( .A1(n4480), .A2(n4309), .ZN(n4475) );
  NAND2_X1 U5428 ( .A1(n4472), .A2(n8777), .ZN(n8916) );
  NAND2_X1 U5429 ( .A1(n6425), .A2(n4529), .ZN(n4528) );
  INV_X1 U5430 ( .A(n9294), .ZN(n4457) );
  OAI21_X1 U5431 ( .B1(n8858), .B2(n4459), .A(n8857), .ZN(n4458) );
  NOR2_X1 U5432 ( .A1(n7424), .A2(n4657), .ZN(n6522) );
  AND2_X1 U5433 ( .A1(n6346), .A2(n6345), .ZN(n6458) );
  NAND2_X1 U5434 ( .A1(n4301), .A2(n8960), .ZN(n4469) );
  INV_X1 U5435 ( .A(n8115), .ZN(n4875) );
  INV_X1 U5436 ( .A(n4877), .ZN(n4876) );
  OAI21_X1 U5437 ( .B1(n8069), .B2(n4305), .A(n4878), .ZN(n4877) );
  INV_X1 U5438 ( .A(n8136), .ZN(n4878) );
  AND2_X1 U5439 ( .A1(n6511), .A2(n6510), .ZN(n6543) );
  NOR2_X1 U5440 ( .A1(n8232), .A2(n4367), .ZN(n4728) );
  NAND2_X1 U5441 ( .A1(n9932), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4735) );
  INV_X1 U5442 ( .A(n4596), .ZN(n4591) );
  NAND2_X1 U5443 ( .A1(n4882), .A2(n5989), .ZN(n4881) );
  AND2_X1 U5444 ( .A1(n5986), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U5445 ( .A1(n4678), .A2(n5602), .ZN(n4677) );
  INV_X1 U5446 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5602) );
  INV_X1 U5447 ( .A(n5601), .ZN(n4678) );
  INV_X1 U5448 ( .A(n8653), .ZN(n4438) );
  NOR2_X1 U5449 ( .A1(n4426), .A2(n4427), .ZN(n4425) );
  INV_X1 U5450 ( .A(n7616), .ZN(n4427) );
  INV_X1 U5451 ( .A(n6169), .ZN(n4422) );
  INV_X1 U5452 ( .A(n8817), .ZN(n4560) );
  INV_X1 U5453 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5049) );
  INV_X1 U5454 ( .A(n4796), .ZN(n4795) );
  OAI21_X1 U5455 ( .B1(n4798), .B2(n4797), .A(n5406), .ZN(n4796) );
  INV_X1 U5456 ( .A(n5009), .ZN(n4797) );
  AND2_X1 U5457 ( .A1(n5369), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5458 ( .A1(n5352), .A2(n4994), .ZN(n4806) );
  INV_X1 U5459 ( .A(n4994), .ZN(n4802) );
  INV_X1 U5460 ( .A(n5337), .ZN(n4770) );
  INV_X1 U5461 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n4954) );
  INV_X1 U5462 ( .A(n4760), .ZN(n4759) );
  OAI21_X1 U5463 ( .B1(n4932), .B2(n4761), .A(n4935), .ZN(n4760) );
  INV_X1 U5464 ( .A(n4934), .ZN(n4761) );
  INV_X1 U5465 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4906) );
  INV_X1 U5466 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4904) );
  AOI21_X1 U5467 ( .B1(n4868), .B2(n4867), .A(n8148), .ZN(n4866) );
  INV_X1 U5468 ( .A(n8091), .ZN(n4867) );
  INV_X1 U5469 ( .A(n7991), .ZN(n4870) );
  NOR3_X1 U5470 ( .A1(n6466), .A2(n6467), .A3(n4385), .ZN(n6486) );
  NOR2_X1 U5471 ( .A1(n6487), .A2(n8298), .ZN(n4385) );
  AOI21_X1 U5472 ( .B1(n8027), .B2(n6488), .A(n6487), .ZN(n4533) );
  NAND2_X1 U5473 ( .A1(n5657), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U5474 ( .A1(n10034), .A2(n4495), .ZN(n8271) );
  OR2_X1 U5475 ( .A1(n10033), .A2(n8530), .ZN(n4495) );
  INV_X1 U5476 ( .A(n4641), .ZN(n4640) );
  INV_X1 U5477 ( .A(n6452), .ZN(n4645) );
  NAND2_X1 U5478 ( .A1(n5594), .A2(n5593), .ZN(n5910) );
  NAND2_X1 U5479 ( .A1(n5592), .A2(n5591), .ZN(n5901) );
  INV_X1 U5480 ( .A(n5894), .ZN(n5592) );
  AND2_X1 U5481 ( .A1(n4312), .A2(n5832), .ZN(n4589) );
  NOR2_X1 U5482 ( .A1(n7868), .A2(n8195), .ZN(n5793) );
  INV_X1 U5483 ( .A(n4535), .ZN(n6397) );
  INV_X1 U5484 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U5485 ( .A1(n4629), .A2(n4627), .ZN(n5719) );
  OAI211_X1 U5486 ( .C1(n5620), .C2(n5619), .A(n4633), .B(n5613), .ZN(n6003)
         );
  OR2_X1 U5487 ( .A1(n6034), .A2(n4634), .ZN(n4633) );
  AND2_X1 U5488 ( .A1(n5988), .A2(n4879), .ZN(n6034) );
  INV_X1 U5489 ( .A(n4881), .ZN(n4879) );
  INV_X1 U5490 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5600) );
  INV_X1 U5491 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5596) );
  OR2_X1 U5492 ( .A1(n8719), .A2(n8723), .ZN(n4817) );
  NAND2_X1 U5493 ( .A1(n8719), .A2(n8723), .ZN(n4816) );
  AND2_X1 U5494 ( .A1(n4439), .A2(n4438), .ZN(n4437) );
  INV_X1 U5495 ( .A(n7296), .ZN(n4431) );
  NAND2_X1 U5496 ( .A1(n4493), .A2(n4488), .ZN(n4487) );
  NOR2_X1 U5497 ( .A1(n9193), .A2(n4455), .ZN(n4454) );
  INV_X1 U5498 ( .A(n4456), .ZN(n4455) );
  NOR2_X1 U5499 ( .A1(n9208), .A2(n9230), .ZN(n4456) );
  OAI21_X1 U5500 ( .B1(n4700), .B2(n4697), .A(n5417), .ZN(n4696) );
  OR2_X1 U5501 ( .A1(n9280), .A2(n9441), .ZN(n5417) );
  INV_X1 U5502 ( .A(n4895), .ZN(n4697) );
  AND2_X1 U5503 ( .A1(n9435), .A2(n9285), .ZN(n9252) );
  NAND2_X1 U5504 ( .A1(n5070), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5398) );
  INV_X1 U5505 ( .A(n5386), .ZN(n5070) );
  NOR2_X1 U5506 ( .A1(n5522), .A2(n4547), .ZN(n4546) );
  INV_X1 U5507 ( .A(n8846), .ZN(n4547) );
  NAND2_X1 U5508 ( .A1(n4544), .A2(n8950), .ZN(n4543) );
  INV_X1 U5509 ( .A(n9329), .ZN(n4544) );
  OR2_X1 U5510 ( .A1(n9338), .A2(n4451), .ZN(n4450) );
  NAND2_X1 U5511 ( .A1(n5067), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U5512 ( .A1(n5066), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5314) );
  INV_X1 U5513 ( .A(n5312), .ZN(n5066) );
  INV_X1 U5514 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5294) );
  OR2_X1 U5515 ( .A1(n5295), .A2(n5294), .ZN(n5312) );
  NOR2_X1 U5516 ( .A1(n4560), .A2(n4559), .ZN(n4558) );
  INV_X1 U5517 ( .A(n8812), .ZN(n4559) );
  OAI21_X1 U5518 ( .B1(n8996), .B2(n4560), .A(n8997), .ZN(n4556) );
  NAND2_X1 U5519 ( .A1(n5065), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5280) );
  INV_X1 U5520 ( .A(n5266), .ZN(n5065) );
  NOR2_X1 U5521 ( .A1(n7557), .A2(n4448), .ZN(n4447) );
  NAND2_X1 U5522 ( .A1(n7492), .A2(n4449), .ZN(n4448) );
  INV_X1 U5523 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5252) );
  OR3_X1 U5524 ( .A1(n8801), .A2(n5515), .A3(n8780), .ZN(n8993) );
  OR2_X1 U5525 ( .A1(n7279), .A2(n7280), .ZN(n7198) );
  NOR2_X1 U5526 ( .A1(n6901), .A2(n7213), .ZN(n6902) );
  XNOR2_X1 U5527 ( .A(n6471), .B(n6470), .ZN(n6469) );
  AOI21_X1 U5528 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n5480) );
  INV_X1 U5529 ( .A(SI_17_), .ZN(n9603) );
  AND2_X1 U5530 ( .A1(n5027), .A2(n5026), .ZN(n5432) );
  AND3_X1 U5531 ( .A1(n5496), .A2(n5495), .A3(n5494), .ZN(n5497) );
  INV_X1 U5532 ( .A(n5322), .ZN(n4776) );
  NAND2_X1 U5533 ( .A1(n4923), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4387) );
  OAI21_X1 U5534 ( .B1(n8770), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4918), .ZN(
        n4919) );
  NAND2_X1 U5535 ( .A1(n4923), .A2(n6614), .ZN(n4918) );
  OAI21_X1 U5536 ( .B1(n4923), .B2(n4713), .A(n4712), .ZN(n4912) );
  NAND2_X1 U5537 ( .A1(n4923), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4712) );
  INV_X1 U5538 ( .A(n4857), .ZN(n4856) );
  NAND2_X1 U5539 ( .A1(n7463), .A2(n4297), .ZN(n4414) );
  NOR2_X1 U5540 ( .A1(n7999), .A2(n8191), .ZN(n4874) );
  INV_X1 U5541 ( .A(n4408), .ZN(n4407) );
  AOI21_X1 U5542 ( .B1(n4408), .B2(n4406), .A(n4338), .ZN(n4405) );
  INV_X1 U5543 ( .A(n8048), .ZN(n4406) );
  OR2_X1 U5544 ( .A1(n7990), .A2(n8441), .ZN(n7991) );
  AND2_X1 U5545 ( .A1(n8079), .A2(n8007), .ZN(n8106) );
  OR2_X1 U5546 ( .A1(n7924), .A2(n4903), .ZN(n4401) );
  NOR2_X1 U5547 ( .A1(n7848), .A2(n4402), .ZN(n7924) );
  OR2_X1 U5548 ( .A1(n7847), .A2(n7923), .ZN(n4402) );
  XNOR2_X1 U5549 ( .A(n7236), .B(n7269), .ZN(n7098) );
  NAND2_X1 U5550 ( .A1(n5590), .A2(n5589), .ZN(n5881) );
  INV_X1 U5551 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U5552 ( .A1(n8011), .A2(n8080), .ZN(n8082) );
  AND2_X1 U5553 ( .A1(n8171), .A2(n4317), .ZN(n4408) );
  NAND2_X1 U5554 ( .A1(n8049), .A2(n8048), .ZN(n4409) );
  AND2_X1 U5555 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  AND4_X1 U5556 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n7232)
         );
  NAND2_X1 U5557 ( .A1(n6788), .A2(n6789), .ZN(n6787) );
  NAND2_X1 U5558 ( .A1(n6922), .A2(n4310), .ZN(n4498) );
  NAND2_X1 U5559 ( .A1(n9951), .A2(n8262), .ZN(n9968) );
  AND2_X1 U5560 ( .A1(n4737), .A2(n4333), .ZN(n10012) );
  NAND2_X1 U5561 ( .A1(n9985), .A2(n8267), .ZN(n10003) );
  NOR2_X1 U5562 ( .A1(n10026), .A2(n8245), .ZN(n10045) );
  INV_X1 U5563 ( .A(n4384), .ZN(n8244) );
  NOR2_X1 U5564 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  NAND2_X1 U5565 ( .A1(n5850), .A2(n4397), .ZN(n4396) );
  NAND2_X1 U5566 ( .A1(n10019), .A2(n8270), .ZN(n10035) );
  NAND2_X1 U5567 ( .A1(n10035), .A2(n10036), .ZN(n10034) );
  XNOR2_X1 U5568 ( .A(n8271), .B(n10051), .ZN(n10055) );
  AND2_X1 U5569 ( .A1(n9738), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4756) );
  NOR2_X1 U5570 ( .A1(n4617), .A2(n5974), .ZN(n4616) );
  INV_X1 U5571 ( .A(n6585), .ZN(n4617) );
  AND2_X1 U5572 ( .A1(n6443), .A2(n6439), .ZN(n4679) );
  AND2_X1 U5573 ( .A1(n6513), .A2(n6512), .ZN(n8334) );
  OR2_X1 U5574 ( .A1(n5916), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U5575 ( .A1(n5927), .A2(n8110), .ZN(n5942) );
  INV_X1 U5576 ( .A(n5928), .ZN(n5927) );
  AND2_X1 U5577 ( .A1(n6439), .A2(n6438), .ZN(n8350) );
  OAI21_X1 U5578 ( .B1(n8373), .B2(n6027), .A(n6434), .ZN(n8360) );
  AOI21_X1 U5579 ( .B1(n4607), .B2(n4609), .A(n4605), .ZN(n4604) );
  INV_X1 U5580 ( .A(n8362), .ZN(n4605) );
  AOI21_X1 U5581 ( .B1(n8401), .B2(n5887), .A(n4294), .ZN(n8384) );
  INV_X1 U5582 ( .A(n4584), .ZN(n4583) );
  OAI21_X1 U5583 ( .B1(n4586), .B2(n4585), .A(n5863), .ZN(n4584) );
  NAND2_X1 U5584 ( .A1(n4652), .A2(n4650), .ZN(n8423) );
  AOI21_X1 U5585 ( .B1(n4653), .B2(n4655), .A(n4651), .ZN(n4650) );
  INV_X1 U5586 ( .A(n6417), .ZN(n4651) );
  INV_X1 U5587 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5585) );
  INV_X1 U5588 ( .A(n5814), .ZN(n5586) );
  NAND2_X1 U5589 ( .A1(n7857), .A2(n7846), .ZN(n4659) );
  INV_X1 U5590 ( .A(n7846), .ZN(n7861) );
  OR2_X1 U5591 ( .A1(n5743), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5757) );
  OR2_X1 U5592 ( .A1(n5703), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U5593 ( .A1(n5581), .A2(n7042), .ZN(n5743) );
  INV_X1 U5594 ( .A(n5729), .ZN(n5581) );
  NAND2_X1 U5595 ( .A1(n7369), .A2(n6521), .ZN(n7407) );
  AND4_X1 U5596 ( .A1(n5692), .A2(n5691), .A3(n5690), .A4(n5689), .ZN(n7482)
         );
  NAND2_X1 U5597 ( .A1(n6390), .A2(n6366), .ZN(n7424) );
  AND2_X1 U5598 ( .A1(n7247), .A2(n10095), .ZN(n6827) );
  NAND2_X1 U5599 ( .A1(n5880), .A2(n5879), .ZN(n8145) );
  AND2_X1 U5600 ( .A1(n5773), .A2(n5772), .ZN(n10100) );
  AND2_X1 U5601 ( .A1(n5701), .A2(n5700), .ZN(n10081) );
  NOR2_X1 U5602 ( .A1(n6840), .A2(n6568), .ZN(n6822) );
  NOR2_X1 U5603 ( .A1(n6833), .A2(n6077), .ZN(n6826) );
  AND2_X1 U5604 ( .A1(n6836), .A2(n6843), .ZN(n6839) );
  AND2_X1 U5605 ( .A1(n6743), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6843) );
  AOI21_X1 U5606 ( .B1(n5613), .B2(n4328), .A(n4849), .ZN(n4848) );
  NAND2_X1 U5607 ( .A1(n6037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6039) );
  INV_X1 U5608 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6035) );
  INV_X1 U5609 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5711) );
  OR2_X1 U5610 ( .A1(n5675), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5695) );
  INV_X1 U5611 ( .A(n4443), .ZN(n4441) );
  OAI21_X1 U5612 ( .B1(n8666), .B2(n6229), .A(n8667), .ZN(n6233) );
  NAND2_X1 U5613 ( .A1(n4811), .A2(n4815), .ZN(n8692) );
  NAND2_X1 U5614 ( .A1(n4293), .A2(n4817), .ZN(n4811) );
  NAND2_X1 U5615 ( .A1(n7614), .A2(n7616), .ZN(n7615) );
  AOI21_X1 U5616 ( .B1(n4836), .B2(n4834), .A(n4833), .ZN(n4832) );
  INV_X1 U5617 ( .A(n6259), .ZN(n4833) );
  INV_X1 U5618 ( .A(n4841), .ZN(n4834) );
  INV_X1 U5619 ( .A(n4836), .ZN(n4835) );
  NAND2_X1 U5620 ( .A1(n5069), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5373) );
  INV_X1 U5621 ( .A(n5362), .ZN(n5069) );
  NAND2_X1 U5622 ( .A1(n4293), .A2(n8719), .ZN(n8722) );
  NAND2_X1 U5623 ( .A1(n7803), .A2(n7804), .ZN(n7802) );
  NAND2_X1 U5624 ( .A1(n5068), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5345) );
  INV_X1 U5625 ( .A(n5343), .ZN(n5068) );
  OR2_X1 U5626 ( .A1(n5345), .A2(n5086), .ZN(n5362) );
  NAND2_X1 U5627 ( .A1(n8665), .A2(n4841), .ZN(n4837) );
  INV_X1 U5628 ( .A(n6132), .ZN(n4828) );
  NAND2_X1 U5629 ( .A1(n4825), .A2(n6132), .ZN(n4827) );
  INV_X1 U5630 ( .A(n8705), .ZN(n6326) );
  INV_X1 U5631 ( .A(n6231), .ZN(n8666) );
  NAND2_X1 U5632 ( .A1(n4306), .A2(n4465), .ZN(n4462) );
  NOR2_X1 U5633 ( .A1(n8885), .A2(n8887), .ZN(n4465) );
  OR2_X1 U5634 ( .A1(n9029), .A2(n9028), .ZN(n4764) );
  OR2_X1 U5635 ( .A1(n9772), .A2(n9771), .ZN(n9774) );
  NAND2_X1 U5636 ( .A1(n9238), .A2(n4454), .ZN(n9191) );
  OR2_X1 U5637 ( .A1(n9193), .A2(n9212), .ZN(n8953) );
  AND2_X1 U5638 ( .A1(n5493), .A2(n5492), .ZN(n9196) );
  AND2_X1 U5639 ( .A1(n8953), .A2(n8870), .ZN(n9188) );
  AND2_X1 U5640 ( .A1(n5085), .A2(n5084), .ZN(n9228) );
  NAND2_X1 U5641 ( .A1(n9238), .A2(n9412), .ZN(n9223) );
  NOR2_X1 U5642 ( .A1(n9221), .A2(n4710), .ZN(n9220) );
  AND2_X1 U5643 ( .A1(n5458), .A2(n5457), .ZN(n9244) );
  OR2_X1 U5644 ( .A1(n9224), .A2(n5488), .ZN(n5458) );
  AND2_X1 U5645 ( .A1(n9420), .A2(n9253), .ZN(n9238) );
  NAND2_X1 U5646 ( .A1(n4571), .A2(n8891), .ZN(n4570) );
  NOR2_X1 U5647 ( .A1(n9259), .A2(n9260), .ZN(n9257) );
  AND2_X1 U5648 ( .A1(n9256), .A2(n9252), .ZN(n9253) );
  NOR2_X1 U5649 ( .A1(n9286), .A2(n9303), .ZN(n9285) );
  AND2_X1 U5650 ( .A1(n5416), .A2(n5415), .ZN(n9291) );
  NAND2_X1 U5651 ( .A1(n4536), .A2(n4539), .ZN(n9300) );
  AND2_X1 U5652 ( .A1(n4540), .A2(n4358), .ZN(n4539) );
  NAND2_X1 U5653 ( .A1(n4545), .A2(n4543), .ZN(n9317) );
  NAND2_X1 U5654 ( .A1(n9343), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U5655 ( .A1(n9317), .A2(n9316), .ZN(n9315) );
  NOR2_X1 U5656 ( .A1(n9372), .A2(n4451), .ZN(n9346) );
  NAND2_X1 U5657 ( .A1(n7893), .A2(n9004), .ZN(n9362) );
  OAI211_X1 U5658 ( .C1(n7627), .C2(n4564), .A(n5521), .B(n4563), .ZN(n7818)
         );
  INV_X1 U5659 ( .A(n4565), .ZN(n4564) );
  NAND2_X1 U5660 ( .A1(n4565), .A2(n8998), .ZN(n4563) );
  AND2_X1 U5661 ( .A1(n8632), .A2(n7706), .ZN(n7821) );
  AOI21_X1 U5662 ( .B1(n7603), .B2(n4683), .A(n4681), .ZN(n4680) );
  NAND2_X1 U5663 ( .A1(n4682), .A2(n5301), .ZN(n4681) );
  OR2_X1 U5664 ( .A1(n8716), .A2(n9041), .ZN(n5301) );
  NOR2_X1 U5665 ( .A1(n8716), .A2(n7630), .ZN(n7706) );
  NAND2_X1 U5666 ( .A1(n4446), .A2(n4447), .ZN(n7630) );
  NOR2_X1 U5667 ( .A1(n7506), .A2(n7947), .ZN(n4446) );
  NAND2_X1 U5668 ( .A1(n7357), .A2(n8812), .ZN(n7487) );
  NAND2_X1 U5669 ( .A1(n4445), .A2(n4447), .ZN(n7604) );
  INV_X1 U5670 ( .A(n7506), .ZN(n4445) );
  NAND2_X1 U5671 ( .A1(n6704), .A2(n8878), .ZN(n5233) );
  NAND2_X1 U5672 ( .A1(n9893), .A2(n9046), .ZN(n8795) );
  AOI21_X1 U5673 ( .B1(n7195), .B2(n5228), .A(n4884), .ZN(n7397) );
  AND2_X1 U5674 ( .A1(n7194), .A2(n5225), .ZN(n5228) );
  INV_X1 U5675 ( .A(n5227), .ZN(n5225) );
  NAND2_X1 U5676 ( .A1(n5226), .A2(n4724), .ZN(n7392) );
  NAND2_X1 U5677 ( .A1(n5119), .A2(n5118), .ZN(n7613) );
  NAND2_X1 U5678 ( .A1(n6661), .A2(n8878), .ZN(n5119) );
  OR2_X1 U5679 ( .A1(n7447), .A2(n7613), .ZN(n7506) );
  NOR2_X1 U5680 ( .A1(n7198), .A2(n7302), .ZN(n7448) );
  OR2_X1 U5681 ( .A1(n8776), .A2(n4551), .ZN(n4550) );
  INV_X1 U5682 ( .A(n4549), .ZN(n4548) );
  AND4_X1 U5683 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n7619)
         );
  NAND2_X1 U5684 ( .A1(n6902), .A2(n7126), .ZN(n6964) );
  NAND2_X1 U5685 ( .A1(n6886), .A2(n5510), .ZN(n6905) );
  NAND2_X1 U5686 ( .A1(n8981), .A2(n6955), .ZN(n6886) );
  AND2_X1 U5687 ( .A1(n8896), .A2(n8859), .ZN(n9301) );
  AOI21_X1 U5688 ( .B1(n4719), .B2(n4718), .A(n4336), .ZN(n4717) );
  NAND2_X1 U5689 ( .A1(n5310), .A2(n5309), .ZN(n7708) );
  AND4_X1 U5690 ( .A1(n5110), .A2(n5109), .A3(n5108), .A4(n5107), .ZN(n8673)
         );
  AND4_X1 U5691 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n7656)
         );
  AND4_X1 U5692 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n7547)
         );
  AND4_X1 U5693 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n7033)
         );
  INV_X1 U5694 ( .A(n9427), .ZN(n9901) );
  AND3_X1 U5695 ( .A1(n6314), .A2(n7131), .A3(n5565), .ZN(n5571) );
  AND2_X1 U5696 ( .A1(n4845), .A2(n5054), .ZN(n4843) );
  NOR2_X1 U5697 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n4846), .ZN(n4845) );
  AND2_X1 U5698 ( .A1(n4844), .A2(n5046), .ZN(n4578) );
  INV_X1 U5699 ( .A(n4846), .ZN(n4844) );
  MUX2_X1 U5700 ( .A(n9554), .B(n5540), .S(P1_IR_REG_24__SCAN_IN), .Z(n5541)
         );
  NAND2_X1 U5701 ( .A1(n4804), .A2(n4994), .ZN(n5370) );
  NAND2_X1 U5702 ( .A1(n4777), .A2(n4778), .ZN(n5323) );
  OAI21_X1 U5703 ( .B1(n5303), .B2(n5302), .A(n4971), .ZN(n5098) );
  OAI21_X1 U5704 ( .B1(n4948), .B2(n4296), .A(n4785), .ZN(n5274) );
  NAND2_X1 U5705 ( .A1(n4948), .A2(n4789), .ZN(n4788) );
  AND2_X1 U5706 ( .A1(n5248), .A2(n5247), .ZN(n5276) );
  XNOR2_X1 U5707 ( .A(n5112), .B(n5111), .ZN(n6661) );
  AND2_X1 U5708 ( .A1(n4688), .A2(n4686), .ZN(n4689) );
  AOI21_X1 U5709 ( .B1(n4930), .B2(n4318), .A(n4687), .ZN(n4686) );
  NAND2_X1 U5710 ( .A1(n8164), .A2(n8015), .ZN(n8038) );
  NAND2_X1 U5711 ( .A1(n4412), .A2(n8105), .ZN(n8055) );
  INV_X1 U5712 ( .A(n4413), .ZN(n4412) );
  INV_X1 U5713 ( .A(n8571), .ZN(n8059) );
  INV_X1 U5714 ( .A(n6359), .ZN(n7114) );
  AND4_X1 U5715 ( .A1(n5763), .A2(n5762), .A3(n5761), .A4(n5760), .ZN(n7577)
         );
  NAND2_X1 U5716 ( .A1(n7519), .A2(n7518), .ZN(n7665) );
  AND3_X1 U5717 ( .A1(n5905), .A2(n5904), .A3(n5903), .ZN(n8387) );
  NAND2_X1 U5718 ( .A1(n5907), .A2(n5906), .ZN(n8074) );
  INV_X1 U5719 ( .A(n4401), .ZN(n7985) );
  OAI21_X1 U5720 ( .B1(n8049), .B2(n4407), .A(n4405), .ZN(n8092) );
  NAND2_X1 U5721 ( .A1(n8092), .A2(n8091), .ZN(n8090) );
  NAND2_X1 U5722 ( .A1(n8090), .A2(n7991), .ZN(n8098) );
  XNOR2_X1 U5723 ( .A(n5683), .B(n7231), .ZN(n7151) );
  OAI21_X1 U5724 ( .B1(n7461), .B2(n4860), .A(n4859), .ZN(n7790) );
  NAND2_X1 U5725 ( .A1(n4399), .A2(n4398), .ZN(n8126) );
  OR2_X1 U5726 ( .A1(n7982), .A2(n7983), .ZN(n4398) );
  NAND2_X1 U5727 ( .A1(n4401), .A2(n4400), .ZN(n4399) );
  INV_X1 U5728 ( .A(n7984), .ZN(n4400) );
  NAND2_X1 U5729 ( .A1(n5812), .A2(n5811), .ZN(n8133) );
  OR2_X1 U5730 ( .A1(n6825), .A2(n6824), .ZN(n8158) );
  AOI21_X1 U5731 ( .B1(n8070), .B2(n8069), .A(n4305), .ZN(n8138) );
  INV_X1 U5732 ( .A(n8177), .ZN(n8155) );
  OR2_X1 U5733 ( .A1(n6825), .A2(n6823), .ZN(n8177) );
  AND2_X1 U5734 ( .A1(n4409), .A2(n4317), .ZN(n8172) );
  NAND2_X1 U5735 ( .A1(n4409), .A2(n4408), .ZN(n8170) );
  NAND2_X1 U5736 ( .A1(n7111), .A2(n7940), .ZN(n8179) );
  NAND2_X1 U5737 ( .A1(n5948), .A2(n5947), .ZN(n8186) );
  INV_X1 U5738 ( .A(n8430), .ZN(n8456) );
  INV_X1 U5739 ( .A(n7661), .ZN(n8198) );
  INV_X1 U5740 ( .A(n7482), .ZN(n8200) );
  NAND4_X1 U5741 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n8201)
         );
  NAND2_X1 U5742 ( .A1(n5657), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5662) );
  OR2_X1 U5743 ( .A1(n5634), .A2(n10118), .ZN(n5659) );
  CLKBUF_X1 U5744 ( .A(n7013), .Z(n8202) );
  OR2_X1 U5745 ( .A1(n6836), .A2(n6626), .ZN(n9736) );
  OR2_X1 U5746 ( .A1(P2_U3150), .A2(n6745), .ZN(n9931) );
  XNOR2_X1 U5747 ( .A(n4498), .B(n4497), .ZN(n7041) );
  INV_X1 U5748 ( .A(n4749), .ZN(n4748) );
  AOI21_X1 U5749 ( .B1(n7041), .B2(P2_REG1_REG_5__SCAN_IN), .A(n4496), .ZN(
        n7068) );
  AND2_X1 U5750 ( .A1(n4498), .A2(n7049), .ZN(n4496) );
  AND2_X1 U5751 ( .A1(n4731), .A2(n4730), .ZN(n9943) );
  INV_X1 U5752 ( .A(n4734), .ZN(n4730) );
  INV_X1 U5753 ( .A(n4737), .ZN(n9995) );
  AND2_X1 U5754 ( .A1(P2_U3893), .A2(n6002), .ZN(n10060) );
  INV_X1 U5755 ( .A(n4743), .ZN(n10063) );
  INV_X1 U5756 ( .A(n9931), .ZN(n10053) );
  INV_X1 U5757 ( .A(n6590), .ZN(n6591) );
  NOR2_X1 U5758 ( .A1(n8444), .A2(n8310), .ZN(n6006) );
  OR2_X1 U5759 ( .A1(n6540), .A2(n8295), .ZN(n6030) );
  NAND2_X1 U5760 ( .A1(n8301), .A2(n8300), .ZN(n8302) );
  NAND2_X1 U5761 ( .A1(n4646), .A2(n6452), .ZN(n8312) );
  NAND2_X1 U5762 ( .A1(n8324), .A2(n6451), .ZN(n4646) );
  NAND2_X1 U5763 ( .A1(n6028), .A2(n6439), .ZN(n8338) );
  NAND2_X1 U5764 ( .A1(n4612), .A2(n4613), .ZN(n8375) );
  AND2_X1 U5765 ( .A1(n4662), .A2(n6422), .ZN(n8400) );
  NAND2_X1 U5766 ( .A1(n8426), .A2(n8425), .ZN(n8424) );
  NAND2_X1 U5767 ( .A1(n8467), .A2(n6412), .ZN(n8436) );
  NAND2_X1 U5768 ( .A1(n5833), .A2(n5832), .ZN(n8438) );
  OR2_X1 U5769 ( .A1(n7247), .A2(n10111), .ZN(n8464) );
  INV_X1 U5770 ( .A(n4592), .ZN(n7932) );
  AOI21_X1 U5771 ( .B1(n4599), .B2(n4598), .A(n4593), .ZN(n4592) );
  INV_X1 U5772 ( .A(n10100), .ZN(n7799) );
  AND2_X1 U5773 ( .A1(n4648), .A2(n6375), .ZN(n7684) );
  NAND2_X1 U5774 ( .A1(n7587), .A2(n6371), .ZN(n7584) );
  INV_X1 U5775 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7429) );
  OAI211_X1 U5776 ( .C1(n6616), .C2(n5680), .A(n5666), .B(n5665), .ZN(n7430)
         );
  INV_X1 U5777 ( .A(n7269), .ZN(n7270) );
  XNOR2_X1 U5778 ( .A(n4656), .B(n6976), .ZN(n6977) );
  NOR2_X1 U5779 ( .A1(n6974), .A2(n4379), .ZN(n7275) );
  OR2_X1 U5780 ( .A1(n8447), .A2(n7248), .ZN(n8452) );
  INV_X1 U5781 ( .A(n8462), .ZN(n8446) );
  INV_X1 U5782 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4671) );
  AOI21_X1 U5783 ( .B1(n8771), .B2(n6500), .A(n4885), .ZN(n8547) );
  INV_X1 U5784 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5785 ( .A1(n5962), .A2(n5961), .ZN(n8553) );
  INV_X1 U5786 ( .A(n8077), .ZN(n8563) );
  AND2_X1 U5787 ( .A1(n5926), .A2(n5925), .ZN(n8567) );
  INV_X1 U5788 ( .A(n8142), .ZN(n8575) );
  INV_X1 U5789 ( .A(n8074), .ZN(n8579) );
  INV_X1 U5790 ( .A(n8145), .ZN(n8586) );
  INV_X1 U5791 ( .A(n8089), .ZN(n8593) );
  INV_X1 U5792 ( .A(n8168), .ZN(n8597) );
  INV_X1 U5793 ( .A(n8133), .ZN(n8603) );
  INV_X1 U5795 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5604) );
  OR2_X1 U5796 ( .A1(n5614), .A2(n5606), .ZN(n5607) );
  INV_X1 U5797 ( .A(n6066), .ZN(n8616) );
  INV_X1 U5798 ( .A(n6045), .ZN(n7959) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7841) );
  XNOR2_X1 U5800 ( .A(n5987), .B(n5986), .ZN(n7843) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7780) );
  XNOR2_X1 U5802 ( .A(n5990), .B(n5989), .ZN(n7782) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U5804 ( .A1(n5993), .A2(n5992), .ZN(n7701) );
  NAND2_X1 U5805 ( .A1(n5889), .A2(n5888), .ZN(n4411) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7626) );
  INV_X1 U5807 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7528) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7381) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7206) );
  INV_X1 U5810 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7086) );
  INV_X1 U5811 ( .A(n9984), .ZN(n8266) );
  INV_X1 U5812 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6985) );
  INV_X1 U5813 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6798) );
  INV_X1 U5814 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6711) );
  INV_X1 U5815 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6663) );
  XNOR2_X1 U5816 ( .A(n5739), .B(n5738), .ZN(n7307) );
  AND2_X1 U5817 ( .A1(n6632), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6603) );
  AND2_X1 U5818 ( .A1(n5404), .A2(n5403), .ZN(n9308) );
  AND2_X1 U5819 ( .A1(n6318), .A2(n8746), .ZN(n6319) );
  INV_X1 U5820 ( .A(n6094), .ZN(n6095) );
  AND2_X1 U5821 ( .A1(n5380), .A2(n5379), .ZN(n9336) );
  NAND2_X1 U5822 ( .A1(n4435), .A2(n4439), .ZN(n8652) );
  OR2_X1 U5823 ( .A1(n8665), .A2(n4441), .ZN(n4435) );
  INV_X1 U5824 ( .A(n4821), .ZN(n4820) );
  NOR2_X1 U5825 ( .A1(n8694), .A2(n6291), .ZN(n8659) );
  OAI21_X1 U5826 ( .B1(n8665), .B2(n6235), .A(n6234), .ZN(n8684) );
  NAND2_X1 U5827 ( .A1(n5421), .A2(n5420), .ZN(n9426) );
  NAND2_X1 U5828 ( .A1(n7953), .A2(n8878), .ZN(n5421) );
  NAND2_X1 U5829 ( .A1(n7030), .A2(n6124), .ZN(n7022) );
  AND4_X1 U5830 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n7654)
         );
  NAND2_X1 U5831 ( .A1(n4442), .A2(n4832), .ZN(n8699) );
  OR2_X1 U5832 ( .A1(n8665), .A2(n4835), .ZN(n4442) );
  AND4_X1 U5833 ( .A1(n5319), .A2(n5318), .A3(n5317), .A4(n5316), .ZN(n8714)
         );
  OAI21_X1 U5834 ( .B1(n4293), .B2(n8719), .A(n8723), .ZN(n8725) );
  AND4_X1 U5835 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n7875)
         );
  NAND2_X1 U5836 ( .A1(n6326), .A2(n6851), .ZN(n8736) );
  NAND2_X1 U5837 ( .A1(n6141), .A2(n6140), .ZN(n7295) );
  INV_X1 U5838 ( .A(n8746), .ZN(n8768) );
  AND4_X1 U5839 ( .A1(n5335), .A2(n5334), .A3(n5333), .A4(n5332), .ZN(n8763)
         );
  INV_X1 U5840 ( .A(n8754), .ZN(n8765) );
  INV_X1 U5841 ( .A(n9244), .ZN(n9417) );
  INV_X1 U5842 ( .A(n9263), .ZN(n9408) );
  NAND2_X1 U5843 ( .A1(n5430), .A2(n5429), .ZN(n9432) );
  INV_X1 U5844 ( .A(n9291), .ZN(n9441) );
  NAND2_X1 U5845 ( .A1(n5146), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5126) );
  NOR2_X1 U5846 ( .A1(n9159), .A2(n9371), .ZN(n9386) );
  NAND2_X1 U5847 ( .A1(n8881), .A2(n8880), .ZN(n9170) );
  INV_X1 U5848 ( .A(n9228), .ZN(n9409) );
  INV_X1 U5849 ( .A(n9420), .ZN(n9246) );
  INV_X1 U5850 ( .A(n9435), .ZN(n9280) );
  AND2_X1 U5851 ( .A1(n5397), .A2(n5396), .ZN(n9443) );
  NAND2_X1 U5852 ( .A1(n9343), .A2(n8846), .ZN(n9330) );
  NAND2_X1 U5853 ( .A1(n5341), .A2(n5340), .ZN(n9379) );
  NAND2_X1 U5854 ( .A1(n4567), .A2(n8929), .ZN(n7704) );
  OAI21_X1 U5855 ( .B1(n7603), .B2(n4685), .A(n4683), .ZN(n7628) );
  NAND2_X1 U5856 ( .A1(n7601), .A2(n5286), .ZN(n7629) );
  NAND2_X1 U5857 ( .A1(n7486), .A2(n8817), .ZN(n7600) );
  NAND2_X1 U5858 ( .A1(n4554), .A2(n4552), .ZN(n7282) );
  OR2_X1 U5859 ( .A1(n9876), .A2(n7136), .ZN(n9869) );
  NAND2_X1 U5860 ( .A1(n4554), .A2(n8777), .ZN(n6961) );
  OR2_X1 U5861 ( .A1(n9876), .A2(n9262), .ZN(n9349) );
  NAND2_X1 U5862 ( .A1(n7197), .A2(n7196), .ZN(n9873) );
  INV_X1 U5863 ( .A(n9374), .ZN(n9865) );
  OR2_X1 U5864 ( .A1(n9876), .A2(n9022), .ZN(n9381) );
  NAND2_X1 U5865 ( .A1(n7135), .A2(n9374), .ZN(n9383) );
  INV_X1 U5866 ( .A(n9381), .ZN(n9863) );
  INV_X1 U5867 ( .A(n9371), .ZN(n9331) );
  NAND2_X1 U5868 ( .A1(n5146), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5134) );
  AOI21_X1 U5869 ( .B1(n4690), .B2(n9430), .A(n5572), .ZN(n4691) );
  NAND2_X1 U5870 ( .A1(n4708), .A2(n4709), .ZN(n9205) );
  NAND2_X1 U5871 ( .A1(n4711), .A2(n4295), .ZN(n9219) );
  OR2_X1 U5872 ( .A1(n9234), .A2(n5444), .ZN(n4711) );
  OAI21_X1 U5873 ( .B1(n4701), .B2(n4703), .A(n4700), .ZN(n9270) );
  NOR2_X1 U5874 ( .A1(n4314), .A2(n4704), .ZN(n9284) );
  INV_X1 U5875 ( .A(n4706), .ZN(n4704) );
  OAI21_X1 U5876 ( .B1(n7891), .B2(n4719), .A(n4718), .ZN(n9342) );
  NOR2_X1 U5877 ( .A1(n7890), .A2(n5336), .ZN(n9360) );
  INV_X1 U5878 ( .A(n7708), .ZN(n8632) );
  AND2_X1 U5879 ( .A1(n5190), .A2(n5189), .ZN(n9870) );
  OR2_X1 U5880 ( .A1(n5155), .A2(n4908), .ZN(n5143) );
  XNOR2_X1 U5881 ( .A(n5544), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9569) );
  INV_X1 U5882 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U5883 ( .A1(n4794), .A2(n5009), .ZN(n5407) );
  INV_X1 U5884 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7840) );
  OR2_X1 U5885 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  INV_X1 U5886 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7778) );
  INV_X1 U5887 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5505) );
  INV_X1 U5888 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7966) );
  INV_X1 U5889 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7530) );
  INV_X1 U5890 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7421) );
  INV_X1 U5891 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7383) );
  INV_X1 U5892 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9669) );
  INV_X1 U5893 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6619) );
  CLKBUF_X1 U5894 ( .A(n7354), .Z(n8278) );
  NOR2_X1 U5895 ( .A1(n4749), .A2(n4348), .ZN(n4746) );
  NAND2_X1 U5896 ( .A1(n4416), .A2(n4371), .ZN(P2_U3180) );
  NAND2_X1 U5897 ( .A1(n4417), .A2(n8169), .ZN(n4416) );
  AND2_X1 U5898 ( .A1(n8167), .A2(n8166), .ZN(n4415) );
  NAND2_X1 U5899 ( .A1(n4504), .A2(n4500), .ZN(P2_U3201) );
  NAND2_X1 U5900 ( .A1(n8276), .A2(n10061), .ZN(n4504) );
  NAND2_X1 U5901 ( .A1(n10128), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U5902 ( .A1(n4623), .A2(n4621), .ZN(n6601) );
  NAND2_X1 U5903 ( .A1(n10117), .A2(n4622), .ZN(n4621) );
  OAI21_X1 U5904 ( .B1(n9402), .B2(n8754), .A(n6580), .ZN(n6581) );
  NAND2_X1 U5905 ( .A1(n4765), .A2(n4762), .ZN(n9035) );
  NAND2_X1 U5906 ( .A1(n4572), .A2(n5570), .ZN(P1_U3519) );
  OAI21_X1 U5907 ( .B1(n5533), .B2(n4573), .A(n9908), .ZN(n4572) );
  AND2_X2 U5908 ( .A1(n7839), .A2(n9022), .ZN(n9025) );
  INV_X2 U5909 ( .A(n5634), .ZN(n5635) );
  AND2_X2 U5910 ( .A1(n4434), .A2(n4436), .ZN(n4293) );
  INV_X2 U5911 ( .A(n6106), .ZN(n6125) );
  AND2_X1 U5912 ( .A1(n8145), .A2(n8413), .ZN(n4294) );
  AND2_X1 U5913 ( .A1(n4710), .A2(n5443), .ZN(n4295) );
  OR2_X1 U5914 ( .A1(n5260), .A2(n4787), .ZN(n4296) );
  AND2_X1 U5915 ( .A1(n4861), .A2(n7789), .ZN(n4297) );
  AND3_X1 U5916 ( .A1(n4439), .A2(n4441), .A3(n4438), .ZN(n4298) );
  INV_X1 U5917 ( .A(n7650), .ZN(n4426) );
  AND2_X1 U5918 ( .A1(n5372), .A2(n5371), .ZN(n9535) );
  AND2_X1 U5919 ( .A1(n4296), .A2(n5273), .ZN(n4299) );
  AND2_X1 U5920 ( .A1(n4709), .A2(n9215), .ZN(n4300) );
  AND2_X1 U5921 ( .A1(n8867), .A2(n4486), .ZN(n4301) );
  AND3_X1 U5922 ( .A1(n8948), .A2(n8960), .A3(n8894), .ZN(n4302) );
  OR2_X1 U5923 ( .A1(n8256), .A2(n4367), .ZN(n4303) );
  AND2_X1 U5924 ( .A1(n6025), .A2(n6420), .ZN(n4304) );
  AND2_X1 U5925 ( .A1(n5476), .A2(n5475), .ZN(n9212) );
  INV_X1 U5926 ( .A(n9212), .ZN(n9400) );
  NAND2_X1 U5927 ( .A1(n4659), .A2(n6401), .ZN(n7915) );
  INV_X2 U5928 ( .A(n5103), .ZN(n6642) );
  NAND2_X2 U5929 ( .A1(n6316), .A2(n6087), .ZN(n6108) );
  INV_X2 U5930 ( .A(n5646), .ZN(n5785) );
  NAND2_X1 U5931 ( .A1(n4635), .A2(n4641), .ZN(n6540) );
  INV_X1 U5932 ( .A(n8766), .ZN(n8830) );
  AND2_X1 U5933 ( .A1(n6316), .A2(n7182), .ZN(n6220) );
  AND2_X1 U5934 ( .A1(n8000), .A2(n8378), .ZN(n4305) );
  OR3_X1 U5935 ( .A1(n8882), .A2(n8975), .A3(n8968), .ZN(n4306) );
  INV_X1 U5936 ( .A(n8425), .ZN(n4585) );
  AND2_X1 U5937 ( .A1(n4855), .A2(n8354), .ZN(n4307) );
  NOR2_X1 U5938 ( .A1(n9394), .A2(n9212), .ZN(n4308) );
  AND2_X1 U5939 ( .A1(n8833), .A2(n8929), .ZN(n4309) );
  INV_X1 U5940 ( .A(n4831), .ZN(n4830) );
  NAND2_X1 U5941 ( .A1(n6152), .A2(n7541), .ZN(n4831) );
  OR2_X1 U5942 ( .A1(n6923), .A2(n6747), .ZN(n4310) );
  NAND2_X1 U5943 ( .A1(n4577), .A2(n5099), .ZN(n4311) );
  INV_X1 U5944 ( .A(n6518), .ZN(n4597) );
  INV_X1 U5945 ( .A(n4775), .ZN(n4774) );
  NAND2_X1 U5946 ( .A1(n4778), .A2(n4776), .ZN(n4775) );
  OR2_X1 U5947 ( .A1(n8168), .A2(n8456), .ZN(n4312) );
  OR2_X1 U5948 ( .A1(n5502), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4313) );
  INV_X1 U5949 ( .A(n6433), .ZN(n4530) );
  AND2_X1 U5950 ( .A1(n9298), .A2(n5393), .ZN(n4314) );
  AND2_X1 U5951 ( .A1(n8701), .A2(n6264), .ZN(n4315) );
  NOR2_X1 U5952 ( .A1(n5769), .A2(n4677), .ZN(n5988) );
  AND2_X1 U5953 ( .A1(n8295), .A2(n4619), .ZN(n4316) );
  NAND2_X1 U5954 ( .A1(n7988), .A2(n8443), .ZN(n4317) );
  AND2_X1 U5955 ( .A1(n4934), .A2(n4931), .ZN(n4318) );
  AND2_X1 U5956 ( .A1(n8167), .A2(n8320), .ZN(n4319) );
  INV_X1 U5957 ( .A(n6519), .ZN(n4520) );
  AND2_X1 U5958 ( .A1(n4866), .A2(n4403), .ZN(n4320) );
  INV_X1 U5959 ( .A(n8437), .ZN(n4587) );
  NOR2_X1 U5960 ( .A1(n8027), .A2(n6584), .ZN(n4321) );
  AND2_X1 U5961 ( .A1(n4600), .A2(n4591), .ZN(n4322) );
  NAND2_X1 U5962 ( .A1(n5467), .A2(n5466), .ZN(n9193) );
  INV_X1 U5963 ( .A(n7075), .ZN(n4752) );
  NOR2_X1 U5964 ( .A1(n8742), .A2(n8743), .ZN(n4323) );
  AND4_X1 U5965 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n7465)
         );
  INV_X1 U5966 ( .A(n7465), .ZN(n4628) );
  NAND2_X1 U5967 ( .A1(n5608), .A2(n8607), .ZN(n5634) );
  AND2_X1 U5968 ( .A1(n8865), .A2(n8901), .ZN(n4324) );
  AND2_X1 U5969 ( .A1(n6021), .A2(n6401), .ZN(n4325) );
  AND2_X1 U5970 ( .A1(n6436), .A2(n6605), .ZN(n4326) );
  AND2_X1 U5971 ( .A1(n4711), .A2(n5443), .ZN(n4327) );
  INV_X1 U5972 ( .A(n4869), .ZN(n4868) );
  OR2_X1 U5973 ( .A1(n8099), .A2(n4870), .ZN(n4869) );
  AND2_X1 U5974 ( .A1(n8965), .A2(n8869), .ZN(n9206) );
  AND2_X1 U5975 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4328) );
  INV_X1 U5976 ( .A(n4644), .ZN(n4643) );
  NOR2_X1 U5977 ( .A1(n6450), .A2(n4645), .ZN(n4644) );
  INV_X1 U5978 ( .A(n4839), .ZN(n4838) );
  NAND3_X1 U5979 ( .A1(n5603), .A2(n5616), .A3(n5618), .ZN(n4329) );
  INV_X1 U5980 ( .A(n9230), .ZN(n9412) );
  NAND2_X1 U5981 ( .A1(n5449), .A2(n5448), .ZN(n9230) );
  AND2_X1 U5982 ( .A1(n4469), .A2(n4807), .ZN(n4330) );
  OR2_X1 U5983 ( .A1(n9426), .A2(n9278), .ZN(n8891) );
  INV_X1 U5984 ( .A(n6597), .ZN(n4672) );
  AND2_X1 U5985 ( .A1(n6176), .A2(n6175), .ZN(n4331) );
  NAND2_X1 U5986 ( .A1(n4807), .A2(n8965), .ZN(n4332) );
  OR2_X1 U5987 ( .A1(n9984), .A2(n8241), .ZN(n4333) );
  AND2_X1 U5988 ( .A1(n8778), .A2(n8777), .ZN(n4334) );
  NOR2_X1 U5989 ( .A1(n6507), .A2(n6508), .ZN(n4335) );
  NOR2_X1 U5990 ( .A1(n9347), .A2(n9464), .ZN(n4336) );
  OR2_X1 U5991 ( .A1(n9257), .A2(n4570), .ZN(n4337) );
  NOR2_X1 U5992 ( .A1(n7989), .A2(n8430), .ZN(n4338) );
  NOR2_X1 U5993 ( .A1(n9412), .A2(n9244), .ZN(n4339) );
  OR2_X1 U5994 ( .A1(n4887), .A2(n4321), .ZN(n4340) );
  AND2_X1 U5995 ( .A1(n4764), .A2(n9027), .ZN(n4341) );
  INV_X1 U5996 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5056) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4908) );
  INV_X1 U5998 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U5999 ( .A(n6469), .B(SI_29_), .ZN(n6342) );
  NAND2_X1 U6000 ( .A1(n7788), .A2(n8197), .ZN(n4342) );
  AND2_X1 U6001 ( .A1(n5988), .A2(n5989), .ZN(n5984) );
  OR2_X1 U6002 ( .A1(n5769), .A2(n5601), .ZN(n4343) );
  AND2_X1 U6003 ( .A1(n8954), .A2(n8956), .ZN(n9010) );
  INV_X1 U6004 ( .A(n9010), .ZN(n4488) );
  AND2_X1 U6005 ( .A1(n6265), .A2(n8700), .ZN(n4344) );
  AND2_X1 U6006 ( .A1(n4936), .A2(SI_7_), .ZN(n4345) );
  AND2_X1 U6007 ( .A1(n6489), .A2(n6588), .ZN(n4346) );
  AND2_X1 U6008 ( .A1(n7663), .A2(n8198), .ZN(n4347) );
  AND2_X1 U6009 ( .A1(n7079), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4348) );
  INV_X1 U6010 ( .A(n4861), .ZN(n4860) );
  NOR2_X1 U6011 ( .A1(n7664), .A2(n4862), .ZN(n4861) );
  AND2_X1 U6012 ( .A1(n4961), .A2(SI_12_), .ZN(n4349) );
  OR2_X1 U6013 ( .A1(n4893), .A2(n4616), .ZN(n4350) );
  AND2_X1 U6014 ( .A1(n8948), .A2(n8960), .ZN(n9009) );
  INV_X1 U6015 ( .A(n9009), .ZN(n4710) );
  NAND2_X1 U6016 ( .A1(n6431), .A2(n6515), .ZN(n4351) );
  INV_X1 U6017 ( .A(n9160), .ZN(n9496) );
  AND2_X1 U6018 ( .A1(n8773), .A2(n8772), .ZN(n9160) );
  NOR2_X1 U6019 ( .A1(n8514), .A2(n8404), .ZN(n4352) );
  AND2_X1 U6020 ( .A1(n6418), .A2(n4585), .ZN(n4353) );
  NAND2_X1 U6021 ( .A1(n4467), .A2(n4576), .ZN(n4354) );
  AND2_X1 U6022 ( .A1(n8633), .A2(n4816), .ZN(n4815) );
  OR2_X1 U6023 ( .A1(n7784), .A2(n7577), .ZN(n6373) );
  INV_X1 U6024 ( .A(n8411), .ZN(n4518) );
  AND2_X1 U6025 ( .A1(n6514), .A2(n6422), .ZN(n4355) );
  NAND2_X1 U6026 ( .A1(n5360), .A2(n5359), .ZN(n9338) );
  AND2_X1 U6027 ( .A1(n4468), .A2(n4382), .ZN(n4356) );
  AND2_X1 U6028 ( .A1(n4468), .A2(n4330), .ZN(n4357) );
  AND2_X1 U6029 ( .A1(n9299), .A2(n9301), .ZN(n4358) );
  AND2_X1 U6030 ( .A1(n6430), .A2(n6434), .ZN(n8376) );
  INV_X1 U6031 ( .A(n8376), .ZN(n4611) );
  AND2_X1 U6032 ( .A1(n6307), .A2(n4897), .ZN(n4359) );
  AND2_X1 U6033 ( .A1(n6422), .A2(n6514), .ZN(n4360) );
  NAND2_X1 U6034 ( .A1(n7929), .A2(n8194), .ZN(n4361) );
  AND2_X1 U6035 ( .A1(n4785), .A2(n5273), .ZN(n4362) );
  AND2_X1 U6036 ( .A1(n4302), .A2(n4324), .ZN(n4363) );
  INV_X1 U6037 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6038 ( .A1(n4876), .A2(n4875), .ZN(n4364) );
  INV_X1 U6039 ( .A(n6010), .ZN(n8226) );
  NAND2_X1 U6040 ( .A1(n7678), .A2(n4600), .ZN(n4599) );
  INV_X1 U6041 ( .A(n6810), .ZN(n4444) );
  NAND2_X1 U6042 ( .A1(n7678), .A2(n5765), .ZN(n7719) );
  AND2_X1 U6043 ( .A1(n8090), .A2(n4868), .ZN(n4365) );
  OR2_X1 U6044 ( .A1(n9372), .A2(n4450), .ZN(n4366) );
  NAND2_X1 U6045 ( .A1(n6024), .A2(n6023), .ZN(n8467) );
  INV_X1 U6046 ( .A(n5160), .ZN(n5103) );
  INV_X1 U6047 ( .A(n5220), .ZN(n5106) );
  OR2_X1 U6048 ( .A1(n9944), .A2(n7681), .ZN(n4367) );
  OAI21_X1 U6049 ( .B1(n5877), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U6050 ( .A1(n7802), .A2(n6184), .ZN(n7871) );
  NAND2_X1 U6051 ( .A1(n5796), .A2(n4599), .ZN(n7912) );
  INV_X1 U6052 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4397) );
  INV_X1 U6053 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5599) );
  AND2_X1 U6054 ( .A1(n8001), .A2(n8367), .ZN(n4368) );
  XNOR2_X1 U6055 ( .A(n6359), .B(n7973), .ZN(n7011) );
  OR2_X1 U6056 ( .A1(n9372), .A2(n9379), .ZN(n4369) );
  NOR2_X1 U6057 ( .A1(n5573), .A2(n9463), .ZN(n4370) );
  NOR2_X1 U6058 ( .A1(n8165), .A2(n4415), .ZN(n4371) );
  AND2_X1 U6059 ( .A1(n5099), .A2(n5046), .ZN(n5324) );
  AND2_X1 U6060 ( .A1(n5923), .A2(n5922), .ZN(n8354) );
  AND2_X1 U6061 ( .A1(n6271), .A2(n6270), .ZN(n4372) );
  AND2_X1 U6062 ( .A1(n8017), .A2(n8015), .ZN(n4373) );
  OR2_X1 U6063 ( .A1(n5809), .A2(n4396), .ZN(n4374) );
  AND2_X2 U6064 ( .A1(n5571), .A2(n6315), .ZN(n9914) );
  INV_X1 U6065 ( .A(n7511), .ZN(n4449) );
  AND2_X2 U6066 ( .A1(n6071), .A2(n6945), .ZN(n10130) );
  NAND2_X1 U6067 ( .A1(n5801), .A2(n5800), .ZN(n7929) );
  INV_X1 U6068 ( .A(n7929), .ZN(n4603) );
  INV_X1 U6069 ( .A(n8798), .ZN(n4724) );
  NAND2_X1 U6070 ( .A1(n7477), .A2(n5684), .ZN(n7372) );
  NAND2_X1 U6071 ( .A1(n4659), .A2(n4325), .ZN(n7916) );
  XNOR2_X1 U6072 ( .A(n6166), .B(n6167), .ZN(n7614) );
  NAND2_X1 U6073 ( .A1(n7461), .A2(n7460), .ZN(n7519) );
  OR2_X1 U6074 ( .A1(n7506), .A2(n7511), .ZN(n4375) );
  NAND2_X1 U6075 ( .A1(n5984), .A2(n5986), .ZN(n6068) );
  AND2_X1 U6076 ( .A1(n7293), .A2(n4830), .ZN(n4376) );
  OR2_X1 U6077 ( .A1(n9735), .A2(n6010), .ZN(n4377) );
  INV_X1 U6078 ( .A(n9906), .ZN(n9908) );
  AND2_X1 U6079 ( .A1(n7293), .A2(n6152), .ZN(n4378) );
  NAND2_X1 U6080 ( .A1(n5615), .A2(n4848), .ZN(n6002) );
  OR2_X1 U6081 ( .A1(n6867), .A2(n6868), .ZN(n6865) );
  INV_X1 U6082 ( .A(n6605), .ZN(n6593) );
  NAND2_X1 U6083 ( .A1(n6569), .A2(n7246), .ZN(n6605) );
  INV_X2 U6084 ( .A(n10117), .ZN(n10116) );
  AND2_X1 U6085 ( .A1(n6079), .A2(n6078), .ZN(n10117) );
  INV_X1 U6086 ( .A(n10033), .ZN(n8252) );
  NAND4_X1 U6087 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n6954)
         );
  INV_X1 U6088 ( .A(n6954), .ZN(n4561) );
  INV_X1 U6089 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U6090 ( .A1(n6803), .A2(n6004), .ZN(n10065) );
  AND2_X1 U6091 ( .A1(n4656), .A2(n6975), .ZN(n4379) );
  INV_X1 U6092 ( .A(n8887), .ZN(n9022) );
  AND2_X1 U6093 ( .A1(n4747), .A2(n4748), .ZN(n4380) );
  INV_X1 U6094 ( .A(n7049), .ZN(n4497) );
  NAND2_X1 U6095 ( .A1(n4739), .A2(n6769), .ZN(n4381) );
  INV_X1 U6096 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4388) );
  INV_X1 U6097 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U6098 ( .A1(n4747), .A2(n4746), .ZN(n4751) );
  OAI21_X1 U6099 ( .B1(n8681), .B2(n4840), .A(n8680), .ZN(n4839) );
  NOR2_X1 U6100 ( .A1(n4372), .A2(n4298), .ZN(n4436) );
  NAND2_X1 U6101 ( .A1(n6235), .A2(n6234), .ZN(n4840) );
  INV_X1 U6102 ( .A(n4595), .ZN(n4594) );
  NAND2_X1 U6103 ( .A1(n4788), .A2(n4952), .ZN(n5261) );
  OR2_X2 U6104 ( .A1(n8454), .A2(n5831), .ZN(n5833) );
  AOI21_X1 U6105 ( .B1(n8361), .B2(n8349), .A(n8350), .ZN(n8352) );
  OAI21_X1 U6106 ( .B1(n8296), .B2(n8295), .A(n8297), .ZN(n8303) );
  NOR2_X1 U6107 ( .A1(n5937), .A2(n4891), .ZN(n8318) );
  OAI22_X1 U6108 ( .A1(n8339), .A2(n5924), .B1(n8059), .B2(n8188), .ZN(n8327)
         );
  NAND2_X1 U6109 ( .A1(n4606), .A2(n4604), .ZN(n8361) );
  NAND2_X2 U6110 ( .A1(n4965), .A2(n4964), .ZN(n5303) );
  NAND2_X1 U6111 ( .A1(n4475), .A2(n8831), .ZN(n4474) );
  NAND3_X1 U6112 ( .A1(n4484), .A2(n4487), .A3(n4483), .ZN(n8883) );
  NAND2_X1 U6113 ( .A1(n4476), .A2(n4473), .ZN(n8840) );
  AOI21_X1 U6114 ( .B1(n4458), .B2(n8860), .A(n4457), .ZN(n8863) );
  INV_X1 U6115 ( .A(n4726), .ZN(n4725) );
  INV_X1 U6116 ( .A(n4501), .ZN(n4500) );
  XNOR2_X1 U6117 ( .A(n5631), .B(n5630), .ZN(n6762) );
  OR2_X1 U6118 ( .A1(n6415), .A2(n4517), .ZN(n4516) );
  OAI21_X1 U6119 ( .B1(n4524), .B2(n4519), .A(n6406), .ZN(n6410) );
  INV_X1 U6120 ( .A(n6400), .ZN(n4525) );
  OAI21_X1 U6121 ( .B1(n4923), .B2(n4388), .A(n4387), .ZN(n4915) );
  NAND3_X1 U6122 ( .A1(n4391), .A2(n4390), .A3(n9624), .ZN(n4389) );
  NAND3_X1 U6123 ( .A1(n4579), .A2(n5597), .A3(n4393), .ZN(n4392) );
  INV_X1 U6124 ( .A(n4394), .ZN(n7108) );
  NAND2_X1 U6125 ( .A1(n4850), .A2(n4394), .ZN(n7235) );
  NAND2_X1 U6126 ( .A1(n4394), .A2(n7148), .ZN(n7150) );
  INV_X1 U6127 ( .A(n4395), .ZN(n5877) );
  NOR2_X2 U6128 ( .A1(n7791), .A2(n7792), .ZN(n7848) );
  NAND2_X1 U6129 ( .A1(n8049), .A2(n4405), .ZN(n4404) );
  OAI21_X1 U6130 ( .B1(n8116), .B2(n4364), .A(n4872), .ZN(n8003) );
  AND2_X2 U6131 ( .A1(n4414), .A2(n4856), .ZN(n7844) );
  NAND2_X2 U6132 ( .A1(n6819), .A2(n4418), .ZN(n7236) );
  NOR2_X2 U6133 ( .A1(n5113), .A2(n4420), .ZN(n5099) );
  NAND4_X1 U6134 ( .A1(n5042), .A2(n5044), .A3(n5043), .A4(n5045), .ZN(n4420)
         );
  NAND4_X1 U6135 ( .A1(n5177), .A2(n5040), .A3(n5151), .A4(n5041), .ZN(n5113)
         );
  OR2_X2 U6136 ( .A1(n8659), .A2(n8658), .ZN(n4421) );
  NAND2_X1 U6137 ( .A1(n7614), .A2(n4425), .ZN(n4424) );
  NAND2_X1 U6138 ( .A1(n7615), .A2(n6169), .ZN(n7649) );
  NAND2_X1 U6139 ( .A1(n5498), .A2(n5497), .ZN(n5502) );
  NAND2_X1 U6140 ( .A1(n8665), .A2(n4437), .ZN(n4434) );
  AND2_X1 U6141 ( .A1(n9238), .A2(n4456), .ZN(n9190) );
  INV_X1 U6142 ( .A(n4766), .ZN(n4463) );
  OAI21_X1 U6143 ( .B1(n4463), .B2(n4462), .A(n4464), .ZN(n4466) );
  AND2_X1 U6144 ( .A1(n4766), .A2(n4306), .ZN(n9021) );
  AND2_X1 U6145 ( .A1(n4843), .A2(n5099), .ZN(n4467) );
  NAND4_X1 U6146 ( .A1(n4576), .A2(n5099), .A3(n4843), .A4(n5076), .ZN(n9555)
         );
  AND2_X2 U6147 ( .A1(n4576), .A2(n5099), .ZN(n5534) );
  NAND2_X1 U6148 ( .A1(n8866), .A2(n4363), .ZN(n4468) );
  OR2_X1 U6149 ( .A1(n8875), .A2(n4485), .ZN(n4483) );
  OR2_X1 U6150 ( .A1(n8874), .A2(n4489), .ZN(n4484) );
  MUX2_X1 U6151 ( .A(n6748), .B(P2_REG1_REG_2__SCAN_IN), .S(n6795), .Z(n6789)
         );
  NAND2_X1 U6152 ( .A1(n4505), .A2(n4929), .ZN(n4930) );
  XNOR2_X2 U6153 ( .A(n4505), .B(n4929), .ZN(n5186) );
  INV_X1 U6154 ( .A(n5153), .ZN(n4914) );
  NAND2_X1 U6155 ( .A1(n6415), .A2(n4510), .ZN(n4508) );
  NOR2_X1 U6156 ( .A1(n4525), .A2(n6605), .ZN(n4524) );
  NAND3_X1 U6157 ( .A1(n4528), .A2(n4527), .A3(n8350), .ZN(n4526) );
  AOI21_X2 U6158 ( .B1(n6490), .B2(n6605), .A(n4531), .ZN(n6505) );
  NAND2_X1 U6159 ( .A1(n4346), .A2(n6593), .ZN(n4532) );
  NAND2_X4 U6160 ( .A1(n5141), .A2(n5058), .ZN(n5155) );
  NAND2_X2 U6161 ( .A1(n9566), .A2(n5509), .ZN(n5141) );
  NAND2_X1 U6162 ( .A1(n9343), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U6163 ( .A1(n4550), .A2(n4548), .ZN(n5514) );
  INV_X1 U6164 ( .A(n8777), .ZN(n4553) );
  NAND2_X1 U6165 ( .A1(n4557), .A2(n4555), .ZN(n5519) );
  INV_X1 U6166 ( .A(n4556), .ZN(n4555) );
  NAND2_X1 U6167 ( .A1(n7357), .A2(n4558), .ZN(n4557) );
  INV_X1 U6168 ( .A(n9235), .ZN(n4571) );
  AND2_X1 U6169 ( .A1(n5052), .A2(n4578), .ZN(n4577) );
  NAND3_X1 U6170 ( .A1(n9624), .A2(n5631), .A3(n5596), .ZN(n5675) );
  NAND2_X1 U6171 ( .A1(n5833), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U6172 ( .A1(n4580), .A2(n4583), .ZN(n8412) );
  NAND2_X1 U6173 ( .A1(n4594), .A2(n4590), .ZN(n8454) );
  NAND2_X1 U6174 ( .A1(n8401), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U6175 ( .A1(n8308), .A2(n5960), .ZN(n4620) );
  NAND2_X1 U6176 ( .A1(n4620), .A2(n4316), .ZN(n8297) );
  AND2_X1 U6177 ( .A1(n4620), .A2(n4619), .ZN(n8296) );
  NAND2_X1 U6178 ( .A1(n8297), .A2(n5974), .ZN(n6586) );
  AND2_X2 U6179 ( .A1(n4629), .A2(n4626), .ZN(n7410) );
  AOI21_X1 U6180 ( .B1(n8367), .B2(n8575), .A(n8352), .ZN(n8339) );
  AOI21_X1 U6181 ( .B1(n8318), .B2(n5950), .A(n5949), .ZN(n8308) );
  OAI22_X1 U6182 ( .A1(n7422), .A2(n5667), .B1(n7974), .B2(n10072), .ZN(n7479)
         );
  NAND2_X1 U6183 ( .A1(n8410), .A2(n5876), .ZN(n8401) );
  NOR2_X1 U6184 ( .A1(n8327), .A2(n5936), .ZN(n5937) );
  NAND2_X1 U6185 ( .A1(n5764), .A2(n7675), .ZN(n7678) );
  NOR2_X2 U6186 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5040) );
  NAND2_X1 U6187 ( .A1(n9345), .A2(n9344), .ZN(n9343) );
  NAND2_X1 U6188 ( .A1(n5663), .A2(n6611), .ZN(n5633) );
  OAI21_X1 U6189 ( .B1(n9183), .B2(n5533), .A(n4691), .ZN(n5577) );
  OAI21_X2 U6190 ( .B1(n5186), .B2(n4931), .A(n4930), .ZN(n5200) );
  NOR2_X2 U6191 ( .A1(n9170), .A2(n9169), .ZN(n9168) );
  OR2_X1 U6192 ( .A1(n8324), .A2(n4643), .ZN(n4635) );
  NAND2_X1 U6193 ( .A1(n8324), .A2(n4639), .ZN(n4638) );
  NAND2_X1 U6194 ( .A1(n7587), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U6195 ( .A1(n6024), .A2(n4653), .ZN(n4652) );
  INV_X1 U6196 ( .A(n6014), .ZN(n6016) );
  CLKBUF_X1 U6197 ( .A(n6014), .Z(n4656) );
  NAND3_X1 U6198 ( .A1(n4658), .A2(n6016), .A3(n7008), .ZN(n4657) );
  NAND2_X1 U6199 ( .A1(n4662), .A2(n4360), .ZN(n6026) );
  NAND2_X1 U6200 ( .A1(n6025), .A2(n4660), .ZN(n4662) );
  NAND2_X1 U6201 ( .A1(n4664), .A2(n4663), .ZN(n7589) );
  NAND3_X1 U6202 ( .A1(n7474), .A2(n6392), .A3(n6367), .ZN(n4664) );
  INV_X1 U6203 ( .A(n7373), .ZN(n6521) );
  NAND2_X1 U6204 ( .A1(n7474), .A2(n6367), .ZN(n7369) );
  NAND2_X1 U6205 ( .A1(n4666), .A2(n4670), .ZN(n6602) );
  NAND3_X1 U6206 ( .A1(n4672), .A2(n4667), .A3(n4669), .ZN(n4666) );
  AND2_X1 U6207 ( .A1(n4672), .A2(n4669), .ZN(n8030) );
  NAND3_X1 U6208 ( .A1(n4675), .A2(n4676), .A3(n4880), .ZN(n5613) );
  AND3_X2 U6209 ( .A1(n4675), .A2(n4676), .A3(n4673), .ZN(n5614) );
  NAND2_X1 U6210 ( .A1(n6028), .A2(n4679), .ZN(n8333) );
  NAND2_X1 U6211 ( .A1(n8333), .A2(n6445), .ZN(n6029) );
  INV_X1 U6212 ( .A(n4680), .ZN(n7703) );
  NAND3_X1 U6213 ( .A1(n5186), .A2(n4930), .A3(n4934), .ZN(n4688) );
  INV_X1 U6214 ( .A(n5533), .ZN(n4690) );
  INV_X1 U6215 ( .A(n9298), .ZN(n4701) );
  INV_X1 U6216 ( .A(n8770), .ZN(n5058) );
  NAND2_X1 U6217 ( .A1(n7891), .A2(n4718), .ZN(n4716) );
  NAND2_X1 U6218 ( .A1(n4716), .A2(n4717), .ZN(n5351) );
  NAND2_X1 U6219 ( .A1(n9486), .A2(n8737), .ZN(n4723) );
  NAND2_X1 U6220 ( .A1(n8794), .A2(n7385), .ZN(n8798) );
  OAI211_X1 U6221 ( .C1(n8231), .C2(n4303), .A(n4727), .B(n4735), .ZN(n4726)
         );
  NAND2_X1 U6222 ( .A1(n8231), .A2(n4728), .ZN(n4727) );
  NAND2_X1 U6223 ( .A1(n4734), .A2(n4733), .ZN(n4729) );
  XNOR2_X1 U6224 ( .A(n8231), .B(n8256), .ZN(n8233) );
  INV_X1 U6225 ( .A(n4736), .ZN(n9942) );
  INV_X1 U6226 ( .A(n6766), .ZN(n4738) );
  NAND2_X1 U6227 ( .A1(n4738), .A2(n6757), .ZN(n4739) );
  NAND3_X1 U6228 ( .A1(n4739), .A2(n6769), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n6994) );
  NAND2_X1 U6229 ( .A1(n4381), .A2(n7432), .ZN(n6993) );
  NAND2_X1 U6230 ( .A1(n4751), .A2(n7161), .ZN(n7172) );
  NAND2_X1 U6231 ( .A1(n4767), .A2(n4769), .ZN(n4985) );
  NAND2_X1 U6232 ( .A1(n5303), .A2(n4771), .ZN(n4767) );
  NAND2_X1 U6233 ( .A1(n5303), .A2(n4781), .ZN(n4777) );
  NAND2_X1 U6234 ( .A1(n4948), .A2(n4362), .ZN(n4783) );
  NAND2_X1 U6235 ( .A1(n4783), .A2(n4784), .ZN(n5288) );
  NAND2_X1 U6236 ( .A1(n4948), .A2(n4947), .ZN(n5243) );
  NAND2_X1 U6237 ( .A1(n5004), .A2(n4795), .ZN(n4793) );
  NAND2_X1 U6238 ( .A1(n5004), .A2(n4798), .ZN(n4794) );
  NAND2_X1 U6239 ( .A1(n5004), .A2(n5003), .ZN(n5395) );
  OAI21_X1 U6240 ( .B1(n5353), .B2(n4803), .A(n4800), .ZN(n5383) );
  OR2_X1 U6241 ( .A1(n5353), .A2(n5352), .ZN(n4804) );
  NAND2_X1 U6242 ( .A1(n8868), .A2(n9025), .ZN(n4807) );
  OAI21_X1 U6243 ( .B1(n4293), .B2(n4810), .A(n4808), .ZN(n8694) );
  NAND2_X1 U6244 ( .A1(n7803), .A2(n4822), .ZN(n4819) );
  NAND2_X1 U6245 ( .A1(n4820), .A2(n4819), .ZN(n7942) );
  OAI211_X2 U6246 ( .C1(n7030), .C2(n4828), .A(n6137), .B(n4827), .ZN(n6141)
         );
  INV_X1 U6247 ( .A(n4825), .ZN(n4829) );
  NAND2_X1 U6248 ( .A1(n7023), .A2(n6132), .ZN(n7091) );
  NAND2_X1 U6249 ( .A1(n7030), .A2(n4829), .ZN(n7023) );
  NAND3_X1 U6250 ( .A1(n5040), .A2(n5151), .A3(n5177), .ZN(n5201) );
  NAND2_X1 U6251 ( .A1(n5534), .A2(n4845), .ZN(n5075) );
  NAND2_X1 U6252 ( .A1(n7235), .A2(n7234), .ZN(n7259) );
  NOR2_X1 U6253 ( .A1(n7151), .A2(n4851), .ZN(n4850) );
  INV_X1 U6254 ( .A(n8055), .ZN(n4855) );
  NAND2_X1 U6255 ( .A1(n4853), .A2(n4852), .ZN(n8078) );
  AOI21_X1 U6256 ( .B1(n8105), .B2(n8188), .A(n4854), .ZN(n4852) );
  NAND2_X1 U6257 ( .A1(n8164), .A2(n4373), .ZN(n8040) );
  OAI21_X1 U6258 ( .B1(n4923), .B2(n4910), .A(n4909), .ZN(n4911) );
  NAND2_X1 U6259 ( .A1(n4923), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4909) );
  XNOR2_X1 U6260 ( .A(n5446), .B(n5445), .ZN(n9572) );
  OAI21_X1 U6261 ( .B1(n5478), .B2(n5477), .A(n9187), .ZN(n9504) );
  NAND2_X1 U6262 ( .A1(n6505), .A2(n7247), .ZN(n6563) );
  XNOR2_X1 U6263 ( .A(n5480), .B(n5479), .ZN(n7963) );
  AND2_X1 U6264 ( .A1(n10114), .A2(n8292), .ZN(n6033) );
  XNOR2_X1 U6265 ( .A(n6032), .B(n6031), .ZN(n8292) );
  NAND2_X1 U6266 ( .A1(n6030), .A2(n6537), .ZN(n6032) );
  AOI21_X1 U6267 ( .B1(n8747), .B2(n4897), .A(n6307), .ZN(n6576) );
  CLKBUF_X1 U6268 ( .A(n8397), .Z(n8511) );
  NAND2_X1 U6269 ( .A1(n6575), .A2(n6319), .ZN(n6340) );
  NAND2_X2 U6270 ( .A1(n7591), .A2(n5737), .ZN(n7572) );
  MUX2_X2 U6271 ( .A(n6081), .B(n6080), .S(n10116), .Z(n6082) );
  MUX2_X2 U6272 ( .A(n9711), .B(n6080), .S(n10130), .Z(n6072) );
  OR2_X1 U6273 ( .A1(n6819), .A2(n6605), .ZN(n6567) );
  INV_X1 U6274 ( .A(n6978), .ZN(n6015) );
  INV_X1 U6275 ( .A(n5559), .ZN(n7957) );
  AND2_X1 U6276 ( .A1(n8226), .A2(n7701), .ZN(n7247) );
  AOI21_X1 U6277 ( .B1(n7259), .B2(n7258), .A(n7257), .ZN(n7261) );
  NAND2_X1 U6278 ( .A1(n5677), .A2(n6762), .ZN(n5632) );
  NAND2_X2 U6279 ( .A1(n6050), .A2(n6049), .ZN(n6821) );
  AOI21_X1 U6280 ( .B1(n6044), .B2(n6045), .A(n6066), .ZN(n6047) );
  NAND2_X2 U6281 ( .A1(n8621), .A2(n6218), .ZN(n8665) );
  NAND2_X1 U6282 ( .A1(n7980), .A2(n5609), .ZN(n5636) );
  NAND2_X1 U6283 ( .A1(n7980), .A2(n8607), .ZN(n5658) );
  INV_X1 U6284 ( .A(n6375), .ZN(n6019) );
  NOR2_X1 U6285 ( .A1(n5227), .A2(n7391), .ZN(n4884) );
  AND2_X1 U6286 ( .A1(n5674), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4885) );
  INV_X1 U6287 ( .A(n8320), .ZN(n8299) );
  AND2_X1 U6288 ( .A1(n5959), .A2(n5958), .ZN(n8320) );
  AND4_X1 U6289 ( .A1(n5848), .A2(n5847), .A3(n5600), .A4(n5599), .ZN(n4886)
         );
  NOR2_X1 U6290 ( .A1(n5573), .A2(n9534), .ZN(n5567) );
  NOR2_X1 U6291 ( .A1(n6538), .A2(n6537), .ZN(n4887) );
  OR2_X1 U6292 ( .A1(n8290), .A2(n8602), .ZN(n4888) );
  OR2_X1 U6293 ( .A1(n8033), .A2(n8543), .ZN(n4889) );
  OR2_X1 U6294 ( .A1(n8033), .A2(n8602), .ZN(n4890) );
  AND2_X1 U6295 ( .A1(n5935), .A2(n8187), .ZN(n4891) );
  OR2_X1 U6296 ( .A1(n8290), .A2(n8543), .ZN(n4892) );
  AND2_X1 U6297 ( .A1(n8290), .A2(n6584), .ZN(n4893) );
  INV_X1 U6298 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5579) );
  INV_X1 U6299 ( .A(n9186), .ZN(n5478) );
  OR2_X1 U6300 ( .A1(n7236), .A2(n7967), .ZN(n4894) );
  AND2_X1 U6301 ( .A1(n5934), .A2(n5933), .ZN(n8342) );
  INV_X1 U6302 ( .A(n8354), .ZN(n8188) );
  OR2_X1 U6303 ( .A1(n9435), .A2(n9291), .ZN(n4895) );
  OR2_X1 U6304 ( .A1(n6013), .A2(n6569), .ZN(n10101) );
  INV_X1 U6305 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4910) );
  AND2_X1 U6306 ( .A1(n4947), .A2(n4946), .ZN(n4896) );
  NAND2_X1 U6307 ( .A1(n6303), .A2(n6302), .ZN(n4897) );
  OR2_X1 U6308 ( .A1(n8830), .A2(n8673), .ZN(n4899) );
  AND2_X1 U6309 ( .A1(n8977), .A2(n8976), .ZN(n4900) );
  AND2_X1 U6310 ( .A1(n6562), .A2(n6561), .ZN(n4901) );
  AND4_X1 U6311 ( .A1(n9188), .A2(n9206), .A3(n9009), .A4(n9008), .ZN(n4902)
         );
  INV_X1 U6312 ( .A(n7588), .ZN(n5737) );
  AND2_X1 U6313 ( .A1(n7923), .A2(n8195), .ZN(n4903) );
  OAI21_X1 U6314 ( .B1(n7718), .B2(n6397), .A(n6382), .ZN(n7857) );
  INV_X1 U6315 ( .A(n9338), .ZN(n9468) );
  AND2_X1 U6316 ( .A1(n5571), .A2(n7132), .ZN(n9544) );
  INV_X1 U6317 ( .A(n9544), .ZN(n9906) );
  OR2_X1 U6318 ( .A1(n6549), .A2(n7782), .ZN(n6550) );
  OR2_X1 U6319 ( .A1(n6551), .A2(n6550), .ZN(n6555) );
  OR2_X1 U6320 ( .A1(n6551), .A2(n6533), .ZN(n6534) );
  NAND2_X1 U6321 ( .A1(n4898), .A2(n4886), .ZN(n5601) );
  INV_X1 U6322 ( .A(n8013), .ZN(n8014) );
  NAND2_X1 U6323 ( .A1(n6106), .A2(n7184), .ZN(n6088) );
  INV_X1 U6324 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5279) );
  INV_X1 U6325 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5120) );
  INV_X1 U6326 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5048) );
  INV_X1 U6327 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6328 ( .A1(n8014), .A2(n8320), .ZN(n8015) );
  INV_X1 U6329 ( .A(n5870), .ZN(n5590) );
  INV_X1 U6330 ( .A(n5908), .ZN(n5594) );
  INV_X1 U6331 ( .A(n8607), .ZN(n5609) );
  NAND2_X1 U6332 ( .A1(n8299), .A2(n8457), .ZN(n8300) );
  INV_X1 U6333 ( .A(n7918), .ZN(n6021) );
  INV_X1 U6334 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7316) );
  INV_X1 U6335 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5578) );
  INV_X1 U6336 ( .A(n10101), .ZN(n6599) );
  INV_X1 U6337 ( .A(n6083), .ZN(n7182) );
  INV_X1 U6338 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5046) );
  INV_X1 U6339 ( .A(SI_22_), .ZN(n5005) );
  INV_X1 U6340 ( .A(SI_14_), .ZN(n4967) );
  INV_X1 U6341 ( .A(n5663), .ZN(n5680) );
  INV_X1 U6342 ( .A(n8232), .ZN(n8256) );
  NAND2_X1 U6343 ( .A1(n5586), .A2(n5585), .ZN(n5825) );
  OR2_X1 U6344 ( .A1(n6074), .A2(n6820), .ZN(n6076) );
  OR2_X1 U6345 ( .A1(n6073), .A2(n6943), .ZN(n6840) );
  XNOR2_X1 U6346 ( .A(n6039), .B(n6038), .ZN(n6045) );
  NAND2_X1 U6347 ( .A1(n5071), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5410) );
  INV_X1 U6348 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5447) );
  OR2_X1 U6349 ( .A1(n7877), .A2(n9043), .ZN(n5272) );
  INV_X1 U6350 ( .A(n9190), .ZN(n9207) );
  INV_X1 U6351 ( .A(n9018), .ZN(n9014) );
  INV_X1 U6352 ( .A(n5563), .ZN(n9013) );
  INV_X1 U6353 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5076) );
  INV_X1 U6354 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U6355 ( .A1(n4981), .A2(n9603), .ZN(n4984) );
  AND2_X1 U6356 ( .A1(n5245), .A2(n5244), .ZN(n5248) );
  XNOR2_X1 U6357 ( .A(n10072), .B(n7236), .ZN(n7147) );
  AND2_X1 U6358 ( .A1(n7996), .A2(n8404), .ZN(n7997) );
  INV_X1 U6359 ( .A(n7843), .ZN(n6569) );
  AND2_X1 U6360 ( .A1(n6746), .A2(n8609), .ZN(n6803) );
  OR2_X1 U6361 ( .A1(n5977), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8031) );
  NOR2_X1 U6362 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND2_X1 U6363 ( .A1(n5941), .A2(n5940), .ZN(n5953) );
  OR2_X1 U6364 ( .A1(n6518), .A2(n6517), .ZN(n7935) );
  OR2_X1 U6365 ( .A1(n6821), .A2(n6054), .ZN(n6833) );
  INV_X1 U6366 ( .A(n8027), .ZN(n8290) );
  INV_X1 U6367 ( .A(n8458), .ZN(n7986) );
  INV_X1 U6368 ( .A(n8194), .ZN(n7983) );
  INV_X1 U6369 ( .A(n7424), .ZN(n7428) );
  NAND2_X1 U6370 ( .A1(n6042), .A2(n6035), .ZN(n6037) );
  AND2_X1 U6371 ( .A1(n9569), .A2(n5557), .ZN(n5558) );
  INV_X1 U6372 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9682) );
  OR2_X1 U6373 ( .A1(n6329), .A2(n9033), .ZN(n8705) );
  INV_X1 U6374 ( .A(n8759), .ZN(n8749) );
  OR2_X1 U6375 ( .A1(n9195), .A2(n5488), .ZN(n5476) );
  OR2_X1 U6376 ( .A1(n9776), .A2(n9775), .ZN(n9778) );
  INV_X1 U6377 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8671) );
  OR2_X1 U6378 ( .A1(n7839), .A2(n7779), .ZN(n5563) );
  OR2_X1 U6379 ( .A1(n9876), .A2(n7446), .ZN(n7196) );
  NAND2_X1 U6380 ( .A1(n9550), .A2(n6322), .ZN(n9374) );
  INV_X1 U6381 ( .A(n9188), .ZN(n5477) );
  INV_X1 U6382 ( .A(n9310), .ZN(n9452) );
  INV_X1 U6383 ( .A(n9473), .ZN(n8737) );
  OR2_X1 U6384 ( .A1(n7708), .A2(n9040), .ZN(n5320) );
  NAND2_X1 U6385 ( .A1(n7491), .A2(n7490), .ZN(n7489) );
  NAND2_X1 U6386 ( .A1(n9013), .A2(n6851), .ZN(n9261) );
  INV_X1 U6387 ( .A(n9895), .ZN(n7450) );
  AND2_X1 U6388 ( .A1(n5460), .A2(n5033), .ZN(n5445) );
  AND2_X1 U6389 ( .A1(n5020), .A2(n5019), .ZN(n5418) );
  AND2_X1 U6390 ( .A1(n4999), .A2(n4998), .ZN(n5369) );
  AND2_X1 U6391 ( .A1(n4984), .A2(n4983), .ZN(n5337) );
  XNOR2_X1 U6392 ( .A(n7147), .B(n8201), .ZN(n7110) );
  INV_X1 U6393 ( .A(n8158), .ZN(n8175) );
  INV_X1 U6394 ( .A(n8162), .ZN(n8169) );
  AND2_X1 U6395 ( .A1(n6503), .A2(n6001), .ZN(n8023) );
  AND4_X1 U6396 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n8427)
         );
  MUX2_X1 U6397 ( .A(n6742), .B(P2_U3893), .S(n6741), .Z(n10052) );
  AND2_X1 U6398 ( .A1(n6803), .A2(n8227), .ZN(n10061) );
  XNOR2_X1 U6399 ( .A(n6592), .B(n6591), .ZN(n8036) );
  AND2_X1 U6400 ( .A1(n6949), .A2(n8462), .ZN(n6946) );
  AND2_X1 U6401 ( .A1(n6823), .A2(n6593), .ZN(n8455) );
  INV_X1 U6402 ( .A(n8449), .ZN(n8393) );
  AND2_X1 U6403 ( .A1(n6833), .A2(n6070), .ZN(n6945) );
  INV_X1 U6404 ( .A(n10114), .ZN(n10106) );
  INV_X1 U6405 ( .A(n10095), .ZN(n10111) );
  OR2_X1 U6406 ( .A1(n7721), .A2(n6599), .ZN(n10114) );
  INV_X1 U6407 ( .A(n6843), .ZN(n6626) );
  AND2_X1 U6408 ( .A1(n6811), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8759) );
  INV_X1 U6409 ( .A(n8762), .ZN(n8751) );
  INV_X1 U6410 ( .A(n6086), .ZN(n9028) );
  INV_X1 U6411 ( .A(n5146), .ZN(n5530) );
  INV_X1 U6412 ( .A(n5331), .ZN(n5488) );
  INV_X1 U6413 ( .A(n9856), .ZN(n9839) );
  OR2_X1 U6414 ( .A1(n9849), .A2(n9848), .ZN(n9858) );
  INV_X1 U6415 ( .A(n7820), .ZN(n9358) );
  INV_X1 U6416 ( .A(n9261), .ZN(n9474) );
  INV_X1 U6417 ( .A(n9482), .ZN(n9258) );
  INV_X1 U6418 ( .A(n9869), .ZN(n9378) );
  INV_X1 U6419 ( .A(n9475), .ZN(n9262) );
  AND2_X1 U6420 ( .A1(n8851), .A2(n8950), .ZN(n9329) );
  AND2_X1 U6421 ( .A1(n7139), .A2(n9028), .ZN(n9427) );
  NAND2_X1 U6422 ( .A1(n7446), .A2(n7450), .ZN(n9905) );
  AND2_X1 U6423 ( .A1(n6316), .A2(n6603), .ZN(n9550) );
  AND2_X1 U6424 ( .A1(n5117), .A2(n5230), .ZN(n9136) );
  AND2_X1 U6425 ( .A1(n6610), .A2(n4288), .ZN(n9571) );
  AND2_X1 U6426 ( .A1(n6817), .A2(n6816), .ZN(n8162) );
  OR2_X1 U6427 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  INV_X1 U6428 ( .A(n8342), .ZN(n8187) );
  INV_X1 U6429 ( .A(n8441), .ZN(n8414) );
  INV_X1 U6430 ( .A(n7577), .ZN(n8197) );
  INV_X1 U6431 ( .A(n10061), .ZN(n9922) );
  NAND2_X1 U6432 ( .A1(n6951), .A2(n6950), .ZN(n8449) );
  INV_X1 U6433 ( .A(n8474), .ZN(n8447) );
  NAND2_X1 U6434 ( .A1(n10130), .A2(n10095), .ZN(n8543) );
  INV_X1 U6435 ( .A(n10130), .ZN(n10128) );
  OR2_X1 U6436 ( .A1(n10117), .A2(n10111), .ZN(n8602) );
  AND3_X1 U6437 ( .A1(n10089), .A2(n10088), .A3(n10087), .ZN(n10122) );
  INV_X1 U6438 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9639) );
  INV_X1 U6439 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7419) );
  INV_X1 U6440 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6707) );
  INV_X1 U6441 ( .A(n6581), .ZN(n6582) );
  INV_X1 U6442 ( .A(n9196), .ZN(n9392) );
  INV_X1 U6443 ( .A(n9308), .ZN(n9449) );
  INV_X1 U6444 ( .A(n8673), .ZN(n9039) );
  OR2_X1 U6445 ( .A1(n9769), .A2(n9032), .ZN(n9847) );
  INV_X1 U6446 ( .A(n9827), .ZN(n9862) );
  INV_X1 U6447 ( .A(n9873), .ZN(n9385) );
  AND2_X1 U6448 ( .A1(n7400), .A2(n7399), .ZN(n9898) );
  NOR2_X1 U6449 ( .A1(n4370), .A2(n5575), .ZN(n5576) );
  NAND2_X1 U6450 ( .A1(n9914), .A2(n9905), .ZN(n9491) );
  NOR2_X1 U6451 ( .A1(n5567), .A2(n5569), .ZN(n5570) );
  NAND2_X1 U6452 ( .A1(n9908), .A2(n9905), .ZN(n9548) );
  AND2_X1 U6453 ( .A1(n9898), .A2(n9897), .ZN(n9911) );
  NAND2_X1 U6454 ( .A1(n9551), .A2(n9550), .ZN(n9883) );
  INV_X1 U6455 ( .A(n5079), .ZN(n9563) );
  INV_X1 U6456 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7955) );
  INV_X1 U6457 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7717) );
  INV_X1 U6458 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7208) );
  INV_X1 U6459 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9684) );
  INV_X2 U6460 ( .A(n9736), .ZN(P2_U3893) );
  AND2_X2 U6461 ( .A1(n6604), .A2(n6603), .ZN(P1_U3973) );
  NAND2_X1 U6462 ( .A1(n7354), .A2(n4904), .ZN(n4905) );
  NAND2_X1 U6463 ( .A1(n4906), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U6464 ( .A1(n4911), .A2(SI_0_), .ZN(n5137) );
  NAND2_X1 U6465 ( .A1(n4912), .A2(SI_1_), .ZN(n4913) );
  OAI21_X2 U6466 ( .B1(n5138), .B2(n5137), .A(n4913), .ZN(n5154) );
  NAND2_X1 U6467 ( .A1(n5154), .A2(n4914), .ZN(n4917) );
  NAND2_X1 U6468 ( .A1(n4915), .A2(SI_2_), .ZN(n4916) );
  NAND2_X1 U6469 ( .A1(n4917), .A2(n4916), .ZN(n5169) );
  INV_X1 U6470 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6615) );
  INV_X1 U6471 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6614) );
  XNOR2_X1 U6472 ( .A(n4919), .B(SI_3_), .ZN(n5168) );
  NAND2_X1 U6473 ( .A1(n5169), .A2(n5168), .ZN(n4922) );
  INV_X1 U6474 ( .A(n4919), .ZN(n4920) );
  NAND2_X1 U6475 ( .A1(n4920), .A2(SI_3_), .ZN(n4921) );
  NAND2_X1 U6476 ( .A1(n4922), .A2(n4921), .ZN(n5181) );
  INV_X1 U6477 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4924) );
  CLKBUF_X3 U6478 ( .A(n4923), .Z(n6610) );
  MUX2_X1 U6479 ( .A(n4924), .B(n6619), .S(n6610), .Z(n4925) );
  XNOR2_X1 U6480 ( .A(n4925), .B(SI_4_), .ZN(n5180) );
  NAND2_X1 U6481 ( .A1(n5181), .A2(n5180), .ZN(n4928) );
  INV_X1 U6482 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6483 ( .A1(n4926), .A2(SI_4_), .ZN(n4927) );
  MUX2_X1 U6484 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8770), .Z(n4929) );
  INV_X1 U6485 ( .A(SI_5_), .ZN(n4931) );
  MUX2_X1 U6486 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6610), .Z(n4933) );
  XNOR2_X1 U6487 ( .A(n4933), .B(SI_6_), .ZN(n5199) );
  INV_X1 U6488 ( .A(n5199), .ZN(n4932) );
  NAND2_X1 U6489 ( .A1(n4933), .A2(SI_6_), .ZN(n4934) );
  MUX2_X1 U6490 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8770), .Z(n4936) );
  XNOR2_X1 U6491 ( .A(n4936), .B(SI_7_), .ZN(n5212) );
  INV_X1 U6492 ( .A(n5212), .ZN(n4935) );
  MUX2_X1 U6493 ( .A(n6663), .B(n9684), .S(n8770), .Z(n4938) );
  INV_X1 U6494 ( .A(SI_8_), .ZN(n4937) );
  NAND2_X1 U6495 ( .A1(n4938), .A2(n4937), .ZN(n4941) );
  INV_X1 U6496 ( .A(n4938), .ZN(n4939) );
  NAND2_X1 U6497 ( .A1(n4939), .A2(SI_8_), .ZN(n4940) );
  NAND2_X1 U6498 ( .A1(n4941), .A2(n4940), .ZN(n5111) );
  INV_X1 U6499 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4942) );
  MUX2_X1 U6500 ( .A(n6707), .B(n4942), .S(n8770), .Z(n4944) );
  INV_X1 U6501 ( .A(SI_9_), .ZN(n4943) );
  NAND2_X1 U6502 ( .A1(n4944), .A2(n4943), .ZN(n4947) );
  INV_X1 U6503 ( .A(n4944), .ZN(n4945) );
  NAND2_X1 U6504 ( .A1(n4945), .A2(SI_9_), .ZN(n4946) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4949) );
  MUX2_X1 U6506 ( .A(n6711), .B(n4949), .S(n6610), .Z(n4950) );
  XNOR2_X1 U6507 ( .A(n4950), .B(SI_10_), .ZN(n5242) );
  INV_X1 U6508 ( .A(n5242), .ZN(n4953) );
  INV_X1 U6509 ( .A(n4950), .ZN(n4951) );
  NAND2_X1 U6510 ( .A1(n4951), .A2(SI_10_), .ZN(n4952) );
  MUX2_X1 U6511 ( .A(n6798), .B(n4954), .S(n6610), .Z(n4956) );
  NAND2_X1 U6512 ( .A1(n4956), .A2(n4955), .ZN(n4959) );
  INV_X1 U6513 ( .A(n4956), .ZN(n4957) );
  NAND2_X1 U6514 ( .A1(n4957), .A2(SI_11_), .ZN(n4958) );
  NAND2_X1 U6515 ( .A1(n4959), .A2(n4958), .ZN(n5260) );
  MUX2_X1 U6516 ( .A(n6985), .B(n9669), .S(n6610), .Z(n4960) );
  XNOR2_X1 U6517 ( .A(n4960), .B(SI_12_), .ZN(n5273) );
  INV_X1 U6518 ( .A(n4960), .ZN(n4961) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8770), .Z(n4963) );
  XNOR2_X1 U6520 ( .A(n4963), .B(SI_13_), .ZN(n5287) );
  INV_X1 U6521 ( .A(n5287), .ZN(n4962) );
  NAND2_X1 U6522 ( .A1(n4963), .A2(SI_13_), .ZN(n4964) );
  MUX2_X1 U6523 ( .A(n7086), .B(n4966), .S(n8770), .Z(n4968) );
  INV_X1 U6524 ( .A(n4968), .ZN(n4969) );
  NAND2_X1 U6525 ( .A1(n4969), .A2(SI_14_), .ZN(n4970) );
  NAND2_X1 U6526 ( .A1(n4971), .A2(n4970), .ZN(n5302) );
  MUX2_X1 U6527 ( .A(n7206), .B(n7208), .S(n8770), .Z(n4972) );
  XNOR2_X1 U6528 ( .A(n4972), .B(SI_15_), .ZN(n5097) );
  INV_X1 U6529 ( .A(n5097), .ZN(n4975) );
  INV_X1 U6530 ( .A(n4972), .ZN(n4973) );
  NAND2_X1 U6531 ( .A1(n4973), .A2(SI_15_), .ZN(n4974) );
  MUX2_X1 U6532 ( .A(n7381), .B(n7383), .S(n6610), .Z(n4977) );
  NAND2_X1 U6533 ( .A1(n4977), .A2(n4976), .ZN(n4980) );
  INV_X1 U6534 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6535 ( .A1(n4978), .A2(SI_16_), .ZN(n4979) );
  NAND2_X1 U6536 ( .A1(n4980), .A2(n4979), .ZN(n5322) );
  MUX2_X1 U6537 ( .A(n7419), .B(n7421), .S(n8770), .Z(n4981) );
  INV_X1 U6538 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6539 ( .A1(n4982), .A2(SI_17_), .ZN(n4983) );
  MUX2_X1 U6540 ( .A(n7528), .B(n7530), .S(n6610), .Z(n4986) );
  XNOR2_X1 U6541 ( .A(n4986), .B(SI_18_), .ZN(n5090) );
  INV_X1 U6542 ( .A(n5090), .ZN(n4989) );
  INV_X1 U6543 ( .A(n4986), .ZN(n4987) );
  NAND2_X1 U6544 ( .A1(n4987), .A2(SI_18_), .ZN(n4988) );
  MUX2_X1 U6545 ( .A(n7626), .B(n7966), .S(n8770), .Z(n4991) );
  INV_X1 U6546 ( .A(SI_19_), .ZN(n4990) );
  NAND2_X1 U6547 ( .A1(n4991), .A2(n4990), .ZN(n4994) );
  INV_X1 U6548 ( .A(n4991), .ZN(n4992) );
  NAND2_X1 U6549 ( .A1(n4992), .A2(SI_19_), .ZN(n4993) );
  NAND2_X1 U6550 ( .A1(n4994), .A2(n4993), .ZN(n5352) );
  MUX2_X1 U6551 ( .A(n7700), .B(n7717), .S(n6610), .Z(n4996) );
  INV_X1 U6552 ( .A(SI_20_), .ZN(n4995) );
  NAND2_X1 U6553 ( .A1(n4996), .A2(n4995), .ZN(n4999) );
  INV_X1 U6554 ( .A(n4996), .ZN(n4997) );
  NAND2_X1 U6555 ( .A1(n4997), .A2(SI_20_), .ZN(n4998) );
  INV_X1 U6556 ( .A(n5383), .ZN(n5000) );
  MUX2_X1 U6557 ( .A(n7780), .B(n7778), .S(n8770), .Z(n5001) );
  XNOR2_X1 U6558 ( .A(n5001), .B(SI_21_), .ZN(n5382) );
  NAND2_X1 U6559 ( .A1(n5000), .A2(n5382), .ZN(n5004) );
  INV_X1 U6560 ( .A(n5001), .ZN(n5002) );
  NAND2_X1 U6561 ( .A1(n5002), .A2(SI_21_), .ZN(n5003) );
  MUX2_X1 U6562 ( .A(n7841), .B(n7840), .S(n6610), .Z(n5006) );
  NAND2_X1 U6563 ( .A1(n5006), .A2(n5005), .ZN(n5009) );
  INV_X1 U6564 ( .A(n5006), .ZN(n5007) );
  NAND2_X1 U6565 ( .A1(n5007), .A2(SI_22_), .ZN(n5008) );
  NAND2_X1 U6566 ( .A1(n5009), .A2(n5008), .ZN(n5394) );
  INV_X1 U6567 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5010) );
  MUX2_X1 U6568 ( .A(n5010), .B(n7952), .S(n8770), .Z(n5012) );
  INV_X1 U6569 ( .A(SI_23_), .ZN(n5011) );
  NAND2_X1 U6570 ( .A1(n5012), .A2(n5011), .ZN(n5015) );
  INV_X1 U6571 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6572 ( .A1(n5013), .A2(SI_23_), .ZN(n5014) );
  MUX2_X1 U6573 ( .A(n9639), .B(n7955), .S(n6610), .Z(n5017) );
  INV_X1 U6574 ( .A(SI_24_), .ZN(n5016) );
  NAND2_X1 U6575 ( .A1(n5017), .A2(n5016), .ZN(n5020) );
  INV_X1 U6576 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6577 ( .A1(n5018), .A2(SI_24_), .ZN(n5019) );
  NAND2_X1 U6578 ( .A1(n5419), .A2(n5418), .ZN(n5021) );
  NAND2_X1 U6579 ( .A1(n5021), .A2(n5020), .ZN(n5433) );
  INV_X1 U6580 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5022) );
  INV_X1 U6581 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9605) );
  MUX2_X1 U6582 ( .A(n5022), .B(n9605), .S(n8770), .Z(n5024) );
  INV_X1 U6583 ( .A(SI_25_), .ZN(n5023) );
  NAND2_X1 U6584 ( .A1(n5024), .A2(n5023), .ZN(n5027) );
  INV_X1 U6585 ( .A(n5024), .ZN(n5025) );
  NAND2_X1 U6586 ( .A1(n5025), .A2(SI_25_), .ZN(n5026) );
  NAND2_X1 U6587 ( .A1(n5433), .A2(n5432), .ZN(n5028) );
  NAND2_X1 U6588 ( .A1(n5028), .A2(n5027), .ZN(n5446) );
  INV_X1 U6589 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5029) );
  MUX2_X1 U6590 ( .A(n5029), .B(n5447), .S(n8770), .Z(n5031) );
  INV_X1 U6591 ( .A(SI_26_), .ZN(n5030) );
  NAND2_X1 U6592 ( .A1(n5031), .A2(n5030), .ZN(n5460) );
  INV_X1 U6593 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6594 ( .A1(n5032), .A2(SI_26_), .ZN(n5033) );
  NAND2_X1 U6595 ( .A1(n5446), .A2(n5445), .ZN(n5464) );
  NAND2_X1 U6596 ( .A1(n5464), .A2(n5460), .ZN(n5039) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5034) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9567) );
  MUX2_X1 U6599 ( .A(n5034), .B(n9567), .S(n6610), .Z(n5036) );
  INV_X1 U6600 ( .A(SI_27_), .ZN(n5035) );
  NAND2_X1 U6601 ( .A1(n5036), .A2(n5035), .ZN(n5459) );
  INV_X1 U6602 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6603 ( .A1(n5037), .A2(SI_27_), .ZN(n5461) );
  AND2_X1 U6604 ( .A1(n5459), .A2(n5461), .ZN(n5038) );
  NOR2_X2 U6605 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5151) );
  NOR2_X1 U6606 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5045) );
  NOR2_X1 U6607 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5044) );
  NOR2_X1 U6608 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5043) );
  NOR2_X1 U6609 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5042) );
  NOR2_X1 U6610 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5047) );
  NAND4_X1 U6611 ( .A1(n5047), .A2(n5092), .A3(n5496), .A4(n5561), .ZN(n5051)
         );
  NAND4_X1 U6612 ( .A1(n5049), .A2(n5495), .A3(n5494), .A4(n5048), .ZN(n5050)
         );
  NOR2_X1 U6613 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  XNOR2_X2 U6614 ( .A(n5055), .B(n5054), .ZN(n5509) );
  NAND2_X1 U6615 ( .A1(n8612), .A2(n8878), .ZN(n5060) );
  OR2_X1 U6616 ( .A1(n5155), .A2(n9567), .ZN(n5059) );
  NAND2_X1 U6617 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5192) );
  INV_X1 U6618 ( .A(n5192), .ZN(n5061) );
  NAND2_X1 U6619 ( .A1(n5061), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5206) );
  INV_X1 U6620 ( .A(n5206), .ZN(n5062) );
  NAND2_X1 U6621 ( .A1(n5062), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5217) );
  INV_X1 U6622 ( .A(n5217), .ZN(n5063) );
  NAND2_X1 U6623 ( .A1(n5063), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5219) );
  INV_X1 U6624 ( .A(n5235), .ZN(n5064) );
  NAND2_X1 U6625 ( .A1(n5064), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5253) );
  INV_X1 U6626 ( .A(n5314), .ZN(n5067) );
  INV_X1 U6627 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5086) );
  INV_X1 U6628 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8704) );
  INV_X1 U6629 ( .A(n5398), .ZN(n5071) );
  INV_X1 U6630 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5422) );
  INV_X1 U6631 ( .A(n5436), .ZN(n5072) );
  NAND2_X1 U6632 ( .A1(n5072), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5451) );
  INV_X1 U6633 ( .A(n5451), .ZN(n5073) );
  NAND2_X1 U6634 ( .A1(n5073), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5453) );
  INV_X1 U6635 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U6636 ( .A1(n5453), .A2(n6577), .ZN(n5074) );
  AND2_X2 U6637 ( .A1(n5080), .A2(n5079), .ZN(n5315) );
  NAND2_X1 U6638 ( .A1(n9209), .A2(n5331), .ZN(n5085) );
  INV_X1 U6639 ( .A(n5080), .ZN(n9559) );
  INV_X1 U6640 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9406) );
  AND2_X2 U6641 ( .A1(n9559), .A2(n9563), .ZN(n5160) );
  NAND2_X1 U6642 ( .A1(n5160), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6643 ( .A1(n5527), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5081) );
  OAI211_X1 U6644 ( .C1(n5530), .C2(n9406), .A(n5082), .B(n5081), .ZN(n5083)
         );
  INV_X1 U6645 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6646 ( .A1(n5345), .A2(n5086), .ZN(n5087) );
  NAND2_X1 U6647 ( .A1(n5362), .A2(n5087), .ZN(n9350) );
  AOI22_X1 U6648 ( .A1(n5146), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5160), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5089) );
  INV_X2 U6649 ( .A(n5106), .ZN(n5527) );
  NAND2_X1 U6650 ( .A1(n5527), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5088) );
  OAI211_X1 U6651 ( .C1(n9350), .C2(n5488), .A(n5089), .B(n5088), .ZN(n9464)
         );
  INV_X1 U6652 ( .A(n9464), .ZN(n8685) );
  XNOR2_X1 U6653 ( .A(n5091), .B(n5090), .ZN(n7527) );
  NAND2_X1 U6654 ( .A1(n7527), .A2(n8878), .ZN(n5096) );
  BUF_X2 U6655 ( .A(n5141), .Z(n8772) );
  INV_X1 U6656 ( .A(n5498), .ZN(n5093) );
  NAND2_X1 U6657 ( .A1(n5339), .A2(n5495), .ZN(n5094) );
  NAND2_X1 U6658 ( .A1(n5094), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5354) );
  XNOR2_X1 U6659 ( .A(n5354), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7761) );
  AOI22_X1 U6660 ( .A1(n5358), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5357), .B2(
        n7761), .ZN(n5095) );
  INV_X1 U6661 ( .A(n9347), .ZN(n9478) );
  XNOR2_X1 U6662 ( .A(n5098), .B(n5097), .ZN(n7205) );
  NAND2_X1 U6663 ( .A1(n7205), .A2(n8878), .ZN(n5102) );
  OR2_X1 U6664 ( .A1(n5099), .A2(n9554), .ZN(n5100) );
  XNOR2_X1 U6665 ( .A(n5100), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U6666 ( .A1(n5358), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5357), .B2(
        n9818), .ZN(n5101) );
  NAND2_X1 U6667 ( .A1(n6642), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6668 ( .A1(n5146), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5109) );
  INV_X1 U6669 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6670 ( .A1(n5314), .A2(n5104), .ZN(n5105) );
  AND2_X1 U6671 ( .A1(n5329), .A2(n5105), .ZN(n8758) );
  NAND2_X1 U6672 ( .A1(n5315), .A2(n8758), .ZN(n5108) );
  NAND2_X1 U6673 ( .A1(n5527), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5107) );
  NOR2_X1 U6674 ( .A1(n5113), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5245) );
  NOR2_X1 U6675 ( .A1(n5245), .A2(n9554), .ZN(n5114) );
  NAND2_X1 U6676 ( .A1(n5114), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5117) );
  INV_X1 U6677 ( .A(n5114), .ZN(n5116) );
  INV_X1 U6678 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6679 ( .A1(n5116), .A2(n5115), .ZN(n5230) );
  AOI22_X1 U6680 ( .A1(n5358), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5357), .B2(
        n9136), .ZN(n5118) );
  NAND2_X1 U6681 ( .A1(n5146), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6682 ( .A1(n6642), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6683 ( .A1(n5219), .A2(n5120), .ZN(n5121) );
  AND2_X1 U6684 ( .A1(n5235), .A2(n5121), .ZN(n7618) );
  NAND2_X1 U6685 ( .A1(n5331), .A2(n7618), .ZN(n5123) );
  NAND2_X1 U6686 ( .A1(n5527), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5122) );
  INV_X1 U6687 ( .A(n7654), .ZN(n9046) );
  NAND2_X1 U6688 ( .A1(n5315), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6689 ( .A1(n5160), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6690 ( .A1(n5220), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5127) );
  INV_X1 U6691 ( .A(SI_0_), .ZN(n5130) );
  NOR2_X1 U6692 ( .A1(n5058), .A2(n5130), .ZN(n5132) );
  INV_X1 U6693 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5131) );
  XNOR2_X1 U6694 ( .A(n5132), .B(n5131), .ZN(n9727) );
  MUX2_X1 U6695 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9727), .S(n8772), .Z(n6810) );
  NAND2_X1 U6696 ( .A1(n6954), .A2(n6810), .ZN(n6883) );
  NAND2_X1 U6697 ( .A1(n5315), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6698 ( .A1(n5220), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5135) );
  XNOR2_X1 U6699 ( .A(n5138), .B(n5137), .ZN(n6611) );
  OR2_X1 U6700 ( .A1(n5182), .A2(n6611), .ZN(n5144) );
  INV_X1 U6701 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6702 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5139) );
  XNOR2_X1 U6703 ( .A(n5140), .B(n5139), .ZN(n6685) );
  OR2_X1 U6704 ( .A1(n5141), .A2(n6685), .ZN(n5142) );
  AND3_X4 U6705 ( .A1(n5144), .A2(n5143), .A3(n5142), .ZN(n8909) );
  NAND2_X1 U6706 ( .A1(n6883), .A2(n6884), .ZN(n6882) );
  INV_X1 U6707 ( .A(n9053), .ZN(n6956) );
  NAND2_X1 U6708 ( .A1(n6956), .A2(n8909), .ZN(n5145) );
  NAND2_X1 U6709 ( .A1(n6882), .A2(n5145), .ZN(n6900) );
  NAND2_X1 U6710 ( .A1(n5315), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6711 ( .A1(n5220), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6712 ( .A1(n5146), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5148) );
  OR2_X1 U6713 ( .A1(n5151), .A2(n9554), .ZN(n5179) );
  INV_X1 U6714 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6715 ( .A1(n5179), .A2(n5152), .ZN(n5165) );
  OAI21_X1 U6716 ( .B1(n5179), .B2(n5152), .A(n5165), .ZN(n6684) );
  XNOR2_X1 U6717 ( .A(n5154), .B(n5153), .ZN(n5651) );
  INV_X1 U6718 ( .A(n5651), .ZN(n6612) );
  OR2_X1 U6719 ( .A1(n5182), .A2(n6612), .ZN(n5157) );
  INV_X1 U6720 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6613) );
  OR2_X1 U6721 ( .A1(n5155), .A2(n6613), .ZN(n5156) );
  NAND2_X1 U6722 ( .A1(n7033), .A2(n7213), .ZN(n5511) );
  INV_X1 U6723 ( .A(n7033), .ZN(n9052) );
  NAND2_X1 U6724 ( .A1(n9052), .A2(n6904), .ZN(n8912) );
  NAND2_X1 U6725 ( .A1(n5511), .A2(n8912), .ZN(n8980) );
  NAND2_X1 U6726 ( .A1(n6900), .A2(n8980), .ZN(n6899) );
  NAND2_X1 U6727 ( .A1(n7033), .A2(n6904), .ZN(n5158) );
  NAND2_X1 U6728 ( .A1(n6899), .A2(n5158), .ZN(n6912) );
  INV_X1 U6729 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6730 ( .A1(n5331), .A2(n5159), .ZN(n5164) );
  NAND2_X1 U6731 ( .A1(n5146), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6732 ( .A1(n5220), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6733 ( .A1(n5160), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6734 ( .A1(n5165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5167) );
  INV_X1 U6735 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6736 ( .A(n5167), .B(n5166), .ZN(n6688) );
  XNOR2_X1 U6737 ( .A(n5169), .B(n5168), .ZN(n6616) );
  OR2_X1 U6738 ( .A1(n5182), .A2(n6616), .ZN(n5171) );
  OR2_X1 U6739 ( .A1(n5155), .A2(n6614), .ZN(n5170) );
  OAI211_X1 U6740 ( .C1(n8772), .C2(n6688), .A(n5171), .B(n5170), .ZN(n7328)
         );
  NAND2_X1 U6741 ( .A1(n6907), .A2(n7328), .ZN(n8777) );
  INV_X1 U6742 ( .A(n6907), .ZN(n9051) );
  NAND2_X1 U6743 ( .A1(n9051), .A2(n7126), .ZN(n8913) );
  NAND2_X1 U6744 ( .A1(n8777), .A2(n8913), .ZN(n6911) );
  NAND2_X1 U6745 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U6746 ( .A1(n6907), .A2(n7126), .ZN(n5172) );
  NAND2_X1 U6747 ( .A1(n6910), .A2(n5172), .ZN(n6967) );
  NAND2_X1 U6748 ( .A1(n5146), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6749 ( .A1(n6642), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5175) );
  OAI21_X1 U6750 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5192), .ZN(n7222) );
  INV_X1 U6751 ( .A(n7222), .ZN(n7027) );
  NAND2_X1 U6752 ( .A1(n5315), .A2(n7027), .ZN(n5174) );
  NAND2_X1 U6753 ( .A1(n5527), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5173) );
  OR2_X1 U6754 ( .A1(n5177), .A2(n9554), .ZN(n5178) );
  NAND2_X1 U6755 ( .A1(n5179), .A2(n5178), .ZN(n5187) );
  XNOR2_X1 U6756 ( .A(n5187), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6690) );
  XNOR2_X1 U6757 ( .A(n5181), .B(n5180), .ZN(n6618) );
  OR2_X1 U6758 ( .A1(n5182), .A2(n6618), .ZN(n5184) );
  OR2_X1 U6759 ( .A1(n5155), .A2(n6619), .ZN(n5183) );
  OAI211_X1 U6760 ( .C1(n6690), .C2(n8772), .A(n5184), .B(n5183), .ZN(n6963)
         );
  NAND2_X1 U6761 ( .A1(n7331), .A2(n6963), .ZN(n8784) );
  INV_X1 U6762 ( .A(n6963), .ZN(n7226) );
  NAND2_X1 U6763 ( .A1(n9050), .A2(n7226), .ZN(n7281) );
  NAND2_X1 U6764 ( .A1(n8784), .A2(n7281), .ZN(n8985) );
  NAND2_X1 U6765 ( .A1(n6967), .A2(n8985), .ZN(n6966) );
  NAND2_X1 U6766 ( .A1(n7331), .A2(n7226), .ZN(n5185) );
  NAND2_X1 U6767 ( .A1(n6966), .A2(n5185), .ZN(n7277) );
  XNOR2_X1 U6768 ( .A(n5186), .B(SI_5_), .ZN(n6620) );
  NAND2_X1 U6769 ( .A1(n6620), .A2(n8878), .ZN(n5190) );
  OAI21_X1 U6770 ( .B1(n5187), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5188) );
  XNOR2_X1 U6771 ( .A(n5188), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9097) );
  AOI22_X1 U6772 ( .A1(n5358), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5357), .B2(
        n9097), .ZN(n5189) );
  NAND2_X1 U6773 ( .A1(n6642), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5197) );
  INV_X1 U6774 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6775 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  AND2_X1 U6776 ( .A1(n5206), .A2(n5193), .ZN(n9866) );
  NAND2_X1 U6777 ( .A1(n5331), .A2(n9866), .ZN(n5196) );
  NAND2_X1 U6778 ( .A1(n5527), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6779 ( .A1(n5146), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5194) );
  NAND4_X1 U6780 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n9049)
         );
  NAND2_X1 U6781 ( .A1(n9870), .A2(n9049), .ZN(n8917) );
  INV_X1 U6782 ( .A(n9049), .ZN(n7298) );
  NAND2_X1 U6783 ( .A1(n7298), .A2(n7280), .ZN(n8785) );
  NAND2_X1 U6784 ( .A1(n8917), .A2(n8785), .ZN(n8986) );
  NAND2_X1 U6785 ( .A1(n7277), .A2(n8986), .ZN(n7276) );
  NAND2_X1 U6786 ( .A1(n9870), .A2(n7298), .ZN(n5198) );
  XNOR2_X1 U6787 ( .A(n5200), .B(n5199), .ZN(n6635) );
  NAND2_X1 U6788 ( .A1(n6635), .A2(n8878), .ZN(n5204) );
  NAND2_X1 U6789 ( .A1(n5201), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5202) );
  XNOR2_X1 U6790 ( .A(n5202), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9110) );
  AOI22_X1 U6791 ( .A1(n5358), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5357), .B2(
        n9110), .ZN(n5203) );
  NAND2_X1 U6792 ( .A1(n5204), .A2(n5203), .ZN(n7302) );
  NAND2_X1 U6793 ( .A1(n6642), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6794 ( .A1(n5146), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5210) );
  INV_X1 U6795 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6796 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  AND2_X1 U6797 ( .A1(n5217), .A2(n5207), .ZN(n7297) );
  NAND2_X1 U6798 ( .A1(n5315), .A2(n7297), .ZN(n5209) );
  NAND2_X1 U6799 ( .A1(n5527), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5208) );
  OR2_X1 U6800 ( .A1(n7302), .A2(n7442), .ZN(n8788) );
  NAND2_X1 U6801 ( .A1(n7302), .A2(n7442), .ZN(n8920) );
  NAND2_X1 U6802 ( .A1(n8788), .A2(n8920), .ZN(n7194) );
  NAND2_X1 U6803 ( .A1(n7613), .A2(n7654), .ZN(n8800) );
  NAND2_X1 U6804 ( .A1(n8795), .A2(n8800), .ZN(n7394) );
  NAND2_X1 U6805 ( .A1(n6640), .A2(n8878), .ZN(n5215) );
  NAND2_X1 U6806 ( .A1(n5113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U6807 ( .A(n5213), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9123) );
  AOI22_X1 U6808 ( .A1(n5358), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5357), .B2(
        n9123), .ZN(n5214) );
  NAND2_X2 U6809 ( .A1(n5215), .A2(n5214), .ZN(n7562) );
  NAND2_X1 U6810 ( .A1(n5146), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6811 ( .A1(n6642), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5223) );
  INV_X1 U6812 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6813 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  AND2_X1 U6814 ( .A1(n5219), .A2(n5218), .ZN(n7561) );
  NAND2_X1 U6815 ( .A1(n5331), .A2(n7561), .ZN(n5222) );
  NAND2_X1 U6816 ( .A1(n5220), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5221) );
  INV_X1 U6817 ( .A(n7619), .ZN(n9047) );
  OR2_X1 U6818 ( .A1(n7562), .A2(n9047), .ZN(n5226) );
  NAND2_X1 U6819 ( .A1(n7562), .A2(n7619), .ZN(n7385) );
  INV_X1 U6820 ( .A(n7442), .ZN(n9048) );
  OR2_X1 U6821 ( .A1(n7302), .A2(n9048), .ZN(n7435) );
  AND2_X1 U6822 ( .A1(n7435), .A2(n5226), .ZN(n7391) );
  OAI21_X1 U6823 ( .B1(n7613), .B2(n9046), .A(n7397), .ZN(n7503) );
  NAND2_X1 U6824 ( .A1(n5230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6825 ( .A(n5231), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7749) );
  AOI22_X1 U6826 ( .A1(n5358), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5357), .B2(
        n7749), .ZN(n5232) );
  NAND2_X1 U6827 ( .A1(n5146), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6828 ( .A1(n6642), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5239) );
  INV_X1 U6829 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6830 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  AND2_X1 U6831 ( .A1(n5253), .A2(n5236), .ZN(n7652) );
  NAND2_X1 U6832 ( .A1(n5331), .A2(n7652), .ZN(n5238) );
  NAND2_X1 U6833 ( .A1(n5527), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6834 ( .A1(n7511), .A2(n7547), .ZN(n8991) );
  NAND2_X1 U6835 ( .A1(n8810), .A2(n8991), .ZN(n7505) );
  NAND2_X1 U6836 ( .A1(n7503), .A2(n7505), .ZN(n7504) );
  INV_X1 U6837 ( .A(n7547), .ZN(n9045) );
  NAND2_X1 U6838 ( .A1(n7504), .A2(n5241), .ZN(n7361) );
  XNOR2_X1 U6839 ( .A(n5243), .B(n5242), .ZN(n6709) );
  NAND2_X1 U6840 ( .A1(n6709), .A2(n8878), .ZN(n5251) );
  NOR2_X1 U6841 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5244) );
  NOR2_X1 U6842 ( .A1(n5248), .A2(n9554), .ZN(n5246) );
  MUX2_X1 U6843 ( .A(n9554), .B(n5246), .S(P1_IR_REG_10__SCAN_IN), .Z(n5249)
         );
  INV_X1 U6844 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5247) );
  NOR2_X1 U6845 ( .A1(n5249), .A2(n5276), .ZN(n9761) );
  AOI22_X1 U6846 ( .A1(n5358), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5357), .B2(
        n9761), .ZN(n5250) );
  NAND2_X1 U6847 ( .A1(n5146), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6848 ( .A1(n6642), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6849 ( .A1(n5253), .A2(n5252), .ZN(n5254) );
  AND2_X1 U6850 ( .A1(n5266), .A2(n5254), .ZN(n7806) );
  NAND2_X1 U6851 ( .A1(n5315), .A2(n7806), .ZN(n5256) );
  NAND2_X1 U6852 ( .A1(n5527), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5255) );
  OR2_X1 U6853 ( .A1(n7557), .A2(n7656), .ZN(n8814) );
  NAND2_X1 U6854 ( .A1(n7557), .A2(n7656), .ZN(n8812) );
  NAND2_X1 U6855 ( .A1(n8814), .A2(n8812), .ZN(n8994) );
  NAND2_X1 U6856 ( .A1(n7361), .A2(n8994), .ZN(n7360) );
  INV_X1 U6857 ( .A(n7656), .ZN(n9044) );
  NAND2_X1 U6858 ( .A1(n7360), .A2(n5259), .ZN(n7491) );
  XNOR2_X1 U6859 ( .A(n5261), .B(n5260), .ZN(n6713) );
  NAND2_X1 U6860 ( .A1(n6713), .A2(n8878), .ZN(n5264) );
  OR2_X1 U6861 ( .A1(n5276), .A2(n9554), .ZN(n5262) );
  XNOR2_X1 U6862 ( .A(n5262), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9149) );
  AOI22_X1 U6863 ( .A1(n5358), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5357), .B2(
        n9149), .ZN(n5263) );
  NAND2_X1 U6864 ( .A1(n6642), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6865 ( .A1(n5146), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5270) );
  INV_X1 U6866 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6867 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  AND2_X1 U6868 ( .A1(n5280), .A2(n5267), .ZN(n7873) );
  NAND2_X1 U6869 ( .A1(n5331), .A2(n7873), .ZN(n5269) );
  NAND2_X1 U6870 ( .A1(n5527), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5268) );
  OR2_X1 U6871 ( .A1(n7877), .A2(n7807), .ZN(n8815) );
  NAND2_X1 U6872 ( .A1(n7877), .A2(n7807), .ZN(n8817) );
  NAND2_X1 U6873 ( .A1(n8815), .A2(n8817), .ZN(n7490) );
  INV_X1 U6874 ( .A(n7807), .ZN(n9043) );
  NAND2_X1 U6875 ( .A1(n7489), .A2(n5272), .ZN(n7603) );
  XNOR2_X1 U6876 ( .A(n5274), .B(n5273), .ZN(n6984) );
  NAND2_X1 U6877 ( .A1(n6984), .A2(n8878), .ZN(n5278) );
  INV_X1 U6878 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6879 ( .A1(n5276), .A2(n5275), .ZN(n5307) );
  NAND2_X1 U6880 ( .A1(n5307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6881 ( .A(n5289), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7756) );
  AOI22_X1 U6882 ( .A1(n5358), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5357), .B2(
        n7756), .ZN(n5277) );
  NAND2_X1 U6883 ( .A1(n6642), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6884 ( .A1(n5527), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6885 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  AND2_X1 U6886 ( .A1(n5295), .A2(n5281), .ZN(n7944) );
  NAND2_X1 U6887 ( .A1(n5315), .A2(n7944), .ZN(n5283) );
  NAND2_X1 U6888 ( .A1(n5146), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5282) );
  OR2_X1 U6889 ( .A1(n7947), .A2(n7875), .ZN(n8819) );
  NAND2_X1 U6890 ( .A1(n7947), .A2(n7875), .ZN(n8928) );
  NAND2_X1 U6891 ( .A1(n8819), .A2(n8928), .ZN(n7602) );
  INV_X1 U6892 ( .A(n7875), .ZN(n9042) );
  XNOR2_X1 U6893 ( .A(n5288), .B(n5287), .ZN(n6971) );
  NAND2_X1 U6894 ( .A1(n6971), .A2(n8878), .ZN(n5293) );
  INV_X1 U6895 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6896 ( .A1(n5289), .A2(n5305), .ZN(n5290) );
  NAND2_X1 U6897 ( .A1(n5290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U6898 ( .A(n5291), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U6899 ( .A1(n5358), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5357), .B2(
        n9794), .ZN(n5292) );
  NAND2_X1 U6900 ( .A1(n6642), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6901 ( .A1(n5146), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6902 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  AND2_X1 U6903 ( .A1(n5312), .A2(n5296), .ZN(n8712) );
  NAND2_X1 U6904 ( .A1(n5331), .A2(n8712), .ZN(n5298) );
  NAND2_X1 U6905 ( .A1(n5527), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5297) );
  OR2_X1 U6906 ( .A1(n8716), .A2(n8626), .ZN(n8834) );
  NAND2_X1 U6907 ( .A1(n8716), .A2(n8626), .ZN(n8929) );
  NAND2_X1 U6908 ( .A1(n8834), .A2(n8929), .ZN(n8998) );
  INV_X1 U6909 ( .A(n8626), .ZN(n9041) );
  XNOR2_X1 U6910 ( .A(n5303), .B(n5302), .ZN(n7039) );
  NAND2_X1 U6911 ( .A1(n7039), .A2(n8878), .ZN(n5310) );
  INV_X1 U6912 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6913 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  OAI21_X1 U6914 ( .B1(n5307), .B2(n5306), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5308) );
  XNOR2_X1 U6915 ( .A(n5308), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U6916 ( .A1(n5358), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5357), .B2(
        n9806), .ZN(n5309) );
  NAND2_X1 U6917 ( .A1(n5146), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6918 ( .A1(n5160), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5318) );
  INV_X1 U6919 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6920 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  AND2_X1 U6921 ( .A1(n5314), .A2(n5313), .ZN(n8625) );
  NAND2_X1 U6922 ( .A1(n5315), .A2(n8625), .ZN(n5317) );
  NAND2_X1 U6923 ( .A1(n5527), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6924 ( .A1(n7708), .A2(n8714), .ZN(n8828) );
  NAND2_X1 U6925 ( .A1(n8835), .A2(n8828), .ZN(n9000) );
  NAND2_X1 U6926 ( .A1(n7703), .A2(n9000), .ZN(n7702) );
  INV_X1 U6927 ( .A(n8714), .ZN(n9040) );
  NAND2_X1 U6928 ( .A1(n7702), .A2(n5320), .ZN(n7814) );
  NAND2_X1 U6929 ( .A1(n7814), .A2(n4899), .ZN(n5321) );
  XNOR2_X1 U6930 ( .A(n5323), .B(n5322), .ZN(n7380) );
  NAND2_X1 U6931 ( .A1(n7380), .A2(n8878), .ZN(n5328) );
  INV_X1 U6932 ( .A(n5324), .ZN(n5325) );
  NAND2_X1 U6933 ( .A1(n5325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5326) );
  XNOR2_X1 U6934 ( .A(n5326), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U6935 ( .A1(n5358), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5357), .B2(
        n9831), .ZN(n5327) );
  NAND2_X1 U6936 ( .A1(n5146), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6937 ( .A1(n5160), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6938 ( .A1(n5329), .A2(n8671), .ZN(n5330) );
  AND2_X1 U6939 ( .A1(n5343), .A2(n5330), .ZN(n8672) );
  NAND2_X1 U6940 ( .A1(n5331), .A2(n8672), .ZN(n5333) );
  NAND2_X1 U6941 ( .A1(n5527), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6942 ( .A1(n8676), .A2(n8763), .ZN(n9361) );
  INV_X1 U6943 ( .A(n8763), .ZN(n9368) );
  XNOR2_X1 U6944 ( .A(n5338), .B(n5337), .ZN(n7418) );
  NAND2_X1 U6945 ( .A1(n7418), .A2(n8878), .ZN(n5341) );
  XNOR2_X1 U6946 ( .A(n5339), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U6947 ( .A1(n5358), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5357), .B2(
        n9840), .ZN(n5340) );
  INV_X1 U6948 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6949 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  NAND2_X1 U6950 ( .A1(n5345), .A2(n5344), .ZN(n9375) );
  OR2_X1 U6951 ( .A1(n5488), .A2(n9375), .ZN(n5349) );
  NAND2_X1 U6952 ( .A1(n5160), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6953 ( .A1(n5146), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6954 ( .A1(n5527), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5346) );
  NAND4_X1 U6955 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n9473)
         );
  NAND2_X1 U6956 ( .A1(n9379), .A2(n9473), .ZN(n5350) );
  INV_X1 U6957 ( .A(n9379), .ZN(n9486) );
  OAI21_X1 U6958 ( .B1(n8685), .B2(n9478), .A(n5351), .ZN(n9328) );
  INV_X1 U6959 ( .A(n9328), .ZN(n5368) );
  XNOR2_X1 U6960 ( .A(n5353), .B(n5352), .ZN(n7625) );
  NAND2_X1 U6961 ( .A1(n7625), .A2(n8878), .ZN(n5360) );
  NAND2_X1 U6962 ( .A1(n5354), .A2(n5496), .ZN(n5355) );
  NAND2_X1 U6963 ( .A1(n5355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5356) );
  XNOR2_X2 U6964 ( .A(n5356), .B(n5494), .ZN(n8887) );
  AOI22_X1 U6965 ( .A1(n5358), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5357), .B2(
        n9022), .ZN(n5359) );
  INV_X1 U6966 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9333) );
  INV_X1 U6967 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6968 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  NAND2_X1 U6969 ( .A1(n5373), .A2(n5363), .ZN(n9332) );
  OR2_X1 U6970 ( .A1(n9332), .A2(n5488), .ZN(n5365) );
  AOI22_X1 U6971 ( .A1(n5146), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5160), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5364) );
  OAI211_X1 U6972 ( .C1(n5106), .C2(n9333), .A(n5365), .B(n5364), .ZN(n9476)
         );
  NAND2_X1 U6973 ( .A1(n9338), .A2(n9476), .ZN(n5367) );
  INV_X1 U6974 ( .A(n9476), .ZN(n9348) );
  AOI21_X2 U6975 ( .B1(n5368), .B2(n5367), .A(n5366), .ZN(n9314) );
  XNOR2_X1 U6976 ( .A(n5370), .B(n5369), .ZN(n7699) );
  NAND2_X1 U6977 ( .A1(n7699), .A2(n8878), .ZN(n5372) );
  OR2_X1 U6978 ( .A1(n5155), .A2(n7717), .ZN(n5371) );
  NAND2_X1 U6979 ( .A1(n5373), .A2(n8704), .ZN(n5374) );
  AND2_X1 U6980 ( .A1(n5386), .A2(n5374), .ZN(n9322) );
  NAND2_X1 U6981 ( .A1(n9322), .A2(n5331), .ZN(n5380) );
  INV_X1 U6982 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6983 ( .A1(n5146), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6984 ( .A1(n6642), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5375) );
  OAI211_X1 U6985 ( .C1(n5377), .C2(n5106), .A(n5376), .B(n5375), .ZN(n5378)
         );
  INV_X1 U6986 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6987 ( .A1(n9535), .A2(n9336), .ZN(n5381) );
  INV_X1 U6988 ( .A(n9336), .ZN(n9465) );
  AOI22_X1 U6989 ( .A1(n9314), .A2(n5381), .B1(n9321), .B2(n9465), .ZN(n9298)
         );
  XNOR2_X1 U6990 ( .A(n5383), .B(n5382), .ZN(n7777) );
  NAND2_X1 U6991 ( .A1(n7777), .A2(n8878), .ZN(n5385) );
  OR2_X1 U6992 ( .A1(n5155), .A2(n7778), .ZN(n5384) );
  INV_X1 U6993 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U6994 ( .A1(n5386), .A2(n9685), .ZN(n5387) );
  NAND2_X1 U6995 ( .A1(n5398), .A2(n5387), .ZN(n9304) );
  OR2_X1 U6996 ( .A1(n9304), .A2(n5488), .ZN(n5392) );
  INV_X1 U6997 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U6998 ( .A1(n5146), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6999 ( .A1(n5527), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U7000 ( .C1(n5103), .C2(n9613), .A(n5389), .B(n5388), .ZN(n5390)
         );
  INV_X1 U7001 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U7002 ( .A1(n5392), .A2(n5391), .ZN(n9440) );
  NAND2_X1 U7003 ( .A1(n9310), .A2(n9440), .ZN(n5393) );
  INV_X1 U7004 ( .A(n9440), .ZN(n8728) );
  XNOR2_X1 U7005 ( .A(n5395), .B(n5394), .ZN(n7838) );
  NAND2_X1 U7006 ( .A1(n7838), .A2(n8878), .ZN(n5397) );
  OR2_X1 U7007 ( .A1(n5155), .A2(n7840), .ZN(n5396) );
  INV_X1 U7008 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U7009 ( .A1(n5398), .A2(n8727), .ZN(n5399) );
  NAND2_X1 U7010 ( .A1(n5410), .A2(n5399), .ZN(n9287) );
  OR2_X1 U7011 ( .A1(n9287), .A2(n5488), .ZN(n5404) );
  INV_X1 U7012 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U7013 ( .A1(n5527), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U7014 ( .A1(n5160), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5400) );
  OAI211_X1 U7015 ( .C1(n5530), .C2(n9447), .A(n5401), .B(n5400), .ZN(n5402)
         );
  INV_X1 U7016 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U7017 ( .A1(n9443), .A2(n9308), .ZN(n5405) );
  XNOR2_X1 U7018 ( .A(n5407), .B(n5406), .ZN(n7950) );
  NAND2_X1 U7019 ( .A1(n7950), .A2(n8878), .ZN(n5409) );
  OR2_X1 U7020 ( .A1(n5155), .A2(n7952), .ZN(n5408) );
  NAND2_X1 U7021 ( .A1(n5410), .A2(n9682), .ZN(n5411) );
  NAND2_X1 U7022 ( .A1(n5423), .A2(n5411), .ZN(n9274) );
  OR2_X1 U7023 ( .A1(n9274), .A2(n5488), .ZN(n5416) );
  INV_X1 U7024 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U7025 ( .A1(n5146), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U7026 ( .A1(n5527), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5412) );
  OAI211_X1 U7027 ( .C1(n5103), .C2(n9671), .A(n5413), .B(n5412), .ZN(n5414)
         );
  INV_X1 U7028 ( .A(n5414), .ZN(n5415) );
  OR2_X1 U7029 ( .A1(n5155), .A2(n7955), .ZN(n5420) );
  NAND2_X1 U7030 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  AND2_X1 U7031 ( .A1(n5436), .A2(n5424), .ZN(n9254) );
  NAND2_X1 U7032 ( .A1(n9254), .A2(n5331), .ZN(n5430) );
  INV_X1 U7033 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U7034 ( .A1(n5527), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U7035 ( .A1(n6642), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5425) );
  OAI211_X1 U7036 ( .C1(n5530), .C2(n5427), .A(n5426), .B(n5425), .ZN(n5428)
         );
  INV_X1 U7037 ( .A(n5428), .ZN(n5429) );
  NOR2_X1 U7038 ( .A1(n9426), .A2(n9432), .ZN(n5431) );
  INV_X1 U7039 ( .A(n9426), .ZN(n9256) );
  OAI22_X2 U7040 ( .A1(n9251), .A2(n5431), .B1(n9256), .B2(n9278), .ZN(n9234)
         );
  XNOR2_X1 U7041 ( .A(n5433), .B(n5432), .ZN(n7958) );
  NAND2_X1 U7042 ( .A1(n7958), .A2(n8878), .ZN(n5435) );
  OR2_X1 U7043 ( .A1(n5155), .A2(n9605), .ZN(n5434) );
  INV_X1 U7044 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U7045 ( .A1(n5436), .A2(n8660), .ZN(n5437) );
  NAND2_X1 U7046 ( .A1(n5451), .A2(n5437), .ZN(n9241) );
  INV_X1 U7047 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U7048 ( .A1(n5527), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7049 ( .A1(n5160), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5438) );
  OAI211_X1 U7050 ( .C1(n5530), .C2(n9423), .A(n5439), .B(n5438), .ZN(n5440)
         );
  INV_X1 U7051 ( .A(n5440), .ZN(n5441) );
  NOR2_X1 U7052 ( .A1(n9420), .A2(n9263), .ZN(n5444) );
  NAND2_X1 U7053 ( .A1(n9420), .A2(n9263), .ZN(n5443) );
  NAND2_X1 U7054 ( .A1(n9572), .A2(n8878), .ZN(n5449) );
  OR2_X1 U7055 ( .A1(n5155), .A2(n5447), .ZN(n5448) );
  INV_X1 U7056 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7057 ( .A1(n5451), .A2(n5450), .ZN(n5452) );
  NAND2_X1 U7058 ( .A1(n5453), .A2(n5452), .ZN(n9224) );
  INV_X1 U7059 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U7060 ( .A1(n6642), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U7061 ( .A1(n5527), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U7062 ( .C1(n5530), .C2(n9415), .A(n5455), .B(n5454), .ZN(n5456)
         );
  INV_X1 U7063 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U7064 ( .A1(n9230), .A2(n9244), .ZN(n8960) );
  NAND2_X1 U7065 ( .A1(n9208), .A2(n9228), .ZN(n8869) );
  OAI21_X1 U7066 ( .B1(n9208), .B2(n9409), .A(n9203), .ZN(n9186) );
  AND2_X1 U7067 ( .A1(n5460), .A2(n5459), .ZN(n5463) );
  INV_X1 U7068 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5465) );
  INV_X1 U7069 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7964) );
  MUX2_X1 U7070 ( .A(n5465), .B(n7964), .S(n6610), .Z(n5482) );
  XNOR2_X1 U7071 ( .A(n5482), .B(SI_28_), .ZN(n5479) );
  NAND2_X1 U7072 ( .A1(n7963), .A2(n8878), .ZN(n5467) );
  OR2_X1 U7073 ( .A1(n5155), .A2(n7964), .ZN(n5466) );
  INV_X1 U7074 ( .A(n5470), .ZN(n5468) );
  NAND2_X1 U7075 ( .A1(n5468), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9176) );
  INV_X1 U7076 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7077 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U7078 ( .A1(n9176), .A2(n5471), .ZN(n9195) );
  INV_X1 U7079 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U7080 ( .A1(n5527), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7081 ( .A1(n6642), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5472) );
  OAI211_X1 U7082 ( .C1(n5530), .C2(n9398), .A(n5473), .B(n5472), .ZN(n5474)
         );
  INV_X1 U7083 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U7084 ( .A1(n9193), .A2(n9212), .ZN(n8870) );
  INV_X1 U7085 ( .A(n9193), .ZN(n9394) );
  NAND2_X1 U7086 ( .A1(n5480), .A2(n5479), .ZN(n5484) );
  INV_X1 U7087 ( .A(SI_28_), .ZN(n5481) );
  NAND2_X1 U7088 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  INV_X1 U7089 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5485) );
  INV_X1 U7090 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9697) );
  MUX2_X1 U7091 ( .A(n5485), .B(n9697), .S(n8770), .Z(n6470) );
  NAND2_X1 U7092 ( .A1(n6342), .A2(n8878), .ZN(n5487) );
  OR2_X1 U7093 ( .A1(n5155), .A2(n9697), .ZN(n5486) );
  OR2_X1 U7094 ( .A1(n9176), .A2(n5488), .ZN(n5493) );
  INV_X1 U7095 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U7096 ( .A1(n6642), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7097 ( .A1(n5527), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5489) );
  OAI211_X1 U7098 ( .C1(n5530), .C2(n5574), .A(n5490), .B(n5489), .ZN(n5491)
         );
  INV_X1 U7099 ( .A(n5491), .ZN(n5492) );
  OR2_X1 U7100 ( .A1(n9178), .A2(n9196), .ZN(n8954) );
  NAND2_X1 U7101 ( .A1(n9178), .A2(n9196), .ZN(n8956) );
  NAND2_X1 U7102 ( .A1(n5502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5503) );
  MUX2_X1 U7103 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5503), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5504) );
  NAND2_X1 U7104 ( .A1(n6085), .A2(n9028), .ZN(n5507) );
  NAND2_X1 U7105 ( .A1(n4313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7106 ( .A1(n7839), .A2(n7779), .ZN(n6958) );
  AND2_X1 U7107 ( .A1(n5507), .A2(n6958), .ZN(n5508) );
  NAND2_X1 U7108 ( .A1(n9013), .A2(n6086), .ZN(n6325) );
  NAND2_X1 U7109 ( .A1(n5508), .A2(n6325), .ZN(n7446) );
  INV_X1 U7110 ( .A(n5509), .ZN(n6851) );
  NAND2_X1 U7111 ( .A1(n6956), .A2(n7184), .ZN(n5510) );
  NAND2_X1 U7112 ( .A1(n6905), .A2(n8912), .ZN(n5512) );
  INV_X1 U7113 ( .A(n6911), .ZN(n8983) );
  INV_X1 U7114 ( .A(n8784), .ZN(n5513) );
  AND2_X1 U7115 ( .A1(n8917), .A2(n7281), .ZN(n8914) );
  NAND2_X1 U7116 ( .A1(n5514), .A2(n8785), .ZN(n7192) );
  INV_X1 U7117 ( .A(n8920), .ZN(n8987) );
  AND2_X1 U7118 ( .A1(n8800), .A2(n7385), .ZN(n8989) );
  INV_X1 U7119 ( .A(n8989), .ZN(n5517) );
  NAND2_X1 U7120 ( .A1(n8810), .A2(n8795), .ZN(n8801) );
  OR2_X1 U7121 ( .A1(n8801), .A2(n8989), .ZN(n8922) );
  INV_X1 U7122 ( .A(n8794), .ZN(n5515) );
  INV_X1 U7123 ( .A(n8788), .ZN(n8780) );
  NAND2_X1 U7124 ( .A1(n8922), .A2(n8993), .ZN(n5516) );
  OAI21_X1 U7125 ( .B1(n7384), .B2(n5517), .A(n5516), .ZN(n5518) );
  NAND2_X1 U7126 ( .A1(n5518), .A2(n8991), .ZN(n7359) );
  INV_X1 U7127 ( .A(n8994), .ZN(n7358) );
  NAND2_X1 U7128 ( .A1(n7359), .A2(n7358), .ZN(n7357) );
  INV_X1 U7129 ( .A(n7490), .ZN(n8996) );
  INV_X1 U7130 ( .A(n7602), .ZN(n8997) );
  NAND2_X1 U7131 ( .A1(n5519), .A2(n8928), .ZN(n7627) );
  INV_X1 U7132 ( .A(n8998), .ZN(n5520) );
  OR2_X1 U7133 ( .A1(n8766), .A2(n8673), .ZN(n8824) );
  NAND2_X1 U7134 ( .A1(n8766), .A2(n8673), .ZN(n8827) );
  NAND2_X1 U7135 ( .A1(n8824), .A2(n8827), .ZN(n9002) );
  INV_X1 U7136 ( .A(n8835), .ZN(n7816) );
  NOR2_X1 U7137 ( .A1(n9002), .A2(n7816), .ZN(n5521) );
  NAND2_X1 U7138 ( .A1(n7818), .A2(n8827), .ZN(n7893) );
  OR2_X1 U7139 ( .A1(n9379), .A2(n8737), .ZN(n8841) );
  NAND2_X1 U7140 ( .A1(n9379), .A2(n8737), .ZN(n8845) );
  NAND3_X1 U7141 ( .A1(n9362), .A2(n9363), .A3(n9361), .ZN(n9366) );
  OR2_X1 U7142 ( .A1(n9347), .A2(n8685), .ZN(n8848) );
  NAND2_X1 U7143 ( .A1(n9347), .A2(n8685), .ZN(n8846) );
  OR2_X1 U7144 ( .A1(n9338), .A2(n9348), .ZN(n8851) );
  NAND2_X1 U7145 ( .A1(n9338), .A2(n9348), .ZN(n8950) );
  INV_X1 U7146 ( .A(n8950), .ZN(n5522) );
  NAND2_X1 U7147 ( .A1(n9321), .A2(n9336), .ZN(n8855) );
  OR2_X1 U7148 ( .A1(n9310), .A2(n8728), .ZN(n8896) );
  NAND2_X1 U7149 ( .A1(n9310), .A2(n8728), .ZN(n8859) );
  OR2_X1 U7150 ( .A1(n9286), .A2(n9308), .ZN(n8775) );
  NAND2_X1 U7151 ( .A1(n9286), .A2(n9308), .ZN(n8774) );
  INV_X1 U7152 ( .A(n8774), .ZN(n5523) );
  NAND2_X1 U7153 ( .A1(n9280), .A2(n9291), .ZN(n8888) );
  NAND2_X1 U7154 ( .A1(n8861), .A2(n8888), .ZN(n9271) );
  OAI21_X1 U7155 ( .B1(n9272), .B2(n9271), .A(n8888), .ZN(n9259) );
  NAND2_X1 U7156 ( .A1(n9426), .A2(n9278), .ZN(n8900) );
  NAND2_X1 U7157 ( .A1(n8891), .A2(n8900), .ZN(n9260) );
  INV_X1 U7158 ( .A(n8891), .ZN(n9236) );
  NAND2_X1 U7159 ( .A1(n9246), .A2(n9263), .ZN(n8901) );
  NAND2_X1 U7160 ( .A1(n8894), .A2(n8901), .ZN(n9235) );
  INV_X1 U7161 ( .A(n8960), .ZN(n8951) );
  NOR2_X1 U7162 ( .A1(n9220), .A2(n8951), .ZN(n9216) );
  INV_X1 U7163 ( .A(n9206), .ZN(n9215) );
  OAI21_X1 U7164 ( .B1(n9216), .B2(n9215), .A(n8869), .ZN(n9189) );
  INV_X1 U7165 ( .A(n8870), .ZN(n8871) );
  AOI21_X1 U7166 ( .B1(n9189), .B2(n8953), .A(n8871), .ZN(n5524) );
  XNOR2_X1 U7167 ( .A(n5524), .B(n4488), .ZN(n5531) );
  OR2_X1 U7168 ( .A1(n7839), .A2(n8887), .ZN(n5525) );
  INV_X1 U7169 ( .A(n7779), .ZN(n8978) );
  NAND2_X1 U7170 ( .A1(n8978), .A2(n9014), .ZN(n8885) );
  NOR2_X2 U7171 ( .A1(n5563), .A2(n6851), .ZN(n9475) );
  INV_X1 U7172 ( .A(n9566), .ZN(n9766) );
  NAND2_X1 U7173 ( .A1(n9766), .A2(P1_B_REG_SCAN_IN), .ZN(n5526) );
  AND2_X1 U7174 ( .A1(n9475), .A2(n5526), .ZN(n9161) );
  INV_X1 U7175 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U7176 ( .A1(n5527), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7177 ( .A1(n5160), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U7178 ( .C1(n5530), .C2(n9390), .A(n5529), .B(n5528), .ZN(n9038)
         );
  OR2_X1 U7179 ( .A1(n6964), .A2(n6963), .ZN(n7279) );
  INV_X1 U7180 ( .A(n7562), .ZN(n7453) );
  NAND2_X1 U7181 ( .A1(n7448), .A2(n7453), .ZN(n7447) );
  INV_X1 U7182 ( .A(n7557), .ZN(n7813) );
  INV_X1 U7183 ( .A(n7877), .ZN(n7492) );
  NAND2_X1 U7184 ( .A1(n8830), .A2(n7821), .ZN(n7895) );
  NAND2_X1 U7185 ( .A1(n9452), .A2(n9320), .ZN(n9303) );
  AOI21_X1 U7186 ( .B1(n9178), .B2(n9191), .A(n9371), .ZN(n5532) );
  NAND2_X1 U7187 ( .A1(n5532), .A2(n9169), .ZN(n9181) );
  INV_X1 U7188 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7189 ( .A1(n5535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5536) );
  MUX2_X1 U7190 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5536), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5537) );
  NAND2_X1 U7191 ( .A1(n5537), .A2(n5543), .ZN(n7962) );
  NAND2_X1 U7192 ( .A1(n7962), .A2(P1_B_REG_SCAN_IN), .ZN(n5542) );
  NOR2_X1 U7193 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5538) );
  AOI21_X1 U7194 ( .B1(n5539), .B2(n5538), .A(n9554), .ZN(n5540) );
  MUX2_X1 U7195 ( .A(P1_B_REG_SCAN_IN), .B(n5542), .S(n7957), .Z(n5545) );
  NAND2_X1 U7196 ( .A1(n5543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5544) );
  INV_X1 U7197 ( .A(n9569), .ZN(n5566) );
  NAND2_X1 U7198 ( .A1(n5566), .A2(n7962), .ZN(n9552) );
  OAI21_X1 U7199 ( .B1(n9551), .B2(P1_D_REG_1__SCAN_IN), .A(n9552), .ZN(n6314)
         );
  INV_X1 U7200 ( .A(n9551), .ZN(n5556) );
  NOR4_X1 U7201 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5554) );
  NOR4_X1 U7202 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5553) );
  INV_X1 U7203 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9881) );
  INV_X1 U7204 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9878) );
  INV_X1 U7205 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9877) );
  INV_X1 U7206 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9880) );
  NAND4_X1 U7207 ( .A1(n9881), .A2(n9878), .A3(n9877), .A4(n9880), .ZN(n5551)
         );
  NOR4_X1 U7208 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5549) );
  NOR4_X1 U7209 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5548) );
  NOR4_X1 U7210 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5547) );
  NOR4_X1 U7211 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5546) );
  NAND4_X1 U7212 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n5550)
         );
  NOR4_X1 U7213 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n5551), .A4(n5550), .ZN(n5552) );
  NAND3_X1 U7214 ( .A1(n5554), .A2(n5553), .A3(n5552), .ZN(n5555) );
  NAND2_X1 U7215 ( .A1(n5556), .A2(n5555), .ZN(n7131) );
  INV_X1 U7216 ( .A(n7962), .ZN(n5557) );
  NAND2_X1 U7217 ( .A1(n5560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5562) );
  OAI211_X1 U7218 ( .C1(n6086), .C2(n5563), .A(n6316), .B(n6632), .ZN(n7130)
         );
  NAND2_X1 U7219 ( .A1(n9895), .A2(n7779), .ZN(n6321) );
  NAND2_X1 U7220 ( .A1(n6321), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5564) );
  NOR2_X1 U7221 ( .A1(n7130), .A2(n5564), .ZN(n5565) );
  NAND2_X1 U7222 ( .A1(n7957), .A2(n5566), .ZN(n9553) );
  INV_X1 U7223 ( .A(n9178), .ZN(n5573) );
  INV_X1 U7224 ( .A(n6958), .ZN(n7139) );
  INV_X1 U7225 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5568) );
  NOR2_X1 U7226 ( .A1(n9908), .A2(n5568), .ZN(n5569) );
  INV_X1 U7227 ( .A(n7132), .ZN(n6315) );
  INV_X1 U7228 ( .A(n9914), .ZN(n5572) );
  NAND2_X1 U7229 ( .A1(n9914), .A2(n9427), .ZN(n9463) );
  NOR2_X1 U7230 ( .A1(n9914), .A2(n5574), .ZN(n5575) );
  NAND2_X1 U7231 ( .A1(n5577), .A2(n5576), .ZN(P1_U3551) );
  INV_X1 U7232 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U7233 ( .A1(n7429), .A2(n5578), .ZN(n5686) );
  INV_X1 U7234 ( .A(n5686), .ZN(n5580) );
  NAND2_X1 U7235 ( .A1(n5580), .A2(n5579), .ZN(n5703) );
  OR2_X2 U7236 ( .A1(n5787), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5802) );
  OR2_X2 U7237 ( .A1(n5825), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5841) );
  OR2_X2 U7238 ( .A1(n5856), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5870) );
  INV_X1 U7239 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5591) );
  OR2_X2 U7240 ( .A1(n5901), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5908) );
  INV_X1 U7241 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7242 ( .A1(n5910), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7243 ( .A1(n5916), .A2(n5595), .ZN(n8355) );
  NAND2_X1 U7244 ( .A1(n6035), .A2(n6038), .ZN(n6040) );
  INV_X1 U7245 ( .A(n6040), .ZN(n5603) );
  NAND2_X1 U7246 ( .A1(n5614), .A2(n5604), .ZN(n8604) );
  XNOR2_X2 U7247 ( .A(n5605), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7980) );
  INV_X1 U7248 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5606) );
  INV_X1 U7249 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8573) );
  INV_X1 U7250 ( .A(n7980), .ZN(n5608) );
  NAND2_X1 U7251 ( .A1(n5635), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7252 ( .A1(n6501), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7253 ( .C1(n8573), .C2(n5646), .A(n5611), .B(n5610), .ZN(n5612)
         );
  INV_X1 U7254 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7255 ( .A1(n5616), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5617) );
  NOR2_X1 U7256 ( .A1(n6040), .A2(n5617), .ZN(n5620) );
  XNOR2_X1 U7257 ( .A(n5618), .B(P2_IR_REG_31__SCAN_IN), .ZN(n5619) );
  INV_X1 U7258 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5618) );
  AND2_X2 U7259 ( .A1(n5694), .A2(n5058), .ZN(n5663) );
  NAND2_X1 U7260 ( .A1(n7838), .A2(n6500), .ZN(n5622) );
  NAND2_X1 U7261 ( .A1(n5674), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5621) );
  INV_X1 U7262 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5623) );
  OR2_X1 U7263 ( .A1(n5646), .A2(n5623), .ZN(n5629) );
  NAND2_X1 U7264 ( .A1(n5624), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5627) );
  INV_X1 U7265 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5625) );
  NAND4_X1 U7266 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n7013)
         );
  INV_X1 U7267 ( .A(n5694), .ZN(n5677) );
  INV_X1 U7268 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7269 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5630) );
  OAI211_X4 U7270 ( .C1(P1_DATAO_REG_1__SCAN_IN), .C2(n5693), .A(n5633), .B(
        n5632), .ZN(n7269) );
  NAND2_X1 U7271 ( .A1(n4292), .A2(n7270), .ZN(n6017) );
  NAND2_X1 U7272 ( .A1(n7013), .A2(n7269), .ZN(n6351) );
  NAND2_X1 U7273 ( .A1(n6017), .A2(n6351), .ZN(n6014) );
  INV_X1 U7274 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U7275 ( .A1(n5635), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7276 ( .A1(n5657), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7277 ( .A1(n5785), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7278 ( .A1(n5058), .A2(SI_0_), .ZN(n5641) );
  XNOR2_X1 U7279 ( .A(n5641), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8620) );
  MUX2_X1 U7280 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8620), .S(n5694), .Z(n7967) );
  NAND2_X1 U7281 ( .A1(n6978), .A2(n7967), .ZN(n6976) );
  NAND2_X1 U7282 ( .A1(n6014), .A2(n6976), .ZN(n5643) );
  NAND2_X1 U7283 ( .A1(n4292), .A2(n7269), .ZN(n5642) );
  NAND2_X1 U7284 ( .A1(n5643), .A2(n5642), .ZN(n7010) );
  INV_X1 U7285 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5644) );
  INV_X1 U7286 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7250) );
  OR2_X1 U7287 ( .A1(n5658), .A2(n7250), .ZN(n5649) );
  INV_X1 U7288 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5645) );
  OR2_X1 U7289 ( .A1(n5646), .A2(n5645), .ZN(n5648) );
  INV_X1 U7290 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U7291 ( .A1(n5663), .A2(n5651), .ZN(n5654) );
  NAND2_X1 U7292 ( .A1(n5674), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7293 ( .A1(n5677), .A2(n6795), .ZN(n5652) );
  NAND2_X1 U7294 ( .A1(n7010), .A2(n7011), .ZN(n5656) );
  INV_X1 U7295 ( .A(n7973), .ZN(n6018) );
  OR2_X1 U7296 ( .A1(n6359), .A2(n6018), .ZN(n5655) );
  NAND2_X1 U7297 ( .A1(n5656), .A2(n5655), .ZN(n7422) );
  NAND2_X1 U7298 ( .A1(n5785), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5661) );
  OR2_X1 U7299 ( .A1(n5858), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7300 ( .A1(n5674), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7301 ( .A1(n5675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5664) );
  XNOR2_X1 U7302 ( .A(n5664), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U7303 ( .A1(n5677), .A2(n6757), .ZN(n5665) );
  NOR2_X1 U7304 ( .A1(n8201), .A2(n7430), .ZN(n5667) );
  INV_X1 U7305 ( .A(n7430), .ZN(n10072) );
  INV_X1 U7306 ( .A(n7479), .ZN(n5682) );
  NAND2_X1 U7307 ( .A1(n6501), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5673) );
  INV_X1 U7308 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6747) );
  OR2_X1 U7309 ( .A1(n6483), .A2(n6747), .ZN(n5672) );
  NAND2_X1 U7310 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5668) );
  AND2_X1 U7311 ( .A1(n5686), .A2(n5668), .ZN(n7476) );
  OR2_X1 U7312 ( .A1(n5858), .A2(n7476), .ZN(n5671) );
  INV_X1 U7313 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5669) );
  OR2_X1 U7314 ( .A1(n5646), .A2(n5669), .ZN(n5670) );
  NAND2_X1 U7315 ( .A1(n5674), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7316 ( .A1(n5695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U7317 ( .A(n5676), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U7318 ( .A1(n5677), .A2(n6923), .ZN(n5678) );
  OAI211_X1 U7319 ( .C1(n6618), .C2(n5680), .A(n5679), .B(n5678), .ZN(n7153)
         );
  NAND2_X1 U7320 ( .A1(n7232), .A2(n7153), .ZN(n6367) );
  INV_X1 U7321 ( .A(n7232), .ZN(n5683) );
  INV_X1 U7322 ( .A(n7153), .ZN(n10076) );
  NAND2_X1 U7323 ( .A1(n5683), .A2(n10076), .ZN(n6387) );
  INV_X1 U7324 ( .A(n7480), .ZN(n5681) );
  NAND2_X1 U7325 ( .A1(n5682), .A2(n5681), .ZN(n7477) );
  OR2_X1 U7326 ( .A1(n5683), .A2(n7153), .ZN(n5684) );
  INV_X1 U7327 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5685) );
  INV_X1 U7328 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7375) );
  OR2_X1 U7329 ( .A1(n5999), .A2(n7375), .ZN(n5691) );
  NAND2_X1 U7330 ( .A1(n5686), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5687) );
  AND2_X1 U7331 ( .A1(n5703), .A2(n5687), .ZN(n7238) );
  OR2_X1 U7332 ( .A1(n5858), .A2(n7238), .ZN(n5690) );
  INV_X1 U7333 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5688) );
  OR2_X1 U7334 ( .A1(n5646), .A2(n5688), .ZN(n5689) );
  NAND2_X1 U7335 ( .A1(n6620), .A2(n6500), .ZN(n5701) );
  INV_X1 U7336 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6629) );
  INV_X1 U7337 ( .A(n5695), .ZN(n5697) );
  INV_X1 U7338 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7339 ( .A1(n5697), .A2(n5696), .ZN(n5710) );
  NAND2_X1 U7340 ( .A1(n5710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5698) );
  XNOR2_X1 U7341 ( .A(n5698), .B(n5711), .ZN(n7049) );
  OAI22_X1 U7342 ( .A1(n5890), .A2(n6629), .B1(n6607), .B2(n7049), .ZN(n5699)
         );
  INV_X1 U7343 ( .A(n5699), .ZN(n5700) );
  NAND2_X1 U7344 ( .A1(n6501), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5709) );
  INV_X1 U7345 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5702) );
  OR2_X1 U7346 ( .A1(n6483), .A2(n5702), .ZN(n5708) );
  NAND2_X1 U7347 ( .A1(n5703), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5704) );
  AND2_X1 U7348 ( .A1(n5729), .A2(n5704), .ZN(n7262) );
  OR2_X1 U7349 ( .A1(n5858), .A2(n7262), .ZN(n5707) );
  INV_X1 U7350 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5705) );
  OR2_X1 U7351 ( .A1(n5646), .A2(n5705), .ZN(n5706) );
  NAND2_X1 U7352 ( .A1(n6635), .A2(n6500), .ZN(n5718) );
  INV_X1 U7353 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6637) );
  INV_X1 U7354 ( .A(n5710), .ZN(n5712) );
  NAND2_X1 U7355 ( .A1(n5712), .A2(n5711), .ZN(n5714) );
  NAND2_X1 U7356 ( .A1(n5714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5713) );
  MUX2_X1 U7357 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5713), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5715) );
  NAND2_X1 U7358 ( .A1(n5715), .A2(n5724), .ZN(n7079) );
  OAI22_X1 U7359 ( .A1(n5890), .A2(n6637), .B1(n6607), .B2(n7079), .ZN(n5716)
         );
  INV_X1 U7360 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7361 ( .A1(n5718), .A2(n5717), .ZN(n10085) );
  NAND2_X1 U7362 ( .A1(n5719), .A2(n10085), .ZN(n5722) );
  INV_X1 U7363 ( .A(n7410), .ZN(n5720) );
  NAND2_X1 U7364 ( .A1(n5720), .A2(n4628), .ZN(n5721) );
  AND2_X2 U7365 ( .A1(n5722), .A2(n5721), .ZN(n7591) );
  NAND2_X1 U7366 ( .A1(n6640), .A2(n6500), .ZN(n5728) );
  INV_X1 U7367 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U7368 ( .A1(n5724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5723) );
  MUX2_X1 U7369 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5723), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5725) );
  NAND2_X1 U7370 ( .A1(n5725), .A2(n5751), .ZN(n7161) );
  OAI22_X1 U7371 ( .A1(n5890), .A2(n9623), .B1(n6607), .B2(n7161), .ZN(n5726)
         );
  INV_X1 U7372 ( .A(n5726), .ZN(n5727) );
  NAND2_X1 U7373 ( .A1(n5728), .A2(n5727), .ZN(n10093) );
  NAND2_X1 U7374 ( .A1(n5635), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5735) );
  INV_X1 U7375 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7056) );
  OR2_X1 U7376 ( .A1(n5999), .A2(n7056), .ZN(n5734) );
  NAND2_X1 U7377 ( .A1(n5729), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5730) );
  AND2_X1 U7378 ( .A1(n5743), .A2(n5730), .ZN(n7596) );
  OR2_X1 U7379 ( .A1(n5858), .A2(n7596), .ZN(n5733) );
  INV_X1 U7380 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5731) );
  OR2_X1 U7381 ( .A1(n5646), .A2(n5731), .ZN(n5732) );
  NAND4_X1 U7382 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n8199)
         );
  OR2_X1 U7383 ( .A1(n10093), .A2(n8199), .ZN(n7573) );
  NAND2_X1 U7384 ( .A1(n10093), .A2(n8199), .ZN(n5736) );
  NAND2_X1 U7385 ( .A1(n7573), .A2(n5736), .ZN(n7588) );
  NAND2_X1 U7386 ( .A1(n7572), .A2(n7573), .ZN(n5750) );
  NAND2_X1 U7387 ( .A1(n6661), .A2(n6500), .ZN(n5742) );
  NAND2_X1 U7388 ( .A1(n5751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5739) );
  INV_X1 U7389 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5738) );
  OAI22_X1 U7390 ( .A1(n5890), .A2(n6663), .B1(n6607), .B2(n7307), .ZN(n5740)
         );
  INV_X1 U7391 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7392 ( .A1(n5742), .A2(n5741), .ZN(n10096) );
  NAND2_X1 U7393 ( .A1(n5635), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5749) );
  INV_X1 U7394 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7581) );
  OR2_X1 U7395 ( .A1(n5999), .A2(n7581), .ZN(n5748) );
  NAND2_X1 U7396 ( .A1(n5743), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5744) );
  AND2_X1 U7397 ( .A1(n5757), .A2(n5744), .ZN(n7580) );
  OR2_X1 U7398 ( .A1(n5858), .A2(n7580), .ZN(n5747) );
  INV_X1 U7399 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5745) );
  OR2_X1 U7400 ( .A1(n5646), .A2(n5745), .ZN(n5746) );
  OR2_X1 U7401 ( .A1(n10096), .A2(n7661), .ZN(n6372) );
  NAND2_X1 U7402 ( .A1(n10096), .A2(n7661), .ZN(n6375) );
  NAND2_X1 U7403 ( .A1(n6372), .A2(n6375), .ZN(n7583) );
  NAND2_X1 U7404 ( .A1(n5750), .A2(n7583), .ZN(n7571) );
  OR2_X1 U7405 ( .A1(n10096), .A2(n8198), .ZN(n7676) );
  NAND2_X1 U7406 ( .A1(n7571), .A2(n7676), .ZN(n5764) );
  NAND2_X1 U7407 ( .A1(n6704), .A2(n6500), .ZN(n5756) );
  OAI21_X1 U7408 ( .B1(n5751), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5753) );
  INV_X1 U7409 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5752) );
  XNOR2_X1 U7410 ( .A(n5753), .B(n5752), .ZN(n8232) );
  OAI22_X1 U7411 ( .A1(n5890), .A2(n6707), .B1(n6607), .B2(n8232), .ZN(n5754)
         );
  INV_X1 U7412 ( .A(n5754), .ZN(n5755) );
  NAND2_X2 U7413 ( .A1(n5756), .A2(n5755), .ZN(n7784) );
  NAND2_X1 U7414 ( .A1(n5635), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5763) );
  INV_X1 U7415 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7681) );
  OR2_X1 U7416 ( .A1(n5999), .A2(n7681), .ZN(n5762) );
  NAND2_X1 U7417 ( .A1(n5757), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5758) );
  AND2_X1 U7418 ( .A1(n5774), .A2(n5758), .ZN(n7680) );
  OR2_X1 U7419 ( .A1(n5858), .A2(n7680), .ZN(n5761) );
  INV_X1 U7420 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5759) );
  OR2_X1 U7421 ( .A1(n5646), .A2(n5759), .ZN(n5760) );
  NAND2_X1 U7422 ( .A1(n7784), .A2(n7577), .ZN(n6376) );
  NAND2_X1 U7423 ( .A1(n6373), .A2(n6376), .ZN(n7675) );
  OR2_X1 U7424 ( .A1(n7784), .A2(n8197), .ZN(n5765) );
  NAND2_X1 U7425 ( .A1(n6709), .A2(n6500), .ZN(n5773) );
  OR2_X1 U7426 ( .A1(n5766), .A2(n5606), .ZN(n5768) );
  MUX2_X1 U7427 ( .A(n5768), .B(P2_IR_REG_31__SCAN_IN), .S(n5767), .Z(n5770)
         );
  NAND2_X1 U7428 ( .A1(n5770), .A2(n5769), .ZN(n9932) );
  OAI22_X1 U7429 ( .A1(n5890), .A2(n6711), .B1(n6607), .B2(n9932), .ZN(n5771)
         );
  INV_X1 U7430 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7431 ( .A1(n6501), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5780) );
  INV_X1 U7432 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8254) );
  OR2_X1 U7433 ( .A1(n6483), .A2(n8254), .ZN(n5779) );
  NAND2_X1 U7434 ( .A1(n5774), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5775) );
  AND2_X1 U7435 ( .A1(n5787), .A2(n5775), .ZN(n7793) );
  OR2_X1 U7436 ( .A1(n5858), .A2(n7793), .ZN(n5778) );
  INV_X1 U7437 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5776) );
  OR2_X1 U7438 ( .A1(n5646), .A2(n5776), .ZN(n5777) );
  NAND4_X1 U7439 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n8196)
         );
  NOR2_X1 U7440 ( .A1(n7799), .A2(n8196), .ZN(n7858) );
  NAND2_X1 U7441 ( .A1(n6713), .A2(n6500), .ZN(n5784) );
  NAND2_X1 U7442 ( .A1(n5769), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5781) );
  XNOR2_X1 U7443 ( .A(n5781), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9950) );
  INV_X1 U7444 ( .A(n9950), .ZN(n8261) );
  OAI22_X1 U7445 ( .A1(n5890), .A2(n6798), .B1(n6607), .B2(n8261), .ZN(n5782)
         );
  INV_X1 U7446 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U7447 ( .A1(n5784), .A2(n5783), .ZN(n7868) );
  NAND2_X1 U7448 ( .A1(n5785), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5792) );
  INV_X1 U7449 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5786) );
  OR2_X1 U7450 ( .A1(n6483), .A2(n5786), .ZN(n5791) );
  INV_X1 U7451 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7866) );
  OR2_X1 U7452 ( .A1(n5999), .A2(n7866), .ZN(n5790) );
  NAND2_X1 U7453 ( .A1(n5787), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5788) );
  AND2_X1 U7454 ( .A1(n5802), .A2(n5788), .ZN(n7865) );
  OR2_X1 U7455 ( .A1(n5858), .A2(n7865), .ZN(n5789) );
  NAND4_X1 U7456 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n8195)
         );
  OR2_X1 U7457 ( .A1(n7858), .A2(n5793), .ZN(n5797) );
  NAND2_X1 U7458 ( .A1(n7799), .A2(n8196), .ZN(n7859) );
  OR2_X1 U7459 ( .A1(n5793), .A2(n7859), .ZN(n5795) );
  NAND2_X1 U7460 ( .A1(n7868), .A2(n8195), .ZN(n5794) );
  AND2_X1 U7461 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7462 ( .A1(n6984), .A2(n6500), .ZN(n5801) );
  NAND2_X1 U7463 ( .A1(n5809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U7464 ( .A(n5798), .B(n4397), .ZN(n8239) );
  OAI22_X1 U7465 ( .A1(n5890), .A2(n6985), .B1(n6607), .B2(n8239), .ZN(n5799)
         );
  INV_X1 U7466 ( .A(n5799), .ZN(n5800) );
  NAND2_X1 U7467 ( .A1(n6501), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5808) );
  INV_X1 U7468 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8263) );
  OR2_X1 U7469 ( .A1(n6483), .A2(n8263), .ZN(n5807) );
  NAND2_X1 U7470 ( .A1(n5802), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5803) );
  AND2_X1 U7471 ( .A1(n5814), .A2(n5803), .ZN(n7927) );
  OR2_X1 U7472 ( .A1(n5858), .A2(n7927), .ZN(n5806) );
  INV_X1 U7473 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5804) );
  OR2_X1 U7474 ( .A1(n5646), .A2(n5804), .ZN(n5805) );
  NAND4_X1 U7475 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n8194)
         );
  NAND2_X1 U7476 ( .A1(n6971), .A2(n6500), .ZN(n5812) );
  INV_X1 U7477 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7006) );
  OR2_X1 U7478 ( .A1(n5851), .A2(n5606), .ZN(n5820) );
  XNOR2_X1 U7479 ( .A(n5820), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9984) );
  OAI22_X1 U7480 ( .A1(n5890), .A2(n7006), .B1(n6607), .B2(n8266), .ZN(n5810)
         );
  INV_X1 U7481 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U7482 ( .A1(n5785), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5819) );
  INV_X1 U7483 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5813) );
  OR2_X1 U7484 ( .A1(n6483), .A2(n5813), .ZN(n5818) );
  INV_X1 U7485 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8243) );
  OR2_X1 U7486 ( .A1(n5999), .A2(n8243), .ZN(n5817) );
  NAND2_X1 U7487 ( .A1(n5814), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5815) );
  AND2_X1 U7488 ( .A1(n5825), .A2(n5815), .ZN(n8131) );
  OR2_X1 U7489 ( .A1(n5858), .A2(n8131), .ZN(n5816) );
  NAND4_X1 U7490 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(n5816), .ZN(n8458)
         );
  NOR2_X1 U7491 ( .A1(n8133), .A2(n8458), .ZN(n6518) );
  NAND2_X1 U7492 ( .A1(n8133), .A2(n8458), .ZN(n6516) );
  NAND2_X1 U7493 ( .A1(n7039), .A2(n6500), .ZN(n5824) );
  NAND2_X1 U7494 ( .A1(n5820), .A2(n5849), .ZN(n5821) );
  NAND2_X1 U7495 ( .A1(n5821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5834) );
  XNOR2_X1 U7496 ( .A(n5834), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10001) );
  INV_X1 U7497 ( .A(n10001), .ZN(n8253) );
  OAI22_X1 U7498 ( .A1(n5890), .A2(n7086), .B1(n6607), .B2(n8253), .ZN(n5822)
         );
  INV_X1 U7499 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U7500 ( .A1(n5785), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5830) );
  INV_X1 U7501 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9680) );
  OR2_X1 U7502 ( .A1(n6483), .A2(n9680), .ZN(n5829) );
  INV_X1 U7503 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8473) );
  OR2_X1 U7504 ( .A1(n5999), .A2(n8473), .ZN(n5828) );
  NAND2_X1 U7505 ( .A1(n5825), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5826) );
  AND2_X1 U7506 ( .A1(n5841), .A2(n5826), .ZN(n8463) );
  OR2_X1 U7507 ( .A1(n5858), .A2(n8463), .ZN(n5827) );
  NAND4_X1 U7508 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n8193)
         );
  AND2_X1 U7509 ( .A1(n8461), .A2(n8193), .ZN(n5831) );
  OR2_X1 U7510 ( .A1(n8461), .A2(n8193), .ZN(n5832) );
  NAND2_X1 U7511 ( .A1(n7205), .A2(n6500), .ZN(n5839) );
  NAND2_X1 U7512 ( .A1(n5834), .A2(n5848), .ZN(n5835) );
  NAND2_X1 U7513 ( .A1(n5835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U7514 ( .A(n5836), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10018) );
  INV_X1 U7515 ( .A(n10018), .ZN(n8269) );
  OAI22_X1 U7516 ( .A1(n5890), .A2(n7206), .B1(n6607), .B2(n8269), .ZN(n5837)
         );
  INV_X1 U7517 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U7518 ( .A1(n5785), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5846) );
  INV_X1 U7519 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8534) );
  OR2_X1 U7520 ( .A1(n6483), .A2(n8534), .ZN(n5845) );
  INV_X1 U7521 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5840) );
  OR2_X1 U7522 ( .A1(n5999), .A2(n5840), .ZN(n5844) );
  NAND2_X1 U7523 ( .A1(n5841), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5842) );
  AND2_X1 U7524 ( .A1(n5856), .A2(n5842), .ZN(n8173) );
  OR2_X1 U7525 ( .A1(n5858), .A2(n8173), .ZN(n5843) );
  NAND2_X1 U7526 ( .A1(n8168), .A2(n8430), .ZN(n6416) );
  NAND2_X1 U7527 ( .A1(n6417), .A2(n6416), .ZN(n8437) );
  NAND2_X1 U7528 ( .A1(n7380), .A2(n6500), .ZN(n5855) );
  AND3_X1 U7529 ( .A1(n5849), .A2(n5848), .A3(n5847), .ZN(n5850) );
  NAND2_X1 U7530 ( .A1(n4374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7531 ( .A(n5852), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10033) );
  OAI22_X1 U7532 ( .A1(n5890), .A2(n7381), .B1(n6607), .B2(n8252), .ZN(n5853)
         );
  INV_X1 U7533 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7534 ( .A1(n6501), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5862) );
  INV_X1 U7535 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8530) );
  OR2_X1 U7536 ( .A1(n6483), .A2(n8530), .ZN(n5861) );
  NAND2_X1 U7537 ( .A1(n5856), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5857) );
  AND2_X1 U7538 ( .A1(n5870), .A2(n5857), .ZN(n8093) );
  OR2_X1 U7539 ( .A1(n8093), .A2(n5858), .ZN(n5860) );
  INV_X1 U7540 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9713) );
  OR2_X1 U7541 ( .A1(n5646), .A2(n9713), .ZN(n5859) );
  NAND2_X1 U7542 ( .A1(n8089), .A2(n8441), .ZN(n6419) );
  NAND2_X1 U7543 ( .A1(n6420), .A2(n6419), .ZN(n8425) );
  NAND2_X1 U7544 ( .A1(n8089), .A2(n8414), .ZN(n5863) );
  NAND2_X1 U7545 ( .A1(n7418), .A2(n6500), .ZN(n5869) );
  NAND2_X1 U7546 ( .A1(n5877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5866) );
  XNOR2_X1 U7547 ( .A(n5866), .B(n5865), .ZN(n8272) );
  OAI22_X1 U7548 ( .A1(n5890), .A2(n7419), .B1(n6607), .B2(n8272), .ZN(n5867)
         );
  INV_X1 U7549 ( .A(n5867), .ZN(n5868) );
  NAND2_X1 U7550 ( .A1(n5870), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7551 ( .A1(n5881), .A2(n5871), .ZN(n8418) );
  NAND2_X1 U7552 ( .A1(n5995), .A2(n8418), .ZN(n5875) );
  INV_X1 U7553 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8526) );
  OR2_X1 U7554 ( .A1(n6483), .A2(n8526), .ZN(n5874) );
  INV_X1 U7555 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8203) );
  OR2_X1 U7556 ( .A1(n5999), .A2(n8203), .ZN(n5873) );
  INV_X1 U7557 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8588) );
  OR2_X1 U7558 ( .A1(n5646), .A2(n8588), .ZN(n5872) );
  OR2_X1 U7559 ( .A1(n8417), .A2(n8427), .ZN(n6426) );
  NAND2_X1 U7560 ( .A1(n8417), .A2(n8427), .ZN(n6422) );
  NAND2_X1 U7561 ( .A1(n6426), .A2(n6422), .ZN(n8411) );
  NAND2_X1 U7562 ( .A1(n8412), .A2(n8411), .ZN(n8410) );
  INV_X1 U7563 ( .A(n8427), .ZN(n8192) );
  NAND2_X1 U7564 ( .A1(n8417), .A2(n8192), .ZN(n5876) );
  NAND2_X1 U7565 ( .A1(n7527), .A2(n6500), .ZN(n5880) );
  XNOR2_X1 U7566 ( .A(n5889), .B(n5888), .ZN(n9738) );
  OAI22_X1 U7567 ( .A1(n5890), .A2(n7528), .B1(n6607), .B2(n9738), .ZN(n5878)
         );
  INV_X1 U7568 ( .A(n5878), .ZN(n5879) );
  NAND2_X1 U7569 ( .A1(n5881), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7570 ( .A1(n5894), .A2(n5882), .ZN(n8405) );
  NAND2_X1 U7571 ( .A1(n8405), .A2(n5995), .ZN(n5886) );
  NAND2_X1 U7572 ( .A1(n5635), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7573 ( .A1(n6501), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7574 ( .A1(n5785), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5883) );
  NAND4_X1 U7575 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n8413)
         );
  OR2_X1 U7576 ( .A1(n8145), .A2(n8413), .ZN(n5887) );
  NAND2_X1 U7577 ( .A1(n7625), .A2(n6500), .ZN(n5893) );
  OAI22_X1 U7578 ( .A1(n5890), .A2(n7626), .B1(n6010), .B2(n6607), .ZN(n5891)
         );
  INV_X1 U7579 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U7580 ( .A1(n5894), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7581 ( .A1(n5901), .A2(n5895), .ZN(n8390) );
  NAND2_X1 U7582 ( .A1(n8390), .A2(n5995), .ZN(n5898) );
  AOI22_X1 U7583 ( .A1(n5785), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6501), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7584 ( .A1(n5635), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7585 ( .A1(n8394), .A2(n8404), .ZN(n6427) );
  AND2_X2 U7586 ( .A1(n6431), .A2(n6427), .ZN(n8395) );
  INV_X1 U7587 ( .A(n8394), .ZN(n8514) );
  NAND2_X1 U7588 ( .A1(n7699), .A2(n6500), .ZN(n5900) );
  NAND2_X1 U7589 ( .A1(n5674), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7590 ( .A1(n5901), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7591 ( .A1(n5908), .A2(n5902), .ZN(n8379) );
  NAND2_X1 U7592 ( .A1(n8379), .A2(n5995), .ZN(n5905) );
  AOI22_X1 U7593 ( .A1(n5635), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6501), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7594 ( .A1(n5785), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7595 ( .A1(n8508), .A2(n8387), .ZN(n6434) );
  INV_X1 U7596 ( .A(n8387), .ZN(n8191) );
  NOR2_X1 U7597 ( .A1(n8508), .A2(n8191), .ZN(n8363) );
  NAND2_X1 U7598 ( .A1(n7777), .A2(n6500), .ZN(n5907) );
  NAND2_X1 U7599 ( .A1(n5674), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7600 ( .A1(n5908), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7601 ( .A1(n5910), .A2(n5909), .ZN(n8368) );
  INV_X1 U7602 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U7603 ( .A1(n5635), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7604 ( .A1(n6501), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5911) );
  OAI211_X1 U7605 ( .C1(n8577), .C2(n5646), .A(n5912), .B(n5911), .ZN(n5913)
         );
  NAND2_X1 U7606 ( .A1(n8074), .A2(n8378), .ZN(n6433) );
  NAND2_X1 U7607 ( .A1(n6436), .A2(n6433), .ZN(n8362) );
  NAND2_X1 U7608 ( .A1(n8579), .A2(n8378), .ZN(n8349) );
  OR2_X1 U7609 ( .A1(n8142), .A2(n8367), .ZN(n6439) );
  NAND2_X1 U7610 ( .A1(n8142), .A2(n8367), .ZN(n6438) );
  NAND2_X1 U7611 ( .A1(n7950), .A2(n6500), .ZN(n5915) );
  NAND2_X1 U7612 ( .A1(n5674), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U7613 ( .A1(n5916), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7614 ( .A1(n5928), .A2(n5917), .ZN(n8343) );
  NAND2_X1 U7615 ( .A1(n8343), .A2(n5995), .ZN(n5923) );
  INV_X1 U7616 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7617 ( .A1(n5785), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7618 ( .A1(n5635), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5918) );
  OAI211_X1 U7619 ( .C1(n5999), .C2(n5920), .A(n5919), .B(n5918), .ZN(n5921)
         );
  INV_X1 U7620 ( .A(n5921), .ZN(n5922) );
  NOR2_X1 U7621 ( .A1(n8571), .A2(n8354), .ZN(n5924) );
  NAND2_X1 U7622 ( .A1(n7953), .A2(n6500), .ZN(n5926) );
  NAND2_X1 U7623 ( .A1(n5674), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5925) );
  INV_X1 U7624 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U7625 ( .A1(n5928), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7626 ( .A1(n5942), .A2(n5929), .ZN(n8331) );
  NAND2_X1 U7627 ( .A1(n8331), .A2(n5995), .ZN(n5934) );
  INV_X1 U7628 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U7629 ( .A1(n5635), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7630 ( .A1(n6501), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U7631 ( .C1(n8565), .C2(n5646), .A(n5931), .B(n5930), .ZN(n5932)
         );
  INV_X1 U7632 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7633 ( .A1(n7958), .A2(n6500), .ZN(n5939) );
  NAND2_X1 U7634 ( .A1(n5674), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5938) );
  INV_X1 U7635 ( .A(n5942), .ZN(n5941) );
  INV_X1 U7636 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7637 ( .A1(n5942), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7638 ( .A1(n5953), .A2(n5943), .ZN(n8322) );
  NAND2_X1 U7639 ( .A1(n8322), .A2(n5995), .ZN(n5948) );
  INV_X1 U7640 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U7641 ( .A1(n6501), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7642 ( .A1(n5635), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5944) );
  OAI211_X1 U7643 ( .C1(n5646), .C2(n8561), .A(n5945), .B(n5944), .ZN(n5946)
         );
  INV_X1 U7644 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U7645 ( .A1(n8077), .A2(n8186), .ZN(n5950) );
  NOR2_X1 U7646 ( .A1(n8077), .A2(n8186), .ZN(n5949) );
  NAND2_X1 U7647 ( .A1(n9572), .A2(n6500), .ZN(n5952) );
  NAND2_X1 U7648 ( .A1(n5674), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5951) );
  OR2_X2 U7649 ( .A1(n5953), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7650 ( .A1(n5953), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7651 ( .A1(n5965), .A2(n5954), .ZN(n8313) );
  NAND2_X1 U7652 ( .A1(n8313), .A2(n5995), .ZN(n5959) );
  INV_X1 U7653 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U7654 ( .A1(n5635), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7655 ( .A1(n6501), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5955) );
  OAI211_X1 U7656 ( .C1(n8557), .C2(n5646), .A(n5956), .B(n5955), .ZN(n5957)
         );
  INV_X1 U7657 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U7658 ( .A1(n8559), .A2(n8320), .ZN(n5960) );
  NAND2_X1 U7659 ( .A1(n8612), .A2(n6500), .ZN(n5962) );
  NAND2_X1 U7660 ( .A1(n5674), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5961) );
  INV_X1 U7661 ( .A(n5965), .ZN(n5964) );
  INV_X1 U7662 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7663 ( .A1(n5964), .A2(n5963), .ZN(n5977) );
  NAND2_X1 U7664 ( .A1(n5965), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7665 ( .A1(n5977), .A2(n5966), .ZN(n8042) );
  NAND2_X1 U7666 ( .A1(n8042), .A2(n5995), .ZN(n5972) );
  INV_X1 U7667 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7668 ( .A1(n5635), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7669 ( .A1(n6501), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5967) );
  OAI211_X1 U7670 ( .C1(n5969), .C2(n5646), .A(n5968), .B(n5967), .ZN(n5970)
         );
  INV_X1 U7671 ( .A(n5970), .ZN(n5971) );
  NAND2_X1 U7672 ( .A1(n8553), .A2(n8185), .ZN(n5973) );
  NAND2_X1 U7673 ( .A1(n7963), .A2(n6500), .ZN(n5976) );
  NAND2_X1 U7674 ( .A1(n5674), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7675 ( .A1(n5977), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7676 ( .A1(n8031), .A2(n5978), .ZN(n8288) );
  NAND2_X1 U7677 ( .A1(n8288), .A2(n5995), .ZN(n5983) );
  NAND2_X1 U7678 ( .A1(n5785), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7679 ( .A1(n6501), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5979) );
  OAI211_X1 U7680 ( .C1(n6483), .C2(n9711), .A(n5980), .B(n5979), .ZN(n5981)
         );
  INV_X1 U7681 ( .A(n5981), .ZN(n5982) );
  XNOR2_X1 U7682 ( .A(n6586), .B(n8020), .ZN(n6009) );
  INV_X1 U7683 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7684 ( .A1(n5985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7685 ( .A1(n8226), .A2(n6569), .ZN(n6074) );
  INV_X1 U7686 ( .A(n5988), .ZN(n5992) );
  NAND2_X1 U7687 ( .A1(n5992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7688 ( .A1(n4343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  MUX2_X1 U7689 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5991), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5993) );
  INV_X1 U7690 ( .A(n7701), .ZN(n6532) );
  NAND2_X1 U7691 ( .A1(n7246), .A2(n6532), .ZN(n5994) );
  INV_X1 U7692 ( .A(n8031), .ZN(n5996) );
  NAND2_X1 U7693 ( .A1(n5996), .A2(n5995), .ZN(n6503) );
  INV_X1 U7694 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U7695 ( .A1(n5635), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7696 ( .A1(n5785), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5997) );
  OAI211_X1 U7697 ( .C1(n5999), .C2(n9620), .A(n5998), .B(n5997), .ZN(n6000)
         );
  INV_X1 U7698 ( .A(n6000), .ZN(n6001) );
  INV_X1 U7699 ( .A(n8023), .ZN(n8184) );
  NAND2_X1 U7700 ( .A1(n8184), .A2(n6593), .ZN(n6345) );
  INV_X1 U7701 ( .A(n6003), .ZN(n6004) );
  OR2_X1 U7702 ( .A1(n6002), .A2(n8227), .ZN(n6005) );
  NAND2_X1 U7703 ( .A1(n6005), .A2(n6607), .ZN(n6823) );
  INV_X1 U7704 ( .A(n6823), .ZN(n6824) );
  NOR2_X1 U7705 ( .A1(n6345), .A2(n6824), .ZN(n6007) );
  NOR2_X2 U7706 ( .A1(n6823), .A2(n6605), .ZN(n8457) );
  NAND2_X1 U7707 ( .A1(n7246), .A2(n7701), .ZN(n6818) );
  NAND2_X1 U7708 ( .A1(n7843), .A2(n6818), .ZN(n6011) );
  NAND2_X1 U7709 ( .A1(n6010), .A2(n6011), .ZN(n6051) );
  INV_X1 U7710 ( .A(n6051), .ZN(n6012) );
  INV_X1 U7711 ( .A(n7247), .ZN(n6013) );
  INV_X1 U7712 ( .A(n7967), .ZN(n6896) );
  NAND2_X1 U7713 ( .A1(n6016), .A2(n6352), .ZN(n6973) );
  NAND2_X1 U7714 ( .A1(n6973), .A2(n6017), .ZN(n7009) );
  INV_X1 U7715 ( .A(n7011), .ZN(n7008) );
  NAND2_X1 U7716 ( .A1(n7009), .A2(n7008), .ZN(n7426) );
  NAND2_X1 U7717 ( .A1(n7114), .A2(n6018), .ZN(n7425) );
  AND2_X1 U7718 ( .A1(n7425), .A2(n6390), .ZN(n6361) );
  NAND2_X1 U7719 ( .A1(n7426), .A2(n6361), .ZN(n7472) );
  NAND2_X1 U7720 ( .A1(n8201), .A2(n10072), .ZN(n6366) );
  NAND2_X1 U7721 ( .A1(n7424), .A2(n6390), .ZN(n7473) );
  NAND3_X1 U7722 ( .A1(n7472), .A2(n7480), .A3(n7473), .ZN(n7474) );
  NAND2_X1 U7723 ( .A1(n8200), .A2(n10081), .ZN(n6386) );
  NAND2_X1 U7724 ( .A1(n7406), .A2(n6386), .ZN(n7373) );
  NAND2_X1 U7725 ( .A1(n7465), .A2(n10085), .ZN(n6350) );
  AND2_X1 U7726 ( .A1(n7406), .A2(n6350), .ZN(n6392) );
  OR2_X1 U7727 ( .A1(n7465), .A2(n10085), .ZN(n6393) );
  NAND2_X1 U7728 ( .A1(n7589), .A2(n7588), .ZN(n7587) );
  INV_X1 U7729 ( .A(n8199), .ZN(n7516) );
  OR2_X1 U7730 ( .A1(n10093), .A2(n7516), .ZN(n6371) );
  NAND2_X1 U7731 ( .A1(n7682), .A2(n6373), .ZN(n7718) );
  INV_X1 U7732 ( .A(n8196), .ZN(n7864) );
  NAND2_X1 U7733 ( .A1(n7799), .A2(n7864), .ZN(n6382) );
  INV_X1 U7734 ( .A(n8195), .ZN(n7914) );
  NAND2_X1 U7735 ( .A1(n7868), .A2(n7914), .ZN(n6401) );
  OR2_X1 U7736 ( .A1(n7868), .A2(n7914), .ZN(n6020) );
  XNOR2_X1 U7737 ( .A(n7929), .B(n7983), .ZN(n7918) );
  OR2_X1 U7738 ( .A1(n7929), .A2(n7983), .ZN(n6403) );
  NAND2_X1 U7739 ( .A1(n7916), .A2(n6403), .ZN(n7936) );
  NOR2_X1 U7740 ( .A1(n8133), .A2(n7986), .ZN(n6022) );
  OAI22_X1 U7741 ( .A1(n7936), .A2(n6022), .B1(n8603), .B2(n8458), .ZN(n8469)
         );
  INV_X1 U7742 ( .A(n8469), .ZN(n6024) );
  NAND2_X1 U7743 ( .A1(n8461), .A2(n8443), .ZN(n6411) );
  NAND2_X1 U7744 ( .A1(n6412), .A2(n6411), .ZN(n8468) );
  INV_X1 U7745 ( .A(n8468), .ZN(n6023) );
  NAND2_X1 U7746 ( .A1(n8423), .A2(n6419), .ZN(n6025) );
  INV_X1 U7747 ( .A(n8413), .ZN(n8386) );
  NAND2_X1 U7748 ( .A1(n8145), .A2(n8386), .ZN(n6514) );
  NAND2_X1 U7749 ( .A1(n6026), .A2(n6515), .ZN(n8396) );
  NAND2_X1 U7750 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  NAND2_X1 U7751 ( .A1(n8397), .A2(n6431), .ZN(n8373) );
  INV_X1 U7752 ( .A(n6430), .ZN(n6027) );
  OAI21_X1 U7753 ( .B1(n8360), .B2(n4530), .A(n6436), .ZN(n8348) );
  NAND2_X1 U7754 ( .A1(n8348), .A2(n6438), .ZN(n6028) );
  NAND2_X1 U7755 ( .A1(n5935), .A2(n8342), .ZN(n6512) );
  NAND2_X1 U7756 ( .A1(n8059), .A2(n8354), .ZN(n8332) );
  AND2_X1 U7757 ( .A1(n6512), .A2(n8332), .ZN(n6445) );
  NAND2_X1 U7758 ( .A1(n6029), .A2(n6513), .ZN(n8324) );
  NAND2_X1 U7759 ( .A1(n8077), .A2(n8329), .ZN(n6451) );
  NOR2_X1 U7760 ( .A1(n8167), .A2(n8320), .ZN(n6450) );
  OR2_X1 U7761 ( .A1(n8553), .A2(n8310), .ZN(n6537) );
  INV_X1 U7762 ( .A(n8020), .ZN(n6031) );
  NOR2_X1 U7763 ( .A1(n8287), .A2(n6033), .ZN(n6080) );
  OR2_X1 U7764 ( .A1(n6042), .A2(n6035), .ZN(n6036) );
  NAND2_X1 U7765 ( .A1(n6037), .A2(n6036), .ZN(n6048) );
  XNOR2_X1 U7766 ( .A(n6048), .B(P2_B_REG_SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7767 ( .A1(n6040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7768 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  INV_X1 U7769 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6628) );
  AND2_X1 U7770 ( .A1(n6045), .A2(n6066), .ZN(n6046) );
  INV_X1 U7771 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U7772 ( .A1(n6047), .A2(n6625), .ZN(n6050) );
  NAND2_X1 U7773 ( .A1(n6066), .A2(n6048), .ZN(n6049) );
  NOR2_X1 U7774 ( .A1(n6821), .A2(n6827), .ZN(n6053) );
  OR2_X1 U7775 ( .A1(n6051), .A2(n7701), .ZN(n6052) );
  MUX2_X1 U7776 ( .A(n6943), .B(n6053), .S(n6940), .Z(n6071) );
  INV_X1 U7777 ( .A(n6943), .ZN(n6054) );
  INV_X1 U7778 ( .A(n6047), .ZN(n6622) );
  NOR2_X1 U7779 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n6058) );
  NOR4_X1 U7780 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6057) );
  NOR4_X1 U7781 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6056) );
  NOR4_X1 U7782 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6055) );
  NAND4_X1 U7783 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n6064)
         );
  NOR4_X1 U7784 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6062) );
  NOR4_X1 U7785 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6061) );
  NOR4_X1 U7786 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6060) );
  NOR4_X1 U7787 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6059) );
  NAND4_X1 U7788 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n6063)
         );
  NOR2_X1 U7789 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  INV_X1 U7790 ( .A(n6048), .ZN(n6623) );
  NAND2_X1 U7791 ( .A1(n6068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7792 ( .A1(n6819), .A2(n6593), .ZN(n6834) );
  AND3_X1 U7793 ( .A1(n6830), .A2(n6839), .A3(n6834), .ZN(n6070) );
  NAND2_X1 U7794 ( .A1(n6072), .A2(n4892), .ZN(P2_U3487) );
  INV_X1 U7795 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7796 ( .A1(n6821), .A2(n6830), .ZN(n6073) );
  INV_X1 U7797 ( .A(n6839), .ZN(n6568) );
  NAND2_X1 U7798 ( .A1(n7782), .A2(n6532), .ZN(n6820) );
  NOR2_X1 U7799 ( .A1(n6593), .A2(n10095), .ZN(n6075) );
  NAND2_X1 U7800 ( .A1(n6076), .A2(n6075), .ZN(n6814) );
  NAND2_X1 U7801 ( .A1(n6814), .A2(n8464), .ZN(n6831) );
  NAND2_X1 U7802 ( .A1(n6822), .A2(n6831), .ZN(n6079) );
  INV_X1 U7803 ( .A(n6567), .ZN(n6937) );
  INV_X1 U7804 ( .A(n6076), .ZN(n6829) );
  NAND2_X1 U7805 ( .A1(n6830), .A2(n6839), .ZN(n6077) );
  OAI21_X1 U7806 ( .B1(n6937), .B2(n6829), .A(n6826), .ZN(n6078) );
  NAND2_X1 U7807 ( .A1(n6082), .A2(n4888), .ZN(P2_U3455) );
  NAND2_X1 U7808 ( .A1(n9053), .A2(n6220), .ZN(n6089) );
  OAI21_X1 U7809 ( .B1(n7182), .B2(n6086), .A(n6085), .ZN(n6087) );
  NAND2_X1 U7810 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  XNOR2_X1 U7811 ( .A(n6090), .B(n6295), .ZN(n6093) );
  NAND2_X1 U7812 ( .A1(n9053), .A2(n6311), .ZN(n6092) );
  OR2_X1 U7813 ( .A1(n6161), .A2(n8909), .ZN(n6091) );
  AND2_X1 U7814 ( .A1(n6092), .A2(n6091), .ZN(n6094) );
  NAND2_X1 U7815 ( .A1(n6093), .A2(n6094), .ZN(n6872) );
  INV_X1 U7816 ( .A(n6093), .ZN(n6096) );
  NAND2_X1 U7817 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  NAND2_X1 U7818 ( .A1(n6872), .A2(n6097), .ZN(n6867) );
  NAND2_X1 U7819 ( .A1(n6954), .A2(n6220), .ZN(n6099) );
  NAND2_X1 U7820 ( .A1(n6106), .A2(n6810), .ZN(n6098) );
  AND2_X1 U7821 ( .A1(n6099), .A2(n6098), .ZN(n6103) );
  INV_X1 U7822 ( .A(n6316), .ZN(n6604) );
  NAND2_X1 U7823 ( .A1(n6604), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7824 ( .A1(n6103), .A2(n6100), .ZN(n6809) );
  NAND2_X1 U7825 ( .A1(n6954), .A2(n6311), .ZN(n6102) );
  AOI22_X1 U7826 ( .A1(n6220), .A2(n6810), .B1(n6604), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7827 ( .A1(n6102), .A2(n6101), .ZN(n6808) );
  NAND2_X1 U7828 ( .A1(n6809), .A2(n6808), .ZN(n6105) );
  NAND2_X1 U7829 ( .A1(n6103), .A2(n6295), .ZN(n6104) );
  NAND2_X1 U7830 ( .A1(n6105), .A2(n6104), .ZN(n6868) );
  NAND2_X1 U7831 ( .A1(n6865), .A2(n6872), .ZN(n6116) );
  OAI22_X1 U7832 ( .A1(n7033), .A2(n6161), .B1(n6904), .B2(n6125), .ZN(n6107)
         );
  XNOR2_X1 U7833 ( .A(n6107), .B(n6295), .ZN(n6111) );
  OR2_X1 U7834 ( .A1(n7033), .A2(n6108), .ZN(n6110) );
  NAND2_X1 U7835 ( .A1(n4291), .A2(n7213), .ZN(n6109) );
  AND2_X1 U7836 ( .A1(n6110), .A2(n6109), .ZN(n6112) );
  NAND2_X1 U7837 ( .A1(n6111), .A2(n6112), .ZN(n6117) );
  INV_X1 U7838 ( .A(n6111), .ZN(n6114) );
  INV_X1 U7839 ( .A(n6112), .ZN(n6113) );
  NAND2_X1 U7840 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  AND2_X1 U7841 ( .A1(n6117), .A2(n6115), .ZN(n6874) );
  NAND2_X1 U7842 ( .A1(n6116), .A2(n6874), .ZN(n6875) );
  NAND2_X1 U7843 ( .A1(n6875), .A2(n6117), .ZN(n7031) );
  OAI22_X1 U7844 ( .A1(n6907), .A2(n6161), .B1(n7126), .B2(n6125), .ZN(n6118)
         );
  XNOR2_X1 U7845 ( .A(n6118), .B(n6295), .ZN(n6123) );
  OR2_X1 U7846 ( .A1(n6907), .A2(n6108), .ZN(n6120) );
  NAND2_X1 U7847 ( .A1(n4291), .A2(n7328), .ZN(n6119) );
  NAND2_X1 U7848 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  XNOR2_X1 U7849 ( .A(n6123), .B(n6121), .ZN(n7032) );
  NAND2_X1 U7850 ( .A1(n7031), .A2(n7032), .ZN(n7030) );
  INV_X1 U7851 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7852 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  INV_X2 U7853 ( .A(n6220), .ZN(n6161) );
  OAI22_X1 U7854 ( .A1(n7331), .A2(n6161), .B1(n7226), .B2(n6125), .ZN(n6127)
         );
  XNOR2_X1 U7855 ( .A(n6127), .B(n6126), .ZN(n6131) );
  OR2_X1 U7856 ( .A1(n7331), .A2(n6108), .ZN(n6129) );
  NAND2_X1 U7857 ( .A1(n4291), .A2(n6963), .ZN(n6128) );
  NAND2_X1 U7858 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  XNOR2_X1 U7859 ( .A(n6131), .B(n6130), .ZN(n7021) );
  NAND2_X1 U7860 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  NAND2_X1 U7861 ( .A1(n9049), .A2(n4291), .ZN(n6133) );
  OAI21_X1 U7862 ( .B1(n9870), .B2(n6125), .A(n6133), .ZN(n6134) );
  XNOR2_X1 U7863 ( .A(n6134), .B(n6295), .ZN(n7089) );
  OR2_X1 U7864 ( .A1(n9870), .A2(n6161), .ZN(n6136) );
  NAND2_X1 U7865 ( .A1(n9049), .A2(n6311), .ZN(n6135) );
  AND2_X1 U7866 ( .A1(n6136), .A2(n6135), .ZN(n6138) );
  NAND2_X1 U7867 ( .A1(n7089), .A2(n6138), .ZN(n6137) );
  INV_X1 U7868 ( .A(n7089), .ZN(n6139) );
  INV_X1 U7869 ( .A(n6138), .ZN(n7088) );
  NAND2_X1 U7870 ( .A1(n6139), .A2(n7088), .ZN(n6140) );
  NAND2_X1 U7871 ( .A1(n7302), .A2(n6219), .ZN(n6143) );
  OR2_X1 U7872 ( .A1(n7442), .A2(n6161), .ZN(n6142) );
  NAND2_X1 U7873 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  XNOR2_X1 U7874 ( .A(n6144), .B(n6295), .ZN(n6147) );
  NAND2_X1 U7875 ( .A1(n7302), .A2(n4291), .ZN(n6146) );
  OR2_X1 U7876 ( .A1(n7442), .A2(n6108), .ZN(n6145) );
  AND2_X1 U7877 ( .A1(n6146), .A2(n6145), .ZN(n6148) );
  NAND2_X1 U7878 ( .A1(n6147), .A2(n6148), .ZN(n6152) );
  INV_X1 U7879 ( .A(n6147), .ZN(n6150) );
  INV_X1 U7880 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7881 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  NAND2_X1 U7882 ( .A1(n6152), .A2(n6151), .ZN(n7296) );
  NAND2_X1 U7883 ( .A1(n7562), .A2(n6219), .ZN(n6154) );
  OR2_X1 U7884 ( .A1(n7619), .A2(n6161), .ZN(n6153) );
  NAND2_X1 U7885 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  XNOR2_X1 U7886 ( .A(n6155), .B(n6295), .ZN(n6157) );
  NOR2_X1 U7887 ( .A1(n7619), .A2(n6108), .ZN(n6156) );
  AOI21_X1 U7888 ( .B1(n7562), .B2(n4291), .A(n6156), .ZN(n6158) );
  NAND2_X1 U7889 ( .A1(n6157), .A2(n6158), .ZN(n7541) );
  INV_X1 U7890 ( .A(n6157), .ZN(n6160) );
  INV_X1 U7891 ( .A(n6158), .ZN(n6159) );
  NAND2_X1 U7892 ( .A1(n6160), .A2(n6159), .ZN(n7543) );
  NAND2_X1 U7893 ( .A1(n7613), .A2(n6219), .ZN(n6163) );
  OR2_X1 U7894 ( .A1(n7654), .A2(n6161), .ZN(n6162) );
  NAND2_X1 U7895 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  XNOR2_X1 U7896 ( .A(n6164), .B(n6295), .ZN(n6167) );
  NOR2_X1 U7897 ( .A1(n7654), .A2(n6108), .ZN(n6165) );
  AOI21_X1 U7898 ( .B1(n7613), .B2(n4291), .A(n6165), .ZN(n7616) );
  INV_X1 U7899 ( .A(n6166), .ZN(n6168) );
  NAND2_X1 U7900 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  NAND2_X1 U7901 ( .A1(n7511), .A2(n6219), .ZN(n6171) );
  OR2_X1 U7902 ( .A1(n7547), .A2(n6161), .ZN(n6170) );
  NAND2_X1 U7903 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  XNOR2_X1 U7904 ( .A(n6172), .B(n6126), .ZN(n6174) );
  NOR2_X1 U7905 ( .A1(n7547), .A2(n6108), .ZN(n6173) );
  AOI21_X1 U7906 ( .B1(n7511), .B2(n4291), .A(n6173), .ZN(n6175) );
  XNOR2_X1 U7907 ( .A(n6174), .B(n6175), .ZN(n7650) );
  INV_X1 U7908 ( .A(n6174), .ZN(n6176) );
  NAND2_X1 U7909 ( .A1(n7557), .A2(n6219), .ZN(n6178) );
  OR2_X1 U7910 ( .A1(n7656), .A2(n6161), .ZN(n6177) );
  NAND2_X1 U7911 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  XNOR2_X1 U7912 ( .A(n6179), .B(n6126), .ZN(n6181) );
  NOR2_X1 U7913 ( .A1(n7656), .A2(n6108), .ZN(n6180) );
  AOI21_X1 U7914 ( .B1(n7557), .B2(n4291), .A(n6180), .ZN(n7804) );
  INV_X1 U7915 ( .A(n6181), .ZN(n6182) );
  NAND2_X1 U7916 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  NAND2_X1 U7917 ( .A1(n7877), .A2(n6219), .ZN(n6186) );
  OR2_X1 U7918 ( .A1(n7807), .A2(n6161), .ZN(n6185) );
  NAND2_X1 U7919 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  XNOR2_X1 U7920 ( .A(n6187), .B(n6126), .ZN(n6189) );
  NOR2_X1 U7921 ( .A1(n7807), .A2(n6108), .ZN(n6188) );
  AOI21_X1 U7922 ( .B1(n7877), .B2(n4291), .A(n6188), .ZN(n6190) );
  XNOR2_X1 U7923 ( .A(n6189), .B(n6190), .ZN(n7872) );
  INV_X1 U7924 ( .A(n6189), .ZN(n6191) );
  NAND2_X1 U7925 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  NAND2_X1 U7926 ( .A1(n7947), .A2(n6219), .ZN(n6194) );
  OR2_X1 U7927 ( .A1(n7875), .A2(n6161), .ZN(n6193) );
  NAND2_X1 U7928 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  XNOR2_X1 U7929 ( .A(n6195), .B(n6126), .ZN(n6197) );
  NOR2_X1 U7930 ( .A1(n7875), .A2(n6108), .ZN(n6196) );
  AOI21_X1 U7931 ( .B1(n7947), .B2(n4291), .A(n6196), .ZN(n6198) );
  XNOR2_X1 U7932 ( .A(n6197), .B(n6198), .ZN(n7943) );
  NAND2_X1 U7933 ( .A1(n7942), .A2(n7943), .ZN(n6201) );
  INV_X1 U7934 ( .A(n6197), .ZN(n6199) );
  NAND2_X1 U7935 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  NAND2_X1 U7936 ( .A1(n6201), .A2(n6200), .ZN(n8710) );
  NAND2_X1 U7937 ( .A1(n8716), .A2(n6219), .ZN(n6203) );
  OR2_X1 U7938 ( .A1(n8626), .A2(n6161), .ZN(n6202) );
  NAND2_X1 U7939 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  XNOR2_X1 U7940 ( .A(n6204), .B(n6126), .ZN(n6206) );
  NOR2_X1 U7941 ( .A1(n8626), .A2(n6108), .ZN(n6205) );
  AOI21_X1 U7942 ( .B1(n8716), .B2(n4291), .A(n6205), .ZN(n6207) );
  XNOR2_X1 U7943 ( .A(n6206), .B(n6207), .ZN(n8711) );
  NAND2_X1 U7944 ( .A1(n8710), .A2(n8711), .ZN(n6210) );
  INV_X1 U7945 ( .A(n6206), .ZN(n6208) );
  NAND2_X1 U7946 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X2 U7947 ( .A1(n6210), .A2(n6209), .ZN(n6217) );
  NAND2_X1 U7948 ( .A1(n7708), .A2(n6219), .ZN(n6212) );
  OR2_X1 U7949 ( .A1(n8714), .A2(n6161), .ZN(n6211) );
  NAND2_X1 U7950 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  XNOR2_X1 U7951 ( .A(n6213), .B(n6126), .ZN(n6215) );
  NOR2_X1 U7952 ( .A1(n8714), .A2(n6108), .ZN(n6214) );
  AOI21_X1 U7953 ( .B1(n7708), .B2(n4291), .A(n6214), .ZN(n8623) );
  INV_X1 U7954 ( .A(n6215), .ZN(n6216) );
  NAND2_X1 U7955 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  NAND2_X1 U7956 ( .A1(n8676), .A2(n6219), .ZN(n6222) );
  OR2_X1 U7957 ( .A1(n8763), .A2(n6161), .ZN(n6221) );
  NAND2_X1 U7958 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  XNOR2_X1 U7959 ( .A(n6223), .B(n6126), .ZN(n8668) );
  NAND2_X1 U7960 ( .A1(n8676), .A2(n4291), .ZN(n6225) );
  OR2_X1 U7961 ( .A1(n8763), .A2(n6108), .ZN(n6224) );
  NAND2_X1 U7962 ( .A1(n6225), .A2(n6224), .ZN(n6230) );
  XNOR2_X1 U7963 ( .A(n6226), .B(n6126), .ZN(n6231) );
  OR2_X1 U7964 ( .A1(n8830), .A2(n6161), .ZN(n6228) );
  OR2_X1 U7965 ( .A1(n8673), .A2(n6108), .ZN(n6227) );
  NAND2_X1 U7966 ( .A1(n6228), .A2(n6227), .ZN(n8756) );
  OAI22_X1 U7967 ( .A1(n8668), .A2(n6230), .B1(n6231), .B2(n8756), .ZN(n6235)
         );
  INV_X1 U7968 ( .A(n8756), .ZN(n6229) );
  INV_X1 U7969 ( .A(n6230), .ZN(n8667) );
  AND2_X1 U7970 ( .A1(n6230), .A2(n8756), .ZN(n6232) );
  AOI22_X1 U7971 ( .A1(n6233), .A2(n8668), .B1(n6232), .B2(n6231), .ZN(n6234)
         );
  NAND2_X1 U7972 ( .A1(n9379), .A2(n6219), .ZN(n6237) );
  NAND2_X1 U7973 ( .A1(n9473), .A2(n4291), .ZN(n6236) );
  NAND2_X1 U7974 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  XNOR2_X1 U7975 ( .A(n6238), .B(n6126), .ZN(n6241) );
  NAND2_X1 U7976 ( .A1(n9379), .A2(n4291), .ZN(n6240) );
  NAND2_X1 U7977 ( .A1(n9473), .A2(n6311), .ZN(n6239) );
  NAND2_X1 U7978 ( .A1(n6240), .A2(n6239), .ZN(n6242) );
  AND2_X1 U7979 ( .A1(n6241), .A2(n6242), .ZN(n8681) );
  INV_X1 U7980 ( .A(n6241), .ZN(n6244) );
  INV_X1 U7981 ( .A(n6242), .ZN(n6243) );
  NAND2_X1 U7982 ( .A1(n6244), .A2(n6243), .ZN(n8680) );
  NAND2_X1 U7983 ( .A1(n9338), .A2(n6219), .ZN(n6246) );
  NAND2_X1 U7984 ( .A1(n9476), .A2(n4291), .ZN(n6245) );
  NAND2_X1 U7985 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  XNOR2_X1 U7986 ( .A(n6247), .B(n6126), .ZN(n8644) );
  NAND2_X1 U7987 ( .A1(n9338), .A2(n4291), .ZN(n6249) );
  NAND2_X1 U7988 ( .A1(n9476), .A2(n6311), .ZN(n6248) );
  NAND2_X1 U7989 ( .A1(n6249), .A2(n6248), .ZN(n6256) );
  NAND2_X1 U7990 ( .A1(n9347), .A2(n4291), .ZN(n6251) );
  NAND2_X1 U7991 ( .A1(n9464), .A2(n6311), .ZN(n6250) );
  NAND2_X1 U7992 ( .A1(n6251), .A2(n6250), .ZN(n8734) );
  NAND2_X1 U7993 ( .A1(n9347), .A2(n6219), .ZN(n6253) );
  NAND2_X1 U7994 ( .A1(n9464), .A2(n4291), .ZN(n6252) );
  NAND2_X1 U7995 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  XNOR2_X1 U7996 ( .A(n6254), .B(n6126), .ZN(n8640) );
  OAI22_X1 U7997 ( .A1(n8644), .A2(n6256), .B1(n8734), .B2(n8640), .ZN(n6260)
         );
  NAND2_X1 U7998 ( .A1(n8640), .A2(n8734), .ZN(n6255) );
  INV_X1 U7999 ( .A(n6256), .ZN(n8643) );
  NAND2_X1 U8000 ( .A1(n6255), .A2(n8643), .ZN(n6258) );
  INV_X1 U8001 ( .A(n6255), .ZN(n6257) );
  AOI22_X1 U8002 ( .A1(n8644), .A2(n6258), .B1(n6257), .B2(n6256), .ZN(n6259)
         );
  OAI22_X1 U8003 ( .A1(n9535), .A2(n6125), .B1(n9336), .B2(n6161), .ZN(n6261)
         );
  XNOR2_X1 U8004 ( .A(n6261), .B(n6295), .ZN(n8701) );
  OR2_X1 U8005 ( .A1(n9535), .A2(n6161), .ZN(n6263) );
  OR2_X1 U8006 ( .A1(n9336), .A2(n6108), .ZN(n6262) );
  NAND2_X1 U8007 ( .A1(n6263), .A2(n6262), .ZN(n8700) );
  INV_X1 U8008 ( .A(n8700), .ZN(n6264) );
  INV_X1 U8009 ( .A(n8701), .ZN(n6265) );
  NAND2_X1 U8010 ( .A1(n9310), .A2(n6219), .ZN(n6267) );
  NAND2_X1 U8011 ( .A1(n9440), .A2(n4291), .ZN(n6266) );
  NAND2_X1 U8012 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  XNOR2_X1 U8013 ( .A(n6268), .B(n6295), .ZN(n6271) );
  AND2_X1 U8014 ( .A1(n9440), .A2(n6311), .ZN(n6269) );
  AOI21_X1 U8015 ( .B1(n9310), .B2(n4291), .A(n6269), .ZN(n6270) );
  XNOR2_X1 U8016 ( .A(n6271), .B(n6270), .ZN(n8653) );
  OAI22_X1 U8017 ( .A1(n9443), .A2(n6125), .B1(n9308), .B2(n6161), .ZN(n6272)
         );
  XNOR2_X1 U8018 ( .A(n6272), .B(n6126), .ZN(n8719) );
  OAI22_X1 U8019 ( .A1(n9443), .A2(n6161), .B1(n9308), .B2(n6108), .ZN(n8723)
         );
  OAI22_X1 U8020 ( .A1(n9435), .A2(n6125), .B1(n9291), .B2(n6161), .ZN(n6273)
         );
  XNOR2_X1 U8021 ( .A(n6273), .B(n6295), .ZN(n6276) );
  OR2_X1 U8022 ( .A1(n9435), .A2(n6161), .ZN(n6275) );
  NAND2_X1 U8023 ( .A1(n9441), .A2(n6311), .ZN(n6274) );
  AND2_X1 U8024 ( .A1(n6275), .A2(n6274), .ZN(n6277) );
  NAND2_X1 U8025 ( .A1(n6276), .A2(n6277), .ZN(n8691) );
  INV_X1 U8026 ( .A(n6276), .ZN(n6279) );
  INV_X1 U8027 ( .A(n6277), .ZN(n6278) );
  NAND2_X1 U8028 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  AND2_X1 U8029 ( .A1(n8691), .A2(n6280), .ZN(n8633) );
  NAND2_X1 U8030 ( .A1(n9426), .A2(n6219), .ZN(n6282) );
  NAND2_X1 U8031 ( .A1(n9432), .A2(n4291), .ZN(n6281) );
  NAND2_X1 U8032 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  XNOR2_X1 U8033 ( .A(n6283), .B(n6295), .ZN(n6285) );
  AND2_X1 U8034 ( .A1(n9432), .A2(n6311), .ZN(n6284) );
  AOI21_X1 U8035 ( .B1(n9426), .B2(n4291), .A(n6284), .ZN(n6286) );
  NAND2_X1 U8036 ( .A1(n6285), .A2(n6286), .ZN(n6290) );
  INV_X1 U8037 ( .A(n6285), .ZN(n6288) );
  INV_X1 U8038 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U8039 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  NAND2_X1 U8040 ( .A1(n6290), .A2(n6289), .ZN(n8690) );
  INV_X1 U8041 ( .A(n6290), .ZN(n6291) );
  OAI22_X1 U8042 ( .A1(n9420), .A2(n6125), .B1(n9263), .B2(n6161), .ZN(n6292)
         );
  XNOR2_X1 U8043 ( .A(n6292), .B(n6126), .ZN(n6299) );
  OAI22_X1 U8044 ( .A1(n9420), .A2(n6161), .B1(n9263), .B2(n6108), .ZN(n6298)
         );
  XNOR2_X1 U8045 ( .A(n6299), .B(n6298), .ZN(n8658) );
  NAND2_X1 U8046 ( .A1(n9230), .A2(n6219), .ZN(n6294) );
  NAND2_X1 U8047 ( .A1(n9417), .A2(n4291), .ZN(n6293) );
  NAND2_X1 U8048 ( .A1(n6294), .A2(n6293), .ZN(n6296) );
  XNOR2_X1 U8049 ( .A(n6296), .B(n6295), .ZN(n6300) );
  NOR2_X1 U8050 ( .A1(n9244), .A2(n6108), .ZN(n6297) );
  AOI21_X1 U8051 ( .B1(n9230), .B2(n4291), .A(n6297), .ZN(n6301) );
  XNOR2_X1 U8052 ( .A(n6300), .B(n6301), .ZN(n8742) );
  NOR2_X1 U8053 ( .A1(n6299), .A2(n6298), .ZN(n8743) );
  INV_X1 U8054 ( .A(n6300), .ZN(n6303) );
  INV_X1 U8055 ( .A(n6301), .ZN(n6302) );
  AOI22_X1 U8056 ( .A1(n9208), .A2(n6219), .B1(n4291), .B2(n9409), .ZN(n6304)
         );
  XNOR2_X1 U8057 ( .A(n6304), .B(n6126), .ZN(n6306) );
  AOI22_X1 U8058 ( .A1(n9208), .A2(n4291), .B1(n6311), .B2(n9409), .ZN(n6305)
         );
  NAND2_X1 U8059 ( .A1(n6306), .A2(n6305), .ZN(n6335) );
  OAI21_X1 U8060 ( .B1(n6306), .B2(n6305), .A(n6335), .ZN(n6574) );
  INV_X1 U8061 ( .A(n6574), .ZN(n6307) );
  NAND2_X1 U8062 ( .A1(n9193), .A2(n6219), .ZN(n6309) );
  NAND2_X1 U8063 ( .A1(n9400), .A2(n4291), .ZN(n6308) );
  NAND2_X1 U8064 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  XNOR2_X1 U8065 ( .A(n6310), .B(n6126), .ZN(n6313) );
  AOI22_X1 U8066 ( .A1(n9193), .A2(n4291), .B1(n6311), .B2(n9400), .ZN(n6312)
         );
  XNOR2_X1 U8067 ( .A(n6313), .B(n6312), .ZN(n6318) );
  INV_X1 U8068 ( .A(n6318), .ZN(n6336) );
  INV_X1 U8069 ( .A(n6314), .ZN(n7134) );
  NAND3_X1 U8070 ( .A1(n6315), .A2(n7134), .A3(n7131), .ZN(n6329) );
  INV_X1 U8071 ( .A(n9550), .ZN(n6631) );
  OR2_X1 U8072 ( .A1(n6329), .A2(n6631), .ZN(n6320) );
  OR2_X1 U8073 ( .A1(n9427), .A2(n9013), .ZN(n6327) );
  NAND3_X1 U8074 ( .A1(n6336), .A2(n8746), .A3(n6335), .ZN(n6317) );
  INV_X1 U8075 ( .A(n6320), .ZN(n6324) );
  OR2_X1 U8076 ( .A1(n6958), .A2(n9018), .ZN(n7136) );
  INV_X1 U8077 ( .A(n7136), .ZN(n6323) );
  INV_X1 U8078 ( .A(n6321), .ZN(n6322) );
  INV_X1 U8079 ( .A(n6325), .ZN(n7140) );
  NAND2_X1 U8080 ( .A1(n9550), .A2(n7140), .ZN(n9033) );
  NAND2_X1 U8081 ( .A1(n6326), .A2(n5509), .ZN(n8762) );
  NAND2_X1 U8082 ( .A1(n9392), .A2(n8751), .ZN(n6334) );
  INV_X1 U8083 ( .A(n9195), .ZN(n6332) );
  NAND3_X1 U8084 ( .A1(n9033), .A2(n6327), .A3(n7136), .ZN(n6328) );
  NAND2_X1 U8085 ( .A1(n6329), .A2(n6328), .ZN(n6331) );
  INV_X1 U8086 ( .A(n7130), .ZN(n6330) );
  NAND2_X1 U8087 ( .A1(n6331), .A2(n6330), .ZN(n6811) );
  AOI22_X1 U8088 ( .A1(n6332), .A2(n8759), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6333) );
  OAI211_X1 U8089 ( .C1(n9228), .C2(n8736), .A(n6334), .B(n6333), .ZN(n6338)
         );
  NOR3_X1 U8090 ( .A1(n6336), .A2(n8768), .A3(n6335), .ZN(n6337) );
  AOI211_X1 U8091 ( .C1(n9193), .C2(n8765), .A(n6338), .B(n6337), .ZN(n6339)
         );
  NAND3_X1 U8092 ( .A1(n6341), .A2(n6340), .A3(n6339), .ZN(P1_U3220) );
  INV_X1 U8093 ( .A(n8298), .ZN(n6584) );
  NAND2_X1 U8094 ( .A1(n6342), .A2(n6500), .ZN(n6344) );
  NAND2_X1 U8095 ( .A1(n5674), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6343) );
  OAI21_X1 U8096 ( .B1(n8033), .B2(n6605), .A(n6588), .ZN(n6346) );
  INV_X1 U8097 ( .A(n6458), .ZN(n6462) );
  MUX2_X1 U8098 ( .A(n8298), .B(n8027), .S(n6605), .Z(n6464) );
  MUX2_X1 U8099 ( .A(n4319), .B(n6450), .S(n6593), .Z(n6347) );
  NOR2_X1 U8100 ( .A1(n8295), .A2(n6347), .ZN(n6461) );
  NAND2_X1 U8101 ( .A1(n6373), .A2(n6372), .ZN(n6349) );
  NAND2_X1 U8102 ( .A1(n6376), .A2(n6375), .ZN(n6348) );
  NOR2_X1 U8103 ( .A1(n6378), .A2(n5737), .ZN(n6394) );
  INV_X1 U8104 ( .A(n6350), .ZN(n6370) );
  MUX2_X1 U8105 ( .A(n6351), .B(n6017), .S(n6593), .Z(n6358) );
  NAND2_X1 U8106 ( .A1(n6978), .A2(n6896), .ZN(n6520) );
  OAI211_X1 U8107 ( .C1(n6352), .C2(n7246), .A(n6520), .B(n6605), .ZN(n6356)
         );
  INV_X1 U8108 ( .A(n6520), .ZN(n6354) );
  NAND2_X1 U8109 ( .A1(n6017), .A2(n6605), .ZN(n6353) );
  NAND2_X1 U8110 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  NAND3_X1 U8111 ( .A1(n6358), .A2(n6357), .A3(n7008), .ZN(n6364) );
  NAND2_X1 U8112 ( .A1(n6359), .A2(n7973), .ZN(n6360) );
  AND2_X1 U8113 ( .A1(n6366), .A2(n6360), .ZN(n6362) );
  MUX2_X1 U8114 ( .A(n6362), .B(n6361), .S(n6605), .Z(n6363) );
  NAND2_X1 U8115 ( .A1(n6364), .A2(n6363), .ZN(n6365) );
  NAND2_X1 U8116 ( .A1(n6365), .A2(n7480), .ZN(n6385) );
  INV_X1 U8117 ( .A(n6366), .ZN(n6368) );
  OAI211_X1 U8118 ( .C1(n6385), .C2(n6368), .A(n6392), .B(n6367), .ZN(n6369)
         );
  OAI211_X1 U8119 ( .C1(n6370), .C2(n6386), .A(n6369), .B(n6393), .ZN(n6381)
         );
  AOI21_X1 U8120 ( .B1(n6372), .B2(n6371), .A(n6378), .ZN(n6374) );
  AOI21_X1 U8121 ( .B1(n7516), .B2(n10093), .A(n6019), .ZN(n6377) );
  OAI211_X1 U8122 ( .C1(n6378), .C2(n6377), .A(n6382), .B(n6376), .ZN(n6379)
         );
  INV_X1 U8123 ( .A(n6382), .ZN(n6383) );
  INV_X1 U8124 ( .A(n6384), .ZN(n6399) );
  INV_X1 U8125 ( .A(n6385), .ZN(n6391) );
  INV_X1 U8126 ( .A(n6386), .ZN(n6389) );
  INV_X1 U8127 ( .A(n6387), .ZN(n6388) );
  AOI211_X1 U8128 ( .C1(n6391), .C2(n6390), .A(n6389), .B(n6388), .ZN(n6396)
         );
  INV_X1 U8129 ( .A(n6392), .ZN(n6395) );
  OAI211_X1 U8130 ( .C1(n6396), .C2(n6395), .A(n6394), .B(n6393), .ZN(n6398)
         );
  AOI21_X1 U8131 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6400) );
  OR2_X1 U8132 ( .A1(n7918), .A2(n7861), .ZN(n6519) );
  INV_X1 U8133 ( .A(n6401), .ZN(n6402) );
  AOI22_X1 U8134 ( .A1(n6403), .A2(n6402), .B1(n7983), .B2(n7929), .ZN(n6404)
         );
  NAND2_X1 U8135 ( .A1(n6519), .A2(n6404), .ZN(n6405) );
  MUX2_X1 U8136 ( .A(n6405), .B(n6404), .S(n6605), .Z(n6406) );
  MUX2_X1 U8137 ( .A(n7986), .B(n8603), .S(n6593), .Z(n6408) );
  INV_X1 U8138 ( .A(n6408), .ZN(n6407) );
  NAND2_X1 U8139 ( .A1(n6407), .A2(n6516), .ZN(n6409) );
  AOI22_X1 U8140 ( .A1(n6410), .A2(n6409), .B1(n6408), .B2(n4597), .ZN(n6414)
         );
  MUX2_X1 U8141 ( .A(n6412), .B(n6411), .S(n6605), .Z(n6413) );
  OAI21_X1 U8142 ( .B1(n6414), .B2(n8468), .A(n6413), .ZN(n6415) );
  MUX2_X1 U8143 ( .A(n6417), .B(n6416), .S(n6605), .Z(n6418) );
  MUX2_X1 U8144 ( .A(n6420), .B(n6419), .S(n6593), .Z(n6421) );
  NAND3_X1 U8145 ( .A1(n6423), .A2(n6427), .A3(n6434), .ZN(n6424) );
  NAND3_X1 U8146 ( .A1(n6424), .A2(n6436), .A3(n6430), .ZN(n6425) );
  NAND2_X1 U8147 ( .A1(n6515), .A2(n6426), .ZN(n6428) );
  OAI211_X1 U8148 ( .C1(n6429), .C2(n6428), .A(n6427), .B(n6514), .ZN(n6432)
         );
  NAND3_X1 U8149 ( .A1(n6432), .A2(n6431), .A3(n6430), .ZN(n6435) );
  NAND3_X1 U8150 ( .A1(n6435), .A2(n6434), .A3(n6433), .ZN(n6437) );
  MUX2_X1 U8151 ( .A(n6439), .B(n6438), .S(n6593), .Z(n6441) );
  INV_X1 U8152 ( .A(n8332), .ZN(n6440) );
  INV_X1 U8153 ( .A(n6442), .ZN(n6443) );
  NAND2_X1 U8154 ( .A1(n6513), .A2(n6443), .ZN(n6444) );
  OAI21_X1 U8155 ( .B1(n6447), .B2(n6444), .A(n6512), .ZN(n6449) );
  INV_X1 U8156 ( .A(n6445), .ZN(n6446) );
  OAI21_X1 U8157 ( .B1(n6447), .B2(n6446), .A(n6513), .ZN(n6448) );
  MUX2_X1 U8158 ( .A(n6449), .B(n6448), .S(n6593), .Z(n6455) );
  NAND2_X1 U8159 ( .A1(n6452), .A2(n6451), .ZN(n8323) );
  INV_X1 U8160 ( .A(n8311), .ZN(n6454) );
  MUX2_X1 U8161 ( .A(n6452), .B(n6451), .S(n6593), .Z(n6453) );
  NOR2_X1 U8162 ( .A1(n8310), .A2(n6593), .ZN(n6457) );
  NOR2_X1 U8163 ( .A1(n8185), .A2(n6605), .ZN(n6456) );
  MUX2_X1 U8164 ( .A(n6457), .B(n6456), .S(n8553), .Z(n6459) );
  NAND2_X1 U8165 ( .A1(n6463), .A2(n8023), .ZN(n6587) );
  INV_X1 U8166 ( .A(n6587), .ZN(n6467) );
  NAND2_X1 U8167 ( .A1(n6465), .A2(n6464), .ZN(n6488) );
  INV_X1 U8168 ( .A(n6488), .ZN(n6466) );
  INV_X1 U8169 ( .A(SI_29_), .ZN(n6468) );
  INV_X1 U8170 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9561) );
  INV_X1 U8171 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6474) );
  MUX2_X1 U8172 ( .A(n9561), .B(n6474), .S(n5058), .Z(n6476) );
  INV_X1 U8173 ( .A(SI_30_), .ZN(n6475) );
  NAND2_X1 U8174 ( .A1(n6476), .A2(n6475), .ZN(n6492) );
  INV_X1 U8175 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U8176 ( .A1(n6477), .A2(SI_30_), .ZN(n6478) );
  NAND2_X1 U8177 ( .A1(n6492), .A2(n6478), .ZN(n6493) );
  NAND2_X1 U8178 ( .A1(n8879), .A2(n6500), .ZN(n6480) );
  NAND2_X1 U8179 ( .A1(n5674), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8180 ( .A1(n6480), .A2(n6479), .ZN(n6541) );
  INV_X1 U8181 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U8182 ( .A1(n5785), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8183 ( .A1(n6501), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6481) );
  OAI211_X1 U8184 ( .C1(n9710), .C2(n6483), .A(n6482), .B(n6481), .ZN(n6484)
         );
  INV_X1 U8185 ( .A(n6484), .ZN(n6485) );
  NAND2_X1 U8186 ( .A1(n6503), .A2(n6485), .ZN(n8183) );
  INV_X1 U8187 ( .A(n8183), .ZN(n6491) );
  OR2_X1 U8188 ( .A1(n6541), .A2(n6491), .ZN(n6489) );
  INV_X1 U8189 ( .A(n6489), .ZN(n6546) );
  NOR2_X1 U8190 ( .A1(n6486), .A2(n6546), .ZN(n6490) );
  AND2_X1 U8191 ( .A1(n6541), .A2(n6491), .ZN(n6508) );
  INV_X1 U8192 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6496) );
  INV_X1 U8193 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U8194 ( .A(n6496), .B(n6495), .S(n5058), .Z(n6497) );
  XNOR2_X1 U8195 ( .A(n6497), .B(SI_31_), .ZN(n6498) );
  INV_X1 U8196 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U8197 ( .A1(n5635), .A2(P2_REG1_REG_31__SCAN_IN), .B1(n6501), .B2(
        P2_REG2_REG_31__SCAN_IN), .ZN(n6502) );
  OAI211_X1 U8198 ( .C1(n5646), .C2(n6504), .A(n6503), .B(n6502), .ZN(n8281)
         );
  AND2_X1 U8199 ( .A1(n8547), .A2(n8281), .ZN(n6507) );
  NOR2_X1 U8200 ( .A1(n8547), .A2(n8281), .ZN(n6551) );
  NOR3_X1 U8201 ( .A1(n6505), .A2(n6551), .A3(n6819), .ZN(n6566) );
  INV_X1 U8202 ( .A(n6551), .ZN(n6506) );
  NOR2_X1 U8203 ( .A1(n6506), .A2(n6010), .ZN(n6536) );
  INV_X1 U8204 ( .A(n6507), .ZN(n6511) );
  INV_X1 U8205 ( .A(n6508), .ZN(n6509) );
  AND2_X1 U8206 ( .A1(n6509), .A2(n6587), .ZN(n6510) );
  INV_X1 U8207 ( .A(n8340), .ZN(n6529) );
  INV_X1 U8208 ( .A(n6516), .ZN(n6517) );
  NAND2_X1 U8209 ( .A1(n6975), .A2(n6520), .ZN(n7968) );
  NAND4_X1 U8210 ( .A1(n6522), .A2(n7480), .A3(n6521), .A4(n7588), .ZN(n6523)
         );
  XNOR2_X1 U8211 ( .A(n7465), .B(n10085), .ZN(n7409) );
  NOR4_X1 U8212 ( .A1(n6523), .A2(n7675), .A3(n7409), .A4(n7583), .ZN(n6524)
         );
  XNOR2_X1 U8213 ( .A(n7799), .B(n8196), .ZN(n7720) );
  NAND4_X1 U8214 ( .A1(n7935), .A2(n4520), .A3(n6524), .A4(n7720), .ZN(n6525)
         );
  NOR4_X1 U8215 ( .A1(n8425), .A2(n8437), .A3(n8468), .A4(n6525), .ZN(n6526)
         );
  NAND4_X1 U8216 ( .A1(n8395), .A2(n4518), .A3(n8402), .A4(n6526), .ZN(n6527)
         );
  NOR3_X1 U8217 ( .A1(n8362), .A2(n4611), .A3(n6527), .ZN(n6528) );
  NAND4_X1 U8218 ( .A1(n6529), .A2(n8334), .A3(n8350), .A4(n6528), .ZN(n6530)
         );
  NOR4_X1 U8219 ( .A1(n8295), .A2(n8311), .A3(n8323), .A4(n6530), .ZN(n6531)
         );
  NAND4_X1 U8220 ( .A1(n6543), .A2(n4346), .A3(n6531), .A4(n8020), .ZN(n6552)
         );
  NAND2_X1 U8221 ( .A1(n6010), .A2(n6532), .ZN(n6549) );
  OR2_X1 U8222 ( .A1(n6549), .A2(n7246), .ZN(n6533) );
  NOR2_X1 U8223 ( .A1(n6552), .A2(n6534), .ZN(n6535) );
  NOR2_X1 U8224 ( .A1(n6536), .A2(n6535), .ZN(n6562) );
  INV_X1 U8225 ( .A(n8020), .ZN(n6538) );
  OR2_X1 U8226 ( .A1(n8295), .A2(n6538), .ZN(n6539) );
  INV_X1 U8227 ( .A(n6588), .ZN(n6544) );
  INV_X1 U8228 ( .A(n8547), .ZN(n6545) );
  INV_X1 U8229 ( .A(n6541), .ZN(n8550) );
  OR2_X1 U8230 ( .A1(n6545), .A2(n8550), .ZN(n6542) );
  OAI211_X1 U8231 ( .C1(n6592), .C2(n6544), .A(n6543), .B(n6542), .ZN(n6548)
         );
  NAND2_X1 U8232 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  NAND2_X1 U8233 ( .A1(n6548), .A2(n6547), .ZN(n6558) );
  INV_X1 U8234 ( .A(n6552), .ZN(n6554) );
  NOR2_X1 U8235 ( .A1(n6010), .A2(n7701), .ZN(n6557) );
  NAND2_X1 U8236 ( .A1(n6557), .A2(n7782), .ZN(n6553) );
  OAI22_X1 U8237 ( .A1(n6558), .A2(n6555), .B1(n6554), .B2(n6553), .ZN(n6556)
         );
  INV_X1 U8238 ( .A(n6556), .ZN(n6560) );
  NAND3_X1 U8239 ( .A1(n6558), .A2(n6557), .A3(n7246), .ZN(n6559) );
  NAND2_X1 U8240 ( .A1(n6563), .A2(n4901), .ZN(n6565) );
  OR2_X1 U8241 ( .A1(n6743), .A2(P2_U3151), .ZN(n7940) );
  INV_X1 U8242 ( .A(n7940), .ZN(n6564) );
  OAI21_X1 U8243 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6573) );
  NOR4_X1 U8244 ( .A1(n6568), .A2(n6004), .A3(n6567), .A4(n6002), .ZN(n6571)
         );
  OAI21_X1 U8245 ( .B1(n7940), .B2(n6569), .A(P2_B_REG_SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8246 ( .A1(n6573), .A2(n6572), .ZN(P2_U3296) );
  OAI21_X1 U8247 ( .B1(n6576), .B2(n6575), .A(n8746), .ZN(n6583) );
  INV_X1 U8248 ( .A(n9208), .ZN(n9402) );
  OAI22_X1 U8249 ( .A1(n9244), .A2(n8736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6577), .ZN(n6579) );
  NOR2_X1 U8250 ( .A1(n9212), .A2(n8762), .ZN(n6578) );
  AOI211_X1 U8251 ( .C1(n9209), .C2(n8759), .A(n6579), .B(n6578), .ZN(n6580)
         );
  NAND2_X1 U8252 ( .A1(n6583), .A2(n6582), .ZN(P1_U3214) );
  NAND2_X1 U8253 ( .A1(n8027), .A2(n8298), .ZN(n6585) );
  XNOR2_X1 U8254 ( .A(n6589), .B(n6590), .ZN(n6598) );
  NAND2_X1 U8255 ( .A1(n8036), .A2(n7721), .ZN(n6596) );
  NAND2_X1 U8256 ( .A1(n6607), .A2(P2_B_REG_SCAN_IN), .ZN(n6594) );
  AND2_X1 U8257 ( .A1(n8455), .A2(n6594), .ZN(n8280) );
  AOI22_X1 U8258 ( .A1(n8457), .A2(n8298), .B1(n8183), .B2(n8280), .ZN(n6595)
         );
  NAND2_X1 U8259 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  NAND2_X1 U8260 ( .A1(n6601), .A2(n4890), .ZN(P2_U3456) );
  NAND2_X1 U8261 ( .A1(n6602), .A2(n4889), .ZN(P2_U3488) );
  NAND2_X1 U8262 ( .A1(n6836), .A2(n6605), .ZN(n6606) );
  NAND2_X1 U8263 ( .A1(n6606), .A2(n6743), .ZN(n6746) );
  NAND2_X1 U8264 ( .A1(n6746), .A2(n6607), .ZN(n6608) );
  NAND2_X1 U8265 ( .A1(n6608), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U8266 ( .A(n9571), .ZN(n9565) );
  NAND2_X1 U8267 ( .A1(n5058), .A2(n4288), .ZN(n9568) );
  OAI222_X1 U8268 ( .A1(n9565), .A2(n6611), .B1(n9568), .B2(n4908), .C1(n4288), 
        .C2(n6685), .ZN(P1_U3354) );
  NOR2_X1 U8269 ( .A1(n5058), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8615) );
  INV_X1 U8270 ( .A(n8615), .ZN(n7954) );
  OAI222_X1 U8271 ( .A1(n6762), .A2(P2_U3151), .B1(n7954), .B2(n4713), .C1(
        n8618), .C2(n6611), .ZN(P2_U3294) );
  INV_X1 U8272 ( .A(n6795), .ZN(n6764) );
  OAI222_X1 U8273 ( .A1(n6764), .A2(P2_U3151), .B1(n8618), .B2(n6612), .C1(
        n4388), .C2(n7954), .ZN(P2_U3293) );
  OAI222_X1 U8274 ( .A1(n9568), .A2(n6613), .B1(n9565), .B2(n6612), .C1(
        P1_U3086), .C2(n6684), .ZN(P1_U3353) );
  OAI222_X1 U8275 ( .A1(n9568), .A2(n6614), .B1(n9565), .B2(n6616), .C1(n4288), 
        .C2(n6688), .ZN(P1_U3352) );
  INV_X1 U8276 ( .A(n6757), .ZN(n6990) );
  OAI222_X1 U8277 ( .A1(n6990), .A2(P2_U3151), .B1(n8618), .B2(n6616), .C1(
        n6615), .C2(n7954), .ZN(P2_U3292) );
  AOI22_X1 U8278 ( .A1(n6923), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n8615), .ZN(n6617) );
  OAI21_X1 U8279 ( .B1(n6618), .B2(n8618), .A(n6617), .ZN(P2_U3291) );
  OAI222_X1 U8280 ( .A1(n6619), .A2(n9568), .B1(P1_U3086), .B2(n6690), .C1(
        n9565), .C2(n6618), .ZN(P1_U3351) );
  INV_X1 U8281 ( .A(n6620), .ZN(n6630) );
  INV_X1 U8282 ( .A(n9568), .ZN(n9570) );
  AOI22_X1 U8283 ( .A1(n9097), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9570), .ZN(n6621) );
  OAI21_X1 U8284 ( .B1(n6630), .B2(n9565), .A(n6621), .ZN(P1_U3350) );
  NAND2_X1 U8285 ( .A1(n6622), .A2(n6839), .ZN(n6648) );
  NOR3_X1 U8286 ( .A1(n8616), .A2(n6626), .A3(n6623), .ZN(n6624) );
  AOI21_X1 U8287 ( .B1(n6648), .B2(n6625), .A(n6624), .ZN(P2_U3376) );
  NOR3_X1 U8288 ( .A1(n7959), .A2(n8616), .A3(n6626), .ZN(n6627) );
  AOI21_X1 U8289 ( .B1(n6648), .B2(n6628), .A(n6627), .ZN(P2_U3377) );
  OAI222_X1 U8290 ( .A1(n7049), .A2(P2_U3151), .B1(n8618), .B2(n6630), .C1(
        n6629), .C2(n7954), .ZN(P2_U3290) );
  OR2_X1 U8291 ( .A1(n6632), .A2(P1_U3086), .ZN(n9024) );
  NAND2_X1 U8292 ( .A1(n6631), .A2(n9024), .ZN(n6682) );
  NAND2_X1 U8293 ( .A1(n6632), .A2(n9013), .ZN(n6633) );
  AND2_X1 U8294 ( .A1(n6633), .A2(n8772), .ZN(n6681) );
  INV_X1 U8295 ( .A(n6681), .ZN(n6634) );
  AND2_X1 U8296 ( .A1(n6682), .A2(n6634), .ZN(n9827) );
  NOR2_X1 U8297 ( .A1(n9827), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8298 ( .A(n6635), .ZN(n6638) );
  AOI22_X1 U8299 ( .A1(n9110), .A2(P1_STATE_REG_SCAN_IN), .B1(n9570), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6636) );
  OAI21_X1 U8300 ( .B1(n6638), .B2(n9565), .A(n6636), .ZN(P1_U3349) );
  OAI222_X1 U8301 ( .A1(n7079), .A2(P2_U3151), .B1(n8618), .B2(n6638), .C1(
        n6637), .C2(n7954), .ZN(P2_U3289) );
  NAND2_X1 U8302 ( .A1(n6954), .A2(P1_U3973), .ZN(n6639) );
  OAI21_X1 U8303 ( .B1(P1_U3973), .B2(n4910), .A(n6639), .ZN(P1_U3554) );
  INV_X1 U8304 ( .A(n6640), .ZN(n6647) );
  AOI22_X1 U8305 ( .A1(n9123), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9570), .ZN(n6641) );
  OAI21_X1 U8306 ( .B1(n6647), .B2(n9565), .A(n6641), .ZN(P1_U3348) );
  NAND2_X1 U8307 ( .A1(n5146), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8308 ( .A1(n6642), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8309 ( .A1(n5527), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6643) );
  AND3_X1 U8310 ( .A1(n6645), .A2(n6644), .A3(n6643), .ZN(n9163) );
  INV_X1 U8311 ( .A(n9163), .ZN(n8974) );
  NAND2_X1 U8312 ( .A1(n8974), .A2(P1_U3973), .ZN(n6646) );
  OAI21_X1 U8313 ( .B1(P1_U3973), .B2(n6495), .A(n6646), .ZN(P1_U3585) );
  OAI222_X1 U8314 ( .A1(n7161), .A2(P2_U3151), .B1(n8618), .B2(n6647), .C1(
        n9623), .C2(n7954), .ZN(P2_U3288) );
  INV_X1 U8315 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U8316 ( .A1(n6715), .A2(n6649), .ZN(P2_U3246) );
  INV_X1 U8317 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6650) );
  NOR2_X1 U8318 ( .A1(n6715), .A2(n6650), .ZN(P2_U3256) );
  INV_X1 U8319 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6651) );
  NOR2_X1 U8320 ( .A1(n6715), .A2(n6651), .ZN(P2_U3253) );
  INV_X1 U8321 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6652) );
  NOR2_X1 U8322 ( .A1(n6715), .A2(n6652), .ZN(P2_U3247) );
  INV_X1 U8323 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6653) );
  NOR2_X1 U8324 ( .A1(n6715), .A2(n6653), .ZN(P2_U3250) );
  INV_X1 U8325 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6654) );
  NOR2_X1 U8326 ( .A1(n6715), .A2(n6654), .ZN(P2_U3249) );
  INV_X1 U8327 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U8328 ( .A1(n6715), .A2(n6655), .ZN(P2_U3255) );
  INV_X1 U8329 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6656) );
  NOR2_X1 U8330 ( .A1(n6715), .A2(n6656), .ZN(P2_U3248) );
  INV_X1 U8331 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6657) );
  NOR2_X1 U8332 ( .A1(n6715), .A2(n6657), .ZN(P2_U3257) );
  INV_X1 U8333 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6658) );
  NOR2_X1 U8334 ( .A1(n6715), .A2(n6658), .ZN(P2_U3252) );
  INV_X1 U8335 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6659) );
  NOR2_X1 U8336 ( .A1(n6715), .A2(n6659), .ZN(P2_U3254) );
  INV_X1 U8337 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U8338 ( .A1(n6715), .A2(n6660), .ZN(P2_U3251) );
  INV_X1 U8339 ( .A(n6661), .ZN(n6664) );
  INV_X1 U8340 ( .A(n9136), .ZN(n6662) );
  OAI222_X1 U8341 ( .A1(n9568), .A2(n9684), .B1(n9565), .B2(n6664), .C1(
        P1_U3086), .C2(n6662), .ZN(P1_U3347) );
  OAI222_X1 U8342 ( .A1(n7307), .A2(P2_U3151), .B1(n8618), .B2(n6664), .C1(
        n6663), .C2(n7954), .ZN(P2_U3287) );
  NAND2_X1 U8343 ( .A1(n6978), .A2(P2_U3893), .ZN(n6665) );
  OAI21_X1 U8344 ( .B1(P2_U3893), .B2(n5131), .A(n6665), .ZN(P2_U3491) );
  INV_X1 U8345 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7509) );
  MUX2_X1 U8346 ( .A(n7509), .B(P1_REG2_REG_9__SCAN_IN), .S(n7749), .Z(n6680)
         );
  XNOR2_X1 U8347 ( .A(n6684), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6855) );
  XNOR2_X1 U8348 ( .A(n6685), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9056) );
  AND2_X1 U8349 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9055) );
  NAND2_X1 U8350 ( .A1(n9056), .A2(n9055), .ZN(n9054) );
  INV_X1 U8351 ( .A(n6685), .ZN(n9060) );
  NAND2_X1 U8352 ( .A1(n9060), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8353 ( .A1(n9054), .A2(n6666), .ZN(n6854) );
  NAND2_X1 U8354 ( .A1(n6855), .A2(n6854), .ZN(n6853) );
  INV_X1 U8355 ( .A(n6684), .ZN(n6859) );
  NAND2_X1 U8356 ( .A1(n6859), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8357 ( .A1(n6853), .A2(n6667), .ZN(n9071) );
  XNOR2_X1 U8358 ( .A(n6688), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U8359 ( .A1(n9071), .A2(n9072), .ZN(n9070) );
  INV_X1 U8360 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7326) );
  OR2_X1 U8361 ( .A1(n6688), .A2(n7326), .ZN(n6668) );
  NAND2_X1 U8362 ( .A1(n9070), .A2(n6668), .ZN(n9086) );
  XNOR2_X1 U8363 ( .A(n6690), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9085) );
  NAND2_X1 U8364 ( .A1(n9086), .A2(n9085), .ZN(n9084) );
  INV_X1 U8365 ( .A(n6690), .ZN(n9083) );
  NAND2_X1 U8366 ( .A1(n9083), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8367 ( .A1(n9084), .A2(n6669), .ZN(n9099) );
  INV_X1 U8368 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6670) );
  MUX2_X1 U8369 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6670), .S(n9097), .Z(n9100)
         );
  NAND2_X1 U8370 ( .A1(n9099), .A2(n9100), .ZN(n9098) );
  NAND2_X1 U8371 ( .A1(n9097), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8372 ( .A1(n9098), .A2(n6671), .ZN(n9112) );
  INV_X1 U8373 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6672) );
  XNOR2_X1 U8374 ( .A(n9110), .B(n6672), .ZN(n9113) );
  NAND2_X1 U8375 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  NAND2_X1 U8376 ( .A1(n9110), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8377 ( .A1(n9111), .A2(n6673), .ZN(n9125) );
  INV_X1 U8378 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6674) );
  MUX2_X1 U8379 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6674), .S(n9123), .Z(n9126)
         );
  NAND2_X1 U8380 ( .A1(n9125), .A2(n9126), .ZN(n9124) );
  NAND2_X1 U8381 ( .A1(n9123), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8382 ( .A1(n9124), .A2(n6675), .ZN(n9141) );
  INV_X1 U8383 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U8384 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6676), .S(n9136), .Z(n9142)
         );
  NAND2_X1 U8385 ( .A1(n9141), .A2(n9142), .ZN(n9140) );
  NAND2_X1 U8386 ( .A1(n9136), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U8387 ( .A1(n9140), .A2(n6677), .ZN(n6679) );
  OR2_X1 U8388 ( .A1(n6679), .A2(n6680), .ZN(n7732) );
  INV_X1 U8389 ( .A(n7732), .ZN(n6678) );
  AOI21_X1 U8390 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6703) );
  NAND2_X1 U8391 ( .A1(n6682), .A2(n6681), .ZN(n9769) );
  OR2_X1 U8392 ( .A1(n5509), .A2(n9566), .ZN(n9032) );
  OR2_X1 U8393 ( .A1(n9769), .A2(n6851), .ZN(n9856) );
  INV_X1 U8394 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U8395 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7655) );
  OAI21_X1 U8396 ( .B1(n9862), .B2(n6683), .A(n7655), .ZN(n6701) );
  INV_X1 U8397 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9642) );
  MUX2_X1 U8398 ( .A(n9642), .B(P1_REG1_REG_3__SCAN_IN), .S(n6688), .Z(n9075)
         );
  XNOR2_X1 U8399 ( .A(n6684), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6858) );
  XNOR2_X1 U8400 ( .A(n6685), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9059) );
  AND2_X1 U8401 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9058) );
  NAND2_X1 U8402 ( .A1(n9059), .A2(n9058), .ZN(n9057) );
  NAND2_X1 U8403 ( .A1(n9060), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U8404 ( .A1(n9057), .A2(n6686), .ZN(n6857) );
  NAND2_X1 U8405 ( .A1(n6858), .A2(n6857), .ZN(n6856) );
  NAND2_X1 U8406 ( .A1(n6859), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6687) );
  NAND2_X1 U8407 ( .A1(n6856), .A2(n6687), .ZN(n9074) );
  NAND2_X1 U8408 ( .A1(n9075), .A2(n9074), .ZN(n9073) );
  INV_X1 U8409 ( .A(n6688), .ZN(n9069) );
  NAND2_X1 U8410 ( .A1(n9069), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U8411 ( .A1(n9073), .A2(n6689), .ZN(n9089) );
  XNOR2_X1 U8412 ( .A(n6690), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U8413 ( .A1(n9089), .A2(n9088), .ZN(n9087) );
  NAND2_X1 U8414 ( .A1(n9083), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U8415 ( .A1(n9087), .A2(n6691), .ZN(n9102) );
  INV_X1 U8416 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7286) );
  MUX2_X1 U8417 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7286), .S(n9097), .Z(n9103)
         );
  NAND2_X1 U8418 ( .A1(n9102), .A2(n9103), .ZN(n9101) );
  NAND2_X1 U8419 ( .A1(n9097), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U8420 ( .A1(n9101), .A2(n6692), .ZN(n9115) );
  INV_X1 U8421 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U8422 ( .A(n9110), .B(n6693), .ZN(n9116) );
  NAND2_X1 U8423 ( .A1(n9115), .A2(n9116), .ZN(n9114) );
  NAND2_X1 U8424 ( .A1(n9110), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U8425 ( .A1(n9114), .A2(n6694), .ZN(n9128) );
  INV_X1 U8426 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9656) );
  MUX2_X1 U8427 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9656), .S(n9123), .Z(n9129)
         );
  NAND2_X1 U8428 ( .A1(n9128), .A2(n9129), .ZN(n9127) );
  NAND2_X1 U8429 ( .A1(n9123), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8430 ( .A1(n9127), .A2(n6695), .ZN(n9138) );
  INV_X1 U8431 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9910) );
  MUX2_X1 U8432 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9910), .S(n9136), .Z(n9139)
         );
  NAND2_X1 U8433 ( .A1(n9138), .A2(n9139), .ZN(n9137) );
  NAND2_X1 U8434 ( .A1(n9136), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8435 ( .A1(n9137), .A2(n6696), .ZN(n6698) );
  INV_X1 U8436 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9912) );
  MUX2_X1 U8437 ( .A(n9912), .B(P1_REG1_REG_9__SCAN_IN), .S(n7749), .Z(n6697)
         );
  OR2_X1 U8438 ( .A1(n6698), .A2(n6697), .ZN(n7751) );
  NAND2_X1 U8439 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  OR2_X1 U8440 ( .A1(n9769), .A2(n9766), .ZN(n9809) );
  AOI21_X1 U8441 ( .B1(n7751), .B2(n6699), .A(n9809), .ZN(n6700) );
  AOI211_X1 U8442 ( .C1(n9839), .C2(n7749), .A(n6701), .B(n6700), .ZN(n6702)
         );
  OAI21_X1 U8443 ( .B1(n6703), .B2(n9847), .A(n6702), .ZN(P1_U3252) );
  INV_X1 U8444 ( .A(n6704), .ZN(n6708) );
  AOI22_X1 U8445 ( .A1(n7749), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9570), .ZN(n6705) );
  OAI21_X1 U8446 ( .B1(n6708), .B2(n9565), .A(n6705), .ZN(P1_U3346) );
  NAND2_X1 U8447 ( .A1(n9736), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n6706) );
  OAI21_X1 U8448 ( .B1(n8404), .B2(n9736), .A(n6706), .ZN(P2_U3510) );
  OAI222_X1 U8449 ( .A1(P2_U3151), .A2(n8232), .B1(n8618), .B2(n6708), .C1(
        n6707), .C2(n7954), .ZN(P2_U3286) );
  INV_X1 U8450 ( .A(n6709), .ZN(n6712) );
  AOI22_X1 U8451 ( .A1(n9761), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9570), .ZN(n6710) );
  OAI21_X1 U8452 ( .B1(n6712), .B2(n9565), .A(n6710), .ZN(P1_U3345) );
  OAI222_X1 U8453 ( .A1(P2_U3151), .A2(n9932), .B1(n8618), .B2(n6712), .C1(
        n6711), .C2(n7954), .ZN(P2_U3285) );
  INV_X1 U8454 ( .A(n6713), .ZN(n6799) );
  AOI22_X1 U8455 ( .A1(n9149), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9570), .ZN(n6714) );
  OAI21_X1 U8456 ( .B1(n6799), .B2(n9565), .A(n6714), .ZN(P1_U3344) );
  INV_X1 U8457 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6716) );
  NOR2_X1 U8458 ( .A1(n6715), .A2(n6716), .ZN(P2_U3261) );
  INV_X1 U8459 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6717) );
  NOR2_X1 U8460 ( .A1(n6715), .A2(n6717), .ZN(P2_U3260) );
  INV_X1 U8461 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6718) );
  NOR2_X1 U8462 ( .A1(n6715), .A2(n6718), .ZN(P2_U3258) );
  INV_X1 U8463 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6719) );
  NOR2_X1 U8464 ( .A1(n6715), .A2(n6719), .ZN(P2_U3234) );
  INV_X1 U8465 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6720) );
  NOR2_X1 U8466 ( .A1(n6715), .A2(n6720), .ZN(P2_U3263) );
  INV_X1 U8467 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6721) );
  NOR2_X1 U8468 ( .A1(n6715), .A2(n6721), .ZN(P2_U3262) );
  INV_X1 U8469 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9608) );
  NOR2_X1 U8470 ( .A1(n6715), .A2(n9608), .ZN(P2_U3245) );
  INV_X1 U8471 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6722) );
  NOR2_X1 U8472 ( .A1(n6715), .A2(n6722), .ZN(P2_U3243) );
  INV_X1 U8473 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6723) );
  NOR2_X1 U8474 ( .A1(n6715), .A2(n6723), .ZN(P2_U3259) );
  INV_X1 U8475 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6724) );
  NOR2_X1 U8476 ( .A1(n6715), .A2(n6724), .ZN(P2_U3241) );
  INV_X1 U8477 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6725) );
  NOR2_X1 U8478 ( .A1(n6715), .A2(n6725), .ZN(P2_U3240) );
  INV_X1 U8479 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U8480 ( .A1(n6715), .A2(n6726), .ZN(P2_U3239) );
  INV_X1 U8481 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6727) );
  NOR2_X1 U8482 ( .A1(n6715), .A2(n6727), .ZN(P2_U3238) );
  INV_X1 U8483 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6728) );
  NOR2_X1 U8484 ( .A1(n6715), .A2(n6728), .ZN(P2_U3237) );
  INV_X1 U8485 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6729) );
  NOR2_X1 U8486 ( .A1(n6715), .A2(n6729), .ZN(P2_U3236) );
  INV_X1 U8487 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6730) );
  NOR2_X1 U8488 ( .A1(n6715), .A2(n6730), .ZN(P2_U3235) );
  INV_X1 U8489 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6731) );
  NOR2_X1 U8490 ( .A1(n6715), .A2(n6731), .ZN(P2_U3242) );
  INV_X1 U8491 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6732) );
  NOR2_X1 U8492 ( .A1(n6715), .A2(n6732), .ZN(P2_U3244) );
  MUX2_X1 U8493 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8227), .Z(n6734) );
  XNOR2_X1 U8494 ( .A(n6734), .B(n6762), .ZN(n9927) );
  MUX2_X1 U8495 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8227), .Z(n6733) );
  INV_X1 U8496 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9624) );
  NOR2_X1 U8497 ( .A1(n6733), .A2(n9624), .ZN(n9926) );
  INV_X1 U8498 ( .A(n6762), .ZN(n9925) );
  INV_X1 U8499 ( .A(n6734), .ZN(n6735) );
  OAI22_X1 U8500 ( .A1(n9927), .A2(n9926), .B1(n9925), .B2(n6735), .ZN(n6781)
         );
  MUX2_X1 U8501 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8227), .Z(n6736) );
  XNOR2_X1 U8502 ( .A(n6736), .B(n6795), .ZN(n6780) );
  AOI22_X1 U8503 ( .A1(n6781), .A2(n6780), .B1(n6736), .B2(n6764), .ZN(n6989)
         );
  MUX2_X1 U8504 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8227), .Z(n6737) );
  XNOR2_X1 U8505 ( .A(n6737), .B(n6757), .ZN(n6988) );
  NAND2_X1 U8506 ( .A1(n6989), .A2(n6988), .ZN(n6987) );
  INV_X1 U8507 ( .A(n6737), .ZN(n6738) );
  NAND2_X1 U8508 ( .A1(n6738), .A2(n6757), .ZN(n6740) );
  MUX2_X1 U8509 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8227), .Z(n6919) );
  XNOR2_X1 U8510 ( .A(n6919), .B(n6923), .ZN(n6739) );
  AOI21_X1 U8511 ( .B1(n6987), .B2(n6740), .A(n6739), .ZN(n6779) );
  NAND3_X1 U8512 ( .A1(n6987), .A2(n6740), .A3(n6739), .ZN(n6920) );
  NAND2_X1 U8513 ( .A1(n6920), .A2(n10060), .ZN(n6778) );
  NOR2_X1 U8514 ( .A1(n8227), .A2(P2_U3151), .ZN(n8613) );
  AND2_X1 U8515 ( .A1(n6746), .A2(n8613), .ZN(n6742) );
  INV_X1 U8516 ( .A(n6002), .ZN(n6741) );
  INV_X1 U8517 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6775) );
  INV_X1 U8518 ( .A(n6743), .ZN(n6744) );
  NOR2_X1 U8519 ( .A1(n6836), .A2(n6744), .ZN(n6745) );
  NOR2_X1 U8520 ( .A1(n6002), .A2(P2_U3151), .ZN(n8609) );
  MUX2_X1 U8521 ( .A(n6747), .B(P2_REG1_REG_4__SCAN_IN), .S(n6923), .Z(n6759)
         );
  NAND2_X1 U8522 ( .A1(n6760), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U8523 ( .A1(n6762), .A2(n6752), .ZN(n6751) );
  NAND2_X1 U8524 ( .A1(n9624), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6749) );
  OR2_X1 U8525 ( .A1(n6749), .A2(n6760), .ZN(n6750) );
  NAND2_X1 U8526 ( .A1(n6751), .A2(n6750), .ZN(n9919) );
  NAND2_X1 U8527 ( .A1(n9919), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6753) );
  NAND2_X1 U8528 ( .A1(n6753), .A2(n6752), .ZN(n6788) );
  NAND2_X1 U8529 ( .A1(n6764), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U8530 ( .A1(n6787), .A2(n6754), .ZN(n6755) );
  XNOR2_X1 U8531 ( .A(n6755), .B(n6990), .ZN(n6991) );
  INV_X1 U8532 ( .A(n6755), .ZN(n6756) );
  OAI22_X1 U8533 ( .A1(n6991), .A2(n10118), .B1(n6757), .B2(n6756), .ZN(n6758)
         );
  OAI21_X1 U8534 ( .B1(n6759), .B2(n6758), .A(n6922), .ZN(n6773) );
  AND2_X1 U8535 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7152) );
  MUX2_X1 U8536 ( .A(n5644), .B(P2_REG2_REG_2__SCAN_IN), .S(n6795), .Z(n6784)
         );
  AND2_X1 U8537 ( .A1(n9624), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U8538 ( .A1(n6760), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6763) );
  OAI21_X1 U8539 ( .B1(n6762), .B2(n6761), .A(n6763), .ZN(n9916) );
  INV_X1 U8540 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9915) );
  OR2_X1 U8541 ( .A1(n9916), .A2(n9915), .ZN(n9918) );
  NAND2_X1 U8542 ( .A1(n9918), .A2(n6763), .ZN(n6783) );
  NAND2_X1 U8543 ( .A1(n6784), .A2(n6783), .ZN(n6782) );
  NAND2_X1 U8544 ( .A1(n6764), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8545 ( .A1(n6782), .A2(n6765), .ZN(n6766) );
  NAND2_X1 U8546 ( .A1(n6766), .A2(n6990), .ZN(n6769) );
  INV_X1 U8547 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7432) );
  NAND2_X1 U8548 ( .A1(n6994), .A2(n6769), .ZN(n6767) );
  INV_X1 U8549 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9619) );
  MUX2_X1 U8550 ( .A(n9619), .B(P2_REG2_REG_4__SCAN_IN), .S(n6923), .Z(n6768)
         );
  NAND2_X1 U8551 ( .A1(n6767), .A2(n6768), .ZN(n6925) );
  INV_X1 U8552 ( .A(n6768), .ZN(n6770) );
  NAND3_X1 U8553 ( .A1(n6994), .A2(n6770), .A3(n6769), .ZN(n6771) );
  AOI21_X1 U8554 ( .B1(n6925), .B2(n6771), .A(n10065), .ZN(n6772) );
  AOI211_X1 U8555 ( .C1(n10061), .C2(n6773), .A(n7152), .B(n6772), .ZN(n6774)
         );
  OAI21_X1 U8556 ( .B1(n6775), .B2(n9931), .A(n6774), .ZN(n6776) );
  AOI21_X1 U8557 ( .B1(n6923), .B2(n10052), .A(n6776), .ZN(n6777) );
  OAI21_X1 U8558 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(P2_U3186) );
  INV_X1 U8559 ( .A(n10060), .ZN(n9739) );
  XNOR2_X1 U8560 ( .A(n6781), .B(n6780), .ZN(n6797) );
  INV_X1 U8561 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6793) );
  INV_X1 U8562 ( .A(n10065), .ZN(n9994) );
  OAI21_X1 U8563 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(n6786) );
  NOR2_X1 U8564 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7250), .ZN(n6785) );
  AOI21_X1 U8565 ( .B1(n9994), .B2(n6786), .A(n6785), .ZN(n6792) );
  OAI21_X1 U8566 ( .B1(n6789), .B2(n6788), .A(n6787), .ZN(n6790) );
  NAND2_X1 U8567 ( .A1(n10061), .A2(n6790), .ZN(n6791) );
  OAI211_X1 U8568 ( .C1(n6793), .C2(n9931), .A(n6792), .B(n6791), .ZN(n6794)
         );
  AOI21_X1 U8569 ( .B1(n6795), .B2(n10052), .A(n6794), .ZN(n6796) );
  OAI21_X1 U8570 ( .B1(n9739), .B2(n6797), .A(n6796), .ZN(P2_U3184) );
  OAI222_X1 U8571 ( .A1(n8261), .A2(P2_U3151), .B1(n8618), .B2(n6799), .C1(
        n6798), .C2(n7954), .ZN(P2_U3284) );
  INV_X1 U8572 ( .A(n10052), .ZN(n9735) );
  INV_X1 U8573 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6948) );
  INV_X1 U8574 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6800) );
  MUX2_X1 U8575 ( .A(n6948), .B(n6800), .S(n8227), .Z(n6801) );
  NOR2_X1 U8576 ( .A1(n6801), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6802) );
  OAI22_X1 U8577 ( .A1(n10060), .A2(n6803), .B1(n9926), .B2(n6802), .ZN(n6804)
         );
  OAI21_X1 U8578 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6805), .A(n6804), .ZN(n6806) );
  AOI21_X1 U8579 ( .B1(n10053), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6806), .ZN(
        n6807) );
  OAI21_X1 U8580 ( .B1(n9624), .B2(n9735), .A(n6807), .ZN(P2_U3182) );
  XOR2_X1 U8581 ( .A(n6809), .B(n6808), .Z(n6848) );
  AOI22_X1 U8582 ( .A1(n8765), .A2(n6810), .B1(n8746), .B2(n6848), .ZN(n6813)
         );
  OR2_X1 U8583 ( .A1(n6811), .A2(P1_U3086), .ZN(n6878) );
  AOI22_X1 U8584 ( .A1(n8751), .A2(n9053), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6878), .ZN(n6812) );
  NAND2_X1 U8585 ( .A1(n6813), .A2(n6812), .ZN(P1_U3232) );
  NAND2_X1 U8586 ( .A1(n6822), .A2(n6829), .ZN(n6817) );
  INV_X1 U8587 ( .A(n6814), .ZN(n6815) );
  NAND2_X1 U8588 ( .A1(n6826), .A2(n6815), .ZN(n6816) );
  XNOR2_X1 U8589 ( .A(n7098), .B(n4292), .ZN(n7097) );
  NAND2_X1 U8590 ( .A1(n6975), .A2(n4894), .ZN(n7096) );
  XOR2_X1 U8591 ( .A(n7097), .B(n7096), .Z(n6847) );
  NAND2_X1 U8592 ( .A1(n6822), .A2(n6937), .ZN(n6825) );
  NAND2_X1 U8593 ( .A1(n6826), .A2(n10095), .ZN(n6828) );
  INV_X1 U8594 ( .A(n8166), .ZN(n8182) );
  OAI22_X1 U8595 ( .A1(n7114), .A2(n8158), .B1(n8182), .B2(n7269), .ZN(n6845)
         );
  NAND2_X1 U8596 ( .A1(n6840), .A2(n6829), .ZN(n6837) );
  INV_X1 U8597 ( .A(n6830), .ZN(n6832) );
  OAI21_X1 U8598 ( .B1(n6833), .B2(n6832), .A(n6831), .ZN(n6835) );
  NAND4_X1 U8599 ( .A1(n6837), .A2(n6836), .A3(n6835), .A4(n6834), .ZN(n6838)
         );
  NAND2_X1 U8600 ( .A1(n6838), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6842) );
  NAND3_X1 U8601 ( .A1(n6840), .A2(n6937), .A3(n6839), .ZN(n6841) );
  AND2_X1 U8602 ( .A1(n6842), .A2(n6841), .ZN(n7111) );
  AND2_X1 U8603 ( .A1(n7111), .A2(n6843), .ZN(n7975) );
  INV_X1 U8604 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U8605 ( .A1(n7975), .A2(n9920), .ZN(n6844) );
  AOI211_X1 U8606 ( .C1(n8155), .C2(n6978), .A(n6845), .B(n6844), .ZN(n6846)
         );
  OAI21_X1 U8607 ( .B1(n8162), .B2(n6847), .A(n6846), .ZN(P2_U3162) );
  INV_X1 U8608 ( .A(n6848), .ZN(n6849) );
  MUX2_X1 U8609 ( .A(n6849), .B(n9055), .S(n9766), .Z(n6852) );
  INV_X1 U8610 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7138) );
  AOI21_X1 U8611 ( .B1(n9766), .B2(n7138), .A(n5509), .ZN(n9765) );
  OAI21_X1 U8612 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9765), .A(P1_U3973), .ZN(
        n6850) );
  AOI21_X1 U8613 ( .B1(n6852), .B2(n6851), .A(n6850), .ZN(n9079) );
  INV_X1 U8614 ( .A(n9847), .ZN(n9842) );
  OAI211_X1 U8615 ( .C1(n6855), .C2(n6854), .A(n9842), .B(n6853), .ZN(n6863)
         );
  AOI22_X1 U8616 ( .A1(n9827), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6862) );
  INV_X1 U8617 ( .A(n9809), .ZN(n9850) );
  OAI211_X1 U8618 ( .C1(n6858), .C2(n6857), .A(n9850), .B(n6856), .ZN(n6861)
         );
  NAND2_X1 U8619 ( .A1(n9839), .A2(n6859), .ZN(n6860) );
  NAND4_X1 U8620 ( .A1(n6863), .A2(n6862), .A3(n6861), .A4(n6860), .ZN(n6864)
         );
  OR2_X1 U8621 ( .A1(n9079), .A2(n6864), .ZN(P1_U3245) );
  INV_X1 U8622 ( .A(n6865), .ZN(n6866) );
  AOI21_X1 U8623 ( .B1(n6868), .B2(n6867), .A(n6866), .ZN(n6871) );
  INV_X1 U8624 ( .A(n8736), .ZN(n8760) );
  AOI22_X1 U8625 ( .A1(n8760), .A2(n6954), .B1(n8751), .B2(n9052), .ZN(n6870)
         );
  AOI22_X1 U8626 ( .A1(n8765), .A2(n7184), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6878), .ZN(n6869) );
  OAI211_X1 U8627 ( .C1(n6871), .C2(n8768), .A(n6870), .B(n6869), .ZN(P1_U3222) );
  INV_X1 U8628 ( .A(n6872), .ZN(n6873) );
  NOR2_X1 U8629 ( .A1(n6874), .A2(n6873), .ZN(n6877) );
  INV_X1 U8630 ( .A(n6875), .ZN(n6876) );
  AOI21_X1 U8631 ( .B1(n6877), .B2(n6865), .A(n6876), .ZN(n6881) );
  AOI22_X1 U8632 ( .A1(n8751), .A2(n9051), .B1(n8760), .B2(n9053), .ZN(n6880)
         );
  AOI22_X1 U8633 ( .A1(n8765), .A2(n7213), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6878), .ZN(n6879) );
  OAI211_X1 U8634 ( .C1(n6881), .C2(n8768), .A(n6880), .B(n6879), .ZN(P1_U3237) );
  OAI21_X1 U8635 ( .B1(n6884), .B2(n6883), .A(n6882), .ZN(n7189) );
  INV_X1 U8636 ( .A(n7189), .ZN(n6890) );
  INV_X1 U8637 ( .A(n7446), .ZN(n7398) );
  OAI22_X1 U8638 ( .A1(n4561), .A2(n9261), .B1(n7033), .B2(n9262), .ZN(n6889)
         );
  INV_X1 U8639 ( .A(n6955), .ZN(n6885) );
  NAND2_X1 U8640 ( .A1(n6885), .A2(n6884), .ZN(n6887) );
  AOI21_X1 U8641 ( .B1(n6887), .B2(n6886), .A(n9258), .ZN(n6888) );
  AOI211_X1 U8642 ( .C1(n7398), .C2(n7189), .A(n6889), .B(n6888), .ZN(n7191)
         );
  OAI211_X1 U8643 ( .C1(n4444), .C2(n8909), .A(n9331), .B(n6901), .ZN(n7187)
         );
  OAI211_X1 U8644 ( .C1(n6890), .C2(n7450), .A(n7191), .B(n7187), .ZN(n7119)
         );
  INV_X1 U8645 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6891) );
  OAI22_X1 U8646 ( .A1(n9463), .A2(n8909), .B1(n9914), .B2(n6891), .ZN(n6892)
         );
  AOI21_X1 U8647 ( .B1(n7119), .B2(n9914), .A(n6892), .ZN(n6893) );
  INV_X1 U8648 ( .A(n6893), .ZN(P1_U3523) );
  INV_X1 U8649 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6898) );
  OAI21_X1 U8650 ( .B1(n8460), .B2(n10114), .A(n7968), .ZN(n6895) );
  NOR2_X1 U8651 ( .A1(n4292), .A2(n8442), .ZN(n6938) );
  INV_X1 U8652 ( .A(n6938), .ZN(n6894) );
  OAI211_X1 U8653 ( .C1(n10111), .C2(n6896), .A(n6895), .B(n6894), .ZN(n8544)
         );
  NAND2_X1 U8654 ( .A1(n8544), .A2(n10116), .ZN(n6897) );
  OAI21_X1 U8655 ( .B1(n6898), .B2(n10116), .A(n6897), .ZN(P2_U3390) );
  OAI21_X1 U8656 ( .B1(n6900), .B2(n8980), .A(n6899), .ZN(n7217) );
  INV_X1 U8657 ( .A(n6901), .ZN(n6903) );
  INV_X1 U8658 ( .A(n6902), .ZN(n6914) );
  OAI211_X1 U8659 ( .C1(n6904), .C2(n6903), .A(n6914), .B(n9331), .ZN(n7215)
         );
  OAI21_X1 U8660 ( .B1(n6904), .B2(n9901), .A(n7215), .ZN(n6908) );
  XNOR2_X1 U8661 ( .A(n6905), .B(n8980), .ZN(n6906) );
  OAI222_X1 U8662 ( .A1(n9261), .A2(n6956), .B1(n9262), .B2(n6907), .C1(n6906), 
        .C2(n9258), .ZN(n7209) );
  AOI211_X1 U8663 ( .C1(n9905), .C2(n7217), .A(n6908), .B(n7209), .ZN(n9885)
         );
  NAND2_X1 U8664 ( .A1(n5572), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6909) );
  OAI21_X1 U8665 ( .B1(n9885), .B2(n5572), .A(n6909), .ZN(P1_U3524) );
  XNOR2_X1 U8666 ( .A(n8776), .B(n6911), .ZN(n7335) );
  OAI21_X1 U8667 ( .B1(n6912), .B2(n6911), .A(n6910), .ZN(n7333) );
  OAI22_X1 U8668 ( .A1(n7033), .A2(n9261), .B1(n7331), .B2(n9262), .ZN(n6915)
         );
  INV_X1 U8669 ( .A(n6964), .ZN(n6913) );
  AOI211_X1 U8670 ( .C1(n7328), .C2(n6914), .A(n9371), .B(n6913), .ZN(n7325)
         );
  AOI211_X1 U8671 ( .C1(n9905), .C2(n7333), .A(n6915), .B(n7325), .ZN(n6916)
         );
  OAI21_X1 U8672 ( .B1(n9258), .B2(n7335), .A(n6916), .ZN(n7128) );
  OAI22_X1 U8673 ( .A1(n9463), .A2(n7126), .B1(n9914), .B2(n9642), .ZN(n6917)
         );
  AOI21_X1 U8674 ( .B1(n7128), .B2(n9914), .A(n6917), .ZN(n6918) );
  INV_X1 U8675 ( .A(n6918), .ZN(P1_U3525) );
  INV_X1 U8676 ( .A(n6919), .ZN(n6921) );
  OAI21_X1 U8677 ( .B1(n6923), .B2(n6921), .A(n6920), .ZN(n7052) );
  MUX2_X1 U8678 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8227), .Z(n7050) );
  XOR2_X1 U8679 ( .A(n7049), .B(n7050), .Z(n7051) );
  XNOR2_X1 U8680 ( .A(n7052), .B(n7051), .ZN(n6936) );
  XNOR2_X1 U8681 ( .A(n7041), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n6934) );
  INV_X1 U8682 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6932) );
  OR2_X1 U8683 ( .A1(n6923), .A2(n9619), .ZN(n6924) );
  NAND2_X1 U8684 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  NAND2_X1 U8685 ( .A1(n6926), .A2(n7049), .ZN(n7074) );
  OAI21_X1 U8686 ( .B1(n6926), .B2(n7049), .A(n7074), .ZN(n6927) );
  NAND2_X1 U8687 ( .A1(n6927), .A2(n7375), .ZN(n6928) );
  NAND2_X1 U8688 ( .A1(n7076), .A2(n6928), .ZN(n6929) );
  NOR2_X1 U8689 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5579), .ZN(n7237) );
  AOI21_X1 U8690 ( .B1(n9994), .B2(n6929), .A(n7237), .ZN(n6931) );
  NAND2_X1 U8691 ( .A1(n10052), .A2(n4497), .ZN(n6930) );
  OAI211_X1 U8692 ( .C1(n6932), .C2(n9931), .A(n6931), .B(n6930), .ZN(n6933)
         );
  AOI21_X1 U8693 ( .B1(n10061), .B2(n6934), .A(n6933), .ZN(n6935) );
  OAI21_X1 U8694 ( .B1(n6936), .B2(n9739), .A(n6935), .ZN(P2_U3187) );
  NOR2_X1 U8695 ( .A1(n6937), .A2(n10095), .ZN(n6939) );
  AOI21_X1 U8696 ( .B1(n7968), .B2(n6939), .A(n6938), .ZN(n6947) );
  INV_X1 U8697 ( .A(n6821), .ZN(n6942) );
  INV_X1 U8698 ( .A(n6940), .ZN(n6941) );
  MUX2_X1 U8699 ( .A(n6943), .B(n6942), .S(n6941), .Z(n6944) );
  NAND2_X1 U8700 ( .A1(n6945), .A2(n6944), .ZN(n6949) );
  MUX2_X1 U8701 ( .A(n6948), .B(n6947), .S(n8474), .Z(n6953) );
  INV_X1 U8702 ( .A(n6949), .ZN(n6951) );
  INV_X1 U8703 ( .A(n8464), .ZN(n6950) );
  AOI22_X1 U8704 ( .A1(n8393), .A2(n7967), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8446), .ZN(n6952) );
  NAND2_X1 U8705 ( .A1(n6953), .A2(n6952), .ZN(P2_U3233) );
  INV_X1 U8706 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6960) );
  AND2_X1 U8707 ( .A1(n6954), .A2(n4444), .ZN(n8908) );
  OR2_X1 U8708 ( .A1(n8908), .A2(n6955), .ZN(n8979) );
  INV_X1 U8709 ( .A(n8979), .ZN(n7141) );
  NOR2_X1 U8710 ( .A1(n9905), .A2(n9482), .ZN(n6957) );
  OAI222_X1 U8711 ( .A1(n4444), .A2(n6958), .B1(n7141), .B2(n6957), .C1(n9262), 
        .C2(n6956), .ZN(n9492) );
  NAND2_X1 U8712 ( .A1(n9492), .A2(n9908), .ZN(n6959) );
  OAI21_X1 U8713 ( .B1(n9544), .B2(n6960), .A(n6959), .ZN(P1_U3453) );
  XNOR2_X1 U8714 ( .A(n6961), .B(n8985), .ZN(n6962) );
  AOI22_X1 U8715 ( .A1(n9051), .A2(n9474), .B1(n9475), .B2(n9049), .ZN(n7025)
         );
  OAI21_X1 U8716 ( .B1(n6962), .B2(n9258), .A(n7025), .ZN(n7220) );
  AOI21_X1 U8717 ( .B1(n6964), .B2(n6963), .A(n9371), .ZN(n6965) );
  AND2_X1 U8718 ( .A1(n6965), .A2(n7279), .ZN(n7221) );
  NOR2_X1 U8719 ( .A1(n7220), .A2(n7221), .ZN(n7124) );
  OAI21_X1 U8720 ( .B1(n6967), .B2(n8985), .A(n6966), .ZN(n7228) );
  INV_X1 U8721 ( .A(n9491), .ZN(n9457) );
  INV_X1 U8722 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6968) );
  OAI22_X1 U8723 ( .A1(n9463), .A2(n7226), .B1(n9914), .B2(n6968), .ZN(n6969)
         );
  AOI21_X1 U8724 ( .B1(n7228), .B2(n9457), .A(n6969), .ZN(n6970) );
  OAI21_X1 U8725 ( .B1(n7124), .B2(n5572), .A(n6970), .ZN(P1_U3526) );
  INV_X1 U8726 ( .A(n6971), .ZN(n7007) );
  AOI22_X1 U8727 ( .A1(n9794), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9570), .ZN(n6972) );
  OAI21_X1 U8728 ( .B1(n7007), .B2(n9565), .A(n6972), .ZN(P1_U3342) );
  INV_X1 U8729 ( .A(n6973), .ZN(n6974) );
  NAND2_X1 U8730 ( .A1(n6977), .A2(n8460), .ZN(n6980) );
  AOI22_X1 U8731 ( .A1(n8457), .A2(n6978), .B1(n6359), .B2(n8455), .ZN(n6979)
         );
  NAND2_X1 U8732 ( .A1(n6980), .A2(n6979), .ZN(n7271) );
  INV_X1 U8733 ( .A(n7271), .ZN(n6981) );
  OAI21_X1 U8734 ( .B1(n7275), .B2(n10106), .A(n6981), .ZN(n7004) );
  OAI22_X1 U8735 ( .A1(n8543), .A2(n7269), .B1(n10130), .B2(n5625), .ZN(n6982)
         );
  AOI21_X1 U8736 ( .B1(n7004), .B2(n10130), .A(n6982), .ZN(n6983) );
  INV_X1 U8737 ( .A(n6983), .ZN(P2_U3460) );
  INV_X1 U8738 ( .A(n6984), .ZN(n6986) );
  OAI222_X1 U8739 ( .A1(P2_U3151), .A2(n8239), .B1(n8618), .B2(n6986), .C1(
        n6985), .C2(n7954), .ZN(P2_U3283) );
  INV_X1 U8740 ( .A(n7756), .ZN(n9779) );
  OAI222_X1 U8741 ( .A1(n9568), .A2(n9669), .B1(n9565), .B2(n6986), .C1(n9779), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  OAI21_X1 U8742 ( .B1(n6989), .B2(n6988), .A(n6987), .ZN(n7001) );
  NOR2_X1 U8743 ( .A1(n9735), .A2(n6990), .ZN(n7000) );
  INV_X1 U8744 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6998) );
  XNOR2_X1 U8745 ( .A(n6991), .B(n10118), .ZN(n6992) );
  AOI22_X1 U8746 ( .A1(n10061), .A2(n6992), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3151), .ZN(n6997) );
  AND2_X1 U8747 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  OR2_X1 U8748 ( .A1(n10065), .A2(n6995), .ZN(n6996) );
  OAI211_X1 U8749 ( .C1(n6998), .C2(n9931), .A(n6997), .B(n6996), .ZN(n6999)
         );
  AOI211_X1 U8750 ( .C1(n10060), .C2(n7001), .A(n7000), .B(n6999), .ZN(n7002)
         );
  INV_X1 U8751 ( .A(n7002), .ZN(P2_U3185) );
  OAI22_X1 U8752 ( .A1(n7269), .A2(n8602), .B1(n10116), .B2(n5623), .ZN(n7003)
         );
  AOI21_X1 U8753 ( .B1(n7004), .B2(n10116), .A(n7003), .ZN(n7005) );
  INV_X1 U8754 ( .A(n7005), .ZN(P2_U3393) );
  OAI222_X1 U8755 ( .A1(n8266), .A2(P2_U3151), .B1(n8618), .B2(n7007), .C1(
        n7006), .C2(n7954), .ZN(P2_U3282) );
  OAI21_X1 U8756 ( .B1(n7009), .B2(n7008), .A(n7426), .ZN(n7249) );
  XNOR2_X1 U8757 ( .A(n7011), .B(n7010), .ZN(n7012) );
  NAND2_X1 U8758 ( .A1(n7012), .A2(n8460), .ZN(n7015) );
  AOI22_X1 U8759 ( .A1(n8457), .A2(n8202), .B1(n8201), .B2(n8455), .ZN(n7014)
         );
  NAND2_X1 U8760 ( .A1(n7015), .A2(n7014), .ZN(n7252) );
  AOI21_X1 U8761 ( .B1(n10114), .B2(n7249), .A(n7252), .ZN(n7020) );
  OAI22_X1 U8762 ( .A1(n7973), .A2(n8602), .B1(n10116), .B2(n5645), .ZN(n7016)
         );
  INV_X1 U8763 ( .A(n7016), .ZN(n7017) );
  OAI21_X1 U8764 ( .B1(n7020), .B2(n10117), .A(n7017), .ZN(P2_U3396) );
  OAI22_X1 U8765 ( .A1(n8543), .A2(n7973), .B1(n10130), .B2(n6748), .ZN(n7018)
         );
  INV_X1 U8766 ( .A(n7018), .ZN(n7019) );
  OAI21_X1 U8767 ( .B1(n7020), .B2(n10128), .A(n7019), .ZN(P2_U3461) );
  AOI21_X1 U8768 ( .B1(n7022), .B2(n7021), .A(n8768), .ZN(n7024) );
  NAND2_X1 U8769 ( .A1(n7024), .A2(n7023), .ZN(n7029) );
  NAND2_X1 U8770 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9080) );
  OAI21_X1 U8771 ( .B1(n8705), .B2(n7025), .A(n9080), .ZN(n7026) );
  AOI21_X1 U8772 ( .B1(n8759), .B2(n7027), .A(n7026), .ZN(n7028) );
  OAI211_X1 U8773 ( .C1(n7226), .C2(n8754), .A(n7029), .B(n7028), .ZN(P1_U3230) );
  OAI21_X1 U8774 ( .B1(n7032), .B2(n7031), .A(n7030), .ZN(n7037) );
  OAI22_X1 U8775 ( .A1(n8754), .A2(n7126), .B1(n7033), .B2(n8736), .ZN(n7036)
         );
  NOR2_X1 U8776 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5159), .ZN(n9065) );
  AOI21_X1 U8777 ( .B1(n8751), .B2(n9050), .A(n9065), .ZN(n7034) );
  OAI21_X1 U8778 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n8749), .A(n7034), .ZN(
        n7035) );
  AOI211_X1 U8779 ( .C1(n7037), .C2(n8746), .A(n7036), .B(n7035), .ZN(n7038)
         );
  INV_X1 U8780 ( .A(n7038), .ZN(P1_U3218) );
  INV_X1 U8781 ( .A(n7039), .ZN(n7087) );
  AOI22_X1 U8782 ( .A1(n9806), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9570), .ZN(n7040) );
  OAI21_X1 U8783 ( .B1(n7087), .B2(n9565), .A(n7040), .ZN(P1_U3341) );
  MUX2_X1 U8784 ( .A(n5702), .B(P2_REG1_REG_6__SCAN_IN), .S(n7079), .Z(n7069)
         );
  NOR2_X1 U8785 ( .A1(n7068), .A2(n7069), .ZN(n7067) );
  AOI21_X1 U8786 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7079), .A(n7067), .ZN(
        n7159) );
  XNOR2_X1 U8787 ( .A(n7159), .B(n7161), .ZN(n7162) );
  INV_X1 U8788 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7055) );
  XNOR2_X1 U8789 ( .A(n7162), .B(n7055), .ZN(n7066) );
  INV_X1 U8790 ( .A(n7161), .ZN(n7057) );
  INV_X1 U8791 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7044) );
  NOR2_X1 U8792 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7042), .ZN(n7467) );
  INV_X1 U8793 ( .A(n7467), .ZN(n7043) );
  OAI21_X1 U8794 ( .B1(n9931), .B2(n7044), .A(n7043), .ZN(n7048) );
  XNOR2_X1 U8795 ( .A(n7079), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7075) );
  OAI21_X1 U8796 ( .B1(n4751), .B2(n7161), .A(n7172), .ZN(n7045) );
  NOR2_X1 U8797 ( .A1(n7045), .A2(n7056), .ZN(n7175) );
  AOI21_X1 U8798 ( .B1(n7056), .B2(n7045), .A(n7175), .ZN(n7046) );
  NOR2_X1 U8799 ( .A1(n7046), .A2(n10065), .ZN(n7047) );
  AOI211_X1 U8800 ( .C1(n10052), .C2(n7057), .A(n7048), .B(n7047), .ZN(n7065)
         );
  AOI22_X1 U8801 ( .A1(n7052), .A2(n7051), .B1(n7050), .B2(n7049), .ZN(n7072)
         );
  MUX2_X1 U8802 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8227), .Z(n7053) );
  NOR2_X1 U8803 ( .A1(n7053), .A2(n7079), .ZN(n7054) );
  AOI21_X1 U8804 ( .B1(n7053), .B2(n7079), .A(n7054), .ZN(n7071) );
  NAND2_X1 U8805 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  INV_X1 U8806 ( .A(n7054), .ZN(n7062) );
  MUX2_X1 U8807 ( .A(n7056), .B(n7055), .S(n8227), .Z(n7058) );
  NAND2_X1 U8808 ( .A1(n7058), .A2(n7057), .ZN(n7165) );
  INV_X1 U8809 ( .A(n7058), .ZN(n7059) );
  NAND2_X1 U8810 ( .A1(n7059), .A2(n7161), .ZN(n7060) );
  NAND2_X1 U8811 ( .A1(n7165), .A2(n7060), .ZN(n7061) );
  AOI21_X1 U8812 ( .B1(n7070), .B2(n7062), .A(n7061), .ZN(n7167) );
  AND3_X1 U8813 ( .A1(n7070), .A2(n7062), .A3(n7061), .ZN(n7063) );
  OAI21_X1 U8814 ( .B1(n7167), .B2(n7063), .A(n10060), .ZN(n7064) );
  OAI211_X1 U8815 ( .C1(n7066), .C2(n9922), .A(n7065), .B(n7064), .ZN(P2_U3189) );
  AOI21_X1 U8816 ( .B1(n7069), .B2(n7068), .A(n7067), .ZN(n7085) );
  OAI21_X1 U8817 ( .B1(n7072), .B2(n7071), .A(n7070), .ZN(n7073) );
  NAND2_X1 U8818 ( .A1(n7073), .A2(n10060), .ZN(n7084) );
  NAND3_X1 U8819 ( .A1(n7076), .A2(n7075), .A3(n7074), .ZN(n7077) );
  NAND2_X1 U8820 ( .A1(n4380), .A2(n7077), .ZN(n7082) );
  INV_X1 U8821 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U8822 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7263) );
  OAI21_X1 U8823 ( .B1(n9931), .B2(n7078), .A(n7263), .ZN(n7081) );
  NOR2_X1 U8824 ( .A1(n9735), .A2(n7079), .ZN(n7080) );
  AOI211_X1 U8825 ( .C1(n9994), .C2(n7082), .A(n7081), .B(n7080), .ZN(n7083)
         );
  OAI211_X1 U8826 ( .C1(n7085), .C2(n9922), .A(n7084), .B(n7083), .ZN(P2_U3188) );
  OAI222_X1 U8827 ( .A1(n8253), .A2(P2_U3151), .B1(n8618), .B2(n7087), .C1(
        n7086), .C2(n7954), .ZN(P2_U3281) );
  XNOR2_X1 U8828 ( .A(n7089), .B(n7088), .ZN(n7090) );
  XNOR2_X1 U8829 ( .A(n7091), .B(n7090), .ZN(n7095) );
  AOI22_X1 U8830 ( .A1(n8760), .A2(n9050), .B1(n8759), .B2(n9866), .ZN(n7092)
         );
  NAND2_X1 U8831 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(n4288), .ZN(n9094) );
  OAI211_X1 U8832 ( .C1(n7442), .C2(n8762), .A(n7092), .B(n9094), .ZN(n7093)
         );
  AOI21_X1 U8833 ( .B1(n7280), .B2(n8765), .A(n7093), .ZN(n7094) );
  OAI21_X1 U8834 ( .B1(n7095), .B2(n8768), .A(n7094), .ZN(P1_U3227) );
  NAND2_X1 U8835 ( .A1(n7097), .A2(n7096), .ZN(n7101) );
  INV_X1 U8836 ( .A(n7098), .ZN(n7099) );
  NAND2_X1 U8837 ( .A1(n7099), .A2(n4292), .ZN(n7100) );
  NAND2_X1 U8838 ( .A1(n7101), .A2(n7100), .ZN(n7971) );
  XNOR2_X1 U8839 ( .A(n7236), .B(n7973), .ZN(n7102) );
  XNOR2_X1 U8840 ( .A(n7102), .B(n7114), .ZN(n7972) );
  NAND2_X1 U8841 ( .A1(n7971), .A2(n7972), .ZN(n7105) );
  INV_X1 U8842 ( .A(n7102), .ZN(n7103) );
  NAND2_X1 U8843 ( .A1(n7103), .A2(n7114), .ZN(n7104) );
  NAND2_X1 U8844 ( .A1(n7105), .A2(n7104), .ZN(n7109) );
  INV_X1 U8845 ( .A(n7109), .ZN(n7107) );
  INV_X1 U8846 ( .A(n7110), .ZN(n7106) );
  AOI211_X1 U8847 ( .C1(n7110), .C2(n7109), .A(n8162), .B(n7108), .ZN(n7116)
         );
  INV_X1 U8848 ( .A(n8179), .ZN(n8130) );
  MUX2_X1 U8849 ( .A(n8130), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7113) );
  AOI22_X1 U8850 ( .A1(n8175), .A2(n5683), .B1(n7430), .B2(n8166), .ZN(n7112)
         );
  OAI211_X1 U8851 ( .C1(n7114), .C2(n8177), .A(n7113), .B(n7112), .ZN(n7115)
         );
  OR2_X1 U8852 ( .A1(n7116), .A2(n7115), .ZN(P2_U3158) );
  INV_X1 U8853 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7117) );
  OAI22_X1 U8854 ( .A1(n9534), .A2(n8909), .B1(n9908), .B2(n7117), .ZN(n7118)
         );
  AOI21_X1 U8855 ( .B1(n7119), .B2(n9908), .A(n7118), .ZN(n7120) );
  INV_X1 U8856 ( .A(n7120), .ZN(P1_U3456) );
  INV_X1 U8857 ( .A(n9548), .ZN(n9528) );
  INV_X1 U8858 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7121) );
  OAI22_X1 U8859 ( .A1(n9534), .A2(n7226), .B1(n9908), .B2(n7121), .ZN(n7122)
         );
  AOI21_X1 U8860 ( .B1(n7228), .B2(n9528), .A(n7122), .ZN(n7123) );
  OAI21_X1 U8861 ( .B1(n7124), .B2(n9906), .A(n7123), .ZN(P1_U3465) );
  INV_X1 U8862 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7125) );
  OAI22_X1 U8863 ( .A1(n9534), .A2(n7126), .B1(n9908), .B2(n7125), .ZN(n7127)
         );
  AOI21_X1 U8864 ( .B1(n7128), .B2(n9908), .A(n7127), .ZN(n7129) );
  INV_X1 U8865 ( .A(n7129), .ZN(P1_U3462) );
  NOR2_X1 U8866 ( .A1(n7130), .A2(n4288), .ZN(n7133) );
  NAND4_X1 U8867 ( .A1(n7134), .A2(n7133), .A3(n7132), .A4(n7131), .ZN(n7135)
         );
  AOI21_X1 U8868 ( .B1(n9863), .B2(n9331), .A(n9378), .ZN(n7146) );
  INV_X1 U8869 ( .A(n9349), .ZN(n7144) );
  INV_X1 U8870 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7137) );
  OAI22_X1 U8871 ( .A1(n9383), .A2(n7138), .B1(n7137), .B2(n9374), .ZN(n7143)
         );
  NOR4_X1 U8872 ( .A1(n9876), .A2(n7141), .A3(n7140), .A4(n7139), .ZN(n7142)
         );
  AOI211_X1 U8873 ( .C1(n7144), .C2(n9053), .A(n7143), .B(n7142), .ZN(n7145)
         );
  OAI21_X1 U8874 ( .B1(n7146), .B2(n4444), .A(n7145), .ZN(P1_U3293) );
  XNOR2_X1 U8875 ( .A(n7236), .B(n10076), .ZN(n7231) );
  NAND2_X1 U8876 ( .A1(n7147), .A2(n8201), .ZN(n7148) );
  INV_X1 U8877 ( .A(n7235), .ZN(n7149) );
  AOI21_X1 U8878 ( .B1(n7151), .B2(n7150), .A(n7149), .ZN(n7158) );
  AOI21_X1 U8879 ( .B1(n8166), .B2(n7153), .A(n7152), .ZN(n7154) );
  OAI21_X1 U8880 ( .B1(n8158), .B2(n7482), .A(n7154), .ZN(n7156) );
  NOR2_X1 U8881 ( .A1(n8130), .A2(n7476), .ZN(n7155) );
  AOI211_X1 U8882 ( .C1(n8155), .C2(n8201), .A(n7156), .B(n7155), .ZN(n7157)
         );
  OAI21_X1 U8883 ( .B1(n7158), .B2(n8162), .A(n7157), .ZN(P2_U3170) );
  INV_X1 U8884 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U8885 ( .A(n10124), .B(P2_REG1_REG_8__SCAN_IN), .S(n7307), .Z(n7164)
         );
  INV_X1 U8886 ( .A(n7159), .ZN(n7160) );
  AOI22_X1 U8887 ( .A1(n7162), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n7161), .B2(
        n7160), .ZN(n7163) );
  NOR2_X1 U8888 ( .A1(n7163), .A2(n7164), .ZN(n7306) );
  AOI21_X1 U8889 ( .B1(n7164), .B2(n7163), .A(n7306), .ZN(n7181) );
  INV_X1 U8890 ( .A(n7165), .ZN(n7166) );
  NOR2_X1 U8891 ( .A1(n7167), .A2(n7166), .ZN(n7169) );
  MUX2_X1 U8892 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8227), .Z(n7308) );
  XNOR2_X1 U8893 ( .A(n7308), .B(n7307), .ZN(n7168) );
  NOR2_X1 U8894 ( .A1(n7169), .A2(n7168), .ZN(n7309) );
  AND2_X1 U8895 ( .A1(n7169), .A2(n7168), .ZN(n7170) );
  OAI21_X1 U8896 ( .B1(n7309), .B2(n7170), .A(n10060), .ZN(n7180) );
  INV_X1 U8897 ( .A(n7307), .ZN(n7315) );
  INV_X1 U8898 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8899 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n7521) );
  OAI21_X1 U8900 ( .B1(n9931), .B2(n7171), .A(n7521), .ZN(n7178) );
  INV_X1 U8901 ( .A(n7172), .ZN(n7174) );
  XNOR2_X1 U8902 ( .A(n7307), .B(n7581), .ZN(n7173) );
  OAI21_X1 U8903 ( .B1(n7175), .B2(n7174), .A(n7173), .ZN(n7314) );
  OR3_X1 U8904 ( .A1(n7175), .A2(n7174), .A3(n7173), .ZN(n7176) );
  AOI21_X1 U8905 ( .B1(n7314), .B2(n7176), .A(n10065), .ZN(n7177) );
  AOI211_X1 U8906 ( .C1(n10052), .C2(n7315), .A(n7178), .B(n7177), .ZN(n7179)
         );
  OAI211_X1 U8907 ( .C1(n7181), .C2(n9922), .A(n7180), .B(n7179), .ZN(P2_U3190) );
  NAND2_X1 U8908 ( .A1(n7182), .A2(n9022), .ZN(n7183) );
  OR2_X1 U8909 ( .A1(n9876), .A2(n7183), .ZN(n7197) );
  INV_X1 U8910 ( .A(n7197), .ZN(n7569) );
  NAND2_X1 U8911 ( .A1(n9378), .A2(n7184), .ZN(n7186) );
  AOI22_X1 U8912 ( .A1(n9876), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9865), .ZN(n7185) );
  OAI211_X1 U8913 ( .C1(n7187), .C2(n9381), .A(n7186), .B(n7185), .ZN(n7188)
         );
  AOI21_X1 U8914 ( .B1(n7569), .B2(n7189), .A(n7188), .ZN(n7190) );
  OAI21_X1 U8915 ( .B1(n7191), .B2(n9876), .A(n7190), .ZN(P1_U3292) );
  XNOR2_X1 U8916 ( .A(n7192), .B(n7194), .ZN(n7193) );
  OAI222_X1 U8917 ( .A1(n9262), .A2(n7619), .B1(n9261), .B2(n7298), .C1(n7193), 
        .C2(n9258), .ZN(n9888) );
  INV_X1 U8918 ( .A(n9888), .ZN(n7204) );
  NAND2_X1 U8919 ( .A1(n7195), .A2(n7194), .ZN(n7436) );
  OAI21_X1 U8920 ( .B1(n7195), .B2(n7194), .A(n7436), .ZN(n9890) );
  INV_X1 U8921 ( .A(n7302), .ZN(n9887) );
  INV_X1 U8922 ( .A(n7198), .ZN(n7278) );
  INV_X1 U8923 ( .A(n7448), .ZN(n7199) );
  OAI211_X1 U8924 ( .C1(n9887), .C2(n7278), .A(n7199), .B(n9331), .ZN(n9886)
         );
  AOI22_X1 U8925 ( .A1(n9876), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7297), .B2(
        n9865), .ZN(n7201) );
  NAND2_X1 U8926 ( .A1(n9378), .A2(n7302), .ZN(n7200) );
  OAI211_X1 U8927 ( .C1(n9886), .C2(n9381), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI21_X1 U8928 ( .B1(n9890), .B2(n9873), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8929 ( .B1(n7204), .B2(n9876), .A(n7203), .ZN(P1_U3287) );
  INV_X1 U8930 ( .A(n7205), .ZN(n7207) );
  OAI222_X1 U8931 ( .A1(P2_U3151), .A2(n8269), .B1(n8618), .B2(n7207), .C1(
        n7206), .C2(n7954), .ZN(P2_U3280) );
  INV_X1 U8932 ( .A(n9818), .ZN(n7758) );
  OAI222_X1 U8933 ( .A1(n9568), .A2(n7208), .B1(n9565), .B2(n7207), .C1(n7758), 
        .C2(n4288), .ZN(P1_U3340) );
  INV_X1 U8934 ( .A(n7209), .ZN(n7219) );
  INV_X1 U8935 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7211) );
  INV_X1 U8936 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7210) );
  OAI22_X1 U8937 ( .A1(n9383), .A2(n7211), .B1(n7210), .B2(n9374), .ZN(n7212)
         );
  AOI21_X1 U8938 ( .B1(n9378), .B2(n7213), .A(n7212), .ZN(n7214) );
  OAI21_X1 U8939 ( .B1(n9381), .B2(n7215), .A(n7214), .ZN(n7216) );
  AOI21_X1 U8940 ( .B1(n9873), .B2(n7217), .A(n7216), .ZN(n7218) );
  OAI21_X1 U8941 ( .B1(n9876), .B2(n7219), .A(n7218), .ZN(P1_U3291) );
  INV_X1 U8942 ( .A(n7220), .ZN(n7230) );
  NAND2_X1 U8943 ( .A1(n9863), .A2(n7221), .ZN(n7225) );
  NOR2_X1 U8944 ( .A1(n9374), .A2(n7222), .ZN(n7223) );
  AOI21_X1 U8945 ( .B1(n9876), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7223), .ZN(
        n7224) );
  OAI211_X1 U8946 ( .C1(n7226), .C2(n9869), .A(n7225), .B(n7224), .ZN(n7227)
         );
  AOI21_X1 U8947 ( .B1(n7228), .B2(n9873), .A(n7227), .ZN(n7229) );
  OAI21_X1 U8948 ( .B1(n7230), .B2(n9876), .A(n7229), .ZN(P1_U3289) );
  INV_X1 U8949 ( .A(n7231), .ZN(n7233) );
  NAND2_X1 U8950 ( .A1(n7233), .A2(n7232), .ZN(n7234) );
  XNOR2_X1 U8951 ( .A(n7236), .B(n10081), .ZN(n7256) );
  XNOR2_X1 U8952 ( .A(n7256), .B(n7482), .ZN(n7258) );
  XNOR2_X1 U8953 ( .A(n7259), .B(n7258), .ZN(n7244) );
  AOI21_X1 U8954 ( .B1(n8175), .B2(n4628), .A(n7237), .ZN(n7242) );
  INV_X1 U8955 ( .A(n10081), .ZN(n7377) );
  NAND2_X1 U8956 ( .A1(n8166), .A2(n7377), .ZN(n7241) );
  INV_X1 U8957 ( .A(n7238), .ZN(n7376) );
  NAND2_X1 U8958 ( .A1(n8179), .A2(n7376), .ZN(n7240) );
  NAND2_X1 U8959 ( .A1(n8155), .A2(n5683), .ZN(n7239) );
  NAND4_X1 U8960 ( .A1(n7242), .A2(n7241), .A3(n7240), .A4(n7239), .ZN(n7243)
         );
  AOI21_X1 U8961 ( .B1(n7244), .B2(n8169), .A(n7243), .ZN(n7245) );
  INV_X1 U8962 ( .A(n7245), .ZN(P2_U3167) );
  AND2_X1 U8963 ( .A1(n7247), .A2(n7246), .ZN(n7590) );
  NOR2_X1 U8964 ( .A1(n7721), .A2(n7590), .ZN(n7248) );
  INV_X1 U8965 ( .A(n7249), .ZN(n7255) );
  OAI22_X1 U8966 ( .A1(n7973), .A2(n8464), .B1(n8462), .B2(n7250), .ZN(n7251)
         );
  NOR2_X1 U8967 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  MUX2_X1 U8968 ( .A(n7253), .B(n5644), .S(n8447), .Z(n7254) );
  OAI21_X1 U8969 ( .B1(n8452), .B2(n7255), .A(n7254), .ZN(P2_U3231) );
  INV_X1 U8970 ( .A(n10085), .ZN(n7268) );
  NOR2_X1 U8971 ( .A1(n7256), .A2(n8200), .ZN(n7257) );
  XNOR2_X1 U8972 ( .A(n10085), .B(n8004), .ZN(n7457) );
  XNOR2_X1 U8973 ( .A(n7457), .B(n7465), .ZN(n7260) );
  NAND2_X1 U8974 ( .A1(n7261), .A2(n7260), .ZN(n7459) );
  OAI211_X1 U8975 ( .C1(n7261), .C2(n7260), .A(n7459), .B(n8169), .ZN(n7267)
         );
  INV_X1 U8976 ( .A(n7262), .ZN(n7415) );
  NAND2_X1 U8977 ( .A1(n8155), .A2(n8200), .ZN(n7264) );
  OAI211_X1 U8978 ( .C1(n7516), .C2(n8158), .A(n7264), .B(n7263), .ZN(n7265)
         );
  AOI21_X1 U8979 ( .B1(n7415), .B2(n8179), .A(n7265), .ZN(n7266) );
  OAI211_X1 U8980 ( .C1(n7268), .C2(n8182), .A(n7267), .B(n7266), .ZN(P2_U3179) );
  AOI22_X1 U8981 ( .A1(n8393), .A2(n7270), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8446), .ZN(n7274) );
  MUX2_X1 U8982 ( .A(n7271), .B(P2_REG2_REG_1__SCAN_IN), .S(n8447), .Z(n7272)
         );
  INV_X1 U8983 ( .A(n7272), .ZN(n7273) );
  OAI211_X1 U8984 ( .C1(n7275), .C2(n8452), .A(n7274), .B(n7273), .ZN(P2_U3232) );
  OAI21_X1 U8985 ( .B1(n7277), .B2(n8986), .A(n7276), .ZN(n9872) );
  AOI211_X1 U8986 ( .C1(n7280), .C2(n7279), .A(n9371), .B(n7278), .ZN(n9864)
         );
  NAND2_X1 U8987 ( .A1(n7282), .A2(n7281), .ZN(n7283) );
  XNOR2_X1 U8988 ( .A(n7283), .B(n8986), .ZN(n7284) );
  AOI222_X1 U8989 ( .A1(n9482), .A2(n7284), .B1(n9048), .B2(n9475), .C1(n9050), 
        .C2(n9474), .ZN(n9875) );
  INV_X1 U8990 ( .A(n9875), .ZN(n7285) );
  AOI211_X1 U8991 ( .C1(n9905), .C2(n9872), .A(n9864), .B(n7285), .ZN(n7292)
         );
  OAI22_X1 U8992 ( .A1(n9463), .A2(n9870), .B1(n9914), .B2(n7286), .ZN(n7287)
         );
  INV_X1 U8993 ( .A(n7287), .ZN(n7288) );
  OAI21_X1 U8994 ( .B1(n7292), .B2(n5572), .A(n7288), .ZN(P1_U3527) );
  INV_X1 U8995 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7289) );
  OAI22_X1 U8996 ( .A1(n9534), .A2(n9870), .B1(n9908), .B2(n7289), .ZN(n7290)
         );
  INV_X1 U8997 ( .A(n7290), .ZN(n7291) );
  OAI21_X1 U8998 ( .B1(n7292), .B2(n9906), .A(n7291), .ZN(P1_U3468) );
  INV_X1 U8999 ( .A(n7293), .ZN(n7294) );
  AOI21_X1 U9000 ( .B1(n7296), .B2(n7295), .A(n7294), .ZN(n7305) );
  NAND2_X1 U9001 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9107) );
  INV_X1 U9002 ( .A(n9107), .ZN(n7301) );
  INV_X1 U9003 ( .A(n7297), .ZN(n7299) );
  OAI22_X1 U9004 ( .A1(n8749), .A2(n7299), .B1(n7298), .B2(n8736), .ZN(n7300)
         );
  AOI211_X1 U9005 ( .C1(n8751), .C2(n9047), .A(n7301), .B(n7300), .ZN(n7304)
         );
  NAND2_X1 U9006 ( .A1(n8765), .A2(n7302), .ZN(n7303) );
  OAI211_X1 U9007 ( .C1(n7305), .C2(n8768), .A(n7304), .B(n7303), .ZN(P1_U3239) );
  AOI21_X1 U9008 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7307), .A(n7306), .ZN(
        n8255) );
  XOR2_X1 U9009 ( .A(n8232), .B(n8255), .Z(n8258) );
  XNOR2_X1 U9010 ( .A(n8258), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7324) );
  INV_X1 U9011 ( .A(n7308), .ZN(n7310) );
  AOI21_X1 U9012 ( .B1(n7315), .B2(n7310), .A(n7309), .ZN(n8213) );
  INV_X1 U9013 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8257) );
  MUX2_X1 U9014 ( .A(n7681), .B(n8257), .S(n8227), .Z(n7311) );
  NOR2_X1 U9015 ( .A1(n7311), .A2(n8256), .ZN(n8212) );
  INV_X1 U9016 ( .A(n8212), .ZN(n7312) );
  NAND2_X1 U9017 ( .A1(n7311), .A2(n8256), .ZN(n8211) );
  NAND2_X1 U9018 ( .A1(n7312), .A2(n8211), .ZN(n7313) );
  XNOR2_X1 U9019 ( .A(n8213), .B(n7313), .ZN(n7322) );
  OAI21_X1 U9020 ( .B1(n7315), .B2(n7581), .A(n7314), .ZN(n8231) );
  XNOR2_X1 U9021 ( .A(n8233), .B(n7681), .ZN(n7320) );
  NOR2_X1 U9022 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7316), .ZN(n7666) );
  INV_X1 U9023 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7317) );
  NOR2_X1 U9024 ( .A1(n9931), .A2(n7317), .ZN(n7318) );
  AOI211_X1 U9025 ( .C1(n8256), .C2(n10052), .A(n7666), .B(n7318), .ZN(n7319)
         );
  OAI21_X1 U9026 ( .B1(n7320), .B2(n10065), .A(n7319), .ZN(n7321) );
  AOI21_X1 U9027 ( .B1(n7322), .B2(n10060), .A(n7321), .ZN(n7323) );
  OAI21_X1 U9028 ( .B1(n7324), .B2(n9922), .A(n7323), .ZN(P2_U3191) );
  OR2_X1 U9029 ( .A1(n9876), .A2(n9258), .ZN(n7820) );
  NOR2_X2 U9030 ( .A1(n9876), .A2(n9261), .ZN(n9354) );
  AOI22_X1 U9031 ( .A1(n7325), .A2(n9863), .B1(n9354), .B2(n9052), .ZN(n7330)
         );
  OAI22_X1 U9032 ( .A1(n9383), .A2(n7326), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9374), .ZN(n7327) );
  AOI21_X1 U9033 ( .B1(n9378), .B2(n7328), .A(n7327), .ZN(n7329) );
  OAI211_X1 U9034 ( .C1(n7331), .C2(n9349), .A(n7330), .B(n7329), .ZN(n7332)
         );
  AOI21_X1 U9035 ( .B1(n9873), .B2(n7333), .A(n7332), .ZN(n7334) );
  OAI21_X1 U9036 ( .B1(n7820), .B2(n7335), .A(n7334), .ZN(P1_U3290) );
  INV_X1 U9037 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10138) );
  INV_X1 U9038 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9846) );
  INV_X1 U9039 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7336) );
  AOI22_X1 U9040 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9846), .B2(n7336), .ZN(n10142) );
  NOR2_X1 U9041 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7337) );
  AOI21_X1 U9042 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7337), .ZN(n10145) );
  NOR2_X1 U9043 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7338) );
  AOI21_X1 U9044 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7338), .ZN(n10148) );
  NOR2_X1 U9045 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7339) );
  AOI21_X1 U9046 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n7339), .ZN(n10151) );
  NOR2_X1 U9047 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7340) );
  AOI21_X1 U9048 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7340), .ZN(n10154) );
  NOR2_X1 U9049 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7341) );
  AOI21_X1 U9050 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7341), .ZN(n10157) );
  NOR2_X1 U9051 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7342) );
  AOI21_X1 U9052 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n7342), .ZN(n10160) );
  NOR2_X1 U9053 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7343) );
  AOI21_X1 U9054 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7343), .ZN(n10163) );
  NOR2_X1 U9055 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7344) );
  AOI21_X1 U9056 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7344), .ZN(n10172) );
  NOR2_X1 U9057 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7345) );
  AOI21_X1 U9058 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7345), .ZN(n10178) );
  NOR2_X1 U9059 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7346) );
  AOI21_X1 U9060 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7346), .ZN(n10175) );
  NOR2_X1 U9061 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7347) );
  AOI21_X1 U9062 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7347), .ZN(n10166) );
  NOR2_X1 U9063 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7348) );
  AOI21_X1 U9064 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7348), .ZN(n10169) );
  AND2_X1 U9065 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7349) );
  NOR2_X1 U9066 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7349), .ZN(n10132) );
  INV_X1 U9067 ( .A(n10132), .ZN(n10133) );
  INV_X1 U9068 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10135) );
  NAND3_X1 U9069 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U9070 ( .A1(n10135), .A2(n10134), .ZN(n10131) );
  NAND2_X1 U9071 ( .A1(n10133), .A2(n10131), .ZN(n10181) );
  NAND2_X1 U9072 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7350) );
  OAI21_X1 U9073 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7350), .ZN(n10180) );
  NOR2_X1 U9074 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  AOI21_X1 U9075 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10179), .ZN(n10184) );
  NAND2_X1 U9076 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7351) );
  OAI21_X1 U9077 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7351), .ZN(n10183) );
  NOR2_X1 U9078 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  AOI21_X1 U9079 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10182), .ZN(n10187) );
  NOR2_X1 U9080 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7352) );
  AOI21_X1 U9081 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7352), .ZN(n10186) );
  NAND2_X1 U9082 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  OAI21_X1 U9083 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10185), .ZN(n10168) );
  NAND2_X1 U9084 ( .A1(n10169), .A2(n10168), .ZN(n10167) );
  OAI21_X1 U9085 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10167), .ZN(n10165) );
  NAND2_X1 U9086 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  OAI21_X1 U9087 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10164), .ZN(n10174) );
  NAND2_X1 U9088 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  OAI21_X1 U9089 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10173), .ZN(n10177) );
  NAND2_X1 U9090 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  OAI21_X1 U9091 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10176), .ZN(n10171) );
  NAND2_X1 U9092 ( .A1(n10172), .A2(n10171), .ZN(n10170) );
  OAI21_X1 U9093 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10170), .ZN(n10162) );
  NAND2_X1 U9094 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  OAI21_X1 U9095 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10161), .ZN(n10159) );
  NAND2_X1 U9096 ( .A1(n10160), .A2(n10159), .ZN(n10158) );
  OAI21_X1 U9097 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10158), .ZN(n10156) );
  NAND2_X1 U9098 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  OAI21_X1 U9099 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10155), .ZN(n10153) );
  NAND2_X1 U9100 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  OAI21_X1 U9101 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10152), .ZN(n10150) );
  NAND2_X1 U9102 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  OAI21_X1 U9103 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10149), .ZN(n10147) );
  NAND2_X1 U9104 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  OAI21_X1 U9105 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10146), .ZN(n10144) );
  NAND2_X1 U9106 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  OAI21_X1 U9107 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10143), .ZN(n10141) );
  NAND2_X1 U9108 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  OAI21_X1 U9109 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10140), .ZN(n10137) );
  NAND2_X1 U9110 ( .A1(n10138), .A2(n10137), .ZN(n7353) );
  NOR2_X1 U9111 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  AOI21_X1 U9112 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7353), .A(n10136), .ZN(
        n7356) );
  XNOR2_X1 U9113 ( .A(n8278), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7355) );
  XNOR2_X1 U9114 ( .A(n7356), .B(n7355), .ZN(ADD_1068_U4) );
  OAI21_X1 U9115 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7550) );
  INV_X1 U9116 ( .A(n7550), .ZN(n7368) );
  OAI21_X1 U9117 ( .B1(n7361), .B2(n8994), .A(n7360), .ZN(n7553) );
  NAND2_X1 U9118 ( .A1(n7553), .A2(n9873), .ZN(n7367) );
  AOI211_X1 U9119 ( .C1(n7557), .C2(n4375), .A(n9371), .B(n7493), .ZN(n7548)
         );
  NOR2_X1 U9120 ( .A1(n7813), .A2(n9869), .ZN(n7365) );
  NAND2_X1 U9121 ( .A1(n9354), .A2(n9045), .ZN(n7363) );
  AOI22_X1 U9122 ( .A1(n9876), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7806), .B2(
        n9865), .ZN(n7362) );
  OAI211_X1 U9123 ( .C1(n7807), .C2(n9349), .A(n7363), .B(n7362), .ZN(n7364)
         );
  AOI211_X1 U9124 ( .C1(n7548), .C2(n9863), .A(n7365), .B(n7364), .ZN(n7366)
         );
  OAI211_X1 U9125 ( .C1(n7368), .C2(n7820), .A(n7367), .B(n7366), .ZN(P1_U3283) );
  INV_X1 U9126 ( .A(n7369), .ZN(n7371) );
  INV_X1 U9127 ( .A(n7407), .ZN(n7370) );
  AOI21_X1 U9128 ( .B1(n7371), .B2(n7373), .A(n7370), .ZN(n10082) );
  XNOR2_X1 U9129 ( .A(n7372), .B(n7373), .ZN(n7374) );
  AOI222_X1 U9130 ( .A1(n8460), .A2(n7374), .B1(n4628), .B2(n8455), .C1(n5683), 
        .C2(n8457), .ZN(n10080) );
  MUX2_X1 U9131 ( .A(n7375), .B(n10080), .S(n8474), .Z(n7379) );
  AOI22_X1 U9132 ( .A1(n8393), .A2(n7377), .B1(n8446), .B2(n7376), .ZN(n7378)
         );
  OAI211_X1 U9133 ( .C1(n10082), .C2(n8452), .A(n7379), .B(n7378), .ZN(
        P2_U3228) );
  INV_X1 U9134 ( .A(n7380), .ZN(n7382) );
  OAI222_X1 U9135 ( .A1(n8252), .A2(P2_U3151), .B1(n8618), .B2(n7382), .C1(
        n7381), .C2(n7954), .ZN(P2_U3279) );
  INV_X1 U9136 ( .A(n9831), .ZN(n7748) );
  OAI222_X1 U9137 ( .A1(n9568), .A2(n7383), .B1(n9565), .B2(n7382), .C1(n4288), 
        .C2(n7748), .ZN(P1_U3339) );
  AND2_X1 U9138 ( .A1(n7384), .A2(n8788), .ZN(n7441) );
  NAND2_X1 U9139 ( .A1(n7441), .A2(n4724), .ZN(n7440) );
  AND2_X1 U9140 ( .A1(n7440), .A2(n7385), .ZN(n7387) );
  INV_X1 U9141 ( .A(n7394), .ZN(n7386) );
  NAND2_X1 U9142 ( .A1(n7387), .A2(n7386), .ZN(n7500) );
  OAI211_X1 U9143 ( .C1(n7387), .C2(n7386), .A(n7500), .B(n9482), .ZN(n7390)
         );
  OAI22_X1 U9144 ( .A1(n7619), .A2(n9261), .B1(n7547), .B2(n9262), .ZN(n7388)
         );
  INV_X1 U9145 ( .A(n7388), .ZN(n7389) );
  AND2_X1 U9146 ( .A1(n7390), .A2(n7389), .ZN(n7400) );
  NAND2_X1 U9147 ( .A1(n7436), .A2(n7391), .ZN(n7393) );
  AND2_X1 U9148 ( .A1(n7393), .A2(n7392), .ZN(n7395) );
  OR2_X1 U9149 ( .A1(n7395), .A2(n7394), .ZN(n7396) );
  NAND2_X1 U9150 ( .A1(n7397), .A2(n7396), .ZN(n9896) );
  NAND2_X1 U9151 ( .A1(n9896), .A2(n7398), .ZN(n7399) );
  AOI21_X1 U9152 ( .B1(n7447), .B2(n7613), .A(n9371), .ZN(n7401) );
  NAND2_X1 U9153 ( .A1(n7401), .A2(n7506), .ZN(n9892) );
  AOI22_X1 U9154 ( .A1(n9876), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7618), .B2(
        n9865), .ZN(n7403) );
  NAND2_X1 U9155 ( .A1(n9378), .A2(n7613), .ZN(n7402) );
  OAI211_X1 U9156 ( .C1(n9892), .C2(n9381), .A(n7403), .B(n7402), .ZN(n7404)
         );
  AOI21_X1 U9157 ( .B1(n9896), .B2(n7569), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9158 ( .B1(n9898), .B2(n9876), .A(n7405), .ZN(P1_U3285) );
  NAND2_X1 U9159 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  XNOR2_X1 U9160 ( .A(n7408), .B(n7409), .ZN(n10086) );
  INV_X1 U9161 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7414) );
  XNOR2_X1 U9162 ( .A(n7410), .B(n7409), .ZN(n7413) );
  NAND2_X1 U9163 ( .A1(n8199), .A2(n8455), .ZN(n7411) );
  OAI21_X1 U9164 ( .B1(n7482), .B2(n8444), .A(n7411), .ZN(n7412) );
  AOI21_X1 U9165 ( .B1(n7413), .B2(n8460), .A(n7412), .ZN(n10089) );
  MUX2_X1 U9166 ( .A(n7414), .B(n10089), .S(n8474), .Z(n7417) );
  AOI22_X1 U9167 ( .A1(n8393), .A2(n10085), .B1(n8446), .B2(n7415), .ZN(n7416)
         );
  OAI211_X1 U9168 ( .C1(n10086), .C2(n8452), .A(n7417), .B(n7416), .ZN(
        P2_U3227) );
  INV_X1 U9169 ( .A(n7418), .ZN(n7420) );
  OAI222_X1 U9170 ( .A1(P2_U3151), .A2(n8272), .B1(n8618), .B2(n7420), .C1(
        n7419), .C2(n7954), .ZN(P2_U3278) );
  INV_X1 U9171 ( .A(n9840), .ZN(n7760) );
  OAI222_X1 U9172 ( .A1(n9568), .A2(n7421), .B1(n9565), .B2(n7420), .C1(n7760), 
        .C2(P1_U3086), .ZN(P1_U3338) );
  XNOR2_X1 U9173 ( .A(n7422), .B(n7424), .ZN(n7423) );
  AOI222_X1 U9174 ( .A1(n8460), .A2(n7423), .B1(n5683), .B2(n8455), .C1(n6359), 
        .C2(n8457), .ZN(n10071) );
  NAND2_X1 U9175 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  XNOR2_X1 U9176 ( .A(n7428), .B(n7427), .ZN(n10074) );
  AOI22_X1 U9177 ( .A1(n8393), .A2(n7430), .B1(n8446), .B2(n7429), .ZN(n7431)
         );
  OAI21_X1 U9178 ( .B1(n7432), .B2(n8474), .A(n7431), .ZN(n7433) );
  AOI21_X1 U9179 ( .B1(n10074), .B2(n8470), .A(n7433), .ZN(n7434) );
  OAI21_X1 U9180 ( .B1(n10071), .B2(n6946), .A(n7434), .ZN(P2_U3230) );
  NAND2_X1 U9181 ( .A1(n7436), .A2(n7435), .ZN(n7437) );
  NAND2_X1 U9182 ( .A1(n7437), .A2(n8798), .ZN(n7439) );
  OR2_X1 U9183 ( .A1(n7437), .A2(n8798), .ZN(n7438) );
  AND2_X1 U9184 ( .A1(n7439), .A2(n7438), .ZN(n7560) );
  OAI21_X1 U9185 ( .B1(n4724), .B2(n7441), .A(n7440), .ZN(n7444) );
  OAI22_X1 U9186 ( .A1(n7442), .A2(n9261), .B1(n7654), .B2(n9262), .ZN(n7443)
         );
  AOI21_X1 U9187 ( .B1(n7444), .B2(n9482), .A(n7443), .ZN(n7445) );
  OAI21_X1 U9188 ( .B1(n7560), .B2(n7446), .A(n7445), .ZN(n7565) );
  INV_X1 U9189 ( .A(n7565), .ZN(n7449) );
  OAI211_X1 U9190 ( .C1(n7448), .C2(n7453), .A(n7447), .B(n9331), .ZN(n7564)
         );
  OAI211_X1 U9191 ( .C1(n7560), .C2(n7450), .A(n7449), .B(n7564), .ZN(n7455)
         );
  OAI22_X1 U9192 ( .A1(n9463), .A2(n7453), .B1(n9914), .B2(n9656), .ZN(n7451)
         );
  AOI21_X1 U9193 ( .B1(n7455), .B2(n9914), .A(n7451), .ZN(n7452) );
  INV_X1 U9194 ( .A(n7452), .ZN(P1_U3529) );
  INV_X1 U9195 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9693) );
  OAI22_X1 U9196 ( .A1(n9534), .A2(n7453), .B1(n9544), .B2(n9693), .ZN(n7454)
         );
  AOI21_X1 U9197 ( .B1(n7455), .B2(n9908), .A(n7454), .ZN(n7456) );
  INV_X1 U9198 ( .A(n7456), .ZN(P1_U3474) );
  XNOR2_X1 U9199 ( .A(n10093), .B(n8016), .ZN(n7517) );
  XNOR2_X1 U9200 ( .A(n7517), .B(n7516), .ZN(n7464) );
  NAND2_X1 U9201 ( .A1(n7457), .A2(n4628), .ZN(n7458) );
  INV_X1 U9202 ( .A(n7464), .ZN(n7460) );
  INV_X1 U9203 ( .A(n7519), .ZN(n7462) );
  AOI21_X1 U9204 ( .B1(n7464), .B2(n7463), .A(n7462), .ZN(n7471) );
  NOR2_X1 U9205 ( .A1(n8177), .A2(n7465), .ZN(n7466) );
  AOI211_X1 U9206 ( .C1(n8175), .C2(n8198), .A(n7467), .B(n7466), .ZN(n7468)
         );
  OAI21_X1 U9207 ( .B1(n7596), .B2(n8130), .A(n7468), .ZN(n7469) );
  AOI21_X1 U9208 ( .B1(n10093), .B2(n8166), .A(n7469), .ZN(n7470) );
  OAI21_X1 U9209 ( .B1(n7471), .B2(n8162), .A(n7470), .ZN(P2_U3153) );
  AND2_X1 U9210 ( .A1(n7473), .A2(n7472), .ZN(n7475) );
  OAI21_X1 U9211 ( .B1(n7475), .B2(n7480), .A(n7474), .ZN(n10079) );
  OAI22_X1 U9212 ( .A1(n8449), .A2(n10076), .B1(n7476), .B2(n8462), .ZN(n7484)
         );
  INV_X1 U9213 ( .A(n7477), .ZN(n7478) );
  AOI21_X1 U9214 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7481) );
  OAI222_X1 U9215 ( .A1(n8442), .A2(n7482), .B1(n8444), .B2(n7974), .C1(n8440), 
        .C2(n7481), .ZN(n10077) );
  MUX2_X1 U9216 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10077), .S(n8474), .Z(n7483)
         );
  AOI211_X1 U9217 ( .C1(n8470), .C2(n10079), .A(n7484), .B(n7483), .ZN(n7485)
         );
  INV_X1 U9218 ( .A(n7485), .ZN(P2_U3229) );
  OAI21_X1 U9219 ( .B1(n8996), .B2(n7487), .A(n7486), .ZN(n7488) );
  NAND2_X1 U9220 ( .A1(n7488), .A2(n9482), .ZN(n7534) );
  OAI21_X1 U9221 ( .B1(n7491), .B2(n7490), .A(n7489), .ZN(n7536) );
  OAI211_X1 U9222 ( .C1(n7493), .C2(n7492), .A(n9331), .B(n7604), .ZN(n7532)
         );
  NAND2_X1 U9223 ( .A1(n9354), .A2(n9044), .ZN(n7495) );
  AOI22_X1 U9224 ( .A1(n9876), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7873), .B2(
        n9865), .ZN(n7494) );
  OAI211_X1 U9225 ( .C1(n7875), .C2(n9349), .A(n7495), .B(n7494), .ZN(n7496)
         );
  AOI21_X1 U9226 ( .B1(n7877), .B2(n9378), .A(n7496), .ZN(n7497) );
  OAI21_X1 U9227 ( .B1(n7532), .B2(n9381), .A(n7497), .ZN(n7498) );
  AOI21_X1 U9228 ( .B1(n7536), .B2(n9873), .A(n7498), .ZN(n7499) );
  OAI21_X1 U9229 ( .B1(n9876), .B2(n7534), .A(n7499), .ZN(P1_U3282) );
  NAND2_X1 U9230 ( .A1(n7500), .A2(n8795), .ZN(n7501) );
  XOR2_X1 U9231 ( .A(n7505), .B(n7501), .Z(n7502) );
  OAI22_X1 U9232 ( .A1(n7502), .A2(n9258), .B1(n7654), .B2(n9261), .ZN(n9902)
         );
  INV_X1 U9233 ( .A(n9902), .ZN(n7515) );
  OAI21_X1 U9234 ( .B1(n7503), .B2(n7505), .A(n7504), .ZN(n9904) );
  XNOR2_X1 U9235 ( .A(n7506), .B(n4449), .ZN(n7507) );
  AOI22_X1 U9236 ( .A1(n7507), .A2(n9331), .B1(n9475), .B2(n9044), .ZN(n9900)
         );
  INV_X1 U9237 ( .A(n7652), .ZN(n7508) );
  OAI22_X1 U9238 ( .A1(n9383), .A2(n7509), .B1(n7508), .B2(n9374), .ZN(n7510)
         );
  AOI21_X1 U9239 ( .B1(n9378), .B2(n7511), .A(n7510), .ZN(n7512) );
  OAI21_X1 U9240 ( .B1(n9900), .B2(n9381), .A(n7512), .ZN(n7513) );
  AOI21_X1 U9241 ( .B1(n9904), .B2(n9873), .A(n7513), .ZN(n7514) );
  OAI21_X1 U9242 ( .B1(n7515), .B2(n9876), .A(n7514), .ZN(P1_U3284) );
  NAND2_X1 U9243 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  INV_X2 U9244 ( .A(n8004), .ZN(n8016) );
  XNOR2_X1 U9245 ( .A(n10096), .B(n8016), .ZN(n7662) );
  XNOR2_X1 U9246 ( .A(n7662), .B(n7661), .ZN(n7520) );
  XNOR2_X1 U9247 ( .A(n7665), .B(n7520), .ZN(n7526) );
  NAND2_X1 U9248 ( .A1(n8155), .A2(n8199), .ZN(n7522) );
  OAI211_X1 U9249 ( .C1(n7577), .C2(n8158), .A(n7522), .B(n7521), .ZN(n7524)
         );
  NOR2_X1 U9250 ( .A1(n8130), .A2(n7580), .ZN(n7523) );
  AOI211_X1 U9251 ( .C1(n10096), .C2(n8166), .A(n7524), .B(n7523), .ZN(n7525)
         );
  OAI21_X1 U9252 ( .B1(n7526), .B2(n8162), .A(n7525), .ZN(P2_U3161) );
  INV_X1 U9253 ( .A(n7527), .ZN(n7529) );
  OAI222_X1 U9254 ( .A1(P2_U3151), .A2(n9738), .B1(n8618), .B2(n7529), .C1(
        n7528), .C2(n7954), .ZN(P2_U3277) );
  INV_X1 U9255 ( .A(n7761), .ZN(n9855) );
  OAI222_X1 U9256 ( .A1(n9568), .A2(n7530), .B1(n9565), .B2(n7529), .C1(n9855), 
        .C2(n4288), .ZN(P1_U3337) );
  OAI22_X1 U9257 ( .A1(n7656), .A2(n9261), .B1(n7875), .B2(n9262), .ZN(n7531)
         );
  INV_X1 U9258 ( .A(n7531), .ZN(n7533) );
  NAND3_X1 U9259 ( .A1(n7534), .A2(n7533), .A3(n7532), .ZN(n7535) );
  AOI21_X1 U9260 ( .B1(n7536), .B2(n9905), .A(n7535), .ZN(n7539) );
  INV_X1 U9261 ( .A(n9534), .ZN(n7696) );
  AOI22_X1 U9262 ( .A1(n7877), .A2(n7696), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9906), .ZN(n7537) );
  OAI21_X1 U9263 ( .B1(n7539), .B2(n9906), .A(n7537), .ZN(P1_U3486) );
  INV_X1 U9264 ( .A(n9463), .ZN(n7694) );
  AOI22_X1 U9265 ( .A1(n7877), .A2(n7694), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n5572), .ZN(n7538) );
  OAI21_X1 U9266 ( .B1(n7539), .B2(n5572), .A(n7538), .ZN(P1_U3533) );
  AOI22_X1 U9267 ( .A1(n8760), .A2(n9048), .B1(n8759), .B2(n7561), .ZN(n7540)
         );
  NAND2_X1 U9268 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(n4288), .ZN(n9120) );
  OAI211_X1 U9269 ( .C1(n7654), .C2(n8762), .A(n7540), .B(n9120), .ZN(n7545)
         );
  AOI21_X1 U9270 ( .B1(n7543), .B2(n7541), .A(n4378), .ZN(n7542) );
  AOI211_X1 U9271 ( .C1(n4376), .C2(n7543), .A(n8768), .B(n7542), .ZN(n7544)
         );
  AOI211_X1 U9272 ( .C1(n7562), .C2(n8765), .A(n7545), .B(n7544), .ZN(n7546)
         );
  INV_X1 U9273 ( .A(n7546), .ZN(P1_U3213) );
  OAI22_X1 U9274 ( .A1(n7547), .A2(n9261), .B1(n7807), .B2(n9262), .ZN(n7549)
         );
  AOI211_X1 U9275 ( .C1(n9482), .C2(n7550), .A(n7549), .B(n7548), .ZN(n7551)
         );
  INV_X1 U9276 ( .A(n7551), .ZN(n7552) );
  AOI21_X1 U9277 ( .B1(n7553), .B2(n9905), .A(n7552), .ZN(n7559) );
  INV_X1 U9278 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7554) );
  OAI22_X1 U9279 ( .A1(n7813), .A2(n9534), .B1(n9544), .B2(n7554), .ZN(n7555)
         );
  INV_X1 U9280 ( .A(n7555), .ZN(n7556) );
  OAI21_X1 U9281 ( .B1(n7559), .B2(n9906), .A(n7556), .ZN(P1_U3483) );
  INV_X1 U9282 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7752) );
  AOI22_X1 U9283 ( .A1(n7557), .A2(n7694), .B1(n5572), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7558) );
  OAI21_X1 U9284 ( .B1(n7559), .B2(n5572), .A(n7558), .ZN(P1_U3532) );
  INV_X1 U9285 ( .A(n7560), .ZN(n7568) );
  AOI22_X1 U9286 ( .A1(n9378), .A2(n7562), .B1(n9865), .B2(n7561), .ZN(n7563)
         );
  OAI21_X1 U9287 ( .B1(n7564), .B2(n9381), .A(n7563), .ZN(n7567) );
  MUX2_X1 U9288 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7565), .S(n9383), .Z(n7566)
         );
  AOI211_X1 U9289 ( .C1(n7569), .C2(n7568), .A(n7567), .B(n7566), .ZN(n7570)
         );
  INV_X1 U9290 ( .A(n7570), .ZN(P1_U3286) );
  INV_X1 U9291 ( .A(n7583), .ZN(n7574) );
  NAND3_X1 U9292 ( .A1(n7572), .A2(n7574), .A3(n7573), .ZN(n7575) );
  NAND2_X1 U9293 ( .A1(n7571), .A2(n7575), .ZN(n7579) );
  NAND2_X1 U9294 ( .A1(n8199), .A2(n8457), .ZN(n7576) );
  OAI21_X1 U9295 ( .B1(n7577), .B2(n8442), .A(n7576), .ZN(n7578) );
  AOI21_X1 U9296 ( .B1(n7579), .B2(n8460), .A(n7578), .ZN(n10099) );
  OAI22_X1 U9297 ( .A1(n8474), .A2(n7581), .B1(n7580), .B2(n8462), .ZN(n7582)
         );
  AOI21_X1 U9298 ( .B1(n8393), .B2(n10096), .A(n7582), .ZN(n7586) );
  XNOR2_X1 U9299 ( .A(n7584), .B(n7583), .ZN(n10094) );
  NAND2_X1 U9300 ( .A1(n10094), .A2(n8470), .ZN(n7585) );
  OAI211_X1 U9301 ( .C1(n10099), .C2(n8447), .A(n7586), .B(n7585), .ZN(
        P2_U3225) );
  OAI21_X1 U9302 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n10090) );
  AND2_X1 U9303 ( .A1(n8474), .A2(n7590), .ZN(n8035) );
  INV_X1 U9304 ( .A(n8035), .ZN(n7729) );
  INV_X1 U9305 ( .A(n7721), .ZN(n7595) );
  OAI21_X1 U9306 ( .B1(n7591), .B2(n5737), .A(n7572), .ZN(n7592) );
  NAND2_X1 U9307 ( .A1(n7592), .A2(n8460), .ZN(n7594) );
  AOI22_X1 U9308 ( .A1(n8457), .A2(n4628), .B1(n8198), .B2(n8455), .ZN(n7593)
         );
  OAI211_X1 U9309 ( .C1(n7595), .C2(n10090), .A(n7594), .B(n7593), .ZN(n10091)
         );
  NAND2_X1 U9310 ( .A1(n10091), .A2(n8474), .ZN(n7599) );
  OAI22_X1 U9311 ( .A1(n8474), .A2(n7056), .B1(n7596), .B2(n8462), .ZN(n7597)
         );
  AOI21_X1 U9312 ( .B1(n8393), .B2(n10093), .A(n7597), .ZN(n7598) );
  OAI211_X1 U9313 ( .C1(n10090), .C2(n7729), .A(n7599), .B(n7598), .ZN(
        P2_U3226) );
  XNOR2_X1 U9314 ( .A(n7600), .B(n7602), .ZN(n7644) );
  OAI21_X1 U9315 ( .B1(n7603), .B2(n7602), .A(n7601), .ZN(n7642) );
  AOI21_X1 U9316 ( .B1(n7604), .B2(n7947), .A(n9371), .ZN(n7605) );
  AND2_X1 U9317 ( .A1(n7605), .A2(n7630), .ZN(n7641) );
  NAND2_X1 U9318 ( .A1(n7641), .A2(n9863), .ZN(n7610) );
  NAND2_X1 U9319 ( .A1(n9354), .A2(n9043), .ZN(n7607) );
  AOI22_X1 U9320 ( .A1(n9876), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7944), .B2(
        n9865), .ZN(n7606) );
  OAI211_X1 U9321 ( .C1(n8626), .C2(n9349), .A(n7607), .B(n7606), .ZN(n7608)
         );
  AOI21_X1 U9322 ( .B1(n7947), .B2(n9378), .A(n7608), .ZN(n7609) );
  NAND2_X1 U9323 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  AOI21_X1 U9324 ( .B1(n7642), .B2(n9873), .A(n7611), .ZN(n7612) );
  OAI21_X1 U9325 ( .B1(n7820), .B2(n7644), .A(n7612), .ZN(P1_U3281) );
  INV_X1 U9326 ( .A(n7613), .ZN(n9893) );
  OAI21_X1 U9327 ( .B1(n7614), .B2(n7616), .A(n7615), .ZN(n7617) );
  NAND2_X1 U9328 ( .A1(n7617), .A2(n8746), .ZN(n7624) );
  NAND2_X1 U9329 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9133) );
  INV_X1 U9330 ( .A(n9133), .ZN(n7622) );
  INV_X1 U9331 ( .A(n7618), .ZN(n7620) );
  OAI22_X1 U9332 ( .A1(n8749), .A2(n7620), .B1(n7619), .B2(n8736), .ZN(n7621)
         );
  AOI211_X1 U9333 ( .C1(n8751), .C2(n9045), .A(n7622), .B(n7621), .ZN(n7623)
         );
  OAI211_X1 U9334 ( .C1(n9893), .C2(n8754), .A(n7624), .B(n7623), .ZN(P1_U3221) );
  INV_X1 U9335 ( .A(n7625), .ZN(n7965) );
  OAI222_X1 U9336 ( .A1(n6010), .A2(P2_U3151), .B1(n8618), .B2(n7965), .C1(
        n7626), .C2(n7954), .ZN(P2_U3276) );
  XNOR2_X1 U9337 ( .A(n7627), .B(n8998), .ZN(n7692) );
  OAI21_X1 U9338 ( .B1(n7629), .B2(n8998), .A(n7628), .ZN(n7690) );
  NAND2_X1 U9339 ( .A1(n8716), .A2(n7630), .ZN(n7631) );
  NAND2_X1 U9340 ( .A1(n7631), .A2(n9331), .ZN(n7632) );
  NOR2_X1 U9341 ( .A1(n7706), .A2(n7632), .ZN(n7689) );
  NAND2_X1 U9342 ( .A1(n7689), .A2(n9863), .ZN(n7637) );
  NAND2_X1 U9343 ( .A1(n9354), .A2(n9042), .ZN(n7634) );
  AOI22_X1 U9344 ( .A1(n9876), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8712), .B2(
        n9865), .ZN(n7633) );
  OAI211_X1 U9345 ( .C1(n8714), .C2(n9349), .A(n7634), .B(n7633), .ZN(n7635)
         );
  AOI21_X1 U9346 ( .B1(n8716), .B2(n9378), .A(n7635), .ZN(n7636) );
  NAND2_X1 U9347 ( .A1(n7637), .A2(n7636), .ZN(n7638) );
  AOI21_X1 U9348 ( .B1(n7690), .B2(n9873), .A(n7638), .ZN(n7639) );
  OAI21_X1 U9349 ( .B1(n7820), .B2(n7692), .A(n7639), .ZN(P1_U3280) );
  OAI22_X1 U9350 ( .A1(n7807), .A2(n9261), .B1(n8626), .B2(n9262), .ZN(n7640)
         );
  AOI211_X1 U9351 ( .C1(n7642), .C2(n9905), .A(n7641), .B(n7640), .ZN(n7643)
         );
  OAI21_X1 U9352 ( .B1(n9258), .B2(n7644), .A(n7643), .ZN(n7645) );
  INV_X1 U9353 ( .A(n7645), .ZN(n7648) );
  AOI22_X1 U9354 ( .A1(n7947), .A2(n7694), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n5572), .ZN(n7646) );
  OAI21_X1 U9355 ( .B1(n7648), .B2(n5572), .A(n7646), .ZN(P1_U3534) );
  AOI22_X1 U9356 ( .A1(n7947), .A2(n7696), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n9906), .ZN(n7647) );
  OAI21_X1 U9357 ( .B1(n7648), .B2(n9906), .A(n7647), .ZN(P1_U3489) );
  XNOR2_X1 U9358 ( .A(n7649), .B(n7650), .ZN(n7651) );
  NAND2_X1 U9359 ( .A1(n7651), .A2(n8746), .ZN(n7660) );
  NAND2_X1 U9360 ( .A1(n8759), .A2(n7652), .ZN(n7653) );
  OAI21_X1 U9361 ( .B1(n8736), .B2(n7654), .A(n7653), .ZN(n7658) );
  OAI21_X1 U9362 ( .B1(n8762), .B2(n7656), .A(n7655), .ZN(n7657) );
  NOR2_X1 U9363 ( .A1(n7658), .A2(n7657), .ZN(n7659) );
  OAI211_X1 U9364 ( .C1(n4449), .C2(n8754), .A(n7660), .B(n7659), .ZN(P1_U3231) );
  AND2_X1 U9365 ( .A1(n7662), .A2(n7661), .ZN(n7664) );
  INV_X1 U9366 ( .A(n7662), .ZN(n7663) );
  XNOR2_X1 U9367 ( .A(n7784), .B(n8016), .ZN(n7787) );
  XNOR2_X1 U9368 ( .A(n7787), .B(n8197), .ZN(n7789) );
  XOR2_X1 U9369 ( .A(n7790), .B(n7789), .Z(n7673) );
  NAND2_X1 U9370 ( .A1(n7784), .A2(n8166), .ZN(n7671) );
  AOI21_X1 U9371 ( .B1(n8175), .B2(n8196), .A(n7666), .ZN(n7670) );
  INV_X1 U9372 ( .A(n7680), .ZN(n7667) );
  NAND2_X1 U9373 ( .A1(n8179), .A2(n7667), .ZN(n7669) );
  NAND2_X1 U9374 ( .A1(n8155), .A2(n8198), .ZN(n7668) );
  NAND4_X1 U9375 ( .A1(n7671), .A2(n7670), .A3(n7669), .A4(n7668), .ZN(n7672)
         );
  AOI21_X1 U9376 ( .B1(n7673), .B2(n8169), .A(n7672), .ZN(n7674) );
  INV_X1 U9377 ( .A(n7674), .ZN(P2_U3171) );
  INV_X1 U9378 ( .A(n7675), .ZN(n7683) );
  NAND3_X1 U9379 ( .A1(n7571), .A2(n7683), .A3(n7676), .ZN(n7677) );
  NAND2_X1 U9380 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  AOI222_X1 U9381 ( .A1(n8460), .A2(n7679), .B1(n8196), .B2(n8455), .C1(n8198), 
        .C2(n8457), .ZN(n7773) );
  OAI22_X1 U9382 ( .A1(n8474), .A2(n7681), .B1(n7680), .B2(n8462), .ZN(n7686)
         );
  OAI21_X1 U9383 ( .B1(n7684), .B2(n7683), .A(n7682), .ZN(n7774) );
  NOR2_X1 U9384 ( .A1(n7774), .A2(n8452), .ZN(n7685) );
  AOI211_X1 U9385 ( .C1(n8393), .C2(n7784), .A(n7686), .B(n7685), .ZN(n7687)
         );
  OAI21_X1 U9386 ( .B1(n7773), .B2(n6946), .A(n7687), .ZN(P2_U3224) );
  OAI22_X1 U9387 ( .A1(n7875), .A2(n9261), .B1(n8714), .B2(n9262), .ZN(n7688)
         );
  AOI211_X1 U9388 ( .C1(n7690), .C2(n9905), .A(n7689), .B(n7688), .ZN(n7691)
         );
  OAI21_X1 U9389 ( .B1(n9258), .B2(n7692), .A(n7691), .ZN(n7693) );
  INV_X1 U9390 ( .A(n7693), .ZN(n7698) );
  AOI22_X1 U9391 ( .A1(n8716), .A2(n7694), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n5572), .ZN(n7695) );
  OAI21_X1 U9392 ( .B1(n7698), .B2(n5572), .A(n7695), .ZN(P1_U3535) );
  AOI22_X1 U9393 ( .A1(n8716), .A2(n7696), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9906), .ZN(n7697) );
  OAI21_X1 U9394 ( .B1(n7698), .B2(n9906), .A(n7697), .ZN(P1_U3492) );
  INV_X1 U9395 ( .A(n7699), .ZN(n7716) );
  OAI222_X1 U9396 ( .A1(P2_U3151), .A2(n7701), .B1(n8618), .B2(n7716), .C1(
        n7700), .C2(n7954), .ZN(P2_U3275) );
  OAI21_X1 U9397 ( .B1(n7703), .B2(n9000), .A(n7702), .ZN(n7832) );
  INV_X1 U9398 ( .A(n7832), .ZN(n7715) );
  AOI21_X1 U9399 ( .B1(n7704), .B2(n9000), .A(n9258), .ZN(n7705) );
  AND2_X1 U9400 ( .A1(n7705), .A2(n7815), .ZN(n7830) );
  INV_X1 U9401 ( .A(n7706), .ZN(n7707) );
  AOI211_X1 U9402 ( .C1(n7708), .C2(n7707), .A(n9371), .B(n7821), .ZN(n7829)
         );
  NAND2_X1 U9403 ( .A1(n7829), .A2(n9863), .ZN(n7712) );
  AOI22_X1 U9404 ( .A1(n9876), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8625), .B2(
        n9865), .ZN(n7709) );
  OAI21_X1 U9405 ( .B1(n9349), .B2(n8673), .A(n7709), .ZN(n7710) );
  AOI21_X1 U9406 ( .B1(n9354), .B2(n9041), .A(n7710), .ZN(n7711) );
  OAI211_X1 U9407 ( .C1(n8632), .C2(n9869), .A(n7712), .B(n7711), .ZN(n7713)
         );
  AOI21_X1 U9408 ( .B1(n7830), .B2(n9383), .A(n7713), .ZN(n7714) );
  OAI21_X1 U9409 ( .B1(n7715), .B2(n9385), .A(n7714), .ZN(P1_U3279) );
  OAI222_X1 U9410 ( .A1(n9568), .A2(n7717), .B1(n4288), .B2(n9018), .C1(n9565), 
        .C2(n7716), .ZN(P1_U3335) );
  XOR2_X1 U9411 ( .A(n7720), .B(n7718), .Z(n7722) );
  INV_X1 U9412 ( .A(n7722), .ZN(n10102) );
  XNOR2_X1 U9413 ( .A(n7719), .B(n7720), .ZN(n7725) );
  NAND2_X1 U9414 ( .A1(n7722), .A2(n7721), .ZN(n7724) );
  AOI22_X1 U9415 ( .A1(n8197), .A2(n8457), .B1(n8455), .B2(n8195), .ZN(n7723)
         );
  OAI211_X1 U9416 ( .C1(n8440), .C2(n7725), .A(n7724), .B(n7723), .ZN(n10104)
         );
  NAND2_X1 U9417 ( .A1(n10104), .A2(n8474), .ZN(n7728) );
  INV_X1 U9418 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9653) );
  OAI22_X1 U9419 ( .A1(n8474), .A2(n9653), .B1(n7793), .B2(n8462), .ZN(n7726)
         );
  AOI21_X1 U9420 ( .B1(n7799), .B2(n8393), .A(n7726), .ZN(n7727) );
  OAI211_X1 U9421 ( .C1(n10102), .C2(n7729), .A(n7728), .B(n7727), .ZN(
        P2_U3223) );
  INV_X1 U9422 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U9423 ( .A1(n9794), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7730) );
  OAI21_X1 U9424 ( .B1(n9794), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7730), .ZN(
        n9787) );
  OR2_X1 U9425 ( .A1(n7749), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U9426 ( .A1(n7732), .A2(n7731), .ZN(n9753) );
  INV_X1 U9427 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7733) );
  MUX2_X1 U9428 ( .A(n7733), .B(P1_REG2_REG_10__SCAN_IN), .S(n9761), .Z(n9754)
         );
  OR2_X1 U9429 ( .A1(n9753), .A2(n9754), .ZN(n9751) );
  NAND2_X1 U9430 ( .A1(n9761), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U9431 ( .A1(n9751), .A2(n7734), .ZN(n9151) );
  INV_X1 U9432 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7735) );
  XNOR2_X1 U9433 ( .A(n9149), .B(n7735), .ZN(n9152) );
  NAND2_X1 U9434 ( .A1(n9151), .A2(n9152), .ZN(n9150) );
  NAND2_X1 U9435 ( .A1(n9149), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U9436 ( .A1(n9150), .A2(n7736), .ZN(n9776) );
  NAND2_X1 U9437 ( .A1(n7756), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7738) );
  OR2_X1 U9438 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7756), .ZN(n7737) );
  NAND2_X1 U9439 ( .A1(n7738), .A2(n7737), .ZN(n9775) );
  OAI21_X1 U9440 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7756), .A(n9778), .ZN(
        n9788) );
  NOR2_X1 U9441 ( .A1(n9787), .A2(n9788), .ZN(n9786) );
  AOI21_X1 U9442 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9794), .A(n9786), .ZN(
        n9803) );
  NAND2_X1 U9443 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9806), .ZN(n7739) );
  OAI21_X1 U9444 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9806), .A(n7739), .ZN(
        n9802) );
  NOR2_X1 U9445 ( .A1(n9803), .A2(n9802), .ZN(n9801) );
  AOI21_X1 U9446 ( .B1(n9806), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9801), .ZN(
        n7740) );
  NOR2_X1 U9447 ( .A1(n7740), .A2(n7758), .ZN(n7741) );
  INV_X1 U9448 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9814) );
  XOR2_X1 U9449 ( .A(n9818), .B(n7740), .Z(n9815) );
  NOR2_X1 U9450 ( .A1(n9814), .A2(n9815), .ZN(n9813) );
  NOR2_X1 U9451 ( .A1(n7741), .A2(n9813), .ZN(n9824) );
  INV_X1 U9452 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7742) );
  AOI22_X1 U9453 ( .A1(n9831), .A2(n7742), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n7748), .ZN(n9823) );
  NOR2_X1 U9454 ( .A1(n9824), .A2(n9823), .ZN(n9822) );
  AOI21_X1 U9455 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9831), .A(n9822), .ZN(
        n9836) );
  INV_X1 U9456 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9376) );
  XNOR2_X1 U9457 ( .A(n9840), .B(n9376), .ZN(n9835) );
  NAND2_X1 U9458 ( .A1(n9836), .A2(n9835), .ZN(n7744) );
  OR2_X1 U9459 ( .A1(n9840), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7743) );
  NAND2_X1 U9460 ( .A1(n7744), .A2(n7743), .ZN(n9849) );
  NAND2_X1 U9461 ( .A1(n7761), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7746) );
  OR2_X1 U9462 ( .A1(n7761), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U9463 ( .A1(n7746), .A2(n7745), .ZN(n9848) );
  NAND2_X1 U9464 ( .A1(n9858), .A2(n7746), .ZN(n7747) );
  XNOR2_X1 U9465 ( .A(n7747), .B(n9333), .ZN(n7765) );
  INV_X1 U9466 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U9467 ( .A1(n9831), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9672), .B2(
        n7748), .ZN(n9830) );
  XNOR2_X1 U9468 ( .A(n9794), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9790) );
  OR2_X1 U9469 ( .A1(n7749), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U9470 ( .A1(n7751), .A2(n7750), .ZN(n9757) );
  MUX2_X1 U9471 ( .A(n7752), .B(P1_REG1_REG_10__SCAN_IN), .S(n9761), .Z(n9758)
         );
  OR2_X1 U9472 ( .A1(n9757), .A2(n9758), .ZN(n9755) );
  NAND2_X1 U9473 ( .A1(n9761), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U9474 ( .A1(n9755), .A2(n7753), .ZN(n9155) );
  INV_X1 U9475 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7754) );
  XNOR2_X1 U9476 ( .A(n9149), .B(n7754), .ZN(n9154) );
  NAND2_X1 U9477 ( .A1(n9155), .A2(n9154), .ZN(n9153) );
  NAND2_X1 U9478 ( .A1(n9149), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U9479 ( .A1(n9153), .A2(n7755), .ZN(n9772) );
  XNOR2_X1 U9480 ( .A(n7756), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n9771) );
  OAI21_X1 U9481 ( .B1(n7756), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9774), .ZN(
        n9791) );
  NOR2_X1 U9482 ( .A1(n9790), .A2(n9791), .ZN(n9789) );
  AOI21_X1 U9483 ( .B1(n9794), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9789), .ZN(
        n9800) );
  XNOR2_X1 U9484 ( .A(n9806), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9799) );
  NOR2_X1 U9485 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  AOI21_X1 U9486 ( .B1(n9806), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9798), .ZN(
        n7757) );
  NOR2_X1 U9487 ( .A1(n7757), .A2(n7758), .ZN(n7759) );
  INV_X1 U9488 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9811) );
  XNOR2_X1 U9489 ( .A(n7758), .B(n7757), .ZN(n9812) );
  NOR2_X1 U9490 ( .A1(n9811), .A2(n9812), .ZN(n9810) );
  NOR2_X1 U9491 ( .A1(n7759), .A2(n9810), .ZN(n9829) );
  NAND2_X1 U9492 ( .A1(n9830), .A2(n9829), .ZN(n9828) );
  OAI21_X1 U9493 ( .B1(n9831), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9828), .ZN(
        n9838) );
  INV_X1 U9494 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9489) );
  XNOR2_X1 U9495 ( .A(n9840), .B(n9489), .ZN(n9837) );
  AOI22_X1 U9496 ( .A1(n9838), .A2(n9837), .B1(n9489), .B2(n7760), .ZN(n9853)
         );
  INV_X1 U9497 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9483) );
  AND2_X1 U9498 ( .A1(n7761), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7762) );
  AOI21_X1 U9499 ( .B1(n9483), .B2(n9855), .A(n7762), .ZN(n9852) );
  NAND2_X1 U9500 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  INV_X1 U9501 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U9502 ( .A1(n9851), .A2(n7763), .ZN(n7764) );
  INV_X1 U9503 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9471) );
  XNOR2_X1 U9504 ( .A(n7764), .B(n9471), .ZN(n7766) );
  AOI22_X1 U9505 ( .A1(n7765), .A2(n9842), .B1(n9850), .B2(n7766), .ZN(n7770)
         );
  INV_X1 U9506 ( .A(n7765), .ZN(n7768) );
  OAI21_X1 U9507 ( .B1(n7766), .B2(n9809), .A(n9856), .ZN(n7767) );
  AOI21_X1 U9508 ( .B1(n7768), .B2(n9842), .A(n7767), .ZN(n7769) );
  MUX2_X1 U9509 ( .A(n7770), .B(n7769), .S(n9022), .Z(n7771) );
  NAND2_X1 U9510 ( .A1(n4288), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8647) );
  OAI211_X1 U9511 ( .C1(n7772), .C2(n9862), .A(n7771), .B(n8647), .ZN(P1_U3262) );
  OAI21_X1 U9512 ( .B1(n10106), .B2(n7774), .A(n7773), .ZN(n7783) );
  INV_X1 U9513 ( .A(n7783), .ZN(n7776) );
  INV_X1 U9514 ( .A(n8602), .ZN(n8554) );
  AOI22_X1 U9515 ( .A1(n8554), .A2(n7784), .B1(n10117), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7775) );
  OAI21_X1 U9516 ( .B1(n7776), .B2(n10117), .A(n7775), .ZN(P2_U3417) );
  INV_X1 U9517 ( .A(n7777), .ZN(n7781) );
  OAI222_X1 U9518 ( .A1(n4288), .A2(n7779), .B1(n9565), .B2(n7781), .C1(n7778), 
        .C2(n9568), .ZN(P1_U3334) );
  OAI222_X1 U9519 ( .A1(P2_U3151), .A2(n7782), .B1(n8618), .B2(n7781), .C1(
        n7780), .C2(n7954), .ZN(P2_U3274) );
  NAND2_X1 U9520 ( .A1(n7783), .A2(n10130), .ZN(n7786) );
  INV_X1 U9521 ( .A(n8543), .ZN(n8481) );
  NAND2_X1 U9522 ( .A1(n7784), .A2(n8481), .ZN(n7785) );
  OAI211_X1 U9523 ( .C1(n10130), .C2(n8257), .A(n7786), .B(n7785), .ZN(
        P2_U3468) );
  XNOR2_X1 U9524 ( .A(n10100), .B(n8016), .ZN(n7792) );
  INV_X1 U9525 ( .A(n7787), .ZN(n7788) );
  XNOR2_X1 U9526 ( .A(n7844), .B(n7864), .ZN(n7791) );
  AOI21_X1 U9527 ( .B1(n7792), .B2(n7791), .A(n7848), .ZN(n7801) );
  INV_X1 U9528 ( .A(n7793), .ZN(n7794) );
  NAND2_X1 U9529 ( .A1(n8179), .A2(n7794), .ZN(n7797) );
  NAND2_X1 U9530 ( .A1(n8155), .A2(n8197), .ZN(n7796) );
  NAND2_X1 U9531 ( .A1(n8175), .A2(n8195), .ZN(n7795) );
  INV_X1 U9532 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9640) );
  OR2_X1 U9533 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9640), .ZN(n9947) );
  NAND4_X1 U9534 ( .A1(n7797), .A2(n7796), .A3(n7795), .A4(n9947), .ZN(n7798)
         );
  AOI21_X1 U9535 ( .B1(n7799), .B2(n8166), .A(n7798), .ZN(n7800) );
  OAI21_X1 U9536 ( .B1(n7801), .B2(n8162), .A(n7800), .ZN(P2_U3157) );
  OAI21_X1 U9537 ( .B1(n7804), .B2(n7803), .A(n7802), .ZN(n7805) );
  NAND2_X1 U9538 ( .A1(n7805), .A2(n8746), .ZN(n7812) );
  NAND2_X1 U9539 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(n4288), .ZN(n9762) );
  INV_X1 U9540 ( .A(n9762), .ZN(n7810) );
  INV_X1 U9541 ( .A(n7806), .ZN(n7808) );
  OAI22_X1 U9542 ( .A1(n8749), .A2(n7808), .B1(n7807), .B2(n8762), .ZN(n7809)
         );
  AOI211_X1 U9543 ( .C1(n8760), .C2(n9045), .A(n7810), .B(n7809), .ZN(n7811)
         );
  OAI211_X1 U9544 ( .C1(n7813), .C2(n8754), .A(n7812), .B(n7811), .ZN(P1_U3217) );
  XOR2_X1 U9545 ( .A(n7814), .B(n9002), .Z(n7889) );
  INV_X1 U9546 ( .A(n7815), .ZN(n7817) );
  OAI21_X1 U9547 ( .B1(n7817), .B2(n7816), .A(n9002), .ZN(n7819) );
  NAND2_X1 U9548 ( .A1(n7819), .A2(n7818), .ZN(n7883) );
  OAI211_X1 U9549 ( .C1(n8830), .C2(n7821), .A(n9331), .B(n7895), .ZN(n7881)
         );
  NAND2_X1 U9550 ( .A1(n9354), .A2(n9040), .ZN(n7823) );
  AOI22_X1 U9551 ( .A1(n9876), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8758), .B2(
        n9865), .ZN(n7822) );
  OAI211_X1 U9552 ( .C1(n8763), .C2(n9349), .A(n7823), .B(n7822), .ZN(n7824)
         );
  AOI21_X1 U9553 ( .B1(n8766), .B2(n9378), .A(n7824), .ZN(n7825) );
  OAI21_X1 U9554 ( .B1(n7881), .B2(n9381), .A(n7825), .ZN(n7826) );
  AOI21_X1 U9555 ( .B1(n7883), .B2(n9358), .A(n7826), .ZN(n7827) );
  OAI21_X1 U9556 ( .B1(n7889), .B2(n9385), .A(n7827), .ZN(P1_U3278) );
  INV_X1 U9557 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7833) );
  OAI22_X1 U9558 ( .A1(n8626), .A2(n9261), .B1(n8673), .B2(n9262), .ZN(n7828)
         );
  OR3_X1 U9559 ( .A1(n7830), .A2(n7829), .A3(n7828), .ZN(n7831) );
  AOI21_X1 U9560 ( .B1(n7832), .B2(n9905), .A(n7831), .ZN(n7835) );
  MUX2_X1 U9561 ( .A(n7833), .B(n7835), .S(n9914), .Z(n7834) );
  OAI21_X1 U9562 ( .B1(n8632), .B2(n9463), .A(n7834), .ZN(P1_U3536) );
  INV_X1 U9563 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7836) );
  MUX2_X1 U9564 ( .A(n7836), .B(n7835), .S(n9544), .Z(n7837) );
  OAI21_X1 U9565 ( .B1(n8632), .B2(n9534), .A(n7837), .ZN(P1_U3495) );
  INV_X1 U9566 ( .A(n7838), .ZN(n7842) );
  OAI222_X1 U9567 ( .A1(n9568), .A2(n7840), .B1(n9565), .B2(n7842), .C1(
        P1_U3086), .C2(n7839), .ZN(P1_U3333) );
  OAI222_X1 U9568 ( .A1(n7843), .A2(P2_U3151), .B1(n8618), .B2(n7842), .C1(
        n7841), .C2(n7954), .ZN(P2_U3273) );
  INV_X1 U9569 ( .A(n7868), .ZN(n10105) );
  INV_X1 U9570 ( .A(n7844), .ZN(n7845) );
  NOR2_X1 U9571 ( .A1(n7845), .A2(n8196), .ZN(n7847) );
  XNOR2_X1 U9572 ( .A(n7846), .B(n8004), .ZN(n7923) );
  INV_X1 U9573 ( .A(n7924), .ZN(n7850) );
  OAI21_X1 U9574 ( .B1(n7848), .B2(n7847), .A(n7923), .ZN(n7849) );
  NAND3_X1 U9575 ( .A1(n7850), .A2(n8169), .A3(n7849), .ZN(n7856) );
  INV_X1 U9576 ( .A(n7865), .ZN(n7854) );
  INV_X1 U9577 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7851) );
  NOR2_X1 U9578 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7851), .ZN(n9958) );
  AOI21_X1 U9579 ( .B1(n8175), .B2(n8194), .A(n9958), .ZN(n7852) );
  OAI21_X1 U9580 ( .B1(n7864), .B2(n8177), .A(n7852), .ZN(n7853) );
  AOI21_X1 U9581 ( .B1(n7854), .B2(n8179), .A(n7853), .ZN(n7855) );
  OAI211_X1 U9582 ( .C1(n10105), .C2(n8182), .A(n7856), .B(n7855), .ZN(
        P2_U3176) );
  XNOR2_X1 U9583 ( .A(n7857), .B(n7861), .ZN(n10107) );
  OR2_X1 U9584 ( .A1(n7719), .A2(n7858), .ZN(n7860) );
  NAND2_X1 U9585 ( .A1(n7860), .A2(n7859), .ZN(n7862) );
  XNOR2_X1 U9586 ( .A(n7862), .B(n7861), .ZN(n7863) );
  OAI222_X1 U9587 ( .A1(n8444), .A2(n7864), .B1(n8442), .B2(n7983), .C1(n7863), 
        .C2(n8440), .ZN(n10109) );
  NAND2_X1 U9588 ( .A1(n10109), .A2(n8474), .ZN(n7870) );
  OAI22_X1 U9589 ( .A1(n8474), .A2(n7866), .B1(n7865), .B2(n8462), .ZN(n7867)
         );
  AOI21_X1 U9590 ( .B1(n7868), .B2(n8393), .A(n7867), .ZN(n7869) );
  OAI211_X1 U9591 ( .C1(n8452), .C2(n10107), .A(n7870), .B(n7869), .ZN(
        P2_U3222) );
  XOR2_X1 U9592 ( .A(n7871), .B(n7872), .Z(n7879) );
  AOI22_X1 U9593 ( .A1(n8760), .A2(n9044), .B1(n8759), .B2(n7873), .ZN(n7874)
         );
  NAND2_X1 U9594 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9146) );
  OAI211_X1 U9595 ( .C1(n7875), .C2(n8762), .A(n7874), .B(n9146), .ZN(n7876)
         );
  AOI21_X1 U9596 ( .B1(n7877), .B2(n8765), .A(n7876), .ZN(n7878) );
  OAI21_X1 U9597 ( .B1(n7879), .B2(n8768), .A(n7878), .ZN(P1_U3236) );
  AOI22_X1 U9598 ( .A1(n9474), .A2(n9040), .B1(n9368), .B2(n9475), .ZN(n7880)
         );
  OAI211_X1 U9599 ( .C1(n8830), .C2(n9901), .A(n7881), .B(n7880), .ZN(n7882)
         );
  AOI21_X1 U9600 ( .B1(n7883), .B2(n9482), .A(n7882), .ZN(n7886) );
  NOR2_X1 U9601 ( .A1(n7886), .A2(n5572), .ZN(n7884) );
  AOI21_X1 U9602 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n5572), .A(n7884), .ZN(
        n7885) );
  OAI21_X1 U9603 ( .B1(n7889), .B2(n9491), .A(n7885), .ZN(P1_U3537) );
  NOR2_X1 U9604 ( .A1(n7886), .A2(n9906), .ZN(n7887) );
  AOI21_X1 U9605 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(n9906), .A(n7887), .ZN(
        n7888) );
  OAI21_X1 U9606 ( .B1(n7889), .B2(n9548), .A(n7888), .ZN(P1_U3498) );
  AOI21_X1 U9607 ( .B1(n9004), .B2(n7891), .A(n7890), .ZN(n7892) );
  INV_X1 U9608 ( .A(n7892), .ZN(n7911) );
  OAI21_X1 U9609 ( .B1(n7893), .B2(n9004), .A(n9362), .ZN(n7906) );
  INV_X1 U9610 ( .A(n8676), .ZN(n7903) );
  INV_X1 U9611 ( .A(n9372), .ZN(n7894) );
  AOI211_X1 U9612 ( .C1(n8676), .C2(n7895), .A(n9371), .B(n7894), .ZN(n7904)
         );
  NAND2_X1 U9613 ( .A1(n7904), .A2(n9863), .ZN(n7899) );
  AOI22_X1 U9614 ( .A1(n9876), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8672), .B2(
        n9865), .ZN(n7896) );
  OAI21_X1 U9615 ( .B1(n9349), .B2(n8737), .A(n7896), .ZN(n7897) );
  AOI21_X1 U9616 ( .B1(n9354), .B2(n9039), .A(n7897), .ZN(n7898) );
  OAI211_X1 U9617 ( .C1(n7903), .C2(n9869), .A(n7899), .B(n7898), .ZN(n7900)
         );
  AOI21_X1 U9618 ( .B1(n9358), .B2(n7906), .A(n7900), .ZN(n7901) );
  OAI21_X1 U9619 ( .B1(n7911), .B2(n9385), .A(n7901), .ZN(P1_U3277) );
  AOI22_X1 U9620 ( .A1(n9039), .A2(n9474), .B1(n9475), .B2(n9473), .ZN(n7902)
         );
  OAI21_X1 U9621 ( .B1(n7903), .B2(n9901), .A(n7902), .ZN(n7905) );
  AOI211_X1 U9622 ( .C1(n9482), .C2(n7906), .A(n7905), .B(n7904), .ZN(n7908)
         );
  MUX2_X1 U9623 ( .A(n9672), .B(n7908), .S(n9914), .Z(n7907) );
  OAI21_X1 U9624 ( .B1(n7911), .B2(n9491), .A(n7907), .ZN(P1_U3538) );
  INV_X1 U9625 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7909) );
  MUX2_X1 U9626 ( .A(n7909), .B(n7908), .S(n9544), .Z(n7910) );
  OAI21_X1 U9627 ( .B1(n7911), .B2(n9548), .A(n7910), .ZN(P1_U3501) );
  XNOR2_X1 U9628 ( .A(n7912), .B(n7918), .ZN(n7913) );
  OAI222_X1 U9629 ( .A1(n8444), .A2(n7914), .B1(n8442), .B2(n7986), .C1(n8440), 
        .C2(n7913), .ZN(n10112) );
  INV_X1 U9630 ( .A(n10112), .ZN(n7922) );
  INV_X1 U9631 ( .A(n7916), .ZN(n7917) );
  AOI21_X1 U9632 ( .B1(n7918), .B2(n7915), .A(n7917), .ZN(n10115) );
  NOR2_X1 U9633 ( .A1(n4603), .A2(n8449), .ZN(n7920) );
  INV_X1 U9634 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8236) );
  OAI22_X1 U9635 ( .A1(n8474), .A2(n8236), .B1(n7927), .B2(n8462), .ZN(n7919)
         );
  AOI211_X1 U9636 ( .C1(n10115), .C2(n8470), .A(n7920), .B(n7919), .ZN(n7921)
         );
  OAI21_X1 U9637 ( .B1(n7922), .B2(n6946), .A(n7921), .ZN(P2_U3221) );
  XNOR2_X1 U9638 ( .A(n7929), .B(n8016), .ZN(n7982) );
  XNOR2_X1 U9639 ( .A(n7982), .B(n7983), .ZN(n7984) );
  XNOR2_X1 U9640 ( .A(n7985), .B(n7984), .ZN(n7931) );
  NAND2_X1 U9641 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n9981) );
  OAI21_X1 U9642 ( .B1(n8158), .B2(n7986), .A(n9981), .ZN(n7925) );
  AOI21_X1 U9643 ( .B1(n8155), .B2(n8195), .A(n7925), .ZN(n7926) );
  OAI21_X1 U9644 ( .B1(n7927), .B2(n8130), .A(n7926), .ZN(n7928) );
  AOI21_X1 U9645 ( .B1(n7929), .B2(n8166), .A(n7928), .ZN(n7930) );
  OAI21_X1 U9646 ( .B1(n7931), .B2(n8162), .A(n7930), .ZN(P2_U3164) );
  XNOR2_X1 U9647 ( .A(n7932), .B(n7935), .ZN(n7933) );
  OAI222_X1 U9648 ( .A1(n8444), .A2(n7983), .B1(n8442), .B2(n8443), .C1(n7933), 
        .C2(n8440), .ZN(n8540) );
  OAI22_X1 U9649 ( .A1(n8603), .A2(n8464), .B1(n8131), .B2(n8462), .ZN(n7934)
         );
  OAI21_X1 U9650 ( .B1(n8540), .B2(n7934), .A(n8474), .ZN(n7938) );
  XOR2_X1 U9651 ( .A(n7936), .B(n7935), .Z(n8541) );
  AOI22_X1 U9652 ( .A1(n8541), .A2(n8470), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6946), .ZN(n7937) );
  NAND2_X1 U9653 ( .A1(n7938), .A2(n7937), .ZN(P2_U3220) );
  INV_X1 U9654 ( .A(n7950), .ZN(n7941) );
  NAND2_X1 U9655 ( .A1(n8615), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7939) );
  OAI211_X1 U9656 ( .C1(n7941), .C2(n8618), .A(n7940), .B(n7939), .ZN(P2_U3272) );
  XOR2_X1 U9657 ( .A(n7942), .B(n7943), .Z(n7949) );
  AOI22_X1 U9658 ( .A1(n8760), .A2(n9043), .B1(n8759), .B2(n7944), .ZN(n7945)
         );
  NAND2_X1 U9659 ( .A1(n4288), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9783) );
  OAI211_X1 U9660 ( .C1(n8626), .C2(n8762), .A(n7945), .B(n9783), .ZN(n7946)
         );
  AOI21_X1 U9661 ( .B1(n7947), .B2(n8765), .A(n7946), .ZN(n7948) );
  OAI21_X1 U9662 ( .B1(n7949), .B2(n8768), .A(n7948), .ZN(P1_U3224) );
  NAND2_X1 U9663 ( .A1(n7950), .A2(n9571), .ZN(n7951) );
  OAI211_X1 U9664 ( .C1(n7952), .C2(n9568), .A(n7951), .B(n9024), .ZN(P1_U3332) );
  INV_X1 U9665 ( .A(n7953), .ZN(n7956) );
  OAI222_X1 U9666 ( .A1(n6048), .A2(P2_U3151), .B1(n8618), .B2(n7956), .C1(
        n9639), .C2(n7954), .ZN(P2_U3271) );
  OAI222_X1 U9667 ( .A1(n7957), .A2(n4288), .B1(n9565), .B2(n7956), .C1(n7955), 
        .C2(n9568), .ZN(P1_U3331) );
  INV_X1 U9668 ( .A(n7958), .ZN(n7961) );
  AOI22_X1 U9669 ( .A1(n7959), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8615), .ZN(n7960) );
  OAI21_X1 U9670 ( .B1(n7961), .B2(n8618), .A(n7960), .ZN(P2_U3270) );
  OAI222_X1 U9671 ( .A1(n7962), .A2(P1_U3086), .B1(n9565), .B2(n7961), .C1(
        n9605), .C2(n9568), .ZN(P1_U3330) );
  INV_X1 U9672 ( .A(n7963), .ZN(n8611) );
  OAI222_X1 U9673 ( .A1(n9568), .A2(n7964), .B1(P1_U3086), .B2(n5509), .C1(
        n9565), .C2(n8611), .ZN(P1_U3327) );
  OAI222_X1 U9674 ( .A1(n9568), .A2(n7966), .B1(n9565), .B2(n7965), .C1(n4288), 
        .C2(n8887), .ZN(P1_U3336) );
  AOI22_X1 U9675 ( .A1(n8169), .A2(n7968), .B1(n7967), .B2(n8166), .ZN(n7970)
         );
  NAND2_X1 U9676 ( .A1(n8175), .A2(n8202), .ZN(n7969) );
  OAI211_X1 U9677 ( .C1(n7975), .C2(n6805), .A(n7970), .B(n7969), .ZN(P2_U3172) );
  XOR2_X1 U9678 ( .A(n7972), .B(n7971), .Z(n7979) );
  OAI22_X1 U9679 ( .A1(n7974), .A2(n8158), .B1(n8182), .B2(n7973), .ZN(n7977)
         );
  NOR2_X1 U9680 ( .A1(n7975), .A2(n7250), .ZN(n7976) );
  AOI211_X1 U9681 ( .C1(n8155), .C2(n8202), .A(n7977), .B(n7976), .ZN(n7978)
         );
  OAI21_X1 U9682 ( .B1(n8162), .B2(n7979), .A(n7978), .ZN(P2_U3177) );
  INV_X1 U9683 ( .A(n8879), .ZN(n9560) );
  AOI22_X1 U9684 ( .A1(n7980), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8615), .ZN(n7981) );
  OAI21_X1 U9685 ( .B1(n9560), .B2(n8618), .A(n7981), .ZN(P2_U3265) );
  XNOR2_X1 U9686 ( .A(n8133), .B(n8016), .ZN(n7987) );
  NAND2_X1 U9687 ( .A1(n7987), .A2(n7986), .ZN(n8122) );
  NOR2_X1 U9688 ( .A1(n7987), .A2(n7986), .ZN(n8124) );
  XNOR2_X1 U9689 ( .A(n8461), .B(n8016), .ZN(n7988) );
  XNOR2_X1 U9690 ( .A(n7988), .B(n8193), .ZN(n8048) );
  XNOR2_X1 U9691 ( .A(n8168), .B(n8016), .ZN(n7989) );
  XNOR2_X1 U9692 ( .A(n7989), .B(n8456), .ZN(n8171) );
  XNOR2_X1 U9693 ( .A(n8089), .B(n8016), .ZN(n7990) );
  XNOR2_X1 U9694 ( .A(n7990), .B(n8414), .ZN(n8091) );
  XNOR2_X1 U9695 ( .A(n8417), .B(n8016), .ZN(n7992) );
  XNOR2_X1 U9696 ( .A(n7992), .B(n8427), .ZN(n8099) );
  INV_X1 U9697 ( .A(n7992), .ZN(n7993) );
  NOR2_X1 U9698 ( .A1(n7993), .A2(n8192), .ZN(n8148) );
  XNOR2_X1 U9699 ( .A(n8145), .B(n8016), .ZN(n7994) );
  XNOR2_X1 U9700 ( .A(n7994), .B(n8413), .ZN(n8147) );
  NAND2_X1 U9701 ( .A1(n7994), .A2(n8386), .ZN(n7995) );
  XNOR2_X1 U9702 ( .A(n8394), .B(n8016), .ZN(n7996) );
  XOR2_X1 U9703 ( .A(n8404), .B(n7996), .Z(n8062) );
  XNOR2_X1 U9704 ( .A(n8508), .B(n8016), .ZN(n7998) );
  XNOR2_X1 U9705 ( .A(n7998), .B(n8387), .ZN(n8115) );
  INV_X1 U9706 ( .A(n7998), .ZN(n7999) );
  XNOR2_X1 U9707 ( .A(n8074), .B(n8016), .ZN(n8000) );
  XOR2_X1 U9708 ( .A(n8378), .B(n8000), .Z(n8069) );
  XNOR2_X1 U9709 ( .A(n8142), .B(n8016), .ZN(n8001) );
  NOR2_X1 U9710 ( .A1(n8001), .A2(n8367), .ZN(n8136) );
  XNOR2_X1 U9711 ( .A(n8059), .B(n8016), .ZN(n8002) );
  NAND2_X1 U9712 ( .A1(n8003), .A2(n8002), .ZN(n8105) );
  XNOR2_X1 U9713 ( .A(n8567), .B(n8004), .ZN(n8005) );
  INV_X1 U9714 ( .A(n8005), .ZN(n8006) );
  NAND2_X1 U9715 ( .A1(n8006), .A2(n8187), .ZN(n8007) );
  NAND2_X1 U9716 ( .A1(n8078), .A2(n8079), .ZN(n8011) );
  XNOR2_X1 U9717 ( .A(n8077), .B(n8016), .ZN(n8008) );
  INV_X1 U9718 ( .A(n8008), .ZN(n8009) );
  NAND2_X1 U9719 ( .A1(n8009), .A2(n8186), .ZN(n8010) );
  NAND2_X1 U9720 ( .A1(n8082), .A2(n8160), .ZN(n8012) );
  XNOR2_X1 U9721 ( .A(n8559), .B(n8016), .ZN(n8013) );
  XNOR2_X1 U9722 ( .A(n8013), .B(n8320), .ZN(n8159) );
  XNOR2_X1 U9723 ( .A(n8553), .B(n8016), .ZN(n8018) );
  XNOR2_X1 U9724 ( .A(n8018), .B(n8310), .ZN(n8039) );
  INV_X1 U9725 ( .A(n8039), .ZN(n8017) );
  NAND2_X1 U9726 ( .A1(n8040), .A2(n8019), .ZN(n8022) );
  XNOR2_X1 U9727 ( .A(n8020), .B(n8016), .ZN(n8021) );
  XNOR2_X1 U9728 ( .A(n8022), .B(n8021), .ZN(n8029) );
  NOR2_X1 U9729 ( .A1(n8023), .A2(n8158), .ZN(n8026) );
  AOI22_X1 U9730 ( .A1(n8288), .A2(n8179), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8024) );
  OAI21_X1 U9731 ( .B1(n8310), .B2(n8177), .A(n8024), .ZN(n8025) );
  AOI211_X1 U9732 ( .C1(n8027), .C2(n8166), .A(n8026), .B(n8025), .ZN(n8028)
         );
  OAI21_X1 U9733 ( .B1(n8029), .B2(n8162), .A(n8028), .ZN(P2_U3160) );
  NOR2_X1 U9734 ( .A1(n8031), .A2(n8462), .ZN(n8282) );
  AOI21_X1 U9735 ( .B1(n8447), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8282), .ZN(
        n8032) );
  OAI21_X1 U9736 ( .B1(n8033), .B2(n8449), .A(n8032), .ZN(n8034) );
  AOI21_X1 U9737 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8037) );
  OAI21_X1 U9738 ( .B1(n8030), .B2(n6946), .A(n8037), .ZN(P2_U3204) );
  INV_X1 U9739 ( .A(n8553), .ZN(n8047) );
  AOI21_X1 U9740 ( .B1(n8038), .B2(n8039), .A(n8162), .ZN(n8041) );
  NAND2_X1 U9741 ( .A1(n8041), .A2(n8040), .ZN(n8046) );
  INV_X1 U9742 ( .A(n8042), .ZN(n8304) );
  AOI22_X1 U9743 ( .A1(n8299), .A2(n8155), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8043) );
  OAI21_X1 U9744 ( .B1(n8304), .B2(n8130), .A(n8043), .ZN(n8044) );
  AOI21_X1 U9745 ( .B1(n8175), .B2(n8298), .A(n8044), .ZN(n8045) );
  OAI211_X1 U9746 ( .C1(n8047), .C2(n8182), .A(n8046), .B(n8045), .ZN(P2_U3154) );
  XOR2_X1 U9747 ( .A(n8049), .B(n8048), .Z(n8054) );
  AOI22_X1 U9748 ( .A1(n8175), .A2(n8456), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8051) );
  NAND2_X1 U9749 ( .A1(n8155), .A2(n8458), .ZN(n8050) );
  OAI211_X1 U9750 ( .C1(n8130), .C2(n8463), .A(n8051), .B(n8050), .ZN(n8052)
         );
  AOI21_X1 U9751 ( .B1(n8461), .B2(n8166), .A(n8052), .ZN(n8053) );
  OAI21_X1 U9752 ( .B1(n8054), .B2(n8162), .A(n8053), .ZN(P2_U3155) );
  AOI21_X1 U9753 ( .B1(n8188), .B2(n8055), .A(n4307), .ZN(n8061) );
  INV_X1 U9754 ( .A(n8367), .ZN(n8189) );
  AOI22_X1 U9755 ( .A1(n8189), .A2(n8155), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8057) );
  NAND2_X1 U9756 ( .A1(n8179), .A2(n8343), .ZN(n8056) );
  OAI211_X1 U9757 ( .C1(n8342), .C2(n8158), .A(n8057), .B(n8056), .ZN(n8058)
         );
  AOI21_X1 U9758 ( .B1(n8059), .B2(n8166), .A(n8058), .ZN(n8060) );
  OAI21_X1 U9759 ( .B1(n8061), .B2(n8162), .A(n8060), .ZN(P2_U3156) );
  XOR2_X1 U9760 ( .A(n8063), .B(n8062), .Z(n8068) );
  AOI22_X1 U9761 ( .A1(n8175), .A2(n8191), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8065) );
  NAND2_X1 U9762 ( .A1(n8179), .A2(n8390), .ZN(n8064) );
  OAI211_X1 U9763 ( .C1(n8386), .C2(n8177), .A(n8065), .B(n8064), .ZN(n8066)
         );
  AOI21_X1 U9764 ( .B1(n8394), .B2(n8166), .A(n8066), .ZN(n8067) );
  OAI21_X1 U9765 ( .B1(n8068), .B2(n8162), .A(n8067), .ZN(P2_U3159) );
  XOR2_X1 U9766 ( .A(n8070), .B(n8069), .Z(n8076) );
  AOI22_X1 U9767 ( .A1(n8189), .A2(n8175), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8072) );
  NAND2_X1 U9768 ( .A1(n8179), .A2(n8368), .ZN(n8071) );
  OAI211_X1 U9769 ( .C1(n8387), .C2(n8177), .A(n8072), .B(n8071), .ZN(n8073)
         );
  AOI21_X1 U9770 ( .B1(n8074), .B2(n8166), .A(n8073), .ZN(n8075) );
  OAI21_X1 U9771 ( .B1(n8076), .B2(n8162), .A(n8075), .ZN(P2_U3163) );
  INV_X1 U9772 ( .A(n8078), .ZN(n8108) );
  INV_X1 U9773 ( .A(n8079), .ZN(n8081) );
  NOR3_X1 U9774 ( .A1(n8108), .A2(n8081), .A3(n8080), .ZN(n8084) );
  INV_X1 U9775 ( .A(n8082), .ZN(n8083) );
  OAI21_X1 U9776 ( .B1(n8084), .B2(n8083), .A(n8169), .ZN(n8088) );
  AOI22_X1 U9777 ( .A1(n8187), .A2(n8155), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8085) );
  OAI21_X1 U9778 ( .B1(n8320), .B2(n8158), .A(n8085), .ZN(n8086) );
  AOI21_X1 U9779 ( .B1(n8322), .B2(n8179), .A(n8086), .ZN(n8087) );
  OAI211_X1 U9780 ( .C1(n8563), .C2(n8182), .A(n8088), .B(n8087), .ZN(P2_U3165) );
  OAI211_X1 U9781 ( .C1(n8092), .C2(n8091), .A(n8090), .B(n8169), .ZN(n8097)
         );
  INV_X1 U9782 ( .A(n8093), .ZN(n8431) );
  AND2_X1 U9783 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10042) );
  AOI21_X1 U9784 ( .B1(n8175), .B2(n8192), .A(n10042), .ZN(n8094) );
  OAI21_X1 U9785 ( .B1(n8430), .B2(n8177), .A(n8094), .ZN(n8095) );
  AOI21_X1 U9786 ( .B1(n8431), .B2(n8179), .A(n8095), .ZN(n8096) );
  OAI211_X1 U9787 ( .C1(n8593), .C2(n8182), .A(n8097), .B(n8096), .ZN(P2_U3166) );
  AOI21_X1 U9788 ( .B1(n8099), .B2(n8098), .A(n4365), .ZN(n8104) );
  AOI22_X1 U9789 ( .A1(n8175), .A2(n8413), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8101) );
  NAND2_X1 U9790 ( .A1(n8179), .A2(n8418), .ZN(n8100) );
  OAI211_X1 U9791 ( .C1(n8441), .C2(n8177), .A(n8101), .B(n8100), .ZN(n8102)
         );
  AOI21_X1 U9792 ( .B1(n8417), .B2(n8166), .A(n8102), .ZN(n8103) );
  OAI21_X1 U9793 ( .B1(n8104), .B2(n8162), .A(n8103), .ZN(P2_U3168) );
  INV_X1 U9794 ( .A(n8105), .ZN(n8107) );
  NOR3_X1 U9795 ( .A1(n4307), .A2(n8107), .A3(n8106), .ZN(n8109) );
  OAI21_X1 U9796 ( .B1(n8109), .B2(n8108), .A(n8169), .ZN(n8114) );
  OAI22_X1 U9797 ( .A1(n8354), .A2(n8177), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8110), .ZN(n8112) );
  NOR2_X1 U9798 ( .A1(n8329), .A2(n8158), .ZN(n8111) );
  AOI211_X1 U9799 ( .C1(n8331), .C2(n8179), .A(n8112), .B(n8111), .ZN(n8113)
         );
  OAI211_X1 U9800 ( .C1(n8567), .C2(n8182), .A(n8114), .B(n8113), .ZN(P2_U3169) );
  XOR2_X1 U9801 ( .A(n8116), .B(n8115), .Z(n8121) );
  INV_X1 U9802 ( .A(n8378), .ZN(n8190) );
  AOI22_X1 U9803 ( .A1(n8190), .A2(n8175), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8118) );
  NAND2_X1 U9804 ( .A1(n8179), .A2(n8379), .ZN(n8117) );
  OAI211_X1 U9805 ( .C1(n8404), .C2(n8177), .A(n8118), .B(n8117), .ZN(n8119)
         );
  AOI21_X1 U9806 ( .B1(n8508), .B2(n8166), .A(n8119), .ZN(n8120) );
  OAI21_X1 U9807 ( .B1(n8121), .B2(n8162), .A(n8120), .ZN(P2_U3173) );
  INV_X1 U9808 ( .A(n8122), .ZN(n8123) );
  NOR2_X1 U9809 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  XNOR2_X1 U9810 ( .A(n8126), .B(n8125), .ZN(n8135) );
  NAND2_X1 U9811 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9998) );
  INV_X1 U9812 ( .A(n9998), .ZN(n8128) );
  NOR2_X1 U9813 ( .A1(n8158), .A2(n8443), .ZN(n8127) );
  AOI211_X1 U9814 ( .C1(n8155), .C2(n8194), .A(n8128), .B(n8127), .ZN(n8129)
         );
  OAI21_X1 U9815 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8132) );
  AOI21_X1 U9816 ( .B1(n8133), .B2(n8166), .A(n8132), .ZN(n8134) );
  OAI21_X1 U9817 ( .B1(n8135), .B2(n8162), .A(n8134), .ZN(P2_U3174) );
  NOR2_X1 U9818 ( .A1(n8136), .A2(n4368), .ZN(n8137) );
  XNOR2_X1 U9819 ( .A(n8138), .B(n8137), .ZN(n8144) );
  AOI22_X1 U9820 ( .A1(n8190), .A2(n8155), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8140) );
  NAND2_X1 U9821 ( .A1(n8179), .A2(n8355), .ZN(n8139) );
  OAI211_X1 U9822 ( .C1(n8354), .C2(n8158), .A(n8140), .B(n8139), .ZN(n8141)
         );
  AOI21_X1 U9823 ( .B1(n8142), .B2(n8166), .A(n8141), .ZN(n8143) );
  OAI21_X1 U9824 ( .B1(n8144), .B2(n8162), .A(n8143), .ZN(P2_U3175) );
  INV_X1 U9825 ( .A(n8146), .ZN(n8150) );
  NOR3_X1 U9826 ( .A1(n4365), .A2(n8148), .A3(n8147), .ZN(n8149) );
  OAI21_X1 U9827 ( .B1(n8150), .B2(n8149), .A(n8169), .ZN(n8154) );
  NOR2_X1 U9828 ( .A1(n8177), .A2(n8427), .ZN(n8152) );
  INV_X1 U9829 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9611) );
  OAI22_X1 U9830 ( .A1(n8158), .A2(n8404), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9611), .ZN(n8151) );
  AOI211_X1 U9831 ( .C1(n8405), .C2(n8179), .A(n8152), .B(n8151), .ZN(n8153)
         );
  OAI211_X1 U9832 ( .C1(n8586), .C2(n8182), .A(n8154), .B(n8153), .ZN(P2_U3178) );
  AOI22_X1 U9833 ( .A1(n8186), .A2(n8155), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8157) );
  NAND2_X1 U9834 ( .A1(n8313), .A2(n8179), .ZN(n8156) );
  OAI211_X1 U9835 ( .C1(n8310), .C2(n8158), .A(n8157), .B(n8156), .ZN(n8165)
         );
  INV_X1 U9836 ( .A(n8159), .ZN(n8161) );
  NAND3_X1 U9837 ( .A1(n8082), .A2(n8161), .A3(n8160), .ZN(n8163) );
  OAI211_X1 U9838 ( .C1(n8172), .C2(n8171), .A(n8170), .B(n8169), .ZN(n8181)
         );
  INV_X1 U9839 ( .A(n8173), .ZN(n8445) );
  NAND2_X1 U9840 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10030) );
  INV_X1 U9841 ( .A(n10030), .ZN(n8174) );
  AOI21_X1 U9842 ( .B1(n8175), .B2(n8414), .A(n8174), .ZN(n8176) );
  OAI21_X1 U9843 ( .B1(n8443), .B2(n8177), .A(n8176), .ZN(n8178) );
  AOI21_X1 U9844 ( .B1(n8445), .B2(n8179), .A(n8178), .ZN(n8180) );
  OAI211_X1 U9845 ( .C1(n8597), .C2(n8182), .A(n8181), .B(n8180), .ZN(P2_U3181) );
  MUX2_X1 U9846 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8281), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9847 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8183), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9848 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8184), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9849 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8298), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8185), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9851 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8299), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9852 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8186), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9853 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8187), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9854 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8188), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9855 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8189), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9856 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8190), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8191), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9858 ( .A(n8413), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9736), .Z(
        P2_U3509) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8192), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8414), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8456), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9862 ( .A(n8193), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9736), .Z(
        P2_U3505) );
  MUX2_X1 U9863 ( .A(n8458), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9736), .Z(
        P2_U3504) );
  MUX2_X1 U9864 ( .A(n8194), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9736), .Z(
        P2_U3503) );
  MUX2_X1 U9865 ( .A(n8195), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9736), .Z(
        P2_U3502) );
  MUX2_X1 U9866 ( .A(n8196), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9736), .Z(
        P2_U3501) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8197), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9868 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8198), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9869 ( .A(n8199), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9736), .Z(
        P2_U3498) );
  MUX2_X1 U9870 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n4628), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8200), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n5683), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9873 ( .A(n8201), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9736), .Z(
        P2_U3494) );
  MUX2_X1 U9874 ( .A(n6359), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9736), .Z(
        P2_U3493) );
  MUX2_X1 U9875 ( .A(n8202), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9736), .Z(
        P2_U3492) );
  INV_X1 U9876 ( .A(n9738), .ZN(n9734) );
  MUX2_X1 U9877 ( .A(n8203), .B(n8526), .S(n8227), .Z(n8222) );
  INV_X1 U9878 ( .A(n8272), .ZN(n10051) );
  XNOR2_X1 U9879 ( .A(n8222), .B(n8272), .ZN(n10058) );
  MUX2_X1 U9880 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8227), .Z(n8204) );
  OR2_X1 U9881 ( .A1(n8204), .A2(n8252), .ZN(n8220) );
  XNOR2_X1 U9882 ( .A(n8204), .B(n10033), .ZN(n10039) );
  MUX2_X1 U9883 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8227), .Z(n8205) );
  OR2_X1 U9884 ( .A1(n8205), .A2(n8269), .ZN(n8219) );
  XNOR2_X1 U9885 ( .A(n8205), .B(n10018), .ZN(n10023) );
  MUX2_X1 U9886 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8227), .Z(n8206) );
  OR2_X1 U9887 ( .A1(n8206), .A2(n8253), .ZN(n8218) );
  XNOR2_X1 U9888 ( .A(n8206), .B(n10001), .ZN(n10007) );
  MUX2_X1 U9889 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8227), .Z(n8207) );
  OR2_X1 U9890 ( .A1(n8207), .A2(n8266), .ZN(n8217) );
  XNOR2_X1 U9891 ( .A(n8207), .B(n9984), .ZN(n9989) );
  INV_X1 U9892 ( .A(n8239), .ZN(n9966) );
  MUX2_X1 U9893 ( .A(n8236), .B(n8263), .S(n8227), .Z(n8208) );
  NAND2_X1 U9894 ( .A1(n9966), .A2(n8208), .ZN(n8216) );
  XNOR2_X1 U9895 ( .A(n8208), .B(n8239), .ZN(n9972) );
  MUX2_X1 U9896 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8227), .Z(n8209) );
  OR2_X1 U9897 ( .A1(n8209), .A2(n8261), .ZN(n8215) );
  XNOR2_X1 U9898 ( .A(n8209), .B(n9950), .ZN(n9955) );
  MUX2_X1 U9899 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8227), .Z(n8210) );
  OR2_X1 U9900 ( .A1(n8210), .A2(n9932), .ZN(n8214) );
  XOR2_X1 U9901 ( .A(n9932), .B(n8210), .Z(n9938) );
  OAI21_X1 U9902 ( .B1(n8213), .B2(n8212), .A(n8211), .ZN(n9939) );
  NAND2_X1 U9903 ( .A1(n9938), .A2(n9939), .ZN(n9937) );
  NAND2_X1 U9904 ( .A1(n8214), .A2(n9937), .ZN(n9954) );
  NAND2_X1 U9905 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  NAND2_X1 U9906 ( .A1(n8215), .A2(n9953), .ZN(n9971) );
  NAND2_X1 U9907 ( .A1(n9972), .A2(n9971), .ZN(n9970) );
  NAND2_X1 U9908 ( .A1(n8216), .A2(n9970), .ZN(n9988) );
  NAND2_X1 U9909 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  NAND2_X1 U9910 ( .A1(n8217), .A2(n9987), .ZN(n10006) );
  NAND2_X1 U9911 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  NAND2_X1 U9912 ( .A1(n8218), .A2(n10005), .ZN(n10022) );
  NAND2_X1 U9913 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  NAND2_X1 U9914 ( .A1(n8219), .A2(n10021), .ZN(n10038) );
  NAND2_X1 U9915 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U9916 ( .A1(n8220), .A2(n10037), .ZN(n10057) );
  NAND2_X1 U9917 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  INV_X1 U9918 ( .A(n10056), .ZN(n8221) );
  AOI21_X1 U9919 ( .B1(n8222), .B2(n10051), .A(n8221), .ZN(n8224) );
  MUX2_X1 U9920 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8227), .Z(n8223) );
  NAND2_X1 U9921 ( .A1(n8224), .A2(n8223), .ZN(n9732) );
  NOR2_X1 U9922 ( .A1(n8224), .A2(n8223), .ZN(n9731) );
  AOI21_X1 U9923 ( .B1(n9734), .B2(n9732), .A(n9731), .ZN(n8230) );
  INV_X1 U9924 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8225) );
  MUX2_X1 U9925 ( .A(n8225), .B(P2_REG2_REG_19__SCAN_IN), .S(n8226), .Z(n8251)
         );
  INV_X1 U9926 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8518) );
  XNOR2_X1 U9927 ( .A(n8226), .B(n8518), .ZN(n8274) );
  INV_X1 U9928 ( .A(n8274), .ZN(n8228) );
  MUX2_X1 U9929 ( .A(n8251), .B(n8228), .S(n8227), .Z(n8229) );
  XNOR2_X1 U9930 ( .A(n8230), .B(n8229), .ZN(n8279) );
  XNOR2_X1 U9931 ( .A(n9932), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U9932 ( .A1(n9950), .A2(n8234), .ZN(n8235) );
  XNOR2_X1 U9933 ( .A(n8234), .B(n9950), .ZN(n9960) );
  OR2_X1 U9934 ( .A1(n8239), .A2(n8236), .ZN(n8238) );
  NAND2_X1 U9935 ( .A1(n8239), .A2(n8236), .ZN(n8237) );
  AND2_X1 U9936 ( .A1(n8238), .A2(n8237), .ZN(n9978) );
  NAND2_X1 U9937 ( .A1(n8239), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8240) );
  INV_X1 U9938 ( .A(n8242), .ZN(n8241) );
  XNOR2_X1 U9939 ( .A(n10001), .B(n8473), .ZN(n10011) );
  NOR2_X1 U9940 ( .A1(n10018), .A2(n8244), .ZN(n8245) );
  NAND2_X1 U9941 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8252), .ZN(n8246) );
  OAI21_X1 U9942 ( .B1(n8252), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8246), .ZN(
        n10044) );
  INV_X1 U9943 ( .A(n8247), .ZN(n8248) );
  INV_X1 U9944 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8250) );
  NOR2_X1 U9945 ( .A1(n9738), .A2(n8250), .ZN(n8249) );
  AOI21_X1 U9946 ( .B1(n8250), .B2(n9738), .A(n8249), .ZN(n9744) );
  INV_X1 U9947 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U9948 ( .A(n9738), .B(n8522), .ZN(n9729) );
  AOI22_X1 U9949 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8252), .B1(n10033), .B2(
        n8530), .ZN(n10036) );
  AOI22_X1 U9950 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8253), .B1(n10001), .B2(
        n9680), .ZN(n10004) );
  NAND2_X1 U9951 ( .A1(n9932), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8259) );
  MUX2_X1 U9952 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8254), .S(n9932), .Z(n9935)
         );
  OAI22_X1 U9953 ( .A1(n8258), .A2(n8257), .B1(n8256), .B2(n8255), .ZN(n9936)
         );
  NAND2_X1 U9954 ( .A1(n9935), .A2(n9936), .ZN(n9934) );
  NAND2_X1 U9955 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  NOR2_X1 U9956 ( .A1(n9966), .A2(n8263), .ZN(n8264) );
  AOI21_X1 U9957 ( .B1(n9966), .B2(n8263), .A(n8264), .ZN(n9969) );
  NAND2_X1 U9958 ( .A1(n9968), .A2(n9969), .ZN(n9967) );
  OAI21_X1 U9959 ( .B1(n9966), .B2(n8263), .A(n9967), .ZN(n8265) );
  NAND2_X1 U9960 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  XOR2_X1 U9961 ( .A(n8266), .B(n8265), .Z(n9986) );
  NAND2_X1 U9962 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U9963 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  NAND2_X1 U9964 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U9965 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  NAND2_X1 U9966 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10055), .ZN(n10054) );
  NAND2_X1 U9967 ( .A1(n8273), .A2(n10054), .ZN(n9728) );
  AOI22_X1 U9968 ( .A1(n9729), .A2(n9728), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9738), .ZN(n8275) );
  XNOR2_X1 U9969 ( .A(n8275), .B(n8274), .ZN(n8276) );
  NAND2_X1 U9970 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8277) );
  NAND2_X1 U9971 ( .A1(n8447), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U9972 ( .A1(n8281), .A2(n8280), .ZN(n8545) );
  INV_X1 U9973 ( .A(n8545), .ZN(n8283) );
  OAI21_X1 U9974 ( .B1(n8283), .B2(n8282), .A(n8474), .ZN(n8285) );
  OAI211_X1 U9975 ( .C1(n8547), .C2(n8449), .A(n8284), .B(n8285), .ZN(P2_U3202) );
  NAND2_X1 U9976 ( .A1(n8447), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8286) );
  OAI211_X1 U9977 ( .C1(n8550), .C2(n8449), .A(n8286), .B(n8285), .ZN(P2_U3203) );
  INV_X1 U9978 ( .A(n8287), .ZN(n8294) );
  AOI22_X1 U9979 ( .A1(n8288), .A2(n8446), .B1(n8447), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8289) );
  OAI21_X1 U9980 ( .B1(n8290), .B2(n8449), .A(n8289), .ZN(n8291) );
  AOI21_X1 U9981 ( .B1(n8292), .B2(n8470), .A(n8291), .ZN(n8293) );
  OAI21_X1 U9982 ( .B1(n8294), .B2(n6946), .A(n8293), .ZN(P2_U3205) );
  XNOR2_X1 U9983 ( .A(n6540), .B(n8295), .ZN(n8479) );
  AOI21_X2 U9984 ( .B1(n8303), .B2(n8460), .A(n8302), .ZN(n8478) );
  OAI21_X1 U9985 ( .B1(n8304), .B2(n8462), .A(n8478), .ZN(n8305) );
  NAND2_X1 U9986 ( .A1(n8305), .A2(n8474), .ZN(n8307) );
  AOI22_X1 U9987 ( .A1(n8553), .A2(n8393), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n6946), .ZN(n8306) );
  OAI211_X1 U9988 ( .C1(n8479), .C2(n8452), .A(n8307), .B(n8306), .ZN(P2_U3206) );
  XNOR2_X1 U9989 ( .A(n8308), .B(n8311), .ZN(n8309) );
  OAI222_X1 U9990 ( .A1(n8442), .A2(n8310), .B1(n8444), .B2(n8329), .C1(n8440), 
        .C2(n8309), .ZN(n8483) );
  INV_X1 U9991 ( .A(n8483), .ZN(n8317) );
  XNOR2_X1 U9992 ( .A(n8312), .B(n8311), .ZN(n8484) );
  AOI22_X1 U9993 ( .A1(n8313), .A2(n8446), .B1(n8447), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8314) );
  OAI21_X1 U9994 ( .B1(n8559), .B2(n8449), .A(n8314), .ZN(n8315) );
  AOI21_X1 U9995 ( .B1(n8484), .B2(n8470), .A(n8315), .ZN(n8316) );
  OAI21_X1 U9996 ( .B1(n8317), .B2(n8447), .A(n8316), .ZN(P2_U3207) );
  NOR2_X1 U9997 ( .A1(n8563), .A2(n8464), .ZN(n8321) );
  XOR2_X1 U9998 ( .A(n8323), .B(n8318), .Z(n8319) );
  OAI222_X1 U9999 ( .A1(n8444), .A2(n8342), .B1(n8442), .B2(n8320), .C1(n8319), 
        .C2(n8440), .ZN(n8487) );
  AOI211_X1 U10000 ( .C1(n8446), .C2(n8322), .A(n8321), .B(n8487), .ZN(n8326)
         );
  XNOR2_X1 U10001 ( .A(n8324), .B(n8323), .ZN(n8488) );
  AOI22_X1 U10002 ( .A1(n8488), .A2(n8470), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n6946), .ZN(n8325) );
  OAI21_X1 U10003 ( .B1(n8326), .B2(n8447), .A(n8325), .ZN(P2_U3208) );
  NOR2_X1 U10004 ( .A1(n8567), .A2(n8464), .ZN(n8330) );
  XNOR2_X1 U10005 ( .A(n8327), .B(n8334), .ZN(n8328) );
  OAI222_X1 U10006 ( .A1(n8444), .A2(n8354), .B1(n8442), .B2(n8329), .C1(n8440), .C2(n8328), .ZN(n8491) );
  AOI211_X1 U10007 ( .C1(n8446), .C2(n8331), .A(n8330), .B(n8491), .ZN(n8337)
         );
  NAND2_X1 U10008 ( .A1(n8333), .A2(n8332), .ZN(n8335) );
  XNOR2_X1 U10009 ( .A(n8335), .B(n8334), .ZN(n8492) );
  AOI22_X1 U10010 ( .A1(n8492), .A2(n8470), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n6946), .ZN(n8336) );
  OAI21_X1 U10011 ( .B1(n8337), .B2(n8447), .A(n8336), .ZN(P2_U3209) );
  XNOR2_X1 U10012 ( .A(n8338), .B(n8340), .ZN(n8496) );
  INV_X1 U10013 ( .A(n8496), .ZN(n8347) );
  XNOR2_X1 U10014 ( .A(n8339), .B(n8340), .ZN(n8341) );
  OAI222_X1 U10015 ( .A1(n8442), .A2(n8342), .B1(n8444), .B2(n8367), .C1(n8440), .C2(n8341), .ZN(n8495) );
  AOI22_X1 U10016 ( .A1(n8343), .A2(n8446), .B1(n8447), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n8344) );
  OAI21_X1 U10017 ( .B1(n8571), .B2(n8449), .A(n8344), .ZN(n8345) );
  AOI21_X1 U10018 ( .B1(n8495), .B2(n8474), .A(n8345), .ZN(n8346) );
  OAI21_X1 U10019 ( .B1(n8347), .B2(n8452), .A(n8346), .ZN(P2_U3210) );
  XOR2_X1 U10020 ( .A(n8350), .B(n8348), .Z(n8500) );
  INV_X1 U10021 ( .A(n8500), .ZN(n8359) );
  AND3_X1 U10022 ( .A1(n8361), .A2(n8350), .A3(n8349), .ZN(n8351) );
  NOR2_X1 U10023 ( .A1(n8352), .A2(n8351), .ZN(n8353) );
  OAI222_X1 U10024 ( .A1(n8444), .A2(n8378), .B1(n8442), .B2(n8354), .C1(n8440), .C2(n8353), .ZN(n8499) );
  AOI22_X1 U10025 ( .A1(n8446), .A2(n8355), .B1(n8447), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8356) );
  OAI21_X1 U10026 ( .B1(n8575), .B2(n8449), .A(n8356), .ZN(n8357) );
  AOI21_X1 U10027 ( .B1(n8499), .B2(n8474), .A(n8357), .ZN(n8358) );
  OAI21_X1 U10028 ( .B1(n8359), .B2(n8452), .A(n8358), .ZN(P2_U3211) );
  XOR2_X1 U10029 ( .A(n8360), .B(n8362), .Z(n8504) );
  INV_X1 U10030 ( .A(n8504), .ZN(n8372) );
  INV_X1 U10031 ( .A(n8361), .ZN(n8365) );
  NOR3_X1 U10032 ( .A1(n8374), .A2(n8363), .A3(n8362), .ZN(n8364) );
  NOR2_X1 U10033 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  OAI222_X1 U10034 ( .A1(n8444), .A2(n8387), .B1(n8442), .B2(n8367), .C1(n8440), .C2(n8366), .ZN(n8503) );
  AOI22_X1 U10035 ( .A1(n8447), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8368), .B2(
        n8446), .ZN(n8369) );
  OAI21_X1 U10036 ( .B1(n8579), .B2(n8449), .A(n8369), .ZN(n8370) );
  AOI21_X1 U10037 ( .B1(n8503), .B2(n8474), .A(n8370), .ZN(n8371) );
  OAI21_X1 U10038 ( .B1(n8452), .B2(n8372), .A(n8371), .ZN(P2_U3212) );
  XNOR2_X1 U10039 ( .A(n8373), .B(n8376), .ZN(n8510) );
  AOI21_X1 U10040 ( .B1(n8376), .B2(n8375), .A(n8374), .ZN(n8377) );
  OAI222_X1 U10041 ( .A1(n8442), .A2(n8378), .B1(n8444), .B2(n8404), .C1(n8440), .C2(n8377), .ZN(n8507) );
  INV_X1 U10042 ( .A(n8508), .ZN(n8381) );
  AOI22_X1 U10043 ( .A1(n8447), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8446), .B2(
        n8379), .ZN(n8380) );
  OAI21_X1 U10044 ( .B1(n8381), .B2(n8449), .A(n8380), .ZN(n8382) );
  AOI21_X1 U10045 ( .B1(n8507), .B2(n8474), .A(n8382), .ZN(n8383) );
  OAI21_X1 U10046 ( .B1(n8510), .B2(n8452), .A(n8383), .ZN(P2_U3213) );
  INV_X1 U10047 ( .A(n8395), .ZN(n8385) );
  XNOR2_X1 U10048 ( .A(n8384), .B(n8385), .ZN(n8389) );
  OAI22_X1 U10049 ( .A1(n8387), .A2(n8442), .B1(n8386), .B2(n8444), .ZN(n8388)
         );
  AOI21_X1 U10050 ( .B1(n8389), .B2(n8460), .A(n8388), .ZN(n8517) );
  INV_X1 U10051 ( .A(n8390), .ZN(n8391) );
  OAI22_X1 U10052 ( .A1(n8474), .A2(n8225), .B1(n8391), .B2(n8462), .ZN(n8392)
         );
  AOI21_X1 U10053 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8399) );
  OR2_X1 U10054 ( .A1(n8396), .A2(n8395), .ZN(n8512) );
  NAND3_X1 U10055 ( .A1(n8512), .A2(n8470), .A3(n8511), .ZN(n8398) );
  OAI211_X1 U10056 ( .C1(n8517), .C2(n8447), .A(n8399), .B(n8398), .ZN(
        P2_U3214) );
  XOR2_X1 U10057 ( .A(n8400), .B(n8402), .Z(n8521) );
  INV_X1 U10058 ( .A(n8521), .ZN(n8409) );
  XOR2_X1 U10059 ( .A(n8402), .B(n8401), .Z(n8403) );
  OAI222_X1 U10060 ( .A1(n8444), .A2(n8427), .B1(n8442), .B2(n8404), .C1(n8403), .C2(n8440), .ZN(n8520) );
  AOI22_X1 U10061 ( .A1(n8447), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8446), .B2(
        n8405), .ZN(n8406) );
  OAI21_X1 U10062 ( .B1(n8586), .B2(n8449), .A(n8406), .ZN(n8407) );
  AOI21_X1 U10063 ( .B1(n8520), .B2(n8474), .A(n8407), .ZN(n8408) );
  OAI21_X1 U10064 ( .B1(n8452), .B2(n8409), .A(n8408), .ZN(P2_U3215) );
  OAI211_X1 U10065 ( .C1(n8412), .C2(n8411), .A(n8410), .B(n8460), .ZN(n8416)
         );
  AOI22_X1 U10066 ( .A1(n8414), .A2(n8457), .B1(n8455), .B2(n8413), .ZN(n8415)
         );
  NAND2_X1 U10067 ( .A1(n8416), .A2(n8415), .ZN(n8524) );
  INV_X1 U10068 ( .A(n8524), .ZN(n8422) );
  OAI21_X1 U10069 ( .B1(n4304), .B2(n4518), .A(n4662), .ZN(n8525) );
  INV_X1 U10070 ( .A(n8417), .ZN(n8590) );
  AOI22_X1 U10071 ( .A1(n8447), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8446), .B2(
        n8418), .ZN(n8419) );
  OAI21_X1 U10072 ( .B1(n8590), .B2(n8449), .A(n8419), .ZN(n8420) );
  AOI21_X1 U10073 ( .B1(n8525), .B2(n8470), .A(n8420), .ZN(n8421) );
  OAI21_X1 U10074 ( .B1(n8422), .B2(n8447), .A(n8421), .ZN(P2_U3216) );
  XNOR2_X1 U10075 ( .A(n8423), .B(n8425), .ZN(n8529) );
  INV_X1 U10076 ( .A(n8529), .ZN(n8435) );
  OAI211_X1 U10077 ( .C1(n8426), .C2(n8425), .A(n8424), .B(n8460), .ZN(n8429)
         );
  OR2_X1 U10078 ( .A1(n8427), .A2(n8442), .ZN(n8428) );
  OAI211_X1 U10079 ( .C1(n8430), .C2(n8444), .A(n8429), .B(n8428), .ZN(n8528)
         );
  AOI22_X1 U10080 ( .A1(n8447), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8446), .B2(
        n8431), .ZN(n8432) );
  OAI21_X1 U10081 ( .B1(n8593), .B2(n8449), .A(n8432), .ZN(n8433) );
  AOI21_X1 U10082 ( .B1(n8528), .B2(n8474), .A(n8433), .ZN(n8434) );
  OAI21_X1 U10083 ( .B1(n8435), .B2(n8452), .A(n8434), .ZN(P2_U3217) );
  XNOR2_X1 U10084 ( .A(n8436), .B(n8437), .ZN(n8533) );
  INV_X1 U10085 ( .A(n8533), .ZN(n8453) );
  XOR2_X1 U10086 ( .A(n8438), .B(n8437), .Z(n8439) );
  OAI222_X1 U10087 ( .A1(n8444), .A2(n8443), .B1(n8442), .B2(n8441), .C1(n8440), .C2(n8439), .ZN(n8532) );
  AOI22_X1 U10088 ( .A1(n8447), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8446), .B2(
        n8445), .ZN(n8448) );
  OAI21_X1 U10089 ( .B1(n8597), .B2(n8449), .A(n8448), .ZN(n8450) );
  AOI21_X1 U10090 ( .B1(n8532), .B2(n8474), .A(n8450), .ZN(n8451) );
  OAI21_X1 U10091 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(P2_U3218) );
  XOR2_X1 U10092 ( .A(n8454), .B(n8468), .Z(n8459) );
  AOI222_X1 U10093 ( .A1(n8460), .A2(n8459), .B1(n8458), .B2(n8457), .C1(n8456), .C2(n8455), .ZN(n8538) );
  INV_X1 U10094 ( .A(n8538), .ZN(n8466) );
  INV_X1 U10095 ( .A(n8461), .ZN(n8539) );
  OAI22_X1 U10096 ( .A1(n8539), .A2(n8464), .B1(n8463), .B2(n8462), .ZN(n8465)
         );
  OAI21_X1 U10097 ( .B1(n8466), .B2(n8465), .A(n8474), .ZN(n8472) );
  NAND2_X1 U10098 ( .A1(n8469), .A2(n8468), .ZN(n8536) );
  NAND3_X1 U10099 ( .A1(n8467), .A2(n8536), .A3(n8470), .ZN(n8471) );
  OAI211_X1 U10100 ( .C1(n8474), .C2(n8473), .A(n8472), .B(n8471), .ZN(
        P2_U3219) );
  NOR2_X1 U10101 ( .A1(n8545), .A2(n10128), .ZN(n8476) );
  AOI21_X1 U10102 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10128), .A(n8476), .ZN(
        n8475) );
  OAI21_X1 U10103 ( .B1(n8547), .B2(n8543), .A(n8475), .ZN(P2_U3490) );
  AOI21_X1 U10104 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10128), .A(n8476), .ZN(
        n8477) );
  OAI21_X1 U10105 ( .B1(n8550), .B2(n8543), .A(n8477), .ZN(P2_U3489) );
  OAI21_X1 U10106 ( .B1(n10106), .B2(n8479), .A(n8478), .ZN(n8551) );
  MUX2_X1 U10107 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8551), .S(n10130), .Z(
        n8480) );
  AOI21_X1 U10108 ( .B1(n8481), .B2(n8553), .A(n8480), .ZN(n8482) );
  INV_X1 U10109 ( .A(n8482), .ZN(P2_U3486) );
  INV_X1 U10110 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8485) );
  AOI21_X1 U10111 ( .B1(n10114), .B2(n8484), .A(n8483), .ZN(n8556) );
  MUX2_X1 U10112 ( .A(n8485), .B(n8556), .S(n10130), .Z(n8486) );
  OAI21_X1 U10113 ( .B1(n8559), .B2(n8543), .A(n8486), .ZN(P2_U3485) );
  INV_X1 U10114 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8489) );
  AOI21_X1 U10115 ( .B1(n10114), .B2(n8488), .A(n8487), .ZN(n8560) );
  MUX2_X1 U10116 ( .A(n8489), .B(n8560), .S(n10130), .Z(n8490) );
  OAI21_X1 U10117 ( .B1(n8563), .B2(n8543), .A(n8490), .ZN(P2_U3484) );
  INV_X1 U10118 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8493) );
  AOI21_X1 U10119 ( .B1(n8492), .B2(n10114), .A(n8491), .ZN(n8564) );
  MUX2_X1 U10120 ( .A(n8493), .B(n8564), .S(n10130), .Z(n8494) );
  OAI21_X1 U10121 ( .B1(n8567), .B2(n8543), .A(n8494), .ZN(P2_U3483) );
  INV_X1 U10122 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8497) );
  AOI21_X1 U10123 ( .B1(n10114), .B2(n8496), .A(n8495), .ZN(n8568) );
  MUX2_X1 U10124 ( .A(n8497), .B(n8568), .S(n10130), .Z(n8498) );
  OAI21_X1 U10125 ( .B1(n8571), .B2(n8543), .A(n8498), .ZN(P2_U3482) );
  INV_X1 U10126 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8501) );
  AOI21_X1 U10127 ( .B1(n10114), .B2(n8500), .A(n8499), .ZN(n8572) );
  MUX2_X1 U10128 ( .A(n8501), .B(n8572), .S(n10130), .Z(n8502) );
  OAI21_X1 U10129 ( .B1(n8575), .B2(n8543), .A(n8502), .ZN(P2_U3481) );
  INV_X1 U10130 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8505) );
  AOI21_X1 U10131 ( .B1(n8504), .B2(n10114), .A(n8503), .ZN(n8576) );
  MUX2_X1 U10132 ( .A(n8505), .B(n8576), .S(n10130), .Z(n8506) );
  OAI21_X1 U10133 ( .B1(n8579), .B2(n8543), .A(n8506), .ZN(P2_U3480) );
  AOI21_X1 U10134 ( .B1(n10095), .B2(n8508), .A(n8507), .ZN(n8509) );
  OAI21_X1 U10135 ( .B1(n10106), .B2(n8510), .A(n8509), .ZN(n8580) );
  MUX2_X1 U10136 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8580), .S(n10130), .Z(
        P2_U3479) );
  NAND3_X1 U10137 ( .A1(n8512), .A2(n8511), .A3(n10114), .ZN(n8513) );
  OAI21_X1 U10138 ( .B1(n8514), .B2(n10111), .A(n8513), .ZN(n8515) );
  INV_X1 U10139 ( .A(n8515), .ZN(n8516) );
  AND2_X1 U10140 ( .A1(n8517), .A2(n8516), .ZN(n8581) );
  MUX2_X1 U10141 ( .A(n8518), .B(n8581), .S(n10130), .Z(n8519) );
  INV_X1 U10142 ( .A(n8519), .ZN(P2_U3478) );
  AOI21_X1 U10143 ( .B1(n8521), .B2(n10114), .A(n8520), .ZN(n8583) );
  MUX2_X1 U10144 ( .A(n8522), .B(n8583), .S(n10130), .Z(n8523) );
  OAI21_X1 U10145 ( .B1(n8586), .B2(n8543), .A(n8523), .ZN(P2_U3477) );
  AOI21_X1 U10146 ( .B1(n10114), .B2(n8525), .A(n8524), .ZN(n8587) );
  MUX2_X1 U10147 ( .A(n8526), .B(n8587), .S(n10130), .Z(n8527) );
  OAI21_X1 U10148 ( .B1(n8590), .B2(n8543), .A(n8527), .ZN(P2_U3476) );
  AOI21_X1 U10149 ( .B1(n10114), .B2(n8529), .A(n8528), .ZN(n8591) );
  MUX2_X1 U10150 ( .A(n8530), .B(n8591), .S(n10130), .Z(n8531) );
  OAI21_X1 U10151 ( .B1(n8593), .B2(n8543), .A(n8531), .ZN(P2_U3475) );
  AOI21_X1 U10152 ( .B1(n10114), .B2(n8533), .A(n8532), .ZN(n8594) );
  MUX2_X1 U10153 ( .A(n8534), .B(n8594), .S(n10130), .Z(n8535) );
  OAI21_X1 U10154 ( .B1(n8597), .B2(n8543), .A(n8535), .ZN(P2_U3474) );
  NAND3_X1 U10155 ( .A1(n8467), .A2(n10114), .A3(n8536), .ZN(n8537) );
  OAI211_X1 U10156 ( .C1(n8539), .C2(n10111), .A(n8538), .B(n8537), .ZN(n8598)
         );
  MUX2_X1 U10157 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8598), .S(n10130), .Z(
        P2_U3473) );
  AOI21_X1 U10158 ( .B1(n8541), .B2(n10114), .A(n8540), .ZN(n8599) );
  MUX2_X1 U10159 ( .A(n5813), .B(n8599), .S(n10130), .Z(n8542) );
  OAI21_X1 U10160 ( .B1(n8603), .B2(n8543), .A(n8542), .ZN(P2_U3472) );
  MUX2_X1 U10161 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8544), .S(n10130), .Z(
        P2_U3459) );
  NOR2_X1 U10162 ( .A1(n8545), .A2(n10117), .ZN(n8548) );
  AOI21_X1 U10163 ( .B1(n10117), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8548), .ZN(
        n8546) );
  OAI21_X1 U10164 ( .B1(n8547), .B2(n8602), .A(n8546), .ZN(P2_U3458) );
  AOI21_X1 U10165 ( .B1(n10117), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8548), .ZN(
        n8549) );
  OAI21_X1 U10166 ( .B1(n8550), .B2(n8602), .A(n8549), .ZN(P2_U3457) );
  MUX2_X1 U10167 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8551), .S(n10116), .Z(
        n8552) );
  AOI21_X1 U10168 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(n8555) );
  INV_X1 U10169 ( .A(n8555), .ZN(P2_U3454) );
  MUX2_X1 U10170 ( .A(n8557), .B(n8556), .S(n10116), .Z(n8558) );
  OAI21_X1 U10171 ( .B1(n8559), .B2(n8602), .A(n8558), .ZN(P2_U3453) );
  MUX2_X1 U10172 ( .A(n8561), .B(n8560), .S(n10116), .Z(n8562) );
  OAI21_X1 U10173 ( .B1(n8563), .B2(n8602), .A(n8562), .ZN(P2_U3452) );
  MUX2_X1 U10174 ( .A(n8565), .B(n8564), .S(n10116), .Z(n8566) );
  OAI21_X1 U10175 ( .B1(n8567), .B2(n8602), .A(n8566), .ZN(P2_U3451) );
  INV_X1 U10176 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8569) );
  MUX2_X1 U10177 ( .A(n8569), .B(n8568), .S(n10116), .Z(n8570) );
  OAI21_X1 U10178 ( .B1(n8571), .B2(n8602), .A(n8570), .ZN(P2_U3450) );
  MUX2_X1 U10179 ( .A(n8573), .B(n8572), .S(n10116), .Z(n8574) );
  OAI21_X1 U10180 ( .B1(n8575), .B2(n8602), .A(n8574), .ZN(P2_U3449) );
  MUX2_X1 U10181 ( .A(n8577), .B(n8576), .S(n10116), .Z(n8578) );
  OAI21_X1 U10182 ( .B1(n8579), .B2(n8602), .A(n8578), .ZN(P2_U3448) );
  MUX2_X1 U10183 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8580), .S(n10116), .Z(
        P2_U3447) );
  INV_X1 U10184 ( .A(n8581), .ZN(n8582) );
  MUX2_X1 U10185 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8582), .S(n10116), .Z(
        P2_U3446) );
  INV_X1 U10186 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8584) );
  MUX2_X1 U10187 ( .A(n8584), .B(n8583), .S(n10116), .Z(n8585) );
  OAI21_X1 U10188 ( .B1(n8586), .B2(n8602), .A(n8585), .ZN(P2_U3444) );
  MUX2_X1 U10189 ( .A(n8588), .B(n8587), .S(n10116), .Z(n8589) );
  OAI21_X1 U10190 ( .B1(n8590), .B2(n8602), .A(n8589), .ZN(P2_U3441) );
  MUX2_X1 U10191 ( .A(n9713), .B(n8591), .S(n10116), .Z(n8592) );
  OAI21_X1 U10192 ( .B1(n8593), .B2(n8602), .A(n8592), .ZN(P2_U3438) );
  INV_X1 U10193 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8595) );
  MUX2_X1 U10194 ( .A(n8595), .B(n8594), .S(n10116), .Z(n8596) );
  OAI21_X1 U10195 ( .B1(n8597), .B2(n8602), .A(n8596), .ZN(P2_U3435) );
  MUX2_X1 U10196 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8598), .S(n10116), .Z(
        P2_U3432) );
  INV_X1 U10197 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U10198 ( .A(n8600), .B(n8599), .S(n10116), .Z(n8601) );
  OAI21_X1 U10199 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(P2_U3429) );
  INV_X1 U10200 ( .A(n8771), .ZN(n9558) );
  NOR4_X1 U10201 ( .A1(n8604), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5606), .ZN(n8605) );
  AOI21_X1 U10202 ( .B1(n8615), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8605), .ZN(
        n8606) );
  OAI21_X1 U10203 ( .B1(n9558), .B2(n8618), .A(n8606), .ZN(P2_U3264) );
  INV_X1 U10204 ( .A(n6342), .ZN(n9562) );
  AOI22_X1 U10205 ( .A1(n8607), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8615), .ZN(n8608) );
  OAI21_X1 U10206 ( .B1(n9562), .B2(n8618), .A(n8608), .ZN(P2_U3266) );
  AOI21_X1 U10207 ( .B1(n8615), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8609), .ZN(
        n8610) );
  OAI21_X1 U10208 ( .B1(n8611), .B2(n8618), .A(n8610), .ZN(P2_U3267) );
  INV_X1 U10209 ( .A(n8612), .ZN(n9564) );
  AOI21_X1 U10210 ( .B1(n8615), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8613), .ZN(
        n8614) );
  OAI21_X1 U10211 ( .B1(n9564), .B2(n8618), .A(n8614), .ZN(P2_U3268) );
  INV_X1 U10212 ( .A(n9572), .ZN(n8619) );
  AOI22_X1 U10213 ( .A1(n8616), .A2(P2_STATE_REG_SCAN_IN), .B1(n8615), .B2(
        P1_DATAO_REG_26__SCAN_IN), .ZN(n8617) );
  OAI21_X1 U10214 ( .B1(n8619), .B2(n8618), .A(n8617), .ZN(P2_U3269) );
  MUX2_X1 U10215 ( .A(n8620), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10216 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8624) );
  NAND2_X1 U10217 ( .A1(n8624), .A2(n8746), .ZN(n8631) );
  NAND2_X1 U10218 ( .A1(n4288), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9807) );
  INV_X1 U10219 ( .A(n9807), .ZN(n8629) );
  INV_X1 U10220 ( .A(n8625), .ZN(n8627) );
  OAI22_X1 U10221 ( .A1(n8749), .A2(n8627), .B1(n8626), .B2(n8736), .ZN(n8628)
         );
  AOI211_X1 U10222 ( .C1(n8751), .C2(n9039), .A(n8629), .B(n8628), .ZN(n8630)
         );
  OAI211_X1 U10223 ( .C1(n8632), .C2(n8754), .A(n8631), .B(n8630), .ZN(
        P1_U3215) );
  INV_X1 U10224 ( .A(n8692), .ZN(n8635) );
  AOI21_X1 U10225 ( .B1(n8725), .B2(n8722), .A(n8633), .ZN(n8634) );
  OAI21_X1 U10226 ( .B1(n8635), .B2(n8634), .A(n8746), .ZN(n8639) );
  OAI22_X1 U10227 ( .A1(n9278), .A2(n8762), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9682), .ZN(n8637) );
  OAI22_X1 U10228 ( .A1(n8749), .A2(n9274), .B1(n9308), .B2(n8736), .ZN(n8636)
         );
  AOI211_X1 U10229 ( .C1(n9280), .C2(n8765), .A(n8637), .B(n8636), .ZN(n8638)
         );
  NAND2_X1 U10230 ( .A1(n8639), .A2(n8638), .ZN(P1_U3216) );
  INV_X1 U10231 ( .A(n8640), .ZN(n8642) );
  XOR2_X1 U10232 ( .A(n8641), .B(n8640), .Z(n8735) );
  NOR2_X1 U10233 ( .A1(n8735), .A2(n8734), .ZN(n8733) );
  AOI21_X1 U10234 ( .B1(n8642), .B2(n8641), .A(n8733), .ZN(n8646) );
  XNOR2_X1 U10235 ( .A(n8644), .B(n8643), .ZN(n8645) );
  XNOR2_X1 U10236 ( .A(n8646), .B(n8645), .ZN(n8651) );
  OAI21_X1 U10237 ( .B1(n8762), .B2(n9336), .A(n8647), .ZN(n8649) );
  OAI22_X1 U10238 ( .A1(n8749), .A2(n9332), .B1(n8685), .B2(n8736), .ZN(n8648)
         );
  AOI211_X1 U10239 ( .C1(n9338), .C2(n8765), .A(n8649), .B(n8648), .ZN(n8650)
         );
  OAI21_X1 U10240 ( .B1(n8651), .B2(n8768), .A(n8650), .ZN(P1_U3219) );
  XOR2_X1 U10241 ( .A(n8653), .B(n8652), .Z(n8657) );
  OAI22_X1 U10242 ( .A1(n8736), .A2(n9336), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9685), .ZN(n8655) );
  OAI22_X1 U10243 ( .A1(n8749), .A2(n9304), .B1(n9308), .B2(n8762), .ZN(n8654)
         );
  AOI211_X1 U10244 ( .C1(n9310), .C2(n8765), .A(n8655), .B(n8654), .ZN(n8656)
         );
  OAI21_X1 U10245 ( .B1(n8657), .B2(n8768), .A(n8656), .ZN(P1_U3223) );
  AOI21_X1 U10246 ( .B1(n8659), .B2(n8658), .A(n8744), .ZN(n8664) );
  OAI22_X1 U10247 ( .A1(n9278), .A2(n8736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8660), .ZN(n8662) );
  OAI22_X1 U10248 ( .A1(n9244), .A2(n8762), .B1(n8749), .B2(n9241), .ZN(n8661)
         );
  AOI211_X1 U10249 ( .C1(n9246), .C2(n8765), .A(n8662), .B(n8661), .ZN(n8663)
         );
  OAI21_X1 U10250 ( .B1(n8664), .B2(n8768), .A(n8663), .ZN(P1_U3225) );
  XNOR2_X1 U10251 ( .A(n8665), .B(n8666), .ZN(n8757) );
  NOR2_X1 U10252 ( .A1(n8757), .A2(n8756), .ZN(n8755) );
  AOI21_X1 U10253 ( .B1(n8666), .B2(n8665), .A(n8755), .ZN(n8670) );
  XNOR2_X1 U10254 ( .A(n8668), .B(n8667), .ZN(n8669) );
  XNOR2_X1 U10255 ( .A(n8670), .B(n8669), .ZN(n8679) );
  NOR2_X1 U10256 ( .A1(n8671), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9826) );
  INV_X1 U10257 ( .A(n8672), .ZN(n8674) );
  OAI22_X1 U10258 ( .A1(n8749), .A2(n8674), .B1(n8673), .B2(n8736), .ZN(n8675)
         );
  AOI211_X1 U10259 ( .C1(n8751), .C2(n9473), .A(n9826), .B(n8675), .ZN(n8678)
         );
  NAND2_X1 U10260 ( .A1(n8676), .A2(n8765), .ZN(n8677) );
  OAI211_X1 U10261 ( .C1(n8679), .C2(n8768), .A(n8678), .B(n8677), .ZN(
        P1_U3226) );
  INV_X1 U10262 ( .A(n8680), .ZN(n8682) );
  NOR2_X1 U10263 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  XNOR2_X1 U10264 ( .A(n8684), .B(n8683), .ZN(n8689) );
  NAND2_X1 U10265 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9844) );
  OAI21_X1 U10266 ( .B1(n8762), .B2(n8685), .A(n9844), .ZN(n8687) );
  OAI22_X1 U10267 ( .A1(n8749), .A2(n9375), .B1(n8763), .B2(n8736), .ZN(n8686)
         );
  AOI211_X1 U10268 ( .C1(n9379), .C2(n8765), .A(n8687), .B(n8686), .ZN(n8688)
         );
  OAI21_X1 U10269 ( .B1(n8689), .B2(n8768), .A(n8688), .ZN(P1_U3228) );
  AND3_X1 U10270 ( .A1(n8692), .A2(n8691), .A3(n8690), .ZN(n8693) );
  OAI21_X1 U10271 ( .B1(n8694), .B2(n8693), .A(n8746), .ZN(n8698) );
  AOI22_X1 U10272 ( .A1(n9408), .A2(n8751), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8697) );
  AOI22_X1 U10273 ( .A1(n9441), .A2(n8760), .B1(n9254), .B2(n8759), .ZN(n8696)
         );
  NAND2_X1 U10274 ( .A1(n9426), .A2(n8765), .ZN(n8695) );
  NAND4_X1 U10275 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(
        P1_U3229) );
  XNOR2_X1 U10276 ( .A(n8701), .B(n8700), .ZN(n8702) );
  XNOR2_X1 U10277 ( .A(n8699), .B(n8702), .ZN(n8709) );
  AND2_X1 U10278 ( .A1(n9476), .A2(n9474), .ZN(n8703) );
  AOI21_X1 U10279 ( .B1(n9440), .B2(n9475), .A(n8703), .ZN(n9318) );
  OAI22_X1 U10280 ( .A1(n9318), .A2(n8705), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8704), .ZN(n8707) );
  NOR2_X1 U10281 ( .A1(n9535), .A2(n8754), .ZN(n8706) );
  AOI211_X1 U10282 ( .C1(n8759), .C2(n9322), .A(n8707), .B(n8706), .ZN(n8708)
         );
  OAI21_X1 U10283 ( .B1(n8709), .B2(n8768), .A(n8708), .ZN(P1_U3233) );
  XOR2_X1 U10284 ( .A(n8710), .B(n8711), .Z(n8718) );
  AOI22_X1 U10285 ( .A1(n8760), .A2(n9042), .B1(n8759), .B2(n8712), .ZN(n8713)
         );
  NAND2_X1 U10286 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9795) );
  OAI211_X1 U10287 ( .C1(n8714), .C2(n8762), .A(n8713), .B(n9795), .ZN(n8715)
         );
  AOI21_X1 U10288 ( .B1(n8716), .B2(n8765), .A(n8715), .ZN(n8717) );
  OAI21_X1 U10289 ( .B1(n8718), .B2(n8768), .A(n8717), .ZN(P1_U3234) );
  XNOR2_X1 U10290 ( .A(n4293), .B(n8719), .ZN(n8721) );
  INV_X1 U10291 ( .A(n8723), .ZN(n8720) );
  NAND2_X1 U10292 ( .A1(n8721), .A2(n8720), .ZN(n8726) );
  INV_X1 U10293 ( .A(n8722), .ZN(n8724) );
  AOI22_X1 U10294 ( .A1(n8726), .A2(n8725), .B1(n8724), .B2(n8723), .ZN(n8732)
         );
  OAI22_X1 U10295 ( .A1(n8736), .A2(n8728), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8727), .ZN(n8730) );
  OAI22_X1 U10296 ( .A1(n9291), .A2(n8762), .B1(n8749), .B2(n9287), .ZN(n8729)
         );
  AOI211_X1 U10297 ( .C1(n9286), .C2(n8765), .A(n8730), .B(n8729), .ZN(n8731)
         );
  OAI21_X1 U10298 ( .B1(n8732), .B2(n8768), .A(n8731), .ZN(P1_U3235) );
  AOI21_X1 U10299 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8741) );
  NAND2_X1 U10300 ( .A1(n4288), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9860) );
  OAI21_X1 U10301 ( .B1(n8762), .B2(n9348), .A(n9860), .ZN(n8739) );
  OAI22_X1 U10302 ( .A1(n8749), .A2(n9350), .B1(n8737), .B2(n8736), .ZN(n8738)
         );
  AOI211_X1 U10303 ( .C1(n9347), .C2(n8765), .A(n8739), .B(n8738), .ZN(n8740)
         );
  OAI21_X1 U10304 ( .B1(n8741), .B2(n8768), .A(n8740), .ZN(P1_U3238) );
  OAI21_X1 U10305 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8745) );
  NAND3_X1 U10306 ( .A1(n8747), .A2(n8746), .A3(n8745), .ZN(n8753) );
  AOI22_X1 U10307 ( .A1(n9408), .A2(n8760), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8748) );
  OAI21_X1 U10308 ( .B1(n9224), .B2(n8749), .A(n8748), .ZN(n8750) );
  AOI21_X1 U10309 ( .B1(n8751), .B2(n9409), .A(n8750), .ZN(n8752) );
  OAI211_X1 U10310 ( .C1(n9412), .C2(n8754), .A(n8753), .B(n8752), .ZN(
        P1_U3240) );
  AOI21_X1 U10311 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8769) );
  AOI22_X1 U10312 ( .A1(n8760), .A2(n9040), .B1(n8759), .B2(n8758), .ZN(n8761)
         );
  NAND2_X1 U10313 ( .A1(n4288), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9819) );
  OAI211_X1 U10314 ( .C1(n8763), .C2(n8762), .A(n8761), .B(n9819), .ZN(n8764)
         );
  AOI21_X1 U10315 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n8767) );
  OAI21_X1 U10316 ( .B1(n8769), .B2(n8768), .A(n8767), .ZN(P1_U3241) );
  MUX2_X1 U10317 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8771), .S(n8770), .Z(
        n8773) );
  NAND2_X1 U10318 ( .A1(n8888), .A2(n8774), .ZN(n8895) );
  NAND2_X1 U10319 ( .A1(n8861), .A2(n8775), .ZN(n8889) );
  MUX2_X1 U10320 ( .A(n8895), .B(n8889), .S(n9025), .Z(n8864) );
  INV_X1 U10321 ( .A(n8913), .ZN(n8783) );
  INV_X1 U10322 ( .A(n8985), .ZN(n8778) );
  NAND2_X1 U10323 ( .A1(n8779), .A2(n8914), .ZN(n8782) );
  AND2_X1 U10324 ( .A1(n8920), .A2(n8785), .ZN(n8781) );
  AOI21_X1 U10325 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8793) );
  NOR2_X1 U10326 ( .A1(n8985), .A2(n8783), .ZN(n8786) );
  NAND2_X1 U10327 ( .A1(n8785), .A2(n8784), .ZN(n8918) );
  AOI21_X1 U10328 ( .B1(n8787), .B2(n8786), .A(n8918), .ZN(n8790) );
  NAND2_X1 U10329 ( .A1(n8788), .A2(n8917), .ZN(n8789) );
  OAI21_X1 U10330 ( .B1(n8790), .B2(n8789), .A(n8920), .ZN(n8791) );
  INV_X1 U10331 ( .A(n8791), .ZN(n8792) );
  MUX2_X1 U10332 ( .A(n8793), .B(n8792), .S(n4486), .Z(n8799) );
  AND2_X1 U10333 ( .A1(n8795), .A2(n8794), .ZN(n8796) );
  MUX2_X1 U10334 ( .A(n8796), .B(n8989), .S(n4486), .Z(n8797) );
  OAI21_X1 U10335 ( .B1(n8799), .B2(n8798), .A(n8797), .ZN(n8805) );
  NAND2_X1 U10336 ( .A1(n8991), .A2(n8800), .ZN(n8802) );
  MUX2_X1 U10337 ( .A(n8802), .B(n8801), .S(n4486), .Z(n8803) );
  INV_X1 U10338 ( .A(n8803), .ZN(n8804) );
  NAND2_X1 U10339 ( .A1(n8805), .A2(n8804), .ZN(n8811) );
  NAND2_X1 U10340 ( .A1(n8817), .A2(n8812), .ZN(n8807) );
  INV_X1 U10341 ( .A(n8991), .ZN(n8806) );
  NOR2_X1 U10342 ( .A1(n8807), .A2(n8806), .ZN(n8923) );
  OAI211_X1 U10343 ( .C1(n8807), .C2(n8814), .A(n8819), .B(n8815), .ZN(n8930)
         );
  AOI21_X1 U10344 ( .B1(n8811), .B2(n8923), .A(n8930), .ZN(n8809) );
  INV_X1 U10345 ( .A(n8928), .ZN(n8808) );
  OR2_X1 U10346 ( .A1(n8809), .A2(n8808), .ZN(n8822) );
  NAND2_X1 U10347 ( .A1(n8811), .A2(n8810), .ZN(n8813) );
  NAND2_X1 U10348 ( .A1(n8813), .A2(n8812), .ZN(n8816) );
  NAND3_X1 U10349 ( .A1(n8816), .A2(n8815), .A3(n8814), .ZN(n8818) );
  NAND3_X1 U10350 ( .A1(n8818), .A2(n8928), .A3(n8817), .ZN(n8820) );
  NAND2_X1 U10351 ( .A1(n8820), .A2(n8819), .ZN(n8821) );
  INV_X1 U10352 ( .A(n8929), .ZN(n8823) );
  NOR2_X1 U10353 ( .A1(n9000), .A2(n8823), .ZN(n8826) );
  AND2_X1 U10354 ( .A1(n8831), .A2(n8824), .ZN(n8906) );
  NAND2_X1 U10355 ( .A1(n8906), .A2(n8835), .ZN(n8825) );
  AND2_X1 U10356 ( .A1(n9361), .A2(n8827), .ZN(n8829) );
  AND2_X1 U10357 ( .A1(n8829), .A2(n8828), .ZN(n8833) );
  INV_X1 U10358 ( .A(n8829), .ZN(n8832) );
  AOI22_X1 U10359 ( .A1(n8832), .A2(n8831), .B1(n9025), .B2(n8830), .ZN(n8838)
         );
  AOI21_X1 U10360 ( .B1(n9361), .B2(n9039), .A(n4486), .ZN(n8837) );
  INV_X1 U10361 ( .A(n8833), .ZN(n8932) );
  NAND2_X1 U10362 ( .A1(n8835), .A2(n8834), .ZN(n8907) );
  NAND2_X1 U10363 ( .A1(n8907), .A2(n9025), .ZN(n8836) );
  OAI22_X1 U10364 ( .A1(n8838), .A2(n8837), .B1(n8932), .B2(n8836), .ZN(n8839)
         );
  OAI21_X1 U10365 ( .B1(n8840), .B2(n8839), .A(n9363), .ZN(n8847) );
  AND2_X1 U10366 ( .A1(n8848), .A2(n8841), .ZN(n8935) );
  NAND2_X1 U10367 ( .A1(n8950), .A2(n8846), .ZN(n8842) );
  AOI21_X1 U10368 ( .B1(n8847), .B2(n8935), .A(n8842), .ZN(n8844) );
  NAND2_X1 U10369 ( .A1(n8855), .A2(n8950), .ZN(n8843) );
  AND2_X1 U10370 ( .A1(n8846), .A2(n8845), .ZN(n8939) );
  NAND2_X1 U10371 ( .A1(n8847), .A2(n8939), .ZN(n8850) );
  NAND2_X1 U10372 ( .A1(n8851), .A2(n8848), .ZN(n8940) );
  NOR2_X1 U10373 ( .A1(n8940), .A2(n9025), .ZN(n8849) );
  NAND2_X1 U10374 ( .A1(n8850), .A2(n8849), .ZN(n8854) );
  NAND2_X1 U10375 ( .A1(n9299), .A2(n8851), .ZN(n8852) );
  NAND2_X1 U10376 ( .A1(n8852), .A2(n9025), .ZN(n8853) );
  NAND2_X1 U10377 ( .A1(n8854), .A2(n8853), .ZN(n8858) );
  NAND2_X1 U10378 ( .A1(n8896), .A2(n9299), .ZN(n8945) );
  NAND2_X1 U10379 ( .A1(n8859), .A2(n8855), .ZN(n8897) );
  MUX2_X1 U10380 ( .A(n8945), .B(n8897), .S(n9025), .Z(n8856) );
  INV_X1 U10381 ( .A(n8856), .ZN(n8857) );
  MUX2_X1 U10382 ( .A(n8859), .B(n8896), .S(n9025), .Z(n8860) );
  INV_X1 U10383 ( .A(n9260), .ZN(n9250) );
  MUX2_X1 U10384 ( .A(n8861), .B(n8888), .S(n9025), .Z(n8862) );
  OAI211_X1 U10385 ( .C1(n8864), .C2(n8863), .A(n9250), .B(n8862), .ZN(n8866)
         );
  MUX2_X1 U10386 ( .A(n8900), .B(n8891), .S(n9025), .Z(n8865) );
  OAI21_X1 U10387 ( .B1(n8867), .B2(n8901), .A(n8960), .ZN(n8868) );
  NAND2_X1 U10388 ( .A1(n8870), .A2(n8869), .ZN(n8904) );
  OAI21_X1 U10389 ( .B1(n4356), .B2(n8904), .A(n8953), .ZN(n8875) );
  INV_X1 U10390 ( .A(n8904), .ZN(n8873) );
  AOI21_X1 U10391 ( .B1(n8953), .B2(n8965), .A(n8871), .ZN(n8872) );
  AOI21_X1 U10392 ( .B1(n4357), .B2(n8873), .A(n8872), .ZN(n8874) );
  NAND2_X1 U10393 ( .A1(n9196), .A2(n4486), .ZN(n8877) );
  MUX2_X1 U10394 ( .A(n4486), .B(n9196), .S(n9178), .Z(n8876) );
  NAND2_X1 U10395 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  OR2_X1 U10396 ( .A1(n5155), .A2(n9561), .ZN(n8880) );
  MUX2_X1 U10397 ( .A(n8883), .B(n4486), .S(n9170), .Z(n8882) );
  NOR2_X1 U10398 ( .A1(n9160), .A2(n9163), .ZN(n8975) );
  INV_X1 U10399 ( .A(n9038), .ZN(n8957) );
  NOR2_X1 U10400 ( .A1(n8957), .A2(n9163), .ZN(n8968) );
  AOI21_X1 U10401 ( .B1(n9025), .B2(n9016), .A(n9021), .ZN(n9037) );
  INV_X1 U10402 ( .A(n8975), .ZN(n8972) );
  INV_X1 U10403 ( .A(n8885), .ZN(n9026) );
  NOR2_X1 U10404 ( .A1(n9024), .A2(n8886), .ZN(n9030) );
  OAI211_X1 U10405 ( .C1(n8972), .C2(n8887), .A(n9026), .B(n9030), .ZN(n9036)
         );
  NAND2_X1 U10406 ( .A1(n8889), .A2(n8888), .ZN(n8890) );
  NAND2_X1 U10407 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  NAND2_X1 U10408 ( .A1(n8892), .A2(n8900), .ZN(n8893) );
  NAND2_X1 U10409 ( .A1(n8894), .A2(n8893), .ZN(n8944) );
  INV_X1 U10410 ( .A(n8895), .ZN(n8899) );
  NAND2_X1 U10411 ( .A1(n8897), .A2(n8896), .ZN(n8898) );
  AND3_X1 U10412 ( .A1(n8900), .A2(n8899), .A3(n8898), .ZN(n8902) );
  OAI21_X1 U10413 ( .B1(n8944), .B2(n8902), .A(n8901), .ZN(n8903) );
  AND2_X1 U10414 ( .A1(n8903), .A2(n8948), .ZN(n8905) );
  AOI21_X1 U10415 ( .B1(n8905), .B2(n8965), .A(n8904), .ZN(n8962) );
  INV_X1 U10416 ( .A(n8906), .ZN(n8938) );
  INV_X1 U10417 ( .A(n8907), .ZN(n8934) );
  INV_X1 U10418 ( .A(n8993), .ZN(n8927) );
  INV_X1 U10419 ( .A(n8908), .ZN(n8911) );
  NAND2_X1 U10420 ( .A1(n9053), .A2(n8909), .ZN(n8910) );
  AND4_X1 U10421 ( .A1(n8912), .A2(n8911), .A3(n8978), .A4(n8910), .ZN(n8915)
         );
  OAI211_X1 U10422 ( .C1(n8916), .C2(n8915), .A(n8914), .B(n8913), .ZN(n8921)
         );
  NAND2_X1 U10423 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  NAND3_X1 U10424 ( .A1(n8921), .A2(n8920), .A3(n8919), .ZN(n8926) );
  INV_X1 U10425 ( .A(n8922), .ZN(n8925) );
  INV_X1 U10426 ( .A(n8923), .ZN(n8924) );
  AOI211_X1 U10427 ( .C1(n8927), .C2(n8926), .A(n8925), .B(n8924), .ZN(n8931)
         );
  OAI211_X1 U10428 ( .C1(n8931), .C2(n8930), .A(n8929), .B(n8928), .ZN(n8933)
         );
  AOI21_X1 U10429 ( .B1(n8934), .B2(n8933), .A(n8932), .ZN(n8937) );
  INV_X1 U10430 ( .A(n8935), .ZN(n8936) );
  AOI211_X1 U10431 ( .C1(n9361), .C2(n8938), .A(n8937), .B(n8936), .ZN(n8943)
         );
  INV_X1 U10432 ( .A(n8939), .ZN(n8942) );
  INV_X1 U10433 ( .A(n8940), .ZN(n8941) );
  OAI21_X1 U10434 ( .B1(n8943), .B2(n8942), .A(n8941), .ZN(n8949) );
  INV_X1 U10435 ( .A(n8944), .ZN(n8947) );
  INV_X1 U10436 ( .A(n8945), .ZN(n8946) );
  NAND3_X1 U10437 ( .A1(n8948), .A2(n8947), .A3(n8946), .ZN(n8961) );
  AOI21_X1 U10438 ( .B1(n8950), .B2(n8949), .A(n8961), .ZN(n8952) );
  OAI21_X1 U10439 ( .B1(n8952), .B2(n8951), .A(n8965), .ZN(n8955) );
  NAND2_X1 U10440 ( .A1(n8954), .A2(n8953), .ZN(n8967) );
  AOI21_X1 U10441 ( .B1(n8962), .B2(n8955), .A(n8967), .ZN(n8958) );
  NAND2_X1 U10442 ( .A1(n9170), .A2(n8957), .ZN(n8976) );
  NAND2_X1 U10443 ( .A1(n8976), .A2(n8956), .ZN(n8970) );
  OAI21_X1 U10444 ( .B1(n8958), .B2(n8970), .A(n8977), .ZN(n8959) );
  AOI21_X1 U10445 ( .B1(n8972), .B2(n8959), .A(n9016), .ZN(n9029) );
  INV_X1 U10446 ( .A(n9170), .ZN(n9500) );
  OAI21_X1 U10447 ( .B1(n8961), .B2(n9317), .A(n8960), .ZN(n8964) );
  INV_X1 U10448 ( .A(n8962), .ZN(n8963) );
  AOI21_X1 U10449 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(n8966) );
  NOR2_X1 U10450 ( .A1(n8967), .A2(n8966), .ZN(n8971) );
  INV_X1 U10451 ( .A(n8968), .ZN(n8969) );
  OAI22_X1 U10452 ( .A1(n8971), .A2(n8970), .B1(n9170), .B2(n8969), .ZN(n8973)
         );
  OAI211_X1 U10453 ( .C1(n9500), .C2(n8974), .A(n8973), .B(n8972), .ZN(n9012)
         );
  INV_X1 U10454 ( .A(n9271), .ZN(n9269) );
  NOR2_X1 U10455 ( .A1(n8979), .A2(n8978), .ZN(n8984) );
  INV_X1 U10456 ( .A(n8980), .ZN(n8982) );
  NAND4_X1 U10457 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n8988)
         );
  NOR4_X1 U10458 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n8990)
         );
  NAND3_X1 U10459 ( .A1(n8991), .A2(n8990), .A3(n8989), .ZN(n8992) );
  NOR3_X1 U10460 ( .A1(n8994), .A2(n8993), .A3(n8992), .ZN(n8995) );
  NAND3_X1 U10461 ( .A1(n8997), .A2(n8996), .A3(n8995), .ZN(n8999) );
  OR3_X1 U10462 ( .A1(n9000), .A2(n8999), .A3(n8998), .ZN(n9001) );
  NOR2_X1 U10463 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  AND4_X1 U10464 ( .A1(n9344), .A2(n9363), .A3(n9004), .A4(n9003), .ZN(n9005)
         );
  AND4_X1 U10465 ( .A1(n9301), .A2(n9316), .A3(n9329), .A4(n9005), .ZN(n9006)
         );
  NAND4_X1 U10466 ( .A1(n9250), .A2(n9269), .A3(n9294), .A4(n9006), .ZN(n9007)
         );
  NOR2_X1 U10467 ( .A1(n9007), .A2(n9235), .ZN(n9008) );
  NAND4_X1 U10468 ( .A1(n8972), .A2(n4900), .A3(n9010), .A4(n4902), .ZN(n9017)
         );
  INV_X1 U10469 ( .A(n9017), .ZN(n9011) );
  AOI21_X1 U10470 ( .B1(n9013), .B2(n9012), .A(n9011), .ZN(n9015) );
  OAI21_X1 U10471 ( .B1(n9015), .B2(n9016), .A(n9014), .ZN(n9023) );
  NOR2_X1 U10472 ( .A1(n9017), .A2(n9016), .ZN(n9019) );
  MUX2_X1 U10473 ( .A(n9019), .B(n9029), .S(n9018), .Z(n9020) );
  AOI21_X1 U10474 ( .B1(n9026), .B2(n9025), .A(n9024), .ZN(n9027) );
  INV_X1 U10475 ( .A(n9030), .ZN(n9031) );
  OAI211_X1 U10476 ( .C1(n9033), .C2(n9032), .A(P1_B_REG_SCAN_IN), .B(n9031), 
        .ZN(n9034) );
  OAI211_X1 U10477 ( .C1(n9037), .C2(n9036), .A(n9035), .B(n9034), .ZN(
        P1_U3242) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9038), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9392), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9400), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9409), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9417), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9408), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9432), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9441), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9449), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9440), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9465), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10489 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9476), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9464), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10491 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9473), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9368), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9039), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9040), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10495 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9041), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9042), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9043), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9044), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9045), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9046), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9047), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9048), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9049), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9050), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9051), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9052), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9053), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10508 ( .C1(n9056), .C2(n9055), .A(n9842), .B(n9054), .ZN(n9064)
         );
  OAI211_X1 U10509 ( .C1(n9059), .C2(n9058), .A(n9850), .B(n9057), .ZN(n9063)
         );
  AOI22_X1 U10510 ( .A1(n9827), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n4288), .ZN(n9062) );
  NAND2_X1 U10511 ( .A1(n9839), .A2(n9060), .ZN(n9061) );
  NAND4_X1 U10512 ( .A1(n9064), .A2(n9063), .A3(n9062), .A4(n9061), .ZN(
        P1_U3244) );
  INV_X1 U10513 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9067) );
  INV_X1 U10514 ( .A(n9065), .ZN(n9066) );
  OAI21_X1 U10515 ( .B1(n9862), .B2(n9067), .A(n9066), .ZN(n9068) );
  AOI21_X1 U10516 ( .B1(n9069), .B2(n9839), .A(n9068), .ZN(n9078) );
  OAI211_X1 U10517 ( .C1(n9072), .C2(n9071), .A(n9842), .B(n9070), .ZN(n9077)
         );
  OAI211_X1 U10518 ( .C1(n9075), .C2(n9074), .A(n9850), .B(n9073), .ZN(n9076)
         );
  NAND3_X1 U10519 ( .A1(n9078), .A2(n9077), .A3(n9076), .ZN(P1_U3246) );
  INV_X1 U10520 ( .A(n9079), .ZN(n9093) );
  INV_X1 U10521 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9081) );
  OAI21_X1 U10522 ( .B1(n9862), .B2(n9081), .A(n9080), .ZN(n9082) );
  AOI21_X1 U10523 ( .B1(n9839), .B2(n9083), .A(n9082), .ZN(n9092) );
  OAI211_X1 U10524 ( .C1(n9086), .C2(n9085), .A(n9842), .B(n9084), .ZN(n9091)
         );
  OAI211_X1 U10525 ( .C1(n9089), .C2(n9088), .A(n9850), .B(n9087), .ZN(n9090)
         );
  NAND4_X1 U10526 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(
        P1_U3247) );
  INV_X1 U10527 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9095) );
  OAI21_X1 U10528 ( .B1(n9862), .B2(n9095), .A(n9094), .ZN(n9096) );
  AOI21_X1 U10529 ( .B1(n9097), .B2(n9839), .A(n9096), .ZN(n9106) );
  OAI211_X1 U10530 ( .C1(n9100), .C2(n9099), .A(n9842), .B(n9098), .ZN(n9105)
         );
  OAI211_X1 U10531 ( .C1(n9103), .C2(n9102), .A(n9850), .B(n9101), .ZN(n9104)
         );
  NAND3_X1 U10532 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(P1_U3248) );
  INV_X1 U10533 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9108) );
  OAI21_X1 U10534 ( .B1(n9862), .B2(n9108), .A(n9107), .ZN(n9109) );
  AOI21_X1 U10535 ( .B1(n9110), .B2(n9839), .A(n9109), .ZN(n9119) );
  OAI211_X1 U10536 ( .C1(n9113), .C2(n9112), .A(n9842), .B(n9111), .ZN(n9118)
         );
  OAI211_X1 U10537 ( .C1(n9116), .C2(n9115), .A(n9850), .B(n9114), .ZN(n9117)
         );
  NAND3_X1 U10538 ( .A1(n9119), .A2(n9118), .A3(n9117), .ZN(P1_U3249) );
  INV_X1 U10539 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9121) );
  OAI21_X1 U10540 ( .B1(n9862), .B2(n9121), .A(n9120), .ZN(n9122) );
  AOI21_X1 U10541 ( .B1(n9123), .B2(n9839), .A(n9122), .ZN(n9132) );
  OAI211_X1 U10542 ( .C1(n9126), .C2(n9125), .A(n9842), .B(n9124), .ZN(n9131)
         );
  OAI211_X1 U10543 ( .C1(n9129), .C2(n9128), .A(n9850), .B(n9127), .ZN(n9130)
         );
  NAND3_X1 U10544 ( .A1(n9132), .A2(n9131), .A3(n9130), .ZN(P1_U3250) );
  INV_X1 U10545 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9134) );
  OAI21_X1 U10546 ( .B1(n9862), .B2(n9134), .A(n9133), .ZN(n9135) );
  AOI21_X1 U10547 ( .B1(n9136), .B2(n9839), .A(n9135), .ZN(n9145) );
  OAI211_X1 U10548 ( .C1(n9139), .C2(n9138), .A(n9850), .B(n9137), .ZN(n9144)
         );
  OAI211_X1 U10549 ( .C1(n9142), .C2(n9141), .A(n9842), .B(n9140), .ZN(n9143)
         );
  NAND3_X1 U10550 ( .A1(n9145), .A2(n9144), .A3(n9143), .ZN(P1_U3251) );
  INV_X1 U10551 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9147) );
  OAI21_X1 U10552 ( .B1(n9862), .B2(n9147), .A(n9146), .ZN(n9148) );
  AOI21_X1 U10553 ( .B1(n9149), .B2(n9839), .A(n9148), .ZN(n9158) );
  OAI211_X1 U10554 ( .C1(n9152), .C2(n9151), .A(n9842), .B(n9150), .ZN(n9157)
         );
  OAI211_X1 U10555 ( .C1(n9155), .C2(n9154), .A(n9153), .B(n9850), .ZN(n9156)
         );
  NAND3_X1 U10556 ( .A1(n9158), .A2(n9157), .A3(n9156), .ZN(P1_U3254) );
  XNOR2_X1 U10557 ( .A(n9496), .B(n9168), .ZN(n9159) );
  NAND2_X1 U10558 ( .A1(n9386), .A2(n9863), .ZN(n9167) );
  NAND2_X1 U10559 ( .A1(n9160), .A2(n9378), .ZN(n9166) );
  INV_X1 U10560 ( .A(n9161), .ZN(n9162) );
  NOR2_X1 U10561 ( .A1(n9163), .A2(n9162), .ZN(n9388) );
  INV_X1 U10562 ( .A(n9388), .ZN(n9164) );
  OR2_X1 U10563 ( .A1(n9876), .A2(n9164), .ZN(n9173) );
  NAND2_X1 U10564 ( .A1(n9876), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9165) );
  NAND4_X1 U10565 ( .A1(n9167), .A2(n9166), .A3(n9173), .A4(n9165), .ZN(
        P1_U3263) );
  AOI211_X1 U10566 ( .C1(n9170), .C2(n9169), .A(n9371), .B(n9168), .ZN(n9389)
         );
  NAND2_X1 U10567 ( .A1(n9389), .A2(n9863), .ZN(n9174) );
  NAND2_X1 U10568 ( .A1(n9170), .A2(n9378), .ZN(n9172) );
  NAND2_X1 U10569 ( .A1(n9876), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9171) );
  NAND4_X1 U10570 ( .A1(n9174), .A2(n9173), .A3(n9172), .A4(n9171), .ZN(
        P1_U3264) );
  INV_X1 U10571 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9175) );
  OAI22_X1 U10572 ( .A1(n9176), .A2(n9374), .B1(n9175), .B2(n9383), .ZN(n9177)
         );
  AOI21_X1 U10573 ( .B1(n9400), .B2(n9354), .A(n9177), .ZN(n9180) );
  NAND2_X1 U10574 ( .A1(n9178), .A2(n9378), .ZN(n9179) );
  OAI211_X1 U10575 ( .C1(n9181), .C2(n9381), .A(n9180), .B(n9179), .ZN(n9182)
         );
  AOI21_X1 U10576 ( .B1(n9183), .B2(n9873), .A(n9182), .ZN(n9184) );
  OAI21_X1 U10577 ( .B1(n9185), .B2(n9876), .A(n9184), .ZN(P1_U3356) );
  XNOR2_X1 U10578 ( .A(n9189), .B(n9188), .ZN(n9397) );
  INV_X1 U10579 ( .A(n9191), .ZN(n9192) );
  AOI211_X1 U10580 ( .C1(n9193), .C2(n9207), .A(n9371), .B(n9192), .ZN(n9396)
         );
  NAND2_X1 U10581 ( .A1(n9396), .A2(n9863), .ZN(n9200) );
  INV_X1 U10582 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9194) );
  OAI22_X1 U10583 ( .A1(n9195), .A2(n9374), .B1(n9194), .B2(n9383), .ZN(n9198)
         );
  NOR2_X1 U10584 ( .A1(n9196), .A2(n9349), .ZN(n9197) );
  AOI211_X1 U10585 ( .C1(n9354), .C2(n9409), .A(n9198), .B(n9197), .ZN(n9199)
         );
  OAI211_X1 U10586 ( .C1(n9394), .C2(n9869), .A(n9200), .B(n9199), .ZN(n9201)
         );
  AOI21_X1 U10587 ( .B1(n9397), .B2(n9358), .A(n9201), .ZN(n9202) );
  OAI21_X1 U10588 ( .B1(n9504), .B2(n9385), .A(n9202), .ZN(P1_U3265) );
  INV_X1 U10589 ( .A(n9203), .ZN(n9204) );
  AOI21_X1 U10590 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9508) );
  AOI211_X1 U10591 ( .C1(n9208), .C2(n9223), .A(n9371), .B(n9190), .ZN(n9404)
         );
  NOR2_X1 U10592 ( .A1(n9402), .A2(n9869), .ZN(n9214) );
  AOI22_X1 U10593 ( .A1(n9209), .A2(n9865), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9876), .ZN(n9211) );
  NAND2_X1 U10594 ( .A1(n9417), .A2(n9354), .ZN(n9210) );
  OAI211_X1 U10595 ( .C1(n9212), .C2(n9349), .A(n9211), .B(n9210), .ZN(n9213)
         );
  AOI211_X1 U10596 ( .C1(n9404), .C2(n9863), .A(n9214), .B(n9213), .ZN(n9218)
         );
  XNOR2_X1 U10597 ( .A(n9216), .B(n9215), .ZN(n9405) );
  NAND2_X1 U10598 ( .A1(n9405), .A2(n9358), .ZN(n9217) );
  OAI211_X1 U10599 ( .C1(n9508), .C2(n9385), .A(n9218), .B(n9217), .ZN(
        P1_U3266) );
  OAI21_X1 U10600 ( .B1(n4327), .B2(n4710), .A(n9219), .ZN(n9512) );
  AOI21_X1 U10601 ( .B1(n9221), .B2(n4710), .A(n9220), .ZN(n9222) );
  INV_X1 U10602 ( .A(n9222), .ZN(n9414) );
  OAI211_X1 U10603 ( .C1(n9412), .C2(n9238), .A(n9331), .B(n9223), .ZN(n9411)
         );
  INV_X1 U10604 ( .A(n9224), .ZN(n9225) );
  AOI22_X1 U10605 ( .A1(n9225), .A2(n9865), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9876), .ZN(n9227) );
  NAND2_X1 U10606 ( .A1(n9408), .A2(n9354), .ZN(n9226) );
  OAI211_X1 U10607 ( .C1(n9228), .C2(n9349), .A(n9227), .B(n9226), .ZN(n9229)
         );
  AOI21_X1 U10608 ( .B1(n9230), .B2(n9378), .A(n9229), .ZN(n9231) );
  OAI21_X1 U10609 ( .B1(n9411), .B2(n9381), .A(n9231), .ZN(n9232) );
  AOI21_X1 U10610 ( .B1(n9414), .B2(n9358), .A(n9232), .ZN(n9233) );
  OAI21_X1 U10611 ( .B1(n9512), .B2(n9385), .A(n9233), .ZN(P1_U3267) );
  XNOR2_X1 U10612 ( .A(n9234), .B(n9235), .ZN(n9516) );
  OAI21_X1 U10613 ( .B1(n9257), .B2(n9236), .A(n9235), .ZN(n9237) );
  NAND2_X1 U10614 ( .A1(n4337), .A2(n9237), .ZN(n9422) );
  INV_X1 U10615 ( .A(n9238), .ZN(n9239) );
  OAI211_X1 U10616 ( .C1(n9420), .C2(n9253), .A(n9239), .B(n9331), .ZN(n9419)
         );
  INV_X1 U10617 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9240) );
  OAI22_X1 U10618 ( .A1(n9241), .A2(n9374), .B1(n9240), .B2(n9383), .ZN(n9242)
         );
  AOI21_X1 U10619 ( .B1(n9354), .B2(n9432), .A(n9242), .ZN(n9243) );
  OAI21_X1 U10620 ( .B1(n9244), .B2(n9349), .A(n9243), .ZN(n9245) );
  AOI21_X1 U10621 ( .B1(n9246), .B2(n9378), .A(n9245), .ZN(n9247) );
  OAI21_X1 U10622 ( .B1(n9419), .B2(n9381), .A(n9247), .ZN(n9248) );
  AOI21_X1 U10623 ( .B1(n9422), .B2(n9358), .A(n9248), .ZN(n9249) );
  OAI21_X1 U10624 ( .B1(n9516), .B2(n9385), .A(n9249), .ZN(P1_U3268) );
  XNOR2_X1 U10625 ( .A(n9251), .B(n9250), .ZN(n9431) );
  INV_X1 U10626 ( .A(n9252), .ZN(n9273) );
  AOI211_X1 U10627 ( .C1(n9426), .C2(n9273), .A(n9371), .B(n9253), .ZN(n9425)
         );
  AOI22_X1 U10628 ( .A1(n9254), .A2(n9865), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9876), .ZN(n9255) );
  OAI21_X1 U10629 ( .B1(n9256), .B2(n9869), .A(n9255), .ZN(n9267) );
  AOI211_X1 U10630 ( .C1(n9260), .C2(n9259), .A(n9258), .B(n9257), .ZN(n9265)
         );
  OAI22_X1 U10631 ( .A1(n9263), .A2(n9262), .B1(n9291), .B2(n9261), .ZN(n9264)
         );
  NOR2_X1 U10632 ( .A1(n9265), .A2(n9264), .ZN(n9429) );
  NOR2_X1 U10633 ( .A1(n9429), .A2(n9876), .ZN(n9266) );
  AOI211_X1 U10634 ( .C1(n9425), .C2(n9863), .A(n9267), .B(n9266), .ZN(n9268)
         );
  OAI21_X1 U10635 ( .B1(n9431), .B2(n9385), .A(n9268), .ZN(P1_U3269) );
  XNOR2_X1 U10636 ( .A(n9270), .B(n9269), .ZN(n9520) );
  XNOR2_X1 U10637 ( .A(n9272), .B(n9271), .ZN(n9437) );
  OAI211_X1 U10638 ( .C1(n9435), .C2(n9285), .A(n9273), .B(n9331), .ZN(n9434)
         );
  INV_X1 U10639 ( .A(n9274), .ZN(n9275) );
  AOI22_X1 U10640 ( .A1(n9275), .A2(n9865), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9876), .ZN(n9277) );
  NAND2_X1 U10641 ( .A1(n9449), .A2(n9354), .ZN(n9276) );
  OAI211_X1 U10642 ( .C1(n9278), .C2(n9349), .A(n9277), .B(n9276), .ZN(n9279)
         );
  AOI21_X1 U10643 ( .B1(n9280), .B2(n9378), .A(n9279), .ZN(n9281) );
  OAI21_X1 U10644 ( .B1(n9434), .B2(n9381), .A(n9281), .ZN(n9282) );
  AOI21_X1 U10645 ( .B1(n9437), .B2(n9358), .A(n9282), .ZN(n9283) );
  OAI21_X1 U10646 ( .B1(n9520), .B2(n9385), .A(n9283), .ZN(P1_U3270) );
  XOR2_X1 U10647 ( .A(n9294), .B(n9284), .Z(n9524) );
  AOI211_X1 U10648 ( .C1(n9286), .C2(n9303), .A(n9371), .B(n9285), .ZN(n9444)
         );
  NOR2_X1 U10649 ( .A1(n9443), .A2(n9869), .ZN(n9293) );
  INV_X1 U10650 ( .A(n9287), .ZN(n9288) );
  AOI22_X1 U10651 ( .A1(n9288), .A2(n9865), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9876), .ZN(n9290) );
  NAND2_X1 U10652 ( .A1(n9354), .A2(n9440), .ZN(n9289) );
  OAI211_X1 U10653 ( .C1(n9291), .C2(n9349), .A(n9290), .B(n9289), .ZN(n9292)
         );
  AOI211_X1 U10654 ( .C1(n9444), .C2(n9863), .A(n9293), .B(n9292), .ZN(n9297)
         );
  XNOR2_X1 U10655 ( .A(n9295), .B(n9294), .ZN(n9446) );
  NAND2_X1 U10656 ( .A1(n9446), .A2(n9358), .ZN(n9296) );
  OAI211_X1 U10657 ( .C1(n9524), .C2(n9385), .A(n9297), .B(n9296), .ZN(
        P1_U3271) );
  XNOR2_X1 U10658 ( .A(n9298), .B(n9301), .ZN(n9527) );
  AND2_X1 U10659 ( .A1(n9315), .A2(n9299), .ZN(n9302) );
  OAI21_X1 U10660 ( .B1(n9302), .B2(n9301), .A(n9300), .ZN(n9454) );
  OAI211_X1 U10661 ( .C1(n9452), .C2(n9320), .A(n9331), .B(n9303), .ZN(n9451)
         );
  INV_X1 U10662 ( .A(n9304), .ZN(n9305) );
  AOI22_X1 U10663 ( .A1(n9305), .A2(n9865), .B1(n9876), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U10664 ( .A1(n9354), .A2(n9465), .ZN(n9306) );
  OAI211_X1 U10665 ( .C1(n9308), .C2(n9349), .A(n9307), .B(n9306), .ZN(n9309)
         );
  AOI21_X1 U10666 ( .B1(n9310), .B2(n9378), .A(n9309), .ZN(n9311) );
  OAI21_X1 U10667 ( .B1(n9451), .B2(n9381), .A(n9311), .ZN(n9312) );
  AOI21_X1 U10668 ( .B1(n9454), .B2(n9358), .A(n9312), .ZN(n9313) );
  OAI21_X1 U10669 ( .B1(n9527), .B2(n9385), .A(n9313), .ZN(P1_U3272) );
  XNOR2_X1 U10670 ( .A(n9314), .B(n9316), .ZN(n9529) );
  INV_X1 U10671 ( .A(n9529), .ZN(n9327) );
  OAI211_X1 U10672 ( .C1(n9317), .C2(n9316), .A(n9315), .B(n9482), .ZN(n9319)
         );
  NAND2_X1 U10673 ( .A1(n9319), .A2(n9318), .ZN(n9459) );
  AOI211_X1 U10674 ( .C1(n9321), .C2(n4366), .A(n9371), .B(n9320), .ZN(n9458)
         );
  NAND2_X1 U10675 ( .A1(n9458), .A2(n9863), .ZN(n9324) );
  AOI22_X1 U10676 ( .A1(n9876), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9322), .B2(
        n9865), .ZN(n9323) );
  OAI211_X1 U10677 ( .C1(n9535), .C2(n9869), .A(n9324), .B(n9323), .ZN(n9325)
         );
  AOI21_X1 U10678 ( .B1(n9383), .B2(n9459), .A(n9325), .ZN(n9326) );
  OAI21_X1 U10679 ( .B1(n9327), .B2(n9385), .A(n9326), .ZN(P1_U3273) );
  XOR2_X1 U10680 ( .A(n9329), .B(n9328), .Z(n9539) );
  XNOR2_X1 U10681 ( .A(n9330), .B(n9329), .ZN(n9470) );
  OAI211_X1 U10682 ( .C1(n9468), .C2(n9346), .A(n4366), .B(n9331), .ZN(n9467)
         );
  OAI22_X1 U10683 ( .A1(n9383), .A2(n9333), .B1(n9332), .B2(n9374), .ZN(n9334)
         );
  AOI21_X1 U10684 ( .B1(n9354), .B2(n9464), .A(n9334), .ZN(n9335) );
  OAI21_X1 U10685 ( .B1(n9336), .B2(n9349), .A(n9335), .ZN(n9337) );
  AOI21_X1 U10686 ( .B1(n9338), .B2(n9378), .A(n9337), .ZN(n9339) );
  OAI21_X1 U10687 ( .B1(n9467), .B2(n9381), .A(n9339), .ZN(n9340) );
  AOI21_X1 U10688 ( .B1(n9470), .B2(n9358), .A(n9340), .ZN(n9341) );
  OAI21_X1 U10689 ( .B1(n9539), .B2(n9385), .A(n9341), .ZN(P1_U3274) );
  XOR2_X1 U10690 ( .A(n9342), .B(n9344), .Z(n9543) );
  OAI21_X1 U10691 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9481) );
  AOI211_X1 U10692 ( .C1(n9347), .C2(n4369), .A(n9371), .B(n9346), .ZN(n9479)
         );
  NAND2_X1 U10693 ( .A1(n9479), .A2(n9863), .ZN(n9356) );
  NOR2_X1 U10694 ( .A1(n9349), .A2(n9348), .ZN(n9353) );
  INV_X1 U10695 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9351) );
  OAI22_X1 U10696 ( .A1(n9383), .A2(n9351), .B1(n9350), .B2(n9374), .ZN(n9352)
         );
  AOI211_X1 U10697 ( .C1(n9354), .C2(n9473), .A(n9353), .B(n9352), .ZN(n9355)
         );
  OAI211_X1 U10698 ( .C1(n9478), .C2(n9869), .A(n9356), .B(n9355), .ZN(n9357)
         );
  AOI21_X1 U10699 ( .B1(n9358), .B2(n9481), .A(n9357), .ZN(n9359) );
  OAI21_X1 U10700 ( .B1(n9543), .B2(n9385), .A(n9359), .ZN(P1_U3275) );
  XNOR2_X1 U10701 ( .A(n9360), .B(n9363), .ZN(n9549) );
  NAND2_X1 U10702 ( .A1(n9362), .A2(n9361), .ZN(n9365) );
  INV_X1 U10703 ( .A(n9363), .ZN(n9364) );
  NAND2_X1 U10704 ( .A1(n9365), .A2(n9364), .ZN(n9367) );
  NAND3_X1 U10705 ( .A1(n9367), .A2(n9366), .A3(n9482), .ZN(n9370) );
  AOI22_X1 U10706 ( .A1(n9474), .A2(n9368), .B1(n9464), .B2(n9475), .ZN(n9369)
         );
  NAND2_X1 U10707 ( .A1(n9370), .A2(n9369), .ZN(n9488) );
  AOI21_X1 U10708 ( .B1(n9379), .B2(n9372), .A(n9371), .ZN(n9373) );
  NAND2_X1 U10709 ( .A1(n9373), .A2(n4369), .ZN(n9485) );
  OAI22_X1 U10710 ( .A1(n9383), .A2(n9376), .B1(n9375), .B2(n9374), .ZN(n9377)
         );
  AOI21_X1 U10711 ( .B1(n9379), .B2(n9378), .A(n9377), .ZN(n9380) );
  OAI21_X1 U10712 ( .B1(n9485), .B2(n9381), .A(n9380), .ZN(n9382) );
  AOI21_X1 U10713 ( .B1(n9488), .B2(n9383), .A(n9382), .ZN(n9384) );
  OAI21_X1 U10714 ( .B1(n9549), .B2(n9385), .A(n9384), .ZN(P1_U3276) );
  INV_X1 U10715 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9694) );
  NOR2_X1 U10716 ( .A1(n9386), .A2(n9388), .ZN(n9493) );
  MUX2_X1 U10717 ( .A(n9694), .B(n9493), .S(n9914), .Z(n9387) );
  OAI21_X1 U10718 ( .B1(n9496), .B2(n9463), .A(n9387), .ZN(P1_U3553) );
  NOR2_X1 U10719 ( .A1(n9389), .A2(n9388), .ZN(n9497) );
  MUX2_X1 U10720 ( .A(n9390), .B(n9497), .S(n9914), .Z(n9391) );
  OAI21_X1 U10721 ( .B1(n9500), .B2(n9463), .A(n9391), .ZN(P1_U3552) );
  AOI22_X1 U10722 ( .A1(n9392), .A2(n9475), .B1(n9409), .B2(n9474), .ZN(n9393)
         );
  OAI21_X1 U10723 ( .B1(n9394), .B2(n9901), .A(n9393), .ZN(n9395) );
  AOI211_X1 U10724 ( .C1(n9397), .C2(n9482), .A(n9396), .B(n9395), .ZN(n9501)
         );
  MUX2_X1 U10725 ( .A(n9398), .B(n9501), .S(n9914), .Z(n9399) );
  OAI21_X1 U10726 ( .B1(n9504), .B2(n9491), .A(n9399), .ZN(P1_U3550) );
  AOI22_X1 U10727 ( .A1(n9400), .A2(n9475), .B1(n9474), .B2(n9417), .ZN(n9401)
         );
  OAI21_X1 U10728 ( .B1(n9402), .B2(n9901), .A(n9401), .ZN(n9403) );
  AOI211_X1 U10729 ( .C1(n9405), .C2(n9482), .A(n9404), .B(n9403), .ZN(n9505)
         );
  MUX2_X1 U10730 ( .A(n9406), .B(n9505), .S(n9914), .Z(n9407) );
  OAI21_X1 U10731 ( .B1(n9508), .B2(n9491), .A(n9407), .ZN(P1_U3549) );
  AOI22_X1 U10732 ( .A1(n9409), .A2(n9475), .B1(n9474), .B2(n9408), .ZN(n9410)
         );
  OAI211_X1 U10733 ( .C1(n9412), .C2(n9901), .A(n9411), .B(n9410), .ZN(n9413)
         );
  AOI21_X1 U10734 ( .B1(n9414), .B2(n9482), .A(n9413), .ZN(n9509) );
  MUX2_X1 U10735 ( .A(n9415), .B(n9509), .S(n9914), .Z(n9416) );
  OAI21_X1 U10736 ( .B1(n9512), .B2(n9491), .A(n9416), .ZN(P1_U3548) );
  AOI22_X1 U10737 ( .A1(n9417), .A2(n9475), .B1(n9474), .B2(n9432), .ZN(n9418)
         );
  OAI211_X1 U10738 ( .C1(n9420), .C2(n9901), .A(n9419), .B(n9418), .ZN(n9421)
         );
  AOI21_X1 U10739 ( .B1(n9422), .B2(n9482), .A(n9421), .ZN(n9513) );
  MUX2_X1 U10740 ( .A(n9423), .B(n9513), .S(n9914), .Z(n9424) );
  OAI21_X1 U10741 ( .B1(n9516), .B2(n9491), .A(n9424), .ZN(P1_U3547) );
  INV_X1 U10742 ( .A(n9905), .ZN(n9430) );
  AOI21_X1 U10743 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(n9428) );
  OAI211_X1 U10744 ( .C1(n9431), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9517)
         );
  MUX2_X1 U10745 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9517), .S(n9914), .Z(
        P1_U3546) );
  INV_X1 U10746 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9438) );
  AOI22_X1 U10747 ( .A1(n9432), .A2(n9475), .B1(n9474), .B2(n9449), .ZN(n9433)
         );
  OAI211_X1 U10748 ( .C1(n9435), .C2(n9901), .A(n9434), .B(n9433), .ZN(n9436)
         );
  AOI21_X1 U10749 ( .B1(n9437), .B2(n9482), .A(n9436), .ZN(n9518) );
  MUX2_X1 U10750 ( .A(n9438), .B(n9518), .S(n9914), .Z(n9439) );
  OAI21_X1 U10751 ( .B1(n9520), .B2(n9491), .A(n9439), .ZN(P1_U3545) );
  AOI22_X1 U10752 ( .A1(n9441), .A2(n9475), .B1(n9474), .B2(n9440), .ZN(n9442)
         );
  OAI21_X1 U10753 ( .B1(n9443), .B2(n9901), .A(n9442), .ZN(n9445) );
  AOI211_X1 U10754 ( .C1(n9446), .C2(n9482), .A(n9445), .B(n9444), .ZN(n9521)
         );
  MUX2_X1 U10755 ( .A(n9447), .B(n9521), .S(n9914), .Z(n9448) );
  OAI21_X1 U10756 ( .B1(n9524), .B2(n9491), .A(n9448), .ZN(P1_U3544) );
  INV_X1 U10757 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9455) );
  AOI22_X1 U10758 ( .A1(n9449), .A2(n9475), .B1(n9474), .B2(n9465), .ZN(n9450)
         );
  OAI211_X1 U10759 ( .C1(n9452), .C2(n9901), .A(n9451), .B(n9450), .ZN(n9453)
         );
  AOI21_X1 U10760 ( .B1(n9454), .B2(n9482), .A(n9453), .ZN(n9525) );
  MUX2_X1 U10761 ( .A(n9455), .B(n9525), .S(n9914), .Z(n9456) );
  OAI21_X1 U10762 ( .B1(n9527), .B2(n9491), .A(n9456), .ZN(P1_U3543) );
  NAND2_X1 U10763 ( .A1(n9529), .A2(n9457), .ZN(n9462) );
  INV_X1 U10764 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9460) );
  NOR2_X1 U10765 ( .A1(n9459), .A2(n9458), .ZN(n9530) );
  MUX2_X1 U10766 ( .A(n9460), .B(n9530), .S(n9914), .Z(n9461) );
  OAI211_X1 U10767 ( .C1(n9535), .C2(n9463), .A(n9462), .B(n9461), .ZN(
        P1_U3542) );
  AOI22_X1 U10768 ( .A1(n9465), .A2(n9475), .B1(n9474), .B2(n9464), .ZN(n9466)
         );
  OAI211_X1 U10769 ( .C1(n9468), .C2(n9901), .A(n9467), .B(n9466), .ZN(n9469)
         );
  AOI21_X1 U10770 ( .B1(n9470), .B2(n9482), .A(n9469), .ZN(n9536) );
  MUX2_X1 U10771 ( .A(n9471), .B(n9536), .S(n9914), .Z(n9472) );
  OAI21_X1 U10772 ( .B1(n9539), .B2(n9491), .A(n9472), .ZN(P1_U3541) );
  AOI22_X1 U10773 ( .A1(n9476), .A2(n9475), .B1(n9474), .B2(n9473), .ZN(n9477)
         );
  OAI21_X1 U10774 ( .B1(n9478), .B2(n9901), .A(n9477), .ZN(n9480) );
  AOI211_X1 U10775 ( .C1(n9482), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9540)
         );
  MUX2_X1 U10776 ( .A(n9483), .B(n9540), .S(n9914), .Z(n9484) );
  OAI21_X1 U10777 ( .B1(n9543), .B2(n9491), .A(n9484), .ZN(P1_U3540) );
  OAI21_X1 U10778 ( .B1(n9486), .B2(n9901), .A(n9485), .ZN(n9487) );
  NOR2_X1 U10779 ( .A1(n9488), .A2(n9487), .ZN(n9545) );
  MUX2_X1 U10780 ( .A(n9489), .B(n9545), .S(n9914), .Z(n9490) );
  OAI21_X1 U10781 ( .B1(n9549), .B2(n9491), .A(n9490), .ZN(P1_U3539) );
  MUX2_X1 U10782 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9492), .S(n9914), .Z(
        P1_U3522) );
  INV_X1 U10783 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9494) );
  MUX2_X1 U10784 ( .A(n9494), .B(n9493), .S(n9908), .Z(n9495) );
  OAI21_X1 U10785 ( .B1(n9496), .B2(n9534), .A(n9495), .ZN(P1_U3521) );
  INV_X1 U10786 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9498) );
  MUX2_X1 U10787 ( .A(n9498), .B(n9497), .S(n9908), .Z(n9499) );
  OAI21_X1 U10788 ( .B1(n9500), .B2(n9534), .A(n9499), .ZN(P1_U3520) );
  INV_X1 U10789 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U10790 ( .A(n9502), .B(n9501), .S(n9908), .Z(n9503) );
  OAI21_X1 U10791 ( .B1(n9504), .B2(n9548), .A(n9503), .ZN(P1_U3518) );
  INV_X1 U10792 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U10793 ( .A(n9506), .B(n9505), .S(n9908), .Z(n9507) );
  OAI21_X1 U10794 ( .B1(n9508), .B2(n9548), .A(n9507), .ZN(P1_U3517) );
  INV_X1 U10795 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9510) );
  MUX2_X1 U10796 ( .A(n9510), .B(n9509), .S(n9908), .Z(n9511) );
  OAI21_X1 U10797 ( .B1(n9512), .B2(n9548), .A(n9511), .ZN(P1_U3516) );
  INV_X1 U10798 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9514) );
  MUX2_X1 U10799 ( .A(n9514), .B(n9513), .S(n9908), .Z(n9515) );
  OAI21_X1 U10800 ( .B1(n9516), .B2(n9548), .A(n9515), .ZN(P1_U3515) );
  MUX2_X1 U10801 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9517), .S(n9544), .Z(
        P1_U3514) );
  MUX2_X1 U10802 ( .A(n9671), .B(n9518), .S(n9544), .Z(n9519) );
  OAI21_X1 U10803 ( .B1(n9520), .B2(n9548), .A(n9519), .ZN(P1_U3513) );
  INV_X1 U10804 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9522) );
  MUX2_X1 U10805 ( .A(n9522), .B(n9521), .S(n9544), .Z(n9523) );
  OAI21_X1 U10806 ( .B1(n9524), .B2(n9548), .A(n9523), .ZN(P1_U3512) );
  MUX2_X1 U10807 ( .A(n9613), .B(n9525), .S(n9544), .Z(n9526) );
  OAI21_X1 U10808 ( .B1(n9527), .B2(n9548), .A(n9526), .ZN(P1_U3511) );
  NAND2_X1 U10809 ( .A1(n9529), .A2(n9528), .ZN(n9533) );
  INV_X1 U10810 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U10811 ( .A(n9531), .B(n9530), .S(n9544), .Z(n9532) );
  OAI211_X1 U10812 ( .C1(n9535), .C2(n9534), .A(n9533), .B(n9532), .ZN(
        P1_U3510) );
  INV_X1 U10813 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9537) );
  MUX2_X1 U10814 ( .A(n9537), .B(n9536), .S(n9544), .Z(n9538) );
  OAI21_X1 U10815 ( .B1(n9539), .B2(n9548), .A(n9538), .ZN(P1_U3509) );
  INV_X1 U10816 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9541) );
  MUX2_X1 U10817 ( .A(n9541), .B(n9540), .S(n9544), .Z(n9542) );
  OAI21_X1 U10818 ( .B1(n9543), .B2(n9548), .A(n9542), .ZN(P1_U3507) );
  INV_X1 U10819 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9546) );
  MUX2_X1 U10820 ( .A(n9546), .B(n9545), .S(n9544), .Z(n9547) );
  OAI21_X1 U10821 ( .B1(n9549), .B2(n9548), .A(n9547), .ZN(P1_U3504) );
  MUX2_X1 U10822 ( .A(n9552), .B(P1_D_REG_1__SCAN_IN), .S(n9883), .Z(P1_U3440)
         );
  MUX2_X1 U10823 ( .A(n9553), .B(P1_D_REG_0__SCAN_IN), .S(n9883), .Z(P1_U3439)
         );
  NOR4_X1 U10824 ( .A1(n9555), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9554), .A4(
        n4288), .ZN(n9556) );
  AOI21_X1 U10825 ( .B1(n9570), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9556), .ZN(
        n9557) );
  OAI21_X1 U10826 ( .B1(n9558), .B2(n9565), .A(n9557), .ZN(P1_U3324) );
  OAI222_X1 U10827 ( .A1(n9568), .A2(n9561), .B1(n9565), .B2(n9560), .C1(n9559), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U10828 ( .A1(n9568), .A2(n9697), .B1(n4288), .B2(n9563), .C1(n9565), .C2(n9562), .ZN(P1_U3326) );
  OAI222_X1 U10829 ( .A1(n9568), .A2(n9567), .B1(P1_U3086), .B2(n9566), .C1(
        n9565), .C2(n9564), .ZN(P1_U3328) );
  AOI222_X1 U10830 ( .A1(n9572), .A2(n9571), .B1(P2_DATAO_REG_26__SCAN_IN), 
        .B2(n9570), .C1(P1_STATE_REG_SCAN_IN), .C2(n9569), .ZN(n9726) );
  NOR2_X1 U10831 ( .A1(keyinput62), .A2(keyinput57), .ZN(n9578) );
  NAND2_X1 U10832 ( .A1(keyinput7), .A2(keyinput34), .ZN(n9576) );
  NOR3_X1 U10833 ( .A1(keyinput0), .A2(keyinput49), .A3(keyinput9), .ZN(n9574)
         );
  NOR3_X1 U10834 ( .A1(keyinput6), .A2(keyinput11), .A3(keyinput1), .ZN(n9573)
         );
  NAND4_X1 U10835 ( .A1(keyinput33), .A2(n9574), .A3(keyinput48), .A4(n9573), 
        .ZN(n9575) );
  NOR4_X1 U10836 ( .A1(keyinput28), .A2(keyinput36), .A3(n9576), .A4(n9575), 
        .ZN(n9577) );
  NAND4_X1 U10837 ( .A1(keyinput15), .A2(keyinput40), .A3(n9578), .A4(n9577), 
        .ZN(n9602) );
  NOR2_X1 U10838 ( .A1(keyinput53), .A2(keyinput13), .ZN(n9579) );
  NAND3_X1 U10839 ( .A1(keyinput39), .A2(keyinput4), .A3(n9579), .ZN(n9584) );
  NAND3_X1 U10840 ( .A1(keyinput42), .A2(keyinput5), .A3(keyinput32), .ZN(
        n9583) );
  NOR2_X1 U10841 ( .A1(keyinput23), .A2(keyinput21), .ZN(n9581) );
  NOR3_X1 U10842 ( .A1(keyinput19), .A2(keyinput24), .A3(keyinput29), .ZN(
        n9580) );
  NAND4_X1 U10843 ( .A1(keyinput58), .A2(n9581), .A3(keyinput2), .A4(n9580), 
        .ZN(n9582) );
  NOR4_X1 U10844 ( .A1(keyinput55), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(
        n9600) );
  NAND2_X1 U10845 ( .A1(keyinput26), .A2(keyinput52), .ZN(n9585) );
  NOR3_X1 U10846 ( .A1(keyinput18), .A2(keyinput60), .A3(n9585), .ZN(n9599) );
  NAND2_X1 U10847 ( .A1(keyinput61), .A2(keyinput46), .ZN(n9589) );
  NOR3_X1 U10848 ( .A1(keyinput38), .A2(keyinput27), .A3(keyinput20), .ZN(
        n9587) );
  NOR3_X1 U10849 ( .A1(keyinput35), .A2(keyinput59), .A3(keyinput47), .ZN(
        n9586) );
  NAND4_X1 U10850 ( .A1(keyinput3), .A2(n9587), .A3(keyinput63), .A4(n9586), 
        .ZN(n9588) );
  NOR4_X1 U10851 ( .A1(keyinput45), .A2(keyinput16), .A3(n9589), .A4(n9588), 
        .ZN(n9598) );
  NOR2_X1 U10852 ( .A1(keyinput22), .A2(keyinput30), .ZN(n9590) );
  NAND3_X1 U10853 ( .A1(keyinput50), .A2(keyinput14), .A3(n9590), .ZN(n9596)
         );
  NAND3_X1 U10854 ( .A1(keyinput54), .A2(keyinput12), .A3(keyinput25), .ZN(
        n9595) );
  NOR3_X1 U10855 ( .A1(keyinput51), .A2(keyinput31), .A3(keyinput43), .ZN(
        n9593) );
  INV_X1 U10856 ( .A(keyinput37), .ZN(n9591) );
  NOR3_X1 U10857 ( .A1(keyinput41), .A2(keyinput8), .A3(n9591), .ZN(n9592) );
  NAND4_X1 U10858 ( .A1(keyinput44), .A2(n9593), .A3(keyinput17), .A4(n9592), 
        .ZN(n9594) );
  NOR4_X1 U10859 ( .A1(keyinput56), .A2(n9596), .A3(n9595), .A4(n9594), .ZN(
        n9597) );
  NAND4_X1 U10860 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9601)
         );
  OAI21_X1 U10861 ( .B1(n9602), .B2(n9601), .A(keyinput10), .ZN(n9724) );
  AOI22_X1 U10862 ( .A1(keyinput23), .A2(n9605), .B1(keyinput10), .B2(n9603), 
        .ZN(n9604) );
  OAI21_X1 U10863 ( .B1(n9605), .B2(keyinput23), .A(n9604), .ZN(n9617) );
  INV_X1 U10864 ( .A(keyinput53), .ZN(n9607) );
  AOI22_X1 U10865 ( .A1(n9608), .A2(keyinput58), .B1(P2_ADDR_REG_15__SCAN_IN), 
        .B2(n9607), .ZN(n9606) );
  OAI221_X1 U10866 ( .B1(n9608), .B2(keyinput58), .C1(n9607), .C2(
        P2_ADDR_REG_15__SCAN_IN), .A(n9606), .ZN(n9616) );
  INV_X1 U10867 ( .A(keyinput4), .ZN(n9610) );
  AOI22_X1 U10868 ( .A1(n9611), .A2(keyinput39), .B1(P2_ADDR_REG_9__SCAN_IN), 
        .B2(n9610), .ZN(n9609) );
  OAI221_X1 U10869 ( .B1(n9611), .B2(keyinput39), .C1(n9610), .C2(
        P2_ADDR_REG_9__SCAN_IN), .A(n9609), .ZN(n9615) );
  AOI22_X1 U10870 ( .A1(n9613), .A2(keyinput13), .B1(n9881), .B2(keyinput19), 
        .ZN(n9612) );
  OAI221_X1 U10871 ( .B1(n9613), .B2(keyinput13), .C1(n9881), .C2(keyinput19), 
        .A(n9612), .ZN(n9614) );
  NOR4_X1 U10872 ( .A1(n9617), .A2(n9616), .A3(n9615), .A4(n9614), .ZN(n9666)
         );
  AOI22_X1 U10873 ( .A1(n9620), .A2(keyinput24), .B1(keyinput29), .B2(n9619), 
        .ZN(n9618) );
  OAI221_X1 U10874 ( .B1(n9620), .B2(keyinput24), .C1(n9619), .C2(keyinput29), 
        .A(n9618), .ZN(n9621) );
  INV_X1 U10875 ( .A(n9621), .ZN(n9636) );
  AOI22_X1 U10876 ( .A1(n5496), .A2(keyinput55), .B1(n9623), .B2(keyinput33), 
        .ZN(n9622) );
  OAI221_X1 U10877 ( .B1(n5496), .B2(keyinput55), .C1(n9623), .C2(keyinput33), 
        .A(n9622), .ZN(n9626) );
  XNOR2_X1 U10878 ( .A(n9624), .B(keyinput32), .ZN(n9625) );
  NOR2_X1 U10879 ( .A1(n9626), .A2(n9625), .ZN(n9635) );
  INV_X1 U10880 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9629) );
  INV_X1 U10881 ( .A(keyinput2), .ZN(n9628) );
  AOI22_X1 U10882 ( .A1(n9629), .A2(keyinput42), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n9628), .ZN(n9627) );
  OAI221_X1 U10883 ( .B1(n9629), .B2(keyinput42), .C1(n9628), .C2(
        P2_ADDR_REG_17__SCAN_IN), .A(n9627), .ZN(n9630) );
  INV_X1 U10884 ( .A(n9630), .ZN(n9634) );
  INV_X1 U10885 ( .A(keyinput5), .ZN(n9632) );
  INV_X1 U10886 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9631) );
  XNOR2_X1 U10887 ( .A(n9632), .B(n9631), .ZN(n9633) );
  AND4_X1 U10888 ( .A1(n9636), .A2(n9635), .A3(n9634), .A4(n9633), .ZN(n9665)
         );
  AOI22_X1 U10889 ( .A1(n9878), .A2(keyinput9), .B1(n5625), .B2(keyinput15), 
        .ZN(n9637) );
  OAI221_X1 U10890 ( .B1(n9878), .B2(keyinput9), .C1(n5625), .C2(keyinput15), 
        .A(n9637), .ZN(n9649) );
  AOI22_X1 U10891 ( .A1(n9640), .A2(keyinput57), .B1(keyinput7), .B2(n9639), 
        .ZN(n9638) );
  OAI221_X1 U10892 ( .B1(n9640), .B2(keyinput57), .C1(n9639), .C2(keyinput7), 
        .A(n9638), .ZN(n9648) );
  INV_X1 U10893 ( .A(keyinput62), .ZN(n9641) );
  XNOR2_X1 U10894 ( .A(n9641), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n9647) );
  XOR2_X1 U10895 ( .A(n9642), .B(keyinput49), .Z(n9645) );
  XNOR2_X1 U10896 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput0), .ZN(n9644) );
  XNOR2_X1 U10897 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput40), .ZN(n9643) );
  NAND3_X1 U10898 ( .A1(n9645), .A2(n9644), .A3(n9643), .ZN(n9646) );
  NOR4_X1 U10899 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(n9664)
         );
  INV_X1 U10900 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9651) );
  AOI22_X1 U10901 ( .A1(n9651), .A2(keyinput48), .B1(n9877), .B2(keyinput52), 
        .ZN(n9650) );
  OAI221_X1 U10902 ( .B1(n9651), .B2(keyinput48), .C1(n9877), .C2(keyinput52), 
        .A(n9650), .ZN(n9662) );
  AOI22_X1 U10903 ( .A1(n5804), .A2(keyinput11), .B1(keyinput1), .B2(n9653), 
        .ZN(n9652) );
  OAI221_X1 U10904 ( .B1(n5804), .B2(keyinput11), .C1(n9653), .C2(keyinput1), 
        .A(n9652), .ZN(n9661) );
  INV_X1 U10905 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U10906 ( .A1(n5920), .A2(keyinput34), .B1(keyinput6), .B2(n9655), 
        .ZN(n9654) );
  OAI221_X1 U10907 ( .B1(n5920), .B2(keyinput34), .C1(n9655), .C2(keyinput6), 
        .A(n9654), .ZN(n9660) );
  XOR2_X1 U10908 ( .A(n9656), .B(keyinput28), .Z(n9658) );
  XNOR2_X1 U10909 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput36), .ZN(n9657) );
  NAND2_X1 U10910 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  NOR4_X1 U10911 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9663)
         );
  NAND4_X1 U10912 ( .A1(n9666), .A2(n9665), .A3(n9664), .A4(n9663), .ZN(n9723)
         );
  AOI22_X1 U10913 ( .A1(n5849), .A2(keyinput61), .B1(keyinput46), .B2(P1_U3086), .ZN(n9667) );
  OAI221_X1 U10914 ( .B1(n5849), .B2(keyinput61), .C1(n4288), .C2(keyinput46), 
        .A(n9667), .ZN(n9678) );
  AOI22_X1 U10915 ( .A1(n7250), .A2(keyinput16), .B1(n9669), .B2(keyinput35), 
        .ZN(n9668) );
  OAI221_X1 U10916 ( .B1(n7250), .B2(keyinput16), .C1(n9669), .C2(keyinput35), 
        .A(n9668), .ZN(n9677) );
  AOI22_X1 U10917 ( .A1(n9672), .A2(keyinput59), .B1(n9671), .B2(keyinput47), 
        .ZN(n9670) );
  OAI221_X1 U10918 ( .B1(n9672), .B2(keyinput59), .C1(n9671), .C2(keyinput47), 
        .A(n9670), .ZN(n9676) );
  XNOR2_X1 U10919 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput51), .ZN(n9674) );
  XNOR2_X1 U10920 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(keyinput63), .ZN(n9673)
         );
  NAND2_X1 U10921 ( .A1(n9674), .A2(n9673), .ZN(n9675) );
  NOR4_X1 U10922 ( .A1(n9678), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(n9721)
         );
  AOI22_X1 U10923 ( .A1(n9680), .A2(keyinput20), .B1(keyinput45), .B2(n5705), 
        .ZN(n9679) );
  OAI221_X1 U10924 ( .B1(n9680), .B2(keyinput20), .C1(n5705), .C2(keyinput45), 
        .A(n9679), .ZN(n9691) );
  AOI22_X1 U10925 ( .A1(n9880), .A2(keyinput38), .B1(keyinput27), .B2(n9682), 
        .ZN(n9681) );
  OAI221_X1 U10926 ( .B1(n9880), .B2(keyinput38), .C1(n9682), .C2(keyinput27), 
        .A(n9681), .ZN(n9690) );
  AOI22_X1 U10927 ( .A1(n9685), .A2(keyinput60), .B1(n9684), .B2(keyinput18), 
        .ZN(n9683) );
  OAI221_X1 U10928 ( .B1(n9685), .B2(keyinput60), .C1(n9684), .C2(keyinput18), 
        .A(n9683), .ZN(n9689) );
  XNOR2_X1 U10929 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput26), .ZN(n9687) );
  XNOR2_X1 U10930 ( .A(keyinput3), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U10931 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  NOR4_X1 U10932 ( .A1(n9691), .A2(n9690), .A3(n9689), .A4(n9688), .ZN(n9720)
         );
  AOI22_X1 U10933 ( .A1(n9694), .A2(keyinput56), .B1(n9693), .B2(keyinput12), 
        .ZN(n9692) );
  OAI221_X1 U10934 ( .B1(n9694), .B2(keyinput56), .C1(n9693), .C2(keyinput12), 
        .A(n9692), .ZN(n9704) );
  INV_X1 U10935 ( .A(SI_7_), .ZN(n9696) );
  AOI22_X1 U10936 ( .A1(n9697), .A2(keyinput21), .B1(keyinput25), .B2(n9696), 
        .ZN(n9695) );
  OAI221_X1 U10937 ( .B1(n9697), .B2(keyinput21), .C1(n9696), .C2(keyinput25), 
        .A(n9695), .ZN(n9703) );
  XOR2_X1 U10938 ( .A(n5159), .B(keyinput8), .Z(n9701) );
  XNOR2_X1 U10939 ( .A(keyinput17), .B(P2_REG0_REG_9__SCAN_IN), .ZN(n9700) );
  XNOR2_X1 U10940 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput54), .ZN(n9699) );
  XNOR2_X1 U10941 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput37), .ZN(n9698) );
  NAND4_X1 U10942 ( .A1(n9701), .A2(n9700), .A3(n9699), .A4(n9698), .ZN(n9702)
         );
  NOR3_X1 U10943 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9719) );
  INV_X1 U10944 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9707) );
  INV_X1 U10945 ( .A(keyinput14), .ZN(n9706) );
  AOI22_X1 U10946 ( .A1(n9707), .A2(keyinput43), .B1(P2_ADDR_REG_8__SCAN_IN), 
        .B2(n9706), .ZN(n9705) );
  OAI221_X1 U10947 ( .B1(n9707), .B2(keyinput43), .C1(n9706), .C2(
        P2_ADDR_REG_8__SCAN_IN), .A(n9705), .ZN(n9717) );
  INV_X1 U10948 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U10949 ( .A1(n9879), .A2(keyinput44), .B1(keyinput31), .B2(n5377), 
        .ZN(n9708) );
  OAI221_X1 U10950 ( .B1(n9879), .B2(keyinput44), .C1(n5377), .C2(keyinput31), 
        .A(n9708), .ZN(n9716) );
  AOI22_X1 U10951 ( .A1(n9711), .A2(keyinput30), .B1(keyinput41), .B2(n9710), 
        .ZN(n9709) );
  OAI221_X1 U10952 ( .B1(n9711), .B2(keyinput30), .C1(n9710), .C2(keyinput41), 
        .A(n9709), .ZN(n9715) );
  AOI22_X1 U10953 ( .A1(n5579), .A2(keyinput50), .B1(keyinput22), .B2(n9713), 
        .ZN(n9712) );
  OAI221_X1 U10954 ( .B1(n5579), .B2(keyinput50), .C1(n9713), .C2(keyinput22), 
        .A(n9712), .ZN(n9714) );
  NOR4_X1 U10955 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n9718)
         );
  NAND4_X1 U10956 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(n9722)
         );
  AOI211_X1 U10957 ( .C1(SI_17_), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9725)
         );
  XNOR2_X1 U10958 ( .A(n9726), .B(n9725), .ZN(P1_U3329) );
  MUX2_X1 U10959 ( .A(n9727), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10960 ( .A(n9729), .B(n9728), .ZN(n9730) );
  AOI22_X1 U10961 ( .A1(n10053), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(n10061), 
        .B2(n9730), .ZN(n9750) );
  INV_X1 U10962 ( .A(n9731), .ZN(n9733) );
  NAND2_X1 U10963 ( .A1(n9733), .A2(n9732), .ZN(n9737) );
  OAI211_X1 U10964 ( .C1(n9737), .C2(n9736), .A(n9735), .B(n9734), .ZN(n9742)
         );
  INV_X1 U10965 ( .A(n9737), .ZN(n9740) );
  OAI21_X1 U10966 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9741) );
  NAND2_X1 U10967 ( .A1(n9742), .A2(n9741), .ZN(n9749) );
  NAND2_X1 U10968 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n9748) );
  AOI21_X1 U10969 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  OR2_X1 U10970 ( .A1(n9746), .A2(n10065), .ZN(n9747) );
  NAND4_X1 U10971 ( .A1(n9750), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(
        P2_U3200) );
  INV_X1 U10972 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9764) );
  INV_X1 U10973 ( .A(n9751), .ZN(n9752) );
  AOI211_X1 U10974 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n9847), .ZN(n9760)
         );
  INV_X1 U10975 ( .A(n9755), .ZN(n9756) );
  AOI211_X1 U10976 ( .C1(n9758), .C2(n9757), .A(n9809), .B(n9756), .ZN(n9759)
         );
  AOI211_X1 U10977 ( .C1(n9839), .C2(n9761), .A(n9760), .B(n9759), .ZN(n9763)
         );
  OAI211_X1 U10978 ( .C1(n9862), .C2(n9764), .A(n9763), .B(n9762), .ZN(
        P1_U3253) );
  XNOR2_X1 U10979 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10980 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10981 ( .B1(n9766), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9765), .ZN(
        n9767) );
  XOR2_X1 U10982 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9767), .Z(n9770) );
  AOI22_X1 U10983 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9827), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n4288), .ZN(n9768) );
  OAI21_X1 U10984 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(P1_U3243) );
  INV_X1 U10985 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U10986 ( .A1(n9772), .A2(n9771), .ZN(n9773) );
  AOI21_X1 U10987 ( .B1(n9774), .B2(n9773), .A(n9809), .ZN(n9782) );
  NAND2_X1 U10988 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  AOI21_X1 U10989 ( .B1(n9778), .B2(n9777), .A(n9847), .ZN(n9781) );
  NOR2_X1 U10990 ( .A1(n9856), .A2(n9779), .ZN(n9780) );
  NOR3_X1 U10991 ( .A1(n9782), .A2(n9781), .A3(n9780), .ZN(n9784) );
  OAI211_X1 U10992 ( .C1(n9862), .C2(n9785), .A(n9784), .B(n9783), .ZN(
        P1_U3255) );
  INV_X1 U10993 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9797) );
  AOI211_X1 U10994 ( .C1(n9788), .C2(n9787), .A(n9786), .B(n9847), .ZN(n9793)
         );
  AOI211_X1 U10995 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9809), .ZN(n9792)
         );
  AOI211_X1 U10996 ( .C1(n9839), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9796)
         );
  OAI211_X1 U10997 ( .C1(n9862), .C2(n9797), .A(n9796), .B(n9795), .ZN(
        P1_U3256) );
  AOI211_X1 U10998 ( .C1(n9800), .C2(n9799), .A(n9798), .B(n9809), .ZN(n9805)
         );
  AOI211_X1 U10999 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9847), .ZN(n9804)
         );
  AOI211_X1 U11000 ( .C1(n9839), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9808)
         );
  OAI211_X1 U11001 ( .C1(n9631), .C2(n9862), .A(n9808), .B(n9807), .ZN(
        P1_U3257) );
  INV_X1 U11002 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9821) );
  AOI211_X1 U11003 ( .C1(n9812), .C2(n9811), .A(n9810), .B(n9809), .ZN(n9817)
         );
  AOI211_X1 U11004 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9847), .ZN(n9816)
         );
  AOI211_X1 U11005 ( .C1(n9839), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9820)
         );
  OAI211_X1 U11006 ( .C1(n9862), .C2(n9821), .A(n9820), .B(n9819), .ZN(
        P1_U3258) );
  AOI211_X1 U11007 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9847), .ZN(n9825)
         );
  AOI211_X1 U11008 ( .C1(n9827), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9826), .B(
        n9825), .ZN(n9834) );
  OAI21_X1 U11009 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9832) );
  AOI22_X1 U11010 ( .A1(n9832), .A2(n9850), .B1(n9831), .B2(n9839), .ZN(n9833)
         );
  NAND2_X1 U11011 ( .A1(n9834), .A2(n9833), .ZN(P1_U3259) );
  XNOR2_X1 U11012 ( .A(n9836), .B(n9835), .ZN(n9843) );
  XNOR2_X1 U11013 ( .A(n9838), .B(n9837), .ZN(n9841) );
  AOI222_X1 U11014 ( .A1(n9843), .A2(n9842), .B1(n9850), .B2(n9841), .C1(n9840), .C2(n9839), .ZN(n9845) );
  OAI211_X1 U11015 ( .C1(n9862), .C2(n9846), .A(n9845), .B(n9844), .ZN(
        P1_U3260) );
  AOI21_X1 U11016 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n9859) );
  OAI211_X1 U11017 ( .C1(n9853), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9854)
         );
  OAI21_X1 U11018 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9857) );
  AOI21_X1 U11019 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9861) );
  OAI211_X1 U11020 ( .C1(n9862), .C2(n10138), .A(n9861), .B(n9860), .ZN(
        P1_U3261) );
  NAND2_X1 U11021 ( .A1(n9864), .A2(n9863), .ZN(n9868) );
  AOI22_X1 U11022 ( .A1(n9876), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9866), .B2(
        n9865), .ZN(n9867) );
  OAI211_X1 U11023 ( .C1(n9870), .C2(n9869), .A(n9868), .B(n9867), .ZN(n9871)
         );
  AOI21_X1 U11024 ( .B1(n9873), .B2(n9872), .A(n9871), .ZN(n9874) );
  OAI21_X1 U11025 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(P1_U3288) );
  AND2_X1 U11026 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9883), .ZN(P1_U3294) );
  INV_X1 U11027 ( .A(n9883), .ZN(n9882) );
  NOR2_X1 U11028 ( .A1(n9882), .A2(n9877), .ZN(P1_U3295) );
  AND2_X1 U11029 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9883), .ZN(P1_U3296) );
  AND2_X1 U11030 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9883), .ZN(P1_U3297) );
  AND2_X1 U11031 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9883), .ZN(P1_U3298) );
  NOR2_X1 U11032 ( .A1(n9882), .A2(n9878), .ZN(P1_U3299) );
  AND2_X1 U11033 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9883), .ZN(P1_U3300) );
  AND2_X1 U11034 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9883), .ZN(P1_U3301) );
  AND2_X1 U11035 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9883), .ZN(P1_U3302) );
  AND2_X1 U11036 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9883), .ZN(P1_U3303) );
  NOR2_X1 U11037 ( .A1(n9882), .A2(n9879), .ZN(P1_U3304) );
  AND2_X1 U11038 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9883), .ZN(P1_U3305) );
  AND2_X1 U11039 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9883), .ZN(P1_U3306) );
  AND2_X1 U11040 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9883), .ZN(P1_U3307) );
  AND2_X1 U11041 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9883), .ZN(P1_U3308) );
  AND2_X1 U11042 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9883), .ZN(P1_U3309) );
  AND2_X1 U11043 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9883), .ZN(P1_U3310) );
  NOR2_X1 U11044 ( .A1(n9882), .A2(n9880), .ZN(P1_U3311) );
  AND2_X1 U11045 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9883), .ZN(P1_U3312) );
  AND2_X1 U11046 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9883), .ZN(P1_U3313) );
  AND2_X1 U11047 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9883), .ZN(P1_U3314) );
  AND2_X1 U11048 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9883), .ZN(P1_U3315) );
  AND2_X1 U11049 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9883), .ZN(P1_U3316) );
  AND2_X1 U11050 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9883), .ZN(P1_U3317) );
  AND2_X1 U11051 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9883), .ZN(P1_U3318) );
  AND2_X1 U11052 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9883), .ZN(P1_U3319) );
  AND2_X1 U11053 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9883), .ZN(P1_U3320) );
  AND2_X1 U11054 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9883), .ZN(P1_U3321) );
  NOR2_X1 U11055 ( .A1(n9882), .A2(n9881), .ZN(P1_U3322) );
  AND2_X1 U11056 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9883), .ZN(P1_U3323) );
  INV_X1 U11057 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9884) );
  AOI22_X1 U11058 ( .A1(n9908), .A2(n9885), .B1(n9884), .B2(n9906), .ZN(
        P1_U3459) );
  OAI21_X1 U11059 ( .B1(n9887), .B2(n9901), .A(n9886), .ZN(n9889) );
  AOI211_X1 U11060 ( .C1(n9905), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9909)
         );
  INV_X1 U11061 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9891) );
  AOI22_X1 U11062 ( .A1(n9908), .A2(n9909), .B1(n9891), .B2(n9906), .ZN(
        P1_U3471) );
  OAI21_X1 U11063 ( .B1(n9893), .B2(n9901), .A(n9892), .ZN(n9894) );
  AOI21_X1 U11064 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9897) );
  INV_X1 U11065 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U11066 ( .A1(n9908), .A2(n9911), .B1(n9899), .B2(n9906), .ZN(
        P1_U3477) );
  OAI21_X1 U11067 ( .B1(n4449), .B2(n9901), .A(n9900), .ZN(n9903) );
  AOI211_X1 U11068 ( .C1(n9905), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9913)
         );
  INV_X1 U11069 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9907) );
  AOI22_X1 U11070 ( .A1(n9908), .A2(n9913), .B1(n9907), .B2(n9906), .ZN(
        P1_U3480) );
  AOI22_X1 U11071 ( .A1(n9914), .A2(n9909), .B1(n6693), .B2(n5572), .ZN(
        P1_U3528) );
  AOI22_X1 U11072 ( .A1(n9914), .A2(n9911), .B1(n9910), .B2(n5572), .ZN(
        P1_U3530) );
  AOI22_X1 U11073 ( .A1(n9914), .A2(n9913), .B1(n9912), .B2(n5572), .ZN(
        P1_U3531) );
  NAND2_X1 U11074 ( .A1(n9916), .A2(n9915), .ZN(n9917) );
  AOI21_X1 U11075 ( .B1(n9918), .B2(n9917), .A(n10065), .ZN(n9924) );
  XOR2_X1 U11076 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9919), .Z(n9921) );
  OAI22_X1 U11077 ( .A1(n9922), .A2(n9921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9920), .ZN(n9923) );
  AOI211_X1 U11078 ( .C1(n10052), .C2(n9925), .A(n9924), .B(n9923), .ZN(n9930)
         );
  XOR2_X1 U11079 ( .A(n9927), .B(n9926), .Z(n9928) );
  NAND2_X1 U11080 ( .A1(n9928), .A2(n10060), .ZN(n9929) );
  OAI211_X1 U11081 ( .C1(n10135), .C2(n9931), .A(n9930), .B(n9929), .ZN(
        P2_U3183) );
  INV_X1 U11082 ( .A(n9932), .ZN(n9933) );
  AOI22_X1 U11083 ( .A1(n10053), .A2(P2_ADDR_REG_10__SCAN_IN), .B1(n10052), 
        .B2(n9933), .ZN(n9949) );
  OAI21_X1 U11084 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9941) );
  OAI21_X1 U11085 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(n9940) );
  AOI22_X1 U11086 ( .A1(n9941), .A2(n10061), .B1(n9940), .B2(n10060), .ZN(
        n9948) );
  AOI21_X1 U11087 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(n9945) );
  OR2_X1 U11088 ( .A1(n9945), .A2(n10065), .ZN(n9946) );
  NAND4_X1 U11089 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(
        P2_U3192) );
  AOI22_X1 U11090 ( .A1(n10053), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10052), 
        .B2(n9950), .ZN(n9965) );
  OAI21_X1 U11091 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n9952), .A(n9951), .ZN(
        n9957) );
  OAI21_X1 U11092 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9956) );
  AOI22_X1 U11093 ( .A1(n9957), .A2(n10061), .B1(n10060), .B2(n9956), .ZN(
        n9964) );
  INV_X1 U11094 ( .A(n9958), .ZN(n9963) );
  AOI21_X1 U11095 ( .B1(n9960), .B2(n7866), .A(n9959), .ZN(n9961) );
  OR2_X1 U11096 ( .A1(n9961), .A2(n10065), .ZN(n9962) );
  NAND4_X1 U11097 ( .A1(n9965), .A2(n9964), .A3(n9963), .A4(n9962), .ZN(
        P2_U3193) );
  AOI22_X1 U11098 ( .A1(n10053), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n10052), 
        .B2(n9966), .ZN(n9983) );
  OAI21_X1 U11099 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9974) );
  OAI21_X1 U11100 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(n9973) );
  AOI22_X1 U11101 ( .A1(n9974), .A2(n10061), .B1(n10060), .B2(n9973), .ZN(
        n9982) );
  INV_X1 U11102 ( .A(n9975), .ZN(n9976) );
  AOI21_X1 U11103 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9979) );
  OR2_X1 U11104 ( .A1(n9979), .A2(n10065), .ZN(n9980) );
  NAND4_X1 U11105 ( .A1(n9983), .A2(n9982), .A3(n9981), .A4(n9980), .ZN(
        P2_U3194) );
  AOI22_X1 U11106 ( .A1(n10053), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(n10052), 
        .B2(n9984), .ZN(n10000) );
  OAI21_X1 U11107 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9986), .A(n9985), .ZN(
        n9991) );
  OAI21_X1 U11108 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(n9990) );
  AOI22_X1 U11109 ( .A1(n9991), .A2(n10061), .B1(n10060), .B2(n9990), .ZN(
        n9999) );
  INV_X1 U11110 ( .A(n9992), .ZN(n9993) );
  NOR2_X1 U11111 ( .A1(n9993), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9996) );
  OAI21_X1 U11112 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9997) );
  NAND4_X1 U11113 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(
        P2_U3195) );
  AOI22_X1 U11114 ( .A1(n10053), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n10052), 
        .B2(n10001), .ZN(n10017) );
  OAI21_X1 U11115 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(n10009) );
  OAI21_X1 U11116 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(n10008) );
  AOI22_X1 U11117 ( .A1(n10009), .A2(n10061), .B1(n10060), .B2(n10008), .ZN(
        n10016) );
  NAND2_X1 U11118 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10015)
         );
  AOI21_X1 U11119 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(n10013) );
  OR2_X1 U11120 ( .A1(n10013), .A2(n10065), .ZN(n10014) );
  NAND4_X1 U11121 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        P2_U3196) );
  AOI22_X1 U11122 ( .A1(n10053), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(n10052), 
        .B2(n10018), .ZN(n10032) );
  OAI21_X1 U11123 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10020), .A(n10019), 
        .ZN(n10025) );
  OAI21_X1 U11124 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n10024) );
  AOI22_X1 U11125 ( .A1(n10025), .A2(n10061), .B1(n10060), .B2(n10024), .ZN(
        n10031) );
  AOI21_X1 U11126 ( .B1(n10027), .B2(n5840), .A(n10026), .ZN(n10028) );
  OR2_X1 U11127 ( .A1(n10065), .A2(n10028), .ZN(n10029) );
  NAND4_X1 U11128 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        P2_U3197) );
  AOI22_X1 U11129 ( .A1(n10053), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(n10052), 
        .B2(n10033), .ZN(n10050) );
  OAI21_X1 U11130 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10041) );
  OAI21_X1 U11131 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(n10040) );
  AOI22_X1 U11132 ( .A1(n10041), .A2(n10061), .B1(n10060), .B2(n10040), .ZN(
        n10049) );
  INV_X1 U11133 ( .A(n10042), .ZN(n10048) );
  AOI21_X1 U11134 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(n10046) );
  OR2_X1 U11135 ( .A1(n10046), .A2(n10065), .ZN(n10047) );
  NAND4_X1 U11136 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        P2_U3198) );
  AOI22_X1 U11137 ( .A1(n10053), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n10052), 
        .B2(n10051), .ZN(n10070) );
  OAI21_X1 U11138 ( .B1(n10055), .B2(P2_REG1_REG_17__SCAN_IN), .A(n10054), 
        .ZN(n10062) );
  OAI21_X1 U11139 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(n10059) );
  AOI22_X1 U11140 ( .A1(n10062), .A2(n10061), .B1(n10060), .B2(n10059), .ZN(
        n10069) );
  NAND2_X1 U11141 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10068)
         );
  AOI21_X1 U11142 ( .B1(n8203), .B2(n10064), .A(n10063), .ZN(n10066) );
  OR2_X1 U11143 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND4_X1 U11144 ( .A1(n10070), .A2(n10069), .A3(n10068), .A4(n10067), .ZN(
        P2_U3199) );
  INV_X1 U11145 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10075) );
  OAI21_X1 U11146 ( .B1(n10072), .B2(n10111), .A(n10071), .ZN(n10073) );
  AOI21_X1 U11147 ( .B1(n10074), .B2(n10114), .A(n10073), .ZN(n10119) );
  AOI22_X1 U11148 ( .A1(n10117), .A2(n10075), .B1(n10119), .B2(n10116), .ZN(
        P2_U3399) );
  NOR2_X1 U11149 ( .A1(n10076), .A2(n10111), .ZN(n10078) );
  AOI211_X1 U11150 ( .C1(n10114), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10120) );
  AOI22_X1 U11151 ( .A1(n10117), .A2(n5669), .B1(n10120), .B2(n10116), .ZN(
        P2_U3402) );
  INV_X1 U11152 ( .A(n10080), .ZN(n10084) );
  OAI22_X1 U11153 ( .A1(n10082), .A2(n10106), .B1(n10081), .B2(n10111), .ZN(
        n10083) );
  NOR2_X1 U11154 ( .A1(n10084), .A2(n10083), .ZN(n10121) );
  AOI22_X1 U11155 ( .A1(n10117), .A2(n5688), .B1(n10121), .B2(n10116), .ZN(
        P2_U3405) );
  NAND2_X1 U11156 ( .A1(n10085), .A2(n10095), .ZN(n10088) );
  OR2_X1 U11157 ( .A1(n10086), .A2(n10106), .ZN(n10087) );
  AOI22_X1 U11158 ( .A1(n10117), .A2(n5705), .B1(n10122), .B2(n10116), .ZN(
        P2_U3408) );
  NOR2_X1 U11159 ( .A1(n10090), .A2(n10101), .ZN(n10092) );
  AOI211_X1 U11160 ( .C1(n10095), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        n10123) );
  AOI22_X1 U11161 ( .A1(n10117), .A2(n5731), .B1(n10123), .B2(n10116), .ZN(
        P2_U3411) );
  NAND2_X1 U11162 ( .A1(n10094), .A2(n10114), .ZN(n10098) );
  NAND2_X1 U11163 ( .A1(n10096), .A2(n10095), .ZN(n10097) );
  AND3_X1 U11164 ( .A1(n10099), .A2(n10098), .A3(n10097), .ZN(n10125) );
  AOI22_X1 U11165 ( .A1(n10117), .A2(n5745), .B1(n10125), .B2(n10116), .ZN(
        P2_U3414) );
  OAI22_X1 U11166 ( .A1(n10102), .A2(n10101), .B1(n10100), .B2(n10111), .ZN(
        n10103) );
  NOR2_X1 U11167 ( .A1(n10104), .A2(n10103), .ZN(n10126) );
  AOI22_X1 U11168 ( .A1(n10117), .A2(n5776), .B1(n10126), .B2(n10116), .ZN(
        P2_U3420) );
  INV_X1 U11169 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10110) );
  OAI22_X1 U11170 ( .A1(n10107), .A2(n10106), .B1(n10105), .B2(n10111), .ZN(
        n10108) );
  NOR2_X1 U11171 ( .A1(n10109), .A2(n10108), .ZN(n10127) );
  AOI22_X1 U11172 ( .A1(n10117), .A2(n10110), .B1(n10127), .B2(n10116), .ZN(
        P2_U3423) );
  NOR2_X1 U11173 ( .A1(n4603), .A2(n10111), .ZN(n10113) );
  AOI211_X1 U11174 ( .C1(n10115), .C2(n10114), .A(n10113), .B(n10112), .ZN(
        n10129) );
  AOI22_X1 U11175 ( .A1(n10117), .A2(n5804), .B1(n10129), .B2(n10116), .ZN(
        P2_U3426) );
  INV_X1 U11176 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U11177 ( .A1(n10130), .A2(n10119), .B1(n10118), .B2(n10128), .ZN(
        P2_U3462) );
  AOI22_X1 U11178 ( .A1(n10130), .A2(n10120), .B1(n6747), .B2(n10128), .ZN(
        P2_U3463) );
  AOI22_X1 U11179 ( .A1(n10130), .A2(n10121), .B1(n5685), .B2(n10128), .ZN(
        P2_U3464) );
  AOI22_X1 U11180 ( .A1(n10130), .A2(n10122), .B1(n5702), .B2(n10128), .ZN(
        P2_U3465) );
  AOI22_X1 U11181 ( .A1(n10130), .A2(n10123), .B1(n7055), .B2(n10128), .ZN(
        P2_U3466) );
  AOI22_X1 U11182 ( .A1(n10130), .A2(n10125), .B1(n10124), .B2(n10128), .ZN(
        P2_U3467) );
  AOI22_X1 U11183 ( .A1(n10130), .A2(n10126), .B1(n8254), .B2(n10128), .ZN(
        P2_U3469) );
  AOI22_X1 U11184 ( .A1(n10130), .A2(n10127), .B1(n5786), .B2(n10128), .ZN(
        P2_U3470) );
  AOI22_X1 U11185 ( .A1(n10130), .A2(n10129), .B1(n8263), .B2(n10128), .ZN(
        P2_U3471) );
  OAI222_X1 U11186 ( .A1(n10135), .A2(n10134), .B1(n10135), .B2(n10133), .C1(
        n10132), .C2(n10131), .ZN(ADD_1068_U5) );
  XOR2_X1 U11187 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11188 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(n10139) );
  XOR2_X1 U11189 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10139), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11190 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(ADD_1068_U56) );
  OAI21_X1 U11191 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(ADD_1068_U57) );
  OAI21_X1 U11192 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(ADD_1068_U58) );
  OAI21_X1 U11193 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(ADD_1068_U59) );
  OAI21_X1 U11194 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(ADD_1068_U60) );
  OAI21_X1 U11195 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(ADD_1068_U61) );
  OAI21_X1 U11196 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(ADD_1068_U62) );
  OAI21_X1 U11197 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(ADD_1068_U63) );
  OAI21_X1 U11198 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(ADD_1068_U50) );
  OAI21_X1 U11199 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(ADD_1068_U51) );
  OAI21_X1 U11200 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(ADD_1068_U47) );
  OAI21_X1 U11201 ( .B1(n10175), .B2(n10174), .A(n10173), .ZN(ADD_1068_U49) );
  OAI21_X1 U11202 ( .B1(n10178), .B2(n10177), .A(n10176), .ZN(ADD_1068_U48) );
  AOI21_X1 U11203 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(ADD_1068_U54) );
  AOI21_X1 U11204 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1068_U53) );
  OAI21_X1 U11205 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(ADD_1068_U52) );
  INV_X2 U4839 ( .A(n9535), .ZN(n9321) );
  CLKBUF_X1 U4811 ( .A(n5636), .Z(n5999) );
  AND3_X1 U4813 ( .A1(n5654), .A2(n5653), .A3(n5652), .ZN(n7973) );
  CLKBUF_X1 U4955 ( .A(n5315), .Z(n5331) );
  CLKBUF_X1 U5794 ( .A(n5694), .Z(n6607) );
endmodule

