

module b21_C_AntiSAT_k_128_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986;

  OR2_X1 U4820 ( .A1(n9441), .A2(n9545), .ZN(n9417) );
  NAND2_X2 U4821 ( .A1(n9282), .A2(n9227), .ZN(n9293) );
  CLKBUF_X2 U4823 ( .A(n5721), .Z(n7858) );
  NAND2_X2 U4824 ( .A1(n6876), .A2(n6954), .ZN(n7920) );
  OR3_X1 U4825 ( .A1(n5539), .A2(n7352), .A3(n7453), .ZN(n6286) );
  CLKBUF_X1 U4826 ( .A(n5143), .Z(n7597) );
  INV_X1 U4827 ( .A(n5843), .ZN(n5703) );
  INV_X1 U4828 ( .A(n5478), .ZN(n5222) );
  INV_X1 U4829 ( .A(n5679), .ZN(n6068) );
  AND2_X1 U4830 ( .A1(n5601), .A2(n4857), .ZN(n4856) );
  INV_X1 U4831 ( .A(n6502), .ZN(n6704) );
  INV_X2 U4832 ( .A(n4333), .ZN(n5505) );
  OR2_X1 U4833 ( .A1(n9264), .A2(n9488), .ZN(n9248) );
  OR2_X1 U4834 ( .A1(n5606), .A2(n5604), .ZN(n5605) );
  BUF_X1 U4835 ( .A(n9747), .Z(n4315) );
  AND4_X1 U4836 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n6829)
         );
  OAI211_X1 U4837 ( .C1(n6210), .C2(n6450), .A(n5106), .B(n5105), .ZN(n6768)
         );
  INV_X1 U4838 ( .A(n6808), .ZN(n9130) );
  NOR2_X2 U4839 ( .A1(n9461), .A2(n4315), .ZN(n6922) );
  XNOR2_X2 U4840 ( .A(n5033), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5043) );
  INV_X2 U4841 ( .A(n6681), .ZN(n6741) );
  AOI21_X2 U4842 ( .B1(n5141), .B2(n4520), .A(n4373), .ZN(n4519) );
  XNOR2_X2 U4843 ( .A(n4901), .B(SI_4_), .ZN(n5141) );
  XNOR2_X2 U4844 ( .A(n5605), .B(n8974), .ZN(n7803) );
  XNOR2_X2 U4845 ( .A(n8880), .B(n8619), .ZN(n8638) );
  INV_X1 U4846 ( .A(n6918), .ZN(n9129) );
  AOI21_X1 U4847 ( .B1(n8059), .B2(n8058), .A(n8057), .ZN(n8066) );
  XNOR2_X1 U4848 ( .A(n7584), .B(n7583), .ZN(n9586) );
  NAND2_X1 U4849 ( .A1(n8621), .A2(n8595), .ZN(n8596) );
  INV_X1 U4850 ( .A(n9365), .ZN(n4873) );
  NAND2_X1 U4851 ( .A1(n6046), .A2(n6045), .ZN(n8886) );
  NOR2_X1 U4852 ( .A1(n9389), .A2(n9219), .ZN(n9390) );
  OAI22_X1 U4853 ( .A1(n8141), .A2(n8140), .B1(n5941), .B2(n5940), .ZN(n8173)
         );
  NAND2_X1 U4854 ( .A1(n5496), .A2(n5495), .ZN(n9505) );
  NAND2_X1 U4855 ( .A1(n5468), .A2(n5467), .ZN(n9510) );
  NOR2_X2 U4856 ( .A1(n9417), .A2(n9539), .ZN(n9405) );
  NAND2_X1 U4857 ( .A1(n7227), .A2(n7316), .ZN(n7315) );
  AOI21_X1 U4858 ( .B1(n6962), .B2(n4344), .A(n4796), .ZN(n7213) );
  NAND2_X1 U4859 ( .A1(n5384), .A2(n5383), .ZN(n9539) );
  NAND2_X1 U4860 ( .A1(n5347), .A2(n5346), .ZN(n9552) );
  OAI21_X1 U4861 ( .B1(n4948), .B2(n4712), .A(n4710), .ZN(n5343) );
  XNOR2_X1 U4862 ( .A(n4631), .B(n5244), .ZN(n6294) );
  NAND2_X1 U4863 ( .A1(n4403), .A2(n4402), .ZN(n6758) );
  AND2_X1 U4864 ( .A1(n7542), .A2(n7637), .ZN(n6916) );
  OR2_X2 U4865 ( .A1(n9667), .A2(n9440), .ZN(n9096) );
  INV_X2 U4866 ( .A(n9837), .ZN(n4316) );
  INV_X2 U4867 ( .A(n9460), .ZN(n9305) );
  NAND2_X1 U4868 ( .A1(n6671), .A2(n7765), .ZN(n6737) );
  INV_X1 U4869 ( .A(n9740), .ZN(n9466) );
  OAI21_X1 U4870 ( .B1(n6226), .B2(n5104), .A(n4612), .ZN(n9747) );
  AND4_X1 U4871 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n6918)
         );
  INV_X2 U4872 ( .A(n9133), .ZN(n6755) );
  NAND2_X2 U4873 ( .A1(n6676), .A2(n5063), .ZN(n5508) );
  AND2_X1 U4874 ( .A1(n5656), .A2(n5655), .ZN(n5659) );
  INV_X2 U4875 ( .A(n6049), .ZN(n7824) );
  CLKBUF_X3 U4876 ( .A(n5703), .Z(n6021) );
  OAI21_X1 U4877 ( .B1(n4522), .B2(n4521), .A(n4519), .ZN(n5160) );
  NAND2_X2 U4878 ( .A1(n6286), .A2(n5063), .ZN(n5478) );
  INV_X1 U4879 ( .A(n5093), .ZN(n5404) );
  AND2_X1 U4880 ( .A1(n8077), .A2(n5042), .ZN(n5093) );
  NAND2_X1 U4881 ( .A1(n7762), .A2(n7792), .ZN(n5063) );
  AND2_X1 U4882 ( .A1(n5025), .A2(n5022), .ZN(n7762) );
  OR2_X1 U4883 ( .A1(n5104), .A2(n6219), .ZN(n5088) );
  NAND2_X1 U4884 ( .A1(n8977), .A2(n5609), .ZN(n8982) );
  NAND2_X1 U4885 ( .A1(n5037), .A2(n9584), .ZN(n5038) );
  CLKBUF_X1 U4886 ( .A(n5036), .Z(n9584) );
  NAND2_X1 U4887 ( .A1(n5036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5033) );
  XNOR2_X1 U4888 ( .A(n5024), .B(n5023), .ZN(n7792) );
  XNOR2_X1 U4889 ( .A(n5649), .B(n5648), .ZN(n8985) );
  INV_X2 U4890 ( .A(n9588), .ZN(n9597) );
  OR2_X1 U4891 ( .A1(n5647), .A2(n4852), .ZN(n5607) );
  NAND2_X1 U4892 ( .A1(n5647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5649) );
  OR2_X1 U4893 ( .A1(n5030), .A2(n5247), .ZN(n4999) );
  INV_X2 U4894 ( .A(n6214), .ZN(n4474) );
  AND2_X1 U4895 ( .A1(n4659), .A2(n5000), .ZN(n4658) );
  NAND2_X1 U4896 ( .A1(n4579), .A2(n4577), .ZN(n4890) );
  AND2_X1 U4897 ( .A1(n4876), .A2(n5557), .ZN(n4659) );
  AND4_X1 U4898 ( .A1(n5016), .A2(n4993), .A3(n8235), .A4(n5023), .ZN(n4997)
         );
  AND2_X1 U4899 ( .A1(n4991), .A2(n4992), .ZN(n4876) );
  AND3_X1 U4900 ( .A1(n4990), .A2(n5055), .A3(n4785), .ZN(n4784) );
  AND2_X1 U4901 ( .A1(n4988), .A2(n4989), .ZN(n4786) );
  INV_X1 U4902 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4581) );
  INV_X1 U4903 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4989) );
  INV_X4 U4904 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4905 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4990) );
  INV_X1 U4906 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4785) );
  INV_X1 U4907 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U4908 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4987) );
  NOR2_X2 U4909 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5099) );
  INV_X4 U4910 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4911 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5023) );
  INV_X1 U4912 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8570) );
  AOI22_X2 U4913 ( .A1(n9431), .A2(n9433), .B1(n9552), .B2(n9424), .ZN(n9416)
         );
  OAI222_X1 U4914 ( .A1(n6866), .A2(n8078), .B1(P2_U3152), .B2(n7803), .C1(
        n7850), .C2(n8987), .ZN(P2_U3328) );
  NAND2_X2 U4915 ( .A1(n5620), .A2(n7803), .ZN(n7854) );
  NAND2_X2 U4916 ( .A1(n7803), .A2(n8982), .ZN(n5843) );
  OR2_X1 U4917 ( .A1(n6681), .A2(n6693), .ZN(n6762) );
  INV_X2 U4918 ( .A(n5417), .ZN(n6181) );
  NOR2_X1 U4919 ( .A1(n7880), .A2(n4530), .ZN(n4529) );
  INV_X1 U4920 ( .A(n7462), .ZN(n4530) );
  OR2_X1 U4921 ( .A1(n9493), .A2(n7530), .ZN(n9253) );
  NAND2_X1 U4922 ( .A1(n5283), .A2(n5282), .ZN(n4948) );
  NOR2_X1 U4923 ( .A1(n5874), .A2(n5633), .ZN(n5650) );
  OR2_X1 U4924 ( .A1(n4787), .A2(n4440), .ZN(n4439) );
  INV_X1 U4925 ( .A(n9030), .ZN(n4440) );
  OR2_X1 U4926 ( .A1(n8109), .A2(n4748), .ZN(n4746) );
  AND2_X1 U4927 ( .A1(n8933), .A2(n8584), .ZN(n4692) );
  AND2_X1 U4928 ( .A1(n7888), .A2(n4821), .ZN(n4820) );
  AOI21_X1 U4929 ( .B1(n4328), .B2(n4395), .A(n4822), .ZN(n4821) );
  AND2_X1 U4930 ( .A1(n8038), .A2(n8036), .ZN(n4822) );
  OR2_X1 U4931 ( .A1(n8875), .A2(n8595), .ZN(n8032) );
  INV_X1 U4932 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4857) );
  AND2_X1 U4933 ( .A1(n5627), .A2(n5788), .ZN(n5804) );
  INV_X1 U4934 ( .A(n9053), .ZN(n4795) );
  CLKBUF_X1 U4935 ( .A(n5090), .Z(n5532) );
  INV_X1 U4936 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4992) );
  OR2_X1 U4937 ( .A1(n7748), .A2(n4698), .ZN(n4697) );
  INV_X1 U4938 ( .A(n5038), .ZN(n5042) );
  NAND2_X1 U4939 ( .A1(n9130), .A2(n6795), .ZN(n7532) );
  INV_X1 U4940 ( .A(n7792), .ZN(n6743) );
  NOR2_X1 U4941 ( .A1(n7797), .A2(n6665), .ZN(n7386) );
  INV_X1 U4942 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U4943 ( .A1(n6061), .A2(n6060), .ZN(n6169) );
  INV_X1 U4944 ( .A(n5424), .ZN(n4732) );
  INV_X1 U4945 ( .A(n4711), .ZN(n4710) );
  OAI21_X1 U4946 ( .B1(n4714), .B2(n4712), .A(n4957), .ZN(n4711) );
  NAND2_X1 U4947 ( .A1(n4713), .A2(n4951), .ZN(n4712) );
  INV_X1 U4948 ( .A(n4704), .ZN(n4703) );
  OR2_X1 U4949 ( .A1(n4930), .A2(n4705), .ZN(n4701) );
  OAI21_X1 U4950 ( .B1(n4707), .B2(n4705), .A(n4941), .ZN(n4704) );
  OAI21_X1 U4951 ( .B1(n4890), .B2(n4540), .A(n5069), .ZN(n4893) );
  NAND2_X1 U4952 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U4953 ( .A1(n7891), .A2(n4743), .ZN(n4742) );
  AND2_X1 U4954 ( .A1(n9850), .A2(n7895), .ZN(n4743) );
  NAND2_X1 U4955 ( .A1(n7274), .A2(n7273), .ZN(n4761) );
  NAND2_X1 U4956 ( .A1(n8163), .A2(n4354), .ZN(n4484) );
  AND2_X1 U4957 ( .A1(n5654), .A2(n4820), .ZN(n4813) );
  OAI21_X1 U4958 ( .B1(n5654), .B2(n4818), .A(n4815), .ZN(n4814) );
  NAND2_X1 U4959 ( .A1(n4818), .A2(n4816), .ZN(n4815) );
  OR2_X1 U4960 ( .A1(n4820), .A2(n5654), .ZN(n4816) );
  INV_X1 U4961 ( .A(n7854), .ZN(n7825) );
  AND2_X1 U4962 ( .A1(n5591), .A2(n5590), .ZN(n5715) );
  NOR2_X1 U4963 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5591) );
  NOR2_X1 U4964 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5590) );
  AND3_X1 U4965 ( .A1(n5715), .A2(n4825), .A3(n8379), .ZN(n5768) );
  NOR2_X1 U4966 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4825) );
  NAND2_X1 U4967 ( .A1(n5635), .A2(n4766), .ZN(n4765) );
  INV_X1 U4968 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5635) );
  INV_X1 U4969 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4766) );
  INV_X1 U4970 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5641) );
  NOR2_X1 U4971 ( .A1(n8706), .A2(n4827), .ZN(n4826) );
  INV_X1 U4972 ( .A(n8005), .ZN(n4827) );
  NOR2_X1 U4973 ( .A1(n8909), .A2(n8914), .ZN(n4563) );
  AOI21_X2 U4974 ( .B1(n8782), .B2(n8587), .A(n8586), .ZN(n8761) );
  NOR2_X1 U4975 ( .A1(n8798), .A2(n8923), .ZN(n8783) );
  OAI21_X1 U4976 ( .B1(n7507), .B2(n7506), .A(n7505), .ZN(n8583) );
  AOI21_X1 U4977 ( .B1(n4529), .B2(n4527), .A(n4366), .ZN(n4526) );
  OR2_X1 U4978 ( .A1(n7476), .A2(n4528), .ZN(n4525) );
  INV_X1 U4979 ( .A(n4529), .ZN(n4528) );
  INV_X1 U4980 ( .A(n7859), .ZN(n5964) );
  NAND2_X1 U4981 ( .A1(n9818), .A2(n7868), .ZN(n4804) );
  NAND2_X1 U4982 ( .A1(n8392), .A2(n9876), .ZN(n7868) );
  NAND2_X1 U4983 ( .A1(n4546), .A2(n4549), .ZN(n4545) );
  OR2_X1 U4984 ( .A1(n8985), .A2(n6214), .ZN(n4544) );
  NAND2_X2 U4985 ( .A1(n4475), .A2(n4473), .ZN(n5767) );
  NOR2_X1 U4986 ( .A1(n4342), .A2(n4409), .ZN(n4473) );
  OR2_X1 U4987 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U4988 ( .A1(n6141), .A2(n8985), .ZN(n5662) );
  INV_X1 U4989 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U4990 ( .A1(n4477), .A2(n4472), .ZN(n6141) );
  INV_X1 U4991 ( .A(n4547), .ZN(n4472) );
  INV_X1 U4992 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5634) );
  AND2_X1 U4993 ( .A1(n6158), .A2(n6157), .ZN(n6193) );
  INV_X1 U4994 ( .A(n4454), .ZN(n4448) );
  NAND2_X1 U4995 ( .A1(n5538), .A2(n5537), .ZN(n8991) );
  AND2_X1 U4996 ( .A1(n7792), .A2(n7383), .ZN(n5568) );
  AND4_X1 U4997 ( .A1(n5579), .A2(n5578), .A3(n5577), .A4(n5576), .ZN(n7530)
         );
  NAND2_X2 U4998 ( .A1(n5043), .A2(n5042), .ZN(n5417) );
  AND2_X1 U4999 ( .A1(n5043), .A2(n5038), .ZN(n5078) );
  AND2_X1 U5000 ( .A1(n9253), .A2(n7727), .ZN(n9271) );
  INV_X1 U5001 ( .A(n4860), .ZN(n4859) );
  OAI21_X1 U5002 ( .B1(n4863), .B2(n4861), .A(n4365), .ZN(n4860) );
  AOI21_X1 U5003 ( .B1(n4621), .B2(n4624), .A(n4368), .ZN(n4619) );
  NAND2_X1 U5004 ( .A1(n4628), .A2(n4317), .ZN(n7336) );
  NAND2_X1 U5005 ( .A1(n4871), .A2(n4870), .ZN(n7312) );
  INV_X1 U5006 ( .A(n7222), .ZN(n4870) );
  INV_X1 U5007 ( .A(n7242), .ZN(n4871) );
  NAND2_X1 U5008 ( .A1(n7677), .A2(n4657), .ZN(n7227) );
  AND2_X1 U5009 ( .A1(n6688), .A2(n9686), .ZN(n9456) );
  NAND2_X1 U5010 ( .A1(n6294), .A2(n5245), .ZN(n4630) );
  NAND2_X1 U5011 ( .A1(n7121), .A2(n7755), .ZN(n9561) );
  AOI21_X1 U5012 ( .B1(n8563), .B2(n9803), .A(n5654), .ZN(n4412) );
  INV_X1 U5013 ( .A(n4770), .ZN(n8992) );
  INV_X1 U5014 ( .A(n7921), .ZN(n4662) );
  NAND2_X1 U5015 ( .A1(n4588), .A2(n4586), .ZN(n7687) );
  NAND2_X1 U5016 ( .A1(n4590), .A2(n4589), .ZN(n4588) );
  INV_X1 U5017 ( .A(n4587), .ZN(n4586) );
  NAND2_X1 U5018 ( .A1(n4591), .A2(n7675), .ZN(n4590) );
  AOI21_X1 U5019 ( .B1(n4610), .B2(n4608), .A(n7689), .ZN(n7693) );
  OAI21_X1 U5020 ( .B1(n4609), .B2(n7681), .A(n4589), .ZN(n4608) );
  INV_X1 U5021 ( .A(n4611), .ZN(n4610) );
  INV_X1 U5022 ( .A(n7718), .ZN(n4716) );
  NOR2_X1 U5023 ( .A1(n4584), .A2(n4319), .ZN(n4717) );
  INV_X1 U5024 ( .A(n7719), .ZN(n4723) );
  INV_X1 U5025 ( .A(n7720), .ZN(n7726) );
  NAND2_X1 U5026 ( .A1(n4601), .A2(n4355), .ZN(n7751) );
  INV_X1 U5027 ( .A(n4908), .ZN(n4617) );
  OR2_X1 U5028 ( .A1(n5995), .A2(n5994), .ZN(n4747) );
  NOR2_X1 U5029 ( .A1(n4361), .A2(n4501), .ZN(n4500) );
  AND2_X1 U5030 ( .A1(n4504), .A2(n4502), .ZN(n4501) );
  INV_X1 U5031 ( .A(n8172), .ZN(n4502) );
  NAND2_X1 U5032 ( .A1(n4500), .A2(n4503), .ZN(n4498) );
  INV_X1 U5033 ( .A(n4504), .ZN(n4503) );
  INV_X1 U5034 ( .A(n7749), .ZN(n4700) );
  INV_X1 U5035 ( .A(SI_15_), .ZN(n4953) );
  INV_X1 U5036 ( .A(n7443), .ZN(n4755) );
  OR2_X1 U5037 ( .A1(n8126), .A2(n5925), .ZN(n4877) );
  AOI21_X1 U5038 ( .B1(n4750), .B2(n4494), .A(n4367), .ZN(n4493) );
  INV_X1 U5039 ( .A(n4496), .ZN(n4494) );
  INV_X1 U5040 ( .A(n4750), .ZN(n4495) );
  AND2_X1 U5041 ( .A1(n8102), .A2(n4345), .ZN(n4504) );
  NOR2_X1 U5042 ( .A1(n4752), .A2(n4497), .ZN(n4496) );
  INV_X1 U5043 ( .A(n5873), .ZN(n4497) );
  NAND2_X1 U5044 ( .A1(n4755), .A2(n5907), .ZN(n4752) );
  NAND2_X1 U5045 ( .A1(n4751), .A2(n5907), .ZN(n4750) );
  INV_X1 U5046 ( .A(n4753), .ZN(n4751) );
  INV_X1 U5047 ( .A(n7803), .ZN(n5621) );
  INV_X1 U5048 ( .A(n8982), .ZN(n5620) );
  NAND2_X1 U5049 ( .A1(n5631), .A2(n5630), .ZN(n5874) );
  INV_X1 U5050 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5630) );
  INV_X1 U5051 ( .A(n5853), .ZN(n5631) );
  NOR2_X1 U5052 ( .A1(n4554), .A2(n8875), .ZN(n4553) );
  OR2_X1 U5053 ( .A1(n8880), .A2(n8886), .ZN(n4554) );
  OR2_X1 U5054 ( .A1(n8891), .A2(n8690), .ZN(n4681) );
  NOR2_X1 U5055 ( .A1(n8687), .A2(n4684), .ZN(n4680) );
  OR2_X1 U5056 ( .A1(n8736), .A2(n8725), .ZN(n4881) );
  INV_X1 U5057 ( .A(n8589), .ZN(n4670) );
  INV_X1 U5058 ( .A(n7997), .ZN(n4811) );
  AOI21_X1 U5059 ( .B1(n4833), .B2(n4839), .A(n7836), .ZN(n4832) );
  OR2_X1 U5060 ( .A1(n8933), .A2(n8803), .ZN(n7982) );
  NOR2_X1 U5061 ( .A1(n4558), .A2(n8581), .ZN(n4557) );
  INV_X1 U5062 ( .A(n4559), .ZN(n4558) );
  NOR2_X1 U5063 ( .A1(n7498), .A2(n8943), .ZN(n4559) );
  INV_X1 U5064 ( .A(n7402), .ZN(n4688) );
  INV_X1 U5065 ( .A(n4846), .ZN(n4845) );
  OAI21_X1 U5066 ( .B1(n4849), .B2(n4847), .A(n4851), .ZN(n4846) );
  OR2_X1 U5067 ( .A1(n7404), .A2(n9907), .ZN(n7954) );
  NAND2_X1 U5068 ( .A1(n6118), .A2(n7909), .ZN(n6700) );
  OAI21_X1 U5069 ( .B1(n8840), .B2(n4534), .A(n4533), .ZN(n4537) );
  AOI21_X1 U5070 ( .B1(n4535), .B2(n4840), .A(n4692), .ZN(n4533) );
  INV_X1 U5071 ( .A(n4535), .ZN(n4534) );
  NAND2_X1 U5072 ( .A1(n6093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6114) );
  INV_X1 U5073 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6091) );
  INV_X1 U5074 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6113) );
  NOR2_X1 U5075 ( .A1(n5599), .A2(n5600), .ZN(n5601) );
  NOR2_X1 U5076 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5598) );
  INV_X1 U5077 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U5078 ( .A1(n4430), .A2(n4427), .ZN(n4426) );
  INV_X1 U5079 ( .A(n5281), .ZN(n4427) );
  AND2_X1 U5080 ( .A1(n5164), .A2(n4340), .ZN(n4780) );
  NAND2_X1 U5081 ( .A1(n6961), .A2(n4799), .ZN(n7196) );
  OR2_X1 U5082 ( .A1(n9036), .A2(n4455), .ZN(n4454) );
  INV_X1 U5083 ( .A(n9045), .ZN(n4455) );
  AND2_X1 U5084 ( .A1(n4389), .A2(n4452), .ZN(n4451) );
  NAND2_X1 U5085 ( .A1(n9045), .A2(n4453), .ZN(n4452) );
  NOR2_X1 U5086 ( .A1(n5478), .A2(n5028), .ZN(n5090) );
  NAND2_X1 U5087 ( .A1(n8998), .A2(n9001), .ZN(n4800) );
  OR2_X1 U5088 ( .A1(n9525), .A2(n9201), .ZN(n7709) );
  NAND2_X1 U5089 ( .A1(n9214), .A2(n4655), .ZN(n4652) );
  NOR2_X1 U5090 ( .A1(n9433), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5091 ( .A1(n9197), .A2(n4568), .ZN(n4566) );
  INV_X1 U5092 ( .A(n7366), .ZN(n4567) );
  OR2_X1 U5093 ( .A1(n7333), .A2(n7421), .ZN(n4568) );
  NAND2_X1 U5094 ( .A1(n6917), .A2(n6916), .ZN(n4648) );
  NAND2_X1 U5095 ( .A1(n9131), .A2(n9718), .ZN(n7764) );
  OAI21_X1 U5096 ( .B1(n5487), .B2(n5486), .A(n5490), .ZN(n5512) );
  NOR2_X1 U5097 ( .A1(n5447), .A2(n4731), .ZN(n4730) );
  INV_X1 U5098 ( .A(n4983), .ZN(n4731) );
  NAND2_X1 U5099 ( .A1(n5019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5021) );
  INV_X1 U5100 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U5101 ( .A1(n5018), .A2(n8235), .ZN(n4801) );
  AND2_X1 U5102 ( .A1(n4961), .A2(n4960), .ZN(n5342) );
  NOR2_X1 U5103 ( .A1(n4952), .A2(n4715), .ZN(n4714) );
  INV_X1 U5104 ( .A(n4947), .ZN(n4715) );
  AND2_X1 U5105 ( .A1(n4947), .A2(n4946), .ZN(n5282) );
  NOR2_X1 U5106 ( .A1(n4934), .A2(n4708), .ZN(n4707) );
  INV_X1 U5107 ( .A(n4929), .ZN(n4708) );
  NAND2_X1 U5108 ( .A1(n5217), .A2(n4886), .ZN(n4930) );
  INV_X1 U5109 ( .A(n4900), .ZN(n4520) );
  INV_X1 U5110 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4580) );
  INV_X1 U5111 ( .A(n6554), .ZN(n4470) );
  NAND2_X1 U5112 ( .A1(n8173), .A2(n8172), .ZN(n4505) );
  XNOR2_X1 U5113 ( .A(n9858), .B(n5679), .ZN(n5667) );
  AND2_X1 U5114 ( .A1(n8155), .A2(n5970), .ZN(n4745) );
  NAND2_X1 U5115 ( .A1(n5982), .A2(n5983), .ZN(n4748) );
  OR2_X1 U5116 ( .A1(n4488), .A2(n4879), .ZN(n4485) );
  AND2_X1 U5117 ( .A1(n4483), .A2(n4486), .ZN(n4481) );
  INV_X1 U5118 ( .A(n8146), .ZN(n4486) );
  NAND2_X1 U5119 ( .A1(n6555), .A2(n4469), .ZN(n4464) );
  OR2_X1 U5120 ( .A1(n4485), .A2(n6025), .ZN(n4483) );
  NAND2_X1 U5121 ( .A1(n4480), .A2(n6017), .ZN(n4479) );
  INV_X1 U5122 ( .A(n4484), .ZN(n4480) );
  AND2_X1 U5123 ( .A1(n5731), .A2(n5714), .ZN(n4758) );
  NOR2_X1 U5124 ( .A1(n5803), .A2(n4516), .ZN(n4515) );
  INV_X1 U5125 ( .A(n7113), .ZN(n4516) );
  NAND2_X1 U5126 ( .A1(n4505), .A2(n4504), .ZN(n8101) );
  AND2_X1 U5127 ( .A1(n5872), .A2(n5852), .ZN(n4760) );
  XNOR2_X1 U5128 ( .A(n5998), .B(n6011), .ZN(n8163) );
  NOR2_X1 U5129 ( .A1(n7105), .A2(n4509), .ZN(n4508) );
  INV_X1 U5130 ( .A(n4511), .ZN(n4509) );
  INV_X1 U5131 ( .A(n4515), .ZN(n4514) );
  NOR2_X1 U5132 ( .A1(n6125), .A2(n9839), .ZN(n6140) );
  NAND2_X1 U5133 ( .A1(n6118), .A2(n8807), .ZN(n6139) );
  AOI21_X1 U5134 ( .B1(n4820), .B2(n4324), .A(n4819), .ZN(n4818) );
  INV_X1 U5135 ( .A(n4823), .ZN(n4819) );
  NOR2_X1 U5136 ( .A1(n8036), .A2(n8037), .ZN(n8600) );
  OR2_X1 U5137 ( .A1(n5843), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U5138 ( .A1(n5621), .A2(n8982), .ZN(n5721) );
  OR2_X1 U5139 ( .A1(n5721), .A2(n5672), .ZN(n5673) );
  NAND2_X1 U5140 ( .A1(n5621), .A2(n5620), .ZN(n5704) );
  NOR2_X1 U5141 ( .A1(n9603), .A2(n4352), .ZN(n9617) );
  INV_X1 U5142 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U5143 ( .A1(n4332), .A2(n8576), .ZN(n8575) );
  AOI21_X1 U5144 ( .B1(n8617), .B2(n8614), .A(n7843), .ZN(n8601) );
  INV_X1 U5145 ( .A(n8875), .ZN(n8621) );
  NAND2_X1 U5146 ( .A1(n8619), .A2(n8819), .ZN(n4421) );
  OR2_X1 U5147 ( .A1(n8891), .A2(n8149), .ZN(n8649) );
  NAND2_X1 U5148 ( .A1(n4523), .A2(n4676), .ZN(n8648) );
  INV_X1 U5149 ( .A(n4677), .ZN(n4676) );
  NAND2_X1 U5150 ( .A1(n8696), .A2(n4678), .ZN(n4523) );
  OAI21_X1 U5151 ( .B1(n8667), .B2(n8593), .A(n4681), .ZN(n4677) );
  NAND2_X1 U5152 ( .A1(n4828), .A2(n4346), .ZN(n8686) );
  NAND2_X1 U5153 ( .A1(n8696), .A2(n4680), .ZN(n4682) );
  OR2_X1 U5154 ( .A1(n8904), .A2(n8591), .ZN(n8005) );
  AOI21_X1 U5155 ( .B1(n8713), .B2(n8592), .A(n4524), .ZN(n8697) );
  NOR2_X1 U5156 ( .A1(n8904), .A2(n8740), .ZN(n4524) );
  NAND2_X1 U5157 ( .A1(n8697), .A2(n8706), .ZN(n8696) );
  INV_X1 U5158 ( .A(n8689), .ZN(n8726) );
  AND2_X1 U5159 ( .A1(n8783), .A2(n8769), .ZN(n8746) );
  INV_X1 U5160 ( .A(n8592), .ZN(n8721) );
  NAND2_X1 U5161 ( .A1(n4807), .A2(n4805), .ZN(n8737) );
  AOI21_X1 U5162 ( .B1(n4808), .B2(n4809), .A(n4806), .ZN(n4805) );
  NAND2_X1 U5163 ( .A1(n8761), .A2(n4343), .ZN(n4671) );
  INV_X1 U5164 ( .A(n4382), .ZN(n4674) );
  INV_X1 U5165 ( .A(n4878), .ZN(n4673) );
  NAND2_X1 U5166 ( .A1(n8810), .A2(n8585), .ZN(n8782) );
  OR2_X1 U5167 ( .A1(n8930), .A2(n8822), .ZN(n8585) );
  OR2_X1 U5168 ( .A1(n8825), .A2(n8930), .ZN(n8798) );
  OR2_X1 U5169 ( .A1(n8938), .A2(n8820), .ZN(n4693) );
  NOR2_X1 U5170 ( .A1(n8833), .A2(n4536), .ZN(n4535) );
  INV_X1 U5171 ( .A(n4693), .ZN(n4536) );
  AND2_X1 U5172 ( .A1(n7982), .A2(n7981), .ZN(n8833) );
  NAND2_X1 U5173 ( .A1(n4840), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U5174 ( .A1(n7509), .A2(n4838), .ZN(n4835) );
  NAND2_X1 U5175 ( .A1(n8840), .A2(n8839), .ZN(n8838) );
  NAND2_X1 U5176 ( .A1(n7509), .A2(n4841), .ZN(n8852) );
  NAND2_X1 U5177 ( .A1(n4525), .A2(n4347), .ZN(n7505) );
  INV_X1 U5178 ( .A(n7968), .ZN(n4532) );
  NAND2_X1 U5179 ( .A1(n7459), .A2(n7968), .ZN(n7509) );
  AND2_X1 U5180 ( .A1(n7971), .A2(n7970), .ZN(n7968) );
  AND2_X1 U5181 ( .A1(n7964), .A2(n7965), .ZN(n7880) );
  OR2_X1 U5182 ( .A1(n7413), .A2(n9907), .ZN(n7479) );
  NOR2_X1 U5183 ( .A1(n7406), .A2(n7942), .ZN(n7457) );
  NAND2_X1 U5184 ( .A1(n6252), .A2(n4539), .ZN(n4538) );
  AND2_X1 U5185 ( .A1(n7000), .A2(n7083), .ZN(n7098) );
  AOI21_X1 U5186 ( .B1(n6995), .B2(n7874), .A(n7933), .ZN(n6935) );
  NAND2_X1 U5187 ( .A1(n6993), .A2(n6932), .ZN(n4675) );
  INV_X1 U5188 ( .A(n9894), .ZN(n7002) );
  NAND2_X1 U5189 ( .A1(n6887), .A2(n6886), .ZN(n9818) );
  AND2_X1 U5190 ( .A1(n7864), .A2(n7891), .ZN(n9815) );
  OR2_X1 U5191 ( .A1(n9867), .A2(n7909), .ZN(n7067) );
  AND2_X1 U5192 ( .A1(n6502), .A2(n8082), .ZN(n6871) );
  INV_X1 U5193 ( .A(n8806), .ZN(n8821) );
  INV_X1 U5194 ( .A(n7279), .ZN(n9900) );
  AND3_X1 U5195 ( .A1(n5719), .A2(n5718), .A3(n5717), .ZN(n9876) );
  NAND2_X1 U5196 ( .A1(n6118), .A2(n7865), .ZN(n9917) );
  INV_X1 U5197 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U5198 ( .A1(n6114), .A2(n6113), .ZN(n6116) );
  OR2_X1 U5199 ( .A1(n5604), .A2(n5641), .ZN(n5636) );
  INV_X1 U5200 ( .A(n4765), .ZN(n4764) );
  NAND2_X1 U5201 ( .A1(n5636), .A2(n5604), .ZN(n4762) );
  INV_X1 U5202 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5593) );
  NOR2_X1 U5203 ( .A1(n4791), .A2(n4444), .ZN(n4442) );
  AOI21_X1 U5204 ( .B1(n4790), .B2(n4789), .A(n4788), .ZN(n4787) );
  INV_X1 U5205 ( .A(n4794), .ZN(n4789) );
  INV_X1 U5206 ( .A(n5484), .ZN(n4788) );
  INV_X1 U5207 ( .A(n9020), .ZN(n4446) );
  INV_X1 U5208 ( .A(n4340), .ZN(n4779) );
  OR2_X1 U5209 ( .A1(n5207), .A2(n5206), .ZN(n5223) );
  INV_X1 U5210 ( .A(n4799), .ZN(n4798) );
  NAND2_X1 U5211 ( .A1(n4436), .A2(n4435), .ZN(n9090) );
  AOI21_X1 U5212 ( .B1(n4774), .B2(n4437), .A(n4434), .ZN(n4435) );
  NAND2_X1 U5213 ( .A1(n6645), .A2(n4437), .ZN(n4436) );
  NAND2_X1 U5214 ( .A1(n5164), .A2(n4778), .ZN(n4437) );
  AND4_X1 U5215 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n9108)
         );
  AOI22_X1 U5216 ( .A1(n6472), .A2(n6471), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6470), .ZN(n6474) );
  NOR2_X1 U5217 ( .A1(n7031), .A2(n7030), .ZN(n7146) );
  AND2_X1 U5218 ( .A1(n9692), .A2(n9691), .ZN(n9694) );
  NAND2_X1 U5219 ( .A1(n7594), .A2(n7593), .ZN(n9237) );
  OR2_X1 U5220 ( .A1(n9244), .A2(n9256), .ZN(n9245) );
  AOI21_X1 U5221 ( .B1(n4322), .B2(n4862), .A(n4371), .ZN(n4632) );
  OR2_X1 U5222 ( .A1(n9505), .A2(n9310), .ZN(n9282) );
  NAND2_X1 U5223 ( .A1(n4866), .A2(n9293), .ZN(n4862) );
  OAI21_X1 U5224 ( .B1(n9307), .B2(n9306), .A(n9226), .ZN(n9292) );
  AOI21_X1 U5225 ( .B1(n4866), .B2(n4864), .A(n4369), .ZN(n4863) );
  INV_X1 U5226 ( .A(n9205), .ZN(n4864) );
  AND2_X1 U5227 ( .A1(n7712), .A2(n9223), .ZN(n9344) );
  AOI21_X1 U5228 ( .B1(n4623), .B2(n4622), .A(n4375), .ZN(n4621) );
  INV_X1 U5229 ( .A(n4872), .ZN(n4622) );
  NAND2_X1 U5230 ( .A1(n9528), .A2(n9394), .ZN(n4872) );
  AND2_X1 U5231 ( .A1(n9399), .A2(n9216), .ZN(n9415) );
  INV_X1 U5232 ( .A(n9196), .ZN(n9437) );
  NAND2_X1 U5233 ( .A1(n4654), .A2(n9212), .ZN(n4653) );
  NAND2_X1 U5234 ( .A1(n7356), .A2(n7321), .ZN(n7337) );
  AOI21_X1 U5235 ( .B1(n7136), .B2(n7646), .A(n7135), .ZN(n7677) );
  AOI21_X1 U5236 ( .B1(n7547), .B2(n7043), .A(n4363), .ZN(n4875) );
  OR2_X1 U5237 ( .A1(n6902), .A2(n7547), .ZN(n7044) );
  INV_X1 U5238 ( .A(n7597), .ZN(n5397) );
  INV_X1 U5239 ( .A(n6210), .ZN(n5396) );
  NAND2_X1 U5240 ( .A1(n9742), .A2(n4334), .ZN(n6913) );
  NAND2_X1 U5241 ( .A1(n4641), .A2(n7532), .ZN(n6807) );
  NOR2_X1 U5242 ( .A1(n6785), .A2(n4642), .ZN(n4640) );
  INV_X1 U5243 ( .A(n6657), .ZN(n4642) );
  NAND2_X1 U5244 ( .A1(n6758), .A2(n6657), .ZN(n7636) );
  INV_X1 U5245 ( .A(n9456), .ZN(n9440) );
  NAND2_X1 U5246 ( .A1(n6176), .A2(n6175), .ZN(n9488) );
  NAND2_X1 U5247 ( .A1(n6152), .A2(n6151), .ZN(n9493) );
  AND2_X1 U5248 ( .A1(n7386), .A2(n7385), .ZN(n7390) );
  AND2_X1 U5249 ( .A1(n6284), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6208) );
  OR2_X1 U5250 ( .A1(n5539), .A2(n5541), .ZN(n6664) );
  AND2_X1 U5251 ( .A1(n6286), .A2(n6208), .ZN(n6240) );
  INV_X1 U5252 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5031) );
  INV_X1 U5253 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5006) );
  INV_X1 U5254 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U5255 ( .A1(n5005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U5256 ( .A1(n5011), .A2(n5010), .ZN(n5013) );
  XNOR2_X1 U5257 ( .A(n5512), .B(n5513), .ZN(n7450) );
  INV_X1 U5258 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5009) );
  OAI21_X1 U5259 ( .B1(n5425), .B2(n4732), .A(n4983), .ZN(n5448) );
  NAND2_X1 U5260 ( .A1(n5015), .A2(n5014), .ZN(n4459) );
  OR2_X1 U5261 ( .A1(n5327), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U5262 ( .A1(n5058), .A2(n5057), .ZN(n4726) );
  NAND2_X1 U5263 ( .A1(n4582), .A2(n4897), .ZN(n5126) );
  NAND2_X1 U5264 ( .A1(n4734), .A2(n4736), .ZN(n6973) );
  INV_X1 U5265 ( .A(n4737), .ZN(n4736) );
  OAI21_X1 U5266 ( .B1(n4335), .B2(n4738), .A(n5787), .ZN(n4737) );
  INV_X1 U5267 ( .A(n8394), .ZN(n6876) );
  NAND2_X1 U5268 ( .A1(n5985), .A2(n5984), .ZN(n8909) );
  NAND2_X1 U5269 ( .A1(n6016), .A2(n6015), .ZN(n8894) );
  NAND2_X1 U5270 ( .A1(n5842), .A2(n5841), .ZN(n8948) );
  INV_X1 U5271 ( .A(n8393), .ZN(n6953) );
  NAND2_X1 U5272 ( .A1(n5944), .A2(n5943), .ZN(n8923) );
  INV_X1 U5273 ( .A(n8804), .ZN(n8819) );
  OAI211_X1 U5274 ( .C1(n8682), .C2(n7824), .A(n6024), .B(n6023), .ZN(n8708)
         );
  NAND2_X1 U5275 ( .A1(n8562), .A2(n9804), .ZN(n4413) );
  OR2_X1 U5276 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  NAND2_X1 U5277 ( .A1(n4376), .A2(n5664), .ZN(n6713) );
  INV_X1 U5278 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8974) );
  AND2_X1 U5279 ( .A1(n6179), .A2(n5575), .ZN(n9267) );
  AND4_X2 U5280 ( .A1(n5098), .A2(n5097), .A3(n5096), .A4(n5095), .ZN(n6674)
         );
  NAND2_X1 U5281 ( .A1(n5393), .A2(n9080), .ZN(n8070) );
  OR2_X1 U5282 ( .A1(n6193), .A2(n9117), .ZN(n4769) );
  NAND2_X1 U5283 ( .A1(n8991), .A2(n6167), .ZN(n4770) );
  AOI21_X1 U5284 ( .B1(n9065), .B2(n9061), .A(n9063), .ZN(n9023) );
  OR2_X1 U5285 ( .A1(n5264), .A2(n5263), .ZN(n4882) );
  AND4_X1 U5286 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n9048)
         );
  AND4_X1 U5287 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n7214)
         );
  AND4_X1 U5288 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n9309)
         );
  AND4_X1 U5289 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n7225)
         );
  INV_X1 U5290 ( .A(n9402), .ZN(n9199) );
  AND2_X1 U5291 ( .A1(n5176), .A2(n4383), .ZN(n4612) );
  NAND2_X1 U5292 ( .A1(n7754), .A2(n7383), .ZN(n4694) );
  INV_X1 U5293 ( .A(n9309), .ZN(n9345) );
  INV_X1 U5294 ( .A(n9108), .ZN(n9424) );
  INV_X1 U5295 ( .A(n7225), .ZN(n9123) );
  INV_X1 U5296 ( .A(n7045), .ZN(n9127) );
  NAND2_X1 U5297 ( .A1(n5094), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U5298 ( .A1(n5077), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5082) );
  AOI21_X1 U5299 ( .B1(n5093), .B2(P1_REG1_REG_0__SCAN_IN), .A(n4318), .ZN(
        n4660) );
  NAND2_X1 U5300 ( .A1(n4637), .A2(n4635), .ZN(n9485) );
  AOI21_X1 U5301 ( .B1(n9273), .B2(n9454), .A(n4636), .ZN(n4635) );
  OR2_X1 U5302 ( .A1(n4638), .A2(n9436), .ZN(n4637) );
  NOR2_X1 U5303 ( .A1(n9234), .A2(n9233), .ZN(n4636) );
  AND2_X1 U5304 ( .A1(n4407), .A2(n4406), .ZN(n9491) );
  AOI22_X1 U5305 ( .A1(n9286), .A2(n9454), .B1(n9258), .B2(n9456), .ZN(n4406)
         );
  NAND2_X1 U5306 ( .A1(n9259), .A2(n9459), .ZN(n4407) );
  AOI21_X1 U5307 ( .B1(n9274), .B2(n9459), .A(n4404), .ZN(n9496) );
  INV_X1 U5308 ( .A(n4405), .ZN(n4404) );
  AOI22_X1 U5309 ( .A1(n9273), .A2(n9456), .B1(n9454), .B2(n9272), .ZN(n4405)
         );
  INV_X1 U5310 ( .A(n9493), .ZN(n9269) );
  NAND2_X1 U5311 ( .A1(n9460), .A2(n6679), .ZN(n9467) );
  AND2_X1 U5312 ( .A1(n9460), .A2(n6680), .ZN(n9429) );
  OAI21_X1 U5313 ( .B1(n7910), .B2(n7911), .A(n4661), .ZN(n7912) );
  NAND2_X1 U5314 ( .A1(n4592), .A2(n7676), .ZN(n4591) );
  OAI21_X1 U5315 ( .B1(n7674), .B2(n7673), .A(n4593), .ZN(n4592) );
  AND2_X1 U5316 ( .A1(n7671), .A2(n7672), .ZN(n4593) );
  OAI21_X1 U5317 ( .B1(n7677), .B2(n4589), .A(n4657), .ZN(n4587) );
  OAI21_X1 U5318 ( .B1(n7688), .B2(n4589), .A(n7690), .ZN(n4611) );
  AOI21_X1 U5319 ( .B1(n7680), .B2(n7679), .A(n7682), .ZN(n4609) );
  NOR2_X1 U5320 ( .A1(n7703), .A2(n4589), .ZN(n4595) );
  OR2_X1 U5321 ( .A1(n9366), .A2(n9217), .ZN(n4596) );
  AOI21_X1 U5322 ( .B1(n7697), .B2(n9415), .A(n7696), .ZN(n4600) );
  NOR2_X1 U5323 ( .A1(n9221), .A2(n7740), .ZN(n4598) );
  NAND2_X1 U5324 ( .A1(n4597), .A2(n4594), .ZN(n7708) );
  OAI21_X1 U5325 ( .B1(n4600), .B2(n4599), .A(n4598), .ZN(n4597) );
  OAI21_X1 U5326 ( .B1(n4600), .B2(n4596), .A(n4595), .ZN(n4594) );
  NAND2_X1 U5327 ( .A1(n7699), .A2(n7698), .ZN(n4599) );
  NAND2_X1 U5328 ( .A1(n9226), .A2(n9282), .ZN(n4718) );
  AOI21_X1 U5329 ( .B1(n4585), .B2(n7712), .A(n4719), .ZN(n4584) );
  NAND2_X1 U5330 ( .A1(n9227), .A2(n4720), .ZN(n4719) );
  OAI21_X1 U5331 ( .B1(n7711), .B2(n9222), .A(n7710), .ZN(n4585) );
  NOR2_X1 U5332 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  INV_X1 U5333 ( .A(n7729), .ZN(n4607) );
  NAND2_X1 U5334 ( .A1(n4606), .A2(n4605), .ZN(n4604) );
  NOR2_X1 U5335 ( .A1(n9281), .A2(n7740), .ZN(n4605) );
  NAND2_X1 U5336 ( .A1(n7724), .A2(n7725), .ZN(n4606) );
  NAND2_X1 U5337 ( .A1(n4603), .A2(n4350), .ZN(n4602) );
  NAND2_X1 U5338 ( .A1(n7726), .A2(n7725), .ZN(n4603) );
  INV_X1 U5339 ( .A(n8109), .ZN(n4744) );
  INV_X1 U5340 ( .A(SI_16_), .ZN(n8251) );
  INV_X1 U5341 ( .A(SI_19_), .ZN(n8237) );
  NOR2_X1 U5342 ( .A1(n7087), .A2(n4850), .ZN(n4849) );
  NOR2_X1 U5343 ( .A1(n5647), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5645) );
  INV_X1 U5344 ( .A(n5361), .ZN(n4453) );
  OAI21_X1 U5345 ( .B1(n7751), .B2(n9258), .A(n7738), .ZN(n7747) );
  NOR2_X1 U5346 ( .A1(n9510), .A2(n9513), .ZN(n4574) );
  INV_X1 U5347 ( .A(n5322), .ZN(n4713) );
  NAND2_X1 U5348 ( .A1(n4706), .A2(n4933), .ZN(n4705) );
  INV_X1 U5349 ( .A(n5265), .ZN(n4706) );
  INV_X1 U5350 ( .A(n5057), .ZN(n4618) );
  AND2_X1 U5351 ( .A1(n4724), .A2(n4616), .ZN(n4615) );
  NOR2_X1 U5352 ( .A1(n5192), .A2(n4725), .ZN(n4724) );
  INV_X1 U5353 ( .A(n4911), .ZN(n4725) );
  NAND2_X1 U5354 ( .A1(n4499), .A2(n4326), .ZN(n6012) );
  INV_X1 U5355 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5807) );
  INV_X1 U5356 ( .A(SI_21_), .ZN(n8297) );
  INV_X1 U5357 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U5358 ( .A1(n6981), .A2(n4415), .ZN(n8504) );
  OR2_X1 U5359 ( .A1(n6982), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4415) );
  OR2_X1 U5360 ( .A1(n8886), .A2(n8594), .ZN(n8020) );
  AND2_X1 U5361 ( .A1(n4679), .A2(n4680), .ZN(n4678) );
  NAND2_X1 U5362 ( .A1(n8790), .A2(n7997), .ZN(n8763) );
  OR2_X1 U5363 ( .A1(n5808), .A2(n5807), .ZN(n5827) );
  NAND2_X1 U5364 ( .A1(n9900), .A2(n8211), .ZN(n7900) );
  NAND2_X1 U5365 ( .A1(n7091), .A2(n4849), .ZN(n4848) );
  NAND2_X1 U5366 ( .A1(n6870), .A2(n9830), .ZN(n7904) );
  NAND2_X1 U5367 ( .A1(n4409), .A2(n4548), .ZN(n4543) );
  OR2_X1 U5368 ( .A1(n5645), .A2(n4550), .ZN(n4549) );
  NAND2_X1 U5369 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n4550) );
  NAND2_X1 U5370 ( .A1(n8812), .A2(n8811), .ZN(n8810) );
  NOR2_X1 U5371 ( .A1(n9854), .A2(n6954), .ZN(n7009) );
  AND2_X1 U5372 ( .A1(n5645), .A2(n5646), .ZN(n4547) );
  AND2_X1 U5373 ( .A1(n4549), .A2(n4548), .ZN(n4477) );
  INV_X1 U5374 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4855) );
  OR2_X1 U5375 ( .A1(n9009), .A2(n9010), .ZN(n4794) );
  OR2_X1 U5376 ( .A1(n5183), .A2(n5184), .ZN(n4799) );
  NOR2_X1 U5377 ( .A1(n4780), .A2(n4775), .ZN(n4774) );
  NOR2_X1 U5378 ( .A1(n4779), .A2(n6826), .ZN(n4775) );
  AOI21_X1 U5379 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n6856), .A(n6855), .ZN(
        n7029) );
  OR2_X1 U5380 ( .A1(n9498), .A2(n9272), .ZN(n9210) );
  NOR2_X1 U5381 ( .A1(n4573), .A2(n9505), .ZN(n4572) );
  INV_X1 U5382 ( .A(n4574), .ZN(n4573) );
  NAND2_X1 U5383 ( .A1(n7781), .A2(n7713), .ZN(n9226) );
  OR2_X1 U5384 ( .A1(n5368), .A2(n5367), .ZN(n5385) );
  OR2_X1 U5385 ( .A1(n4339), .A2(n7222), .ZN(n4869) );
  NOR2_X1 U5386 ( .A1(n7046), .A2(n4647), .ZN(n4646) );
  INV_X1 U5387 ( .A(n7542), .ZN(n4647) );
  AND2_X1 U5388 ( .A1(n7671), .A2(n7768), .ZN(n4649) );
  NAND2_X1 U5389 ( .A1(n9337), .A2(n4574), .ZN(n9311) );
  OR2_X1 U5390 ( .A1(n9382), .A2(n9528), .ZN(n9373) );
  AND2_X1 U5391 ( .A1(n7580), .A2(n7579), .ZN(n7595) );
  AND2_X1 U5392 ( .A1(n7574), .A2(n7573), .ZN(n7591) );
  AND2_X1 U5393 ( .A1(n6170), .A2(n6065), .ZN(n6168) );
  AND2_X1 U5394 ( .A1(n6060), .A2(n5518), .ZN(n6058) );
  AND2_X1 U5395 ( .A1(n4980), .A2(n4979), .ZN(n5409) );
  NAND2_X1 U5396 ( .A1(n5175), .A2(n5174), .ZN(n4909) );
  NAND2_X1 U5397 ( .A1(n6214), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4400) );
  INV_X1 U5398 ( .A(n8640), .ZN(n8594) );
  INV_X1 U5399 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5893) );
  AND2_X1 U5400 ( .A1(n5906), .A2(n4757), .ZN(n4753) );
  OR2_X1 U5401 ( .A1(n5887), .A2(n5886), .ZN(n4757) );
  NAND2_X1 U5402 ( .A1(n4756), .A2(n4755), .ZN(n4754) );
  AOI21_X1 U5403 ( .B1(n4515), .B2(n4513), .A(n4512), .ZN(n4511) );
  INV_X1 U5404 ( .A(n5821), .ZN(n4512) );
  INV_X1 U5405 ( .A(n6972), .ZN(n4513) );
  OR2_X1 U5406 ( .A1(n6845), .A2(n4739), .ZN(n4738) );
  INV_X1 U5407 ( .A(n5766), .ZN(n4739) );
  INV_X1 U5408 ( .A(n4738), .ZN(n4735) );
  AOI21_X1 U5409 ( .B1(n4493), .B2(n4495), .A(n4374), .ZN(n4490) );
  OR2_X1 U5410 ( .A1(n5999), .A2(n8165), .ZN(n6007) );
  NAND2_X1 U5411 ( .A1(n8163), .A2(n8162), .ZN(n8161) );
  NAND2_X1 U5412 ( .A1(n6139), .A2(n6509), .ZN(n7066) );
  NAND2_X1 U5413 ( .A1(n4740), .A2(n4335), .ZN(n6837) );
  OR2_X1 U5414 ( .A1(n5894), .A2(n5893), .ZN(n5915) );
  INV_X1 U5415 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5914) );
  OR2_X1 U5416 ( .A1(n5915), .A2(n5914), .ZN(n5917) );
  NAND2_X1 U5417 ( .A1(n7435), .A2(n4496), .ZN(n4492) );
  INV_X1 U5418 ( .A(n9850), .ZN(n7865) );
  NAND2_X1 U5419 ( .A1(n4377), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6092) );
  NOR2_X1 U5420 ( .A1(n9604), .A2(n4416), .ZN(n9603) );
  NAND2_X1 U5421 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n4416) );
  NOR2_X1 U5422 ( .A1(n8404), .A2(n8403), .ZN(n8402) );
  NOR2_X1 U5423 ( .A1(n8430), .A2(n8431), .ZN(n8429) );
  AND2_X1 U5424 ( .A1(n8482), .A2(n8483), .ZN(n8480) );
  NOR2_X1 U5425 ( .A1(n6526), .A2(n6525), .ZN(n6601) );
  OR2_X1 U5426 ( .A1(n8496), .A2(n8495), .ZN(n8498) );
  NAND2_X1 U5427 ( .A1(n6729), .A2(n6730), .ZN(n6981) );
  INV_X1 U5428 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U5429 ( .A1(n8510), .A2(n8509), .ZN(n8531) );
  NAND2_X1 U5430 ( .A1(n8531), .A2(n4410), .ZN(n8534) );
  NAND2_X1 U5431 ( .A1(n8518), .A2(n8508), .ZN(n4410) );
  NAND2_X1 U5432 ( .A1(n4553), .A2(n8869), .ZN(n4552) );
  NOR2_X1 U5433 ( .A1(n8655), .A2(n4551), .ZN(n8620) );
  INV_X1 U5434 ( .A(n4553), .ZN(n4551) );
  OR2_X1 U5435 ( .A1(n8655), .A2(n4554), .ZN(n8630) );
  AND2_X1 U5436 ( .A1(n6071), .A2(n6048), .ZN(n8656) );
  NOR2_X1 U5437 ( .A1(n8698), .A2(n8894), .ZN(n8681) );
  NAND2_X1 U5438 ( .A1(n8746), .A2(n4560), .ZN(n8698) );
  NOR2_X1 U5439 ( .A1(n8899), .A2(n4562), .ZN(n4560) );
  NAND2_X1 U5440 ( .A1(n4671), .A2(n4668), .ZN(n8590) );
  NOR2_X1 U5441 ( .A1(n4337), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U5442 ( .A1(n4881), .A2(n4670), .ZN(n4669) );
  NAND2_X1 U5443 ( .A1(n4378), .A2(n8001), .ZN(n4808) );
  NAND2_X1 U5444 ( .A1(n8764), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U5445 ( .A1(n8764), .A2(n8001), .ZN(n4809) );
  NAND2_X1 U5446 ( .A1(n8763), .A2(n8764), .ZN(n8762) );
  NAND2_X1 U5447 ( .A1(n8746), .A2(n8752), .ZN(n8747) );
  OR2_X1 U5448 ( .A1(n5946), .A2(n5945), .ZN(n5957) );
  AND2_X1 U5449 ( .A1(n7989), .A2(n7997), .ZN(n8791) );
  NAND2_X1 U5450 ( .A1(n4831), .A2(n4829), .ZN(n8801) );
  AOI21_X1 U5451 ( .B1(n4832), .B2(n4834), .A(n4830), .ZN(n4829) );
  INV_X1 U5452 ( .A(n7982), .ZN(n4830) );
  AND2_X1 U5453 ( .A1(n7495), .A2(n4555), .ZN(n8842) );
  NOR2_X1 U5454 ( .A1(n8938), .A2(n4556), .ZN(n4555) );
  INV_X1 U5455 ( .A(n4557), .ZN(n4556) );
  AND2_X1 U5456 ( .A1(n8850), .A2(n7974), .ZN(n8582) );
  NAND2_X1 U5457 ( .A1(n7495), .A2(n9916), .ZN(n7494) );
  INV_X1 U5458 ( .A(n8206), .ZN(n7506) );
  NOR2_X1 U5459 ( .A1(n7479), .A2(n8948), .ZN(n7495) );
  NAND2_X1 U5460 ( .A1(n4691), .A2(n7402), .ZN(n4686) );
  NOR2_X1 U5461 ( .A1(n4689), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U5462 ( .A1(n4844), .A2(n4842), .ZN(n7406) );
  AOI21_X1 U5463 ( .B1(n4845), .B2(n4847), .A(n4843), .ZN(n4842) );
  INV_X1 U5464 ( .A(n7946), .ZN(n4843) );
  NAND2_X1 U5465 ( .A1(n7098), .A2(n9900), .ZN(n7291) );
  OR2_X1 U5466 ( .A1(n7291), .A2(n7394), .ZN(n7413) );
  NAND2_X1 U5467 ( .A1(n7281), .A2(n4690), .ZN(n7403) );
  AND2_X1 U5468 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  NAND2_X1 U5469 ( .A1(n7088), .A2(n7087), .ZN(n7281) );
  AND2_X1 U5470 ( .A1(n7951), .A2(n7937), .ZN(n7931) );
  NAND2_X1 U5471 ( .A1(n4803), .A2(n4802), .ZN(n6995) );
  NAND2_X1 U5472 ( .A1(n6928), .A2(n7926), .ZN(n4802) );
  NOR2_X1 U5473 ( .A1(n7001), .A2(n7002), .ZN(n7000) );
  NAND2_X1 U5474 ( .A1(n4542), .A2(n4541), .ZN(n7001) );
  NOR2_X1 U5475 ( .A1(n9830), .A2(n9885), .ZN(n4541) );
  INV_X1 U5476 ( .A(n9826), .ZN(n4542) );
  AND3_X1 U5477 ( .A1(n5739), .A2(n5738), .A3(n5737), .ZN(n6930) );
  NAND2_X1 U5478 ( .A1(n7903), .A2(n7869), .ZN(n9820) );
  AND2_X1 U5479 ( .A1(n7920), .A2(n7921), .ZN(n4663) );
  OR2_X1 U5480 ( .A1(n7859), .A2(n6216), .ZN(n5665) );
  INV_X1 U5481 ( .A(n4665), .ZN(n6702) );
  NAND2_X1 U5482 ( .A1(n6143), .A2(n6509), .ZN(n8804) );
  NAND2_X1 U5483 ( .A1(n6142), .A2(n6509), .ZN(n8806) );
  NAND2_X1 U5484 ( .A1(n6704), .A2(n8082), .ZN(n7021) );
  NAND2_X1 U5485 ( .A1(n7813), .A2(n7812), .ZN(n8875) );
  NAND2_X1 U5486 ( .A1(n6067), .A2(n6066), .ZN(n8880) );
  NAND2_X1 U5487 ( .A1(n5653), .A2(n5652), .ZN(n8933) );
  AND3_X1 U5488 ( .A1(n5772), .A2(n5771), .A3(n5770), .ZN(n7083) );
  INV_X1 U5489 ( .A(n9915), .ZN(n9886) );
  INV_X1 U5490 ( .A(n9917), .ZN(n9868) );
  NAND2_X1 U5491 ( .A1(n6139), .A2(n7865), .ZN(n9915) );
  NAND2_X1 U5492 ( .A1(n7123), .A2(n7895), .ZN(n9850) );
  NAND2_X1 U5493 ( .A1(n7465), .A2(n9867), .ZN(n9921) );
  OR2_X1 U5494 ( .A1(n6507), .A2(n6117), .ZN(n9839) );
  OR2_X1 U5495 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  NAND2_X1 U5496 ( .A1(n5648), .A2(n5646), .ZN(n4852) );
  INV_X1 U5497 ( .A(n6084), .ZN(n6089) );
  XNOR2_X1 U5498 ( .A(n5640), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U5499 ( .A1(n5627), .A2(n5601), .ZN(n5639) );
  AND3_X1 U5500 ( .A1(n5837), .A2(n5822), .A3(n5628), .ZN(n5629) );
  NOR2_X1 U5501 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4824) );
  NAND2_X1 U5502 ( .A1(n6962), .A2(n6963), .ZN(n6961) );
  NAND2_X1 U5503 ( .A1(n4425), .A2(n4428), .ZN(n8998) );
  AND2_X1 U5504 ( .A1(n4429), .A2(n5320), .ZN(n4428) );
  OR2_X1 U5505 ( .A1(n4320), .A2(n4430), .ZN(n4429) );
  NAND2_X1 U5506 ( .A1(n4336), .A2(n5321), .ZN(n8999) );
  INV_X1 U5507 ( .A(n5508), .ZN(n6188) );
  NAND2_X1 U5508 ( .A1(n9009), .A2(n9010), .ZN(n4793) );
  NAND2_X1 U5509 ( .A1(n9013), .A2(n4794), .ZN(n4792) );
  AND2_X1 U5510 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  INV_X1 U5511 ( .A(n9510), .ZN(n9206) );
  INV_X1 U5512 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U5513 ( .A1(n4433), .A2(n4320), .ZN(n7422) );
  OR2_X1 U5514 ( .A1(n5288), .A2(n5287), .ZN(n5312) );
  OR2_X1 U5515 ( .A1(n5223), .A2(n6401), .ZN(n5252) );
  OAI21_X1 U5516 ( .B1(n6482), .B2(n6481), .A(n6484), .ZN(n6483) );
  AND2_X1 U5517 ( .A1(n4449), .A2(n4388), .ZN(n9081) );
  NOR2_X1 U5518 ( .A1(n4454), .A2(n5392), .ZN(n4450) );
  NOR2_X1 U5519 ( .A1(n5312), .A2(n9002), .ZN(n5331) );
  OR2_X1 U5520 ( .A1(n9476), .A2(n9188), .ZN(n7790) );
  INV_X1 U5521 ( .A(n4697), .ZN(n7757) );
  AND4_X1 U5522 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n6832)
         );
  NOR2_X1 U5523 ( .A1(n6439), .A2(n6438), .ZN(n6437) );
  NOR2_X1 U5524 ( .A1(n6354), .A2(n6355), .ZN(n6353) );
  INV_X1 U5525 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9084) );
  AND3_X1 U5526 ( .A1(n7604), .A2(n7603), .A3(n7602), .ZN(n9233) );
  XNOR2_X1 U5527 ( .A(n4639), .B(n9232), .ZN(n4638) );
  NAND2_X1 U5528 ( .A1(n9255), .A2(n9230), .ZN(n4639) );
  AND2_X1 U5529 ( .A1(n7730), .A2(n9230), .ZN(n9256) );
  OR2_X1 U5530 ( .A1(n9493), .A2(n9286), .ZN(n4398) );
  AND2_X1 U5531 ( .A1(n9337), .A2(n4570), .ZN(n9278) );
  NOR2_X1 U5532 ( .A1(n9498), .A2(n4571), .ZN(n4570) );
  INV_X1 U5533 ( .A(n4572), .ZN(n4571) );
  AND4_X1 U5534 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n9330)
         );
  NAND2_X1 U5535 ( .A1(n9337), .A2(n9326), .ZN(n9321) );
  AOI21_X1 U5536 ( .B1(n9354), .B2(n9353), .A(n9222), .ZN(n9343) );
  AND2_X1 U5537 ( .A1(n9358), .A2(n9341), .ZN(n9337) );
  AND2_X1 U5538 ( .A1(n5413), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5428) );
  AND2_X1 U5539 ( .A1(n9220), .A2(n7701), .ZN(n9368) );
  NAND2_X1 U5540 ( .A1(n9421), .A2(n9439), .ZN(n4417) );
  AND2_X1 U5541 ( .A1(n4323), .A2(n9216), .ZN(n4651) );
  NAND2_X1 U5542 ( .A1(n4567), .A2(n4325), .ZN(n9441) );
  NAND2_X1 U5543 ( .A1(n4567), .A2(n4566), .ZN(n9443) );
  NOR2_X1 U5544 ( .A1(n7366), .A2(n4568), .ZN(n7343) );
  NAND2_X1 U5545 ( .A1(n5286), .A2(n5285), .ZN(n7421) );
  NOR2_X1 U5546 ( .A1(n7366), .A2(n7421), .ZN(n7367) );
  INV_X1 U5547 ( .A(n7310), .ZN(n7553) );
  AND2_X1 U5548 ( .A1(n7675), .A2(n7625), .ZN(n7552) );
  AND4_X1 U5549 ( .A1(n5212), .A2(n5211), .A3(n5210), .A4(n5209), .ZN(n7239)
         );
  NAND2_X1 U5550 ( .A1(n4645), .A2(n4649), .ZN(n7134) );
  NAND2_X1 U5551 ( .A1(n4648), .A2(n4646), .ZN(n4645) );
  NOR2_X1 U5552 ( .A1(n7052), .A2(n7127), .ZN(n7246) );
  NAND2_X1 U5553 ( .A1(n4648), .A2(n7542), .ZN(n7770) );
  NAND2_X1 U5554 ( .A1(n6786), .A2(n7541), .ZN(n6917) );
  AND4_X1 U5555 ( .A1(n5053), .A2(n5052), .A3(n5051), .A4(n5050), .ZN(n9095)
         );
  NAND2_X1 U5556 ( .A1(n6798), .A2(n6797), .ZN(n9471) );
  NAND2_X1 U5557 ( .A1(n6807), .A2(n7538), .ZN(n9452) );
  OR2_X1 U5558 ( .A1(n6815), .A2(n6819), .ZN(n9463) );
  NOR2_X1 U5559 ( .A1(n6762), .A2(n6768), .ZN(n6763) );
  INV_X1 U5560 ( .A(n7535), .ZN(n4402) );
  INV_X1 U5561 ( .A(n6756), .ZN(n4403) );
  OR2_X1 U5562 ( .A1(n5404), .A2(n5116), .ZN(n5120) );
  INV_X1 U5563 ( .A(n6491), .ZN(n6746) );
  NAND2_X1 U5564 ( .A1(n7599), .A2(n7598), .ZN(n9480) );
  AND2_X1 U5565 ( .A1(n5205), .A2(n5204), .ZN(n9774) );
  OR2_X1 U5566 ( .A1(n9561), .A2(n5568), .ZN(n9773) );
  AND2_X1 U5567 ( .A1(n7568), .A2(n6174), .ZN(n7566) );
  XNOR2_X1 U5568 ( .A(n6169), .B(n6168), .ZN(n8984) );
  AOI21_X1 U5569 ( .B1(n4730), .B2(n4732), .A(n4729), .ZN(n4728) );
  INV_X1 U5570 ( .A(n5446), .ZN(n4729) );
  AND2_X1 U5571 ( .A1(n5465), .A2(n5452), .ZN(n5463) );
  XNOR2_X1 U5572 ( .A(n5558), .B(n5557), .ZN(n6284) );
  OR2_X1 U5573 ( .A1(n5021), .A2(n5020), .ZN(n5022) );
  NAND2_X1 U5574 ( .A1(n4458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5024) );
  NOR2_X1 U5575 ( .A1(n4457), .A2(n4801), .ZN(n4456) );
  INV_X1 U5576 ( .A(n5015), .ZN(n4457) );
  NAND2_X1 U5577 ( .A1(n4709), .A2(n4951), .ZN(n5323) );
  NAND2_X1 U5578 ( .A1(n4948), .A2(n4714), .ZN(n4709) );
  NAND2_X1 U5579 ( .A1(n4702), .A2(n4933), .ZN(n5266) );
  NAND2_X1 U5580 ( .A1(n4930), .A2(n4707), .ZN(n4702) );
  AND2_X1 U5581 ( .A1(n5250), .A2(n5284), .ZN(n6470) );
  AND2_X1 U5582 ( .A1(n5202), .A2(n4991), .ZN(n5218) );
  OR2_X1 U5583 ( .A1(n4783), .A2(n5054), .ZN(n5194) );
  NAND2_X1 U5584 ( .A1(n4909), .A2(n4908), .ZN(n5058) );
  NAND2_X1 U5585 ( .A1(n4583), .A2(n4894), .ZN(n5103) );
  NAND2_X1 U5586 ( .A1(n6837), .A2(n5766), .ZN(n6846) );
  NAND2_X1 U5587 ( .A1(n4754), .A2(n4757), .ZN(n7521) );
  NAND2_X1 U5588 ( .A1(n5892), .A2(n5891), .ZN(n8581) );
  NAND2_X1 U5589 ( .A1(n4510), .A2(n4511), .ZN(n7106) );
  OR2_X1 U5590 ( .A1(n6973), .A2(n4514), .ZN(n4510) );
  NAND2_X1 U5591 ( .A1(n4465), .A2(n4469), .ZN(n6589) );
  INV_X1 U5592 ( .A(n6555), .ZN(n4471) );
  AND2_X1 U5593 ( .A1(n4505), .A2(n4345), .ZN(n8103) );
  INV_X1 U5594 ( .A(n8210), .ZN(n7407) );
  AND2_X1 U5595 ( .A1(n5681), .A2(n5669), .ZN(n6498) );
  INV_X1 U5596 ( .A(n5667), .ZN(n4460) );
  NAND2_X1 U5597 ( .A1(n8101), .A2(n4745), .ZN(n4749) );
  NAND2_X1 U5598 ( .A1(n4761), .A2(n5852), .ZN(n7437) );
  NAND2_X1 U5599 ( .A1(n6028), .A2(n6027), .ZN(n8119) );
  NAND2_X1 U5600 ( .A1(n4484), .A2(n4485), .ZN(n6026) );
  OAI211_X1 U5601 ( .C1(n4466), .C2(n4463), .A(n5732), .B(n4461), .ZN(n6636)
         );
  INV_X1 U5602 ( .A(n4758), .ZN(n4463) );
  NAND2_X1 U5603 ( .A1(n4462), .A2(n4758), .ZN(n4461) );
  NAND2_X1 U5604 ( .A1(n4478), .A2(n4482), .ZN(n8147) );
  AND2_X1 U5605 ( .A1(n4483), .A2(n4479), .ZN(n4478) );
  INV_X1 U5606 ( .A(n9876), .ZN(n9830) );
  NAND2_X1 U5607 ( .A1(n4759), .A2(n5714), .ZN(n6630) );
  AND2_X1 U5608 ( .A1(n4517), .A2(n4518), .ZN(n7114) );
  NAND2_X1 U5609 ( .A1(n6973), .A2(n6972), .ZN(n4517) );
  AND2_X1 U5610 ( .A1(n8101), .A2(n5970), .ZN(n8154) );
  NAND2_X1 U5611 ( .A1(n7435), .A2(n5873), .ZN(n7444) );
  NAND2_X1 U5612 ( .A1(n5876), .A2(n5875), .ZN(n8943) );
  NAND2_X1 U5613 ( .A1(n4507), .A2(n4506), .ZN(n7274) );
  AOI21_X1 U5614 ( .B1(n4508), .B2(n4514), .A(n4372), .ZN(n4506) );
  INV_X1 U5615 ( .A(n8175), .ZN(n8167) );
  INV_X1 U5616 ( .A(n8174), .ZN(n8166) );
  AND3_X1 U5617 ( .A1(n5755), .A2(n5754), .A3(n5753), .ZN(n9894) );
  INV_X1 U5618 ( .A(n8204), .ZN(n8180) );
  INV_X1 U5619 ( .A(n8191), .ZN(n8202) );
  NAND2_X1 U5620 ( .A1(n4818), .A2(n8807), .ZN(n4817) );
  XNOR2_X1 U5621 ( .A(n6092), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U5622 ( .A1(n6078), .A2(n6077), .ZN(n8619) );
  NAND4_X1 U5623 ( .A1(n5710), .A2(n5709), .A3(n5708), .A4(n5707), .ZN(n8393)
         );
  NAND3_X1 U5624 ( .A1(n5696), .A2(n5695), .A3(n5694), .ZN(n8394) );
  AND2_X1 U5625 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  OR2_X1 U5626 ( .A1(n5843), .A2(n5671), .ZN(n5675) );
  OR2_X1 U5627 ( .A1(n7854), .A2(n9925), .ZN(n5674) );
  INV_X2 U5628 ( .A(P2_U3966), .ZN(n8395) );
  OR2_X1 U5629 ( .A1(n8456), .A2(n8455), .ZN(n8458) );
  NAND2_X1 U5630 ( .A1(n8458), .A2(n6519), .ZN(n8469) );
  OAI21_X1 U5631 ( .B1(n5928), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5942) );
  AOI21_X1 U5632 ( .B1(n4423), .B2(n8824), .A(n4420), .ZN(n8878) );
  NAND2_X1 U5633 ( .A1(n4422), .A2(n4421), .ZN(n4420) );
  XNOR2_X1 U5634 ( .A(n8617), .B(n8616), .ZN(n4423) );
  NAND2_X1 U5635 ( .A1(n8618), .A2(n8821), .ZN(n4422) );
  INV_X1 U5636 ( .A(n8886), .ZN(n8659) );
  NAND2_X1 U5637 ( .A1(n6030), .A2(n6029), .ZN(n8891) );
  AND2_X1 U5638 ( .A1(n4682), .A2(n8593), .ZN(n8663) );
  AND2_X1 U5639 ( .A1(n4828), .A2(n4338), .ZN(n8688) );
  INV_X1 U5640 ( .A(n4682), .ZN(n8679) );
  NAND2_X1 U5641 ( .A1(n8696), .A2(n4683), .ZN(n8680) );
  NAND2_X1 U5642 ( .A1(n8720), .A2(n8005), .ZN(n8705) );
  NAND2_X1 U5643 ( .A1(n8746), .A2(n4563), .ZN(n8715) );
  NOR2_X1 U5644 ( .A1(n4667), .A2(n4666), .ZN(n8732) );
  OR2_X1 U5645 ( .A1(n4337), .A2(n8589), .ZN(n4666) );
  INV_X1 U5646 ( .A(n4671), .ZN(n4667) );
  OAI21_X1 U5647 ( .B1(n4672), .B2(n4382), .A(n4878), .ZN(n8745) );
  INV_X1 U5648 ( .A(n8761), .ZN(n4672) );
  NAND2_X1 U5649 ( .A1(n5966), .A2(n5965), .ZN(n8920) );
  NAND2_X1 U5650 ( .A1(n5931), .A2(n5930), .ZN(n8930) );
  AND2_X1 U5651 ( .A1(n8838), .A2(n4535), .ZN(n8831) );
  NAND2_X1 U5652 ( .A1(n8838), .A2(n4693), .ZN(n8832) );
  AND2_X1 U5653 ( .A1(n4835), .A2(n4833), .ZN(n8818) );
  NAND2_X1 U5654 ( .A1(n4835), .A2(n4836), .ZN(n8851) );
  NAND2_X1 U5655 ( .A1(n4525), .A2(n4526), .ZN(n7463) );
  NAND2_X1 U5656 ( .A1(n4531), .A2(n7462), .ZN(n7488) );
  NAND2_X1 U5657 ( .A1(n7476), .A2(n7877), .ZN(n4531) );
  NAND2_X1 U5658 ( .A1(n5826), .A2(n5825), .ZN(n9907) );
  NAND2_X1 U5659 ( .A1(n5792), .A2(n4359), .ZN(n7279) );
  NAND2_X1 U5660 ( .A1(n4804), .A2(n6888), .ZN(n6934) );
  INV_X2 U5661 ( .A(n4316), .ZN(n8846) );
  OR2_X1 U5662 ( .A1(n6710), .A2(n5678), .ZN(n9833) );
  INV_X1 U5663 ( .A(n9831), .ZN(n8848) );
  OR2_X1 U5664 ( .A1(n7067), .A2(n9839), .ZN(n9827) );
  INV_X2 U5665 ( .A(n9937), .ZN(n9939) );
  AND2_X1 U5666 ( .A1(n6127), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9847) );
  CLKBUF_X1 U5667 ( .A(n6141), .Z(n6142) );
  XNOR2_X1 U5668 ( .A(n6095), .B(n6094), .ZN(n7355) );
  NAND2_X1 U5669 ( .A1(n6116), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  INV_X1 U5670 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7258) );
  INV_X1 U5671 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7125) );
  INV_X1 U5672 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7063) );
  INV_X1 U5673 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5637) );
  OAI21_X1 U5674 ( .B1(n5928), .B2(n4763), .A(n4762), .ZN(n5638) );
  NAND2_X1 U5675 ( .A1(n5636), .A2(n4764), .ZN(n4763) );
  INV_X1 U5676 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8315) );
  INV_X1 U5677 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6655) );
  INV_X1 U5678 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6618) );
  INV_X1 U5679 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6614) );
  INV_X1 U5680 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6496) );
  INV_X1 U5681 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6296) );
  INV_X1 U5682 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6244) );
  OR2_X1 U5683 ( .A1(n5627), .A2(n5604), .ZN(n5789) );
  INV_X1 U5684 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6227) );
  INV_X1 U5685 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6225) );
  INV_X1 U5686 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U5687 ( .A(n5661), .B(n5660), .ZN(n9599) );
  AND4_X1 U5688 ( .A1(n5191), .A2(n5190), .A3(n5189), .A4(n5188), .ZN(n7045)
         );
  OR2_X1 U5689 ( .A1(n6234), .A2(n5104), .ZN(n4565) );
  NAND2_X1 U5690 ( .A1(n5399), .A2(n5398), .ZN(n9533) );
  NAND2_X1 U5691 ( .A1(n5427), .A2(n5426), .ZN(n9525) );
  NAND2_X1 U5692 ( .A1(n4438), .A2(n4787), .ZN(n9029) );
  NAND2_X1 U5693 ( .A1(n5341), .A2(n9105), .ZN(n9037) );
  NOR2_X1 U5694 ( .A1(n4776), .A2(n4777), .ZN(n9092) );
  NAND2_X1 U5695 ( .A1(n4773), .A2(n4772), .ZN(n4777) );
  AOI21_X1 U5696 ( .B1(n4782), .B2(n4779), .A(n6826), .ZN(n4772) );
  NAND2_X1 U5697 ( .A1(n5165), .A2(n4781), .ZN(n6825) );
  OAI21_X1 U5698 ( .B1(n9037), .B2(n9036), .A(n5361), .ZN(n9044) );
  OAI21_X1 U5699 ( .B1(n8070), .B2(n5408), .A(n8067), .ZN(n4424) );
  AND4_X1 U5700 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n7430)
         );
  NOR2_X1 U5701 ( .A1(n4431), .A2(n5280), .ZN(n7423) );
  INV_X1 U5702 ( .A(n4433), .ZN(n4431) );
  NAND2_X1 U5703 ( .A1(n5003), .A2(n5002), .ZN(n9519) );
  NAND2_X1 U5704 ( .A1(n4797), .A2(n7261), .ZN(n4796) );
  NAND2_X1 U5705 ( .A1(n5238), .A2(n4351), .ZN(n4797) );
  INV_X1 U5706 ( .A(n9678), .ZN(n9117) );
  AND2_X1 U5707 ( .A1(n5566), .A2(n5565), .ZN(n9683) );
  INV_X1 U5708 ( .A(n9056), .ZN(n9115) );
  NAND2_X1 U5709 ( .A1(n4408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5001) );
  OR2_X1 U5710 ( .A1(n5406), .A2(n5405), .ZN(n9402) );
  INV_X1 U5711 ( .A(n6832), .ZN(n9457) );
  BUF_X1 U5712 ( .A(P1_U4006), .Z(n9132) );
  CLKBUF_X1 U5713 ( .A(n5570), .Z(n9686) );
  NAND2_X1 U5714 ( .A1(n6391), .A2(n6258), .ZN(n6452) );
  NOR2_X1 U5715 ( .A1(n6266), .A2(n6267), .ZN(n6306) );
  NOR2_X1 U5716 ( .A1(n6314), .A2(n6313), .ZN(n6334) );
  AOI21_X1 U5717 ( .B1(n7153), .B2(n7148), .A(n7147), .ZN(n7150) );
  AOI21_X1 U5718 ( .B1(n9699), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9694), .ZN(
        n9167) );
  INV_X1 U5719 ( .A(n9480), .ZN(n9192) );
  OR2_X1 U5720 ( .A1(n9320), .A2(n4862), .ZN(n4634) );
  OAI21_X1 U5721 ( .B1(n9320), .B2(n4865), .A(n4863), .ZN(n9291) );
  AND2_X1 U5722 ( .A1(n4867), .A2(n4868), .ZN(n9304) );
  NAND2_X1 U5723 ( .A1(n9320), .A2(n9205), .ZN(n4867) );
  INV_X1 U5724 ( .A(n9519), .ZN(n9341) );
  OAI21_X1 U5725 ( .B1(n4873), .B2(n4624), .A(n4621), .ZN(n9336) );
  NAND2_X1 U5726 ( .A1(n4625), .A2(n4623), .ZN(n9350) );
  AND2_X1 U5727 ( .A1(n4625), .A2(n4321), .ZN(n9352) );
  NAND2_X1 U5728 ( .A1(n4873), .A2(n4872), .ZN(n4625) );
  AND2_X1 U5729 ( .A1(n4650), .A2(n4323), .ZN(n9423) );
  AOI21_X1 U5730 ( .B1(n9214), .B2(n9213), .A(n9212), .ZN(n9434) );
  NAND2_X1 U5731 ( .A1(n4650), .A2(n4653), .ZN(n9432) );
  NAND2_X1 U5732 ( .A1(n7312), .A2(n7311), .ZN(n7360) );
  INV_X1 U5733 ( .A(n7677), .ZN(n7137) );
  INV_X1 U5734 ( .A(n9774), .ZN(n7127) );
  NAND2_X1 U5735 ( .A1(n7044), .A2(n7043), .ZN(n7126) );
  NAND2_X1 U5736 ( .A1(n9742), .A2(n6802), .ZN(n6915) );
  NAND2_X1 U5737 ( .A1(n5561), .A2(n9749), .ZN(n9465) );
  INV_X1 U5738 ( .A(n9467), .ZN(n9374) );
  AND2_X2 U5739 ( .A1(n7390), .A2(n7388), .ZN(n9802) );
  INV_X1 U5740 ( .A(n9486), .ZN(n4576) );
  INV_X1 U5741 ( .A(n9485), .ZN(n4399) );
  AND2_X2 U5742 ( .A1(n7390), .A2(n7389), .ZN(n9784) );
  INV_X1 U5743 ( .A(n6208), .ZN(n6241) );
  MUX2_X1 U5744 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5035), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5037) );
  XNOR2_X1 U5745 ( .A(n7567), .B(n7566), .ZN(n9589) );
  NAND2_X1 U5746 ( .A1(n5013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U5747 ( .A1(n5013), .A2(n5012), .ZN(n7453) );
  OR2_X1 U5748 ( .A1(n5011), .A2(n5010), .ZN(n5012) );
  XNOR2_X1 U5749 ( .A(n5008), .B(n5009), .ZN(n7352) );
  INV_X1 U5750 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7255) );
  INV_X1 U5751 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7122) );
  INV_X1 U5752 ( .A(n5061), .ZN(n7121) );
  INV_X1 U5753 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8304) );
  INV_X1 U5754 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U5755 ( .A1(n5364), .A2(n5018), .ZN(n5027) );
  INV_X1 U5756 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8298) );
  INV_X1 U5757 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6561) );
  INV_X1 U5758 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6295) );
  INV_X1 U5759 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6222) );
  INV_X1 U5760 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6218) );
  INV_X1 U5761 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U5762 ( .A1(n4522), .A2(n4900), .ZN(n5142) );
  XNOR2_X1 U5763 ( .A(n5126), .B(n5125), .ZN(n6234) );
  NAND2_X1 U5764 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U5765 ( .A1(n4770), .A2(n4348), .ZN(n4768) );
  AOI21_X1 U5766 ( .B1(n5588), .B2(n5587), .A(n5586), .ZN(n5589) );
  OAI21_X1 U5767 ( .B1(n9281), .B2(n9056), .A(n5585), .ZN(n5586) );
  NOR2_X1 U5768 ( .A1(n9491), .A2(n9305), .ZN(n9260) );
  NOR2_X1 U5769 ( .A1(n9496), .A2(n9305), .ZN(n9275) );
  INV_X1 U5770 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5247) );
  AND2_X2 U5771 ( .A1(n6286), .A2(n6677), .ZN(n4333) );
  INV_X1 U5772 ( .A(n8839), .ZN(n4840) );
  CLKBUF_X3 U5773 ( .A(n4474), .Z(n4409) );
  OR2_X1 U5774 ( .A1(n8914), .A2(n8111), .ZN(n8001) );
  INV_X1 U5775 ( .A(n4624), .ZN(n4623) );
  NAND2_X1 U5776 ( .A1(n9351), .A2(n4321), .ZN(n4624) );
  OR2_X1 U5777 ( .A1(n7311), .A2(n4339), .ZN(n4317) );
  AND2_X1 U5778 ( .A1(n5078), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4318) );
  AND3_X1 U5779 ( .A1(n4718), .A2(n9227), .A3(n7740), .ZN(n4319) );
  AND2_X1 U5780 ( .A1(n4432), .A2(n7425), .ZN(n4320) );
  OR2_X1 U5781 ( .A1(n9528), .A2(n9394), .ZN(n4321) );
  INV_X1 U5782 ( .A(n9293), .ZN(n4861) );
  INV_X1 U5783 ( .A(n7877), .ZN(n4527) );
  AND2_X1 U5784 ( .A1(n4859), .A2(n9210), .ZN(n4322) );
  NAND2_X1 U5785 ( .A1(n7920), .A2(n7921), .ZN(n6947) );
  INV_X1 U5786 ( .A(n7284), .ZN(n4847) );
  INV_X1 U5787 ( .A(n5662), .ZN(n6252) );
  NAND2_X1 U5788 ( .A1(n4792), .A2(n4793), .ZN(n9052) );
  AND2_X1 U5789 ( .A1(n4653), .A2(n9215), .ZN(n4323) );
  NOR2_X1 U5790 ( .A1(n8038), .A2(n4395), .ZN(n4324) );
  NAND2_X1 U5791 ( .A1(n6006), .A2(n6005), .ZN(n8899) );
  AND2_X1 U5792 ( .A1(n4566), .A2(n4569), .ZN(n4325) );
  INV_X1 U5793 ( .A(n5164), .ZN(n4782) );
  AND2_X1 U5794 ( .A1(n4498), .A2(n4360), .ZN(n4326) );
  INV_X1 U5795 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5646) );
  INV_X1 U5796 ( .A(n9421), .ZN(n9545) );
  AND2_X1 U5797 ( .A1(n5366), .A2(n5365), .ZN(n9421) );
  OR2_X1 U5798 ( .A1(n8938), .A2(n8135), .ZN(n4327) );
  NAND2_X1 U5799 ( .A1(n7847), .A2(n8867), .ZN(n4328) );
  INV_X1 U5800 ( .A(n7547), .ZN(n6901) );
  AND2_X1 U5801 ( .A1(n6796), .A2(n6675), .ZN(n4329) );
  AND2_X1 U5802 ( .A1(n9487), .A2(n4380), .ZN(n4330) );
  INV_X1 U5803 ( .A(n7740), .ZN(n4589) );
  NAND2_X1 U5804 ( .A1(n7495), .A2(n4557), .ZN(n4331) );
  NAND2_X1 U5805 ( .A1(n9858), .A2(n6697), .ZN(n4665) );
  OR2_X1 U5806 ( .A1(n8655), .A2(n4552), .ZN(n4332) );
  NAND2_X1 U5808 ( .A1(n4630), .A2(n5251), .ZN(n9651) );
  BUF_X1 U5809 ( .A(n4333), .Z(n5229) );
  XNOR2_X1 U5810 ( .A(n5026), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5061) );
  AND2_X1 U5811 ( .A1(n4441), .A2(n4439), .ZN(n5538) );
  NAND2_X1 U5812 ( .A1(n5099), .A2(n4987), .ZN(n5054) );
  NAND2_X1 U5813 ( .A1(n7283), .A2(n7279), .ZN(n7284) );
  INV_X1 U5814 ( .A(n4469), .ZN(n4468) );
  OR2_X1 U5815 ( .A1(n5698), .A2(n5697), .ZN(n4469) );
  AND2_X1 U5816 ( .A1(n6803), .A2(n6802), .ZN(n4334) );
  AND2_X1 U5817 ( .A1(n6839), .A2(n4741), .ZN(n4335) );
  INV_X1 U5818 ( .A(n5704), .ZN(n6049) );
  INV_X1 U5819 ( .A(n9433), .ZN(n4654) );
  NAND2_X1 U5820 ( .A1(n4824), .A2(n5715), .ZN(n5735) );
  AND2_X1 U5821 ( .A1(n7422), .A2(n7424), .ZN(n4336) );
  AND2_X1 U5822 ( .A1(n8755), .A2(n4673), .ZN(n4337) );
  NAND2_X1 U5823 ( .A1(n8899), .A2(n8726), .ZN(n4338) );
  NAND2_X1 U5824 ( .A1(n7313), .A2(n7359), .ZN(n4339) );
  NAND4_X1 U5825 ( .A1(n5676), .A2(n5675), .A3(n5674), .A4(n5673), .ZN(n6502)
         );
  NAND2_X1 U5826 ( .A1(n5151), .A2(n5150), .ZN(n4340) );
  OR2_X1 U5827 ( .A1(n8894), .A2(n8708), .ZN(n8593) );
  INV_X1 U5828 ( .A(n7713), .ZN(n4722) );
  INV_X1 U5829 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U5830 ( .A1(n7919), .A2(n4665), .ZN(n6873) );
  OR2_X1 U5831 ( .A1(n6210), .A2(n6415), .ZN(n4341) );
  NAND2_X1 U5832 ( .A1(n5997), .A2(n5996), .ZN(n8904) );
  AND2_X1 U5833 ( .A1(n4547), .A2(n8985), .ZN(n4342) );
  INV_X1 U5834 ( .A(n8880), .ZN(n8636) );
  NAND2_X1 U5835 ( .A1(n5442), .A2(n4445), .ZN(n4443) );
  AND2_X1 U5836 ( .A1(n8755), .A2(n4674), .ZN(n4343) );
  AND2_X1 U5837 ( .A1(n5238), .A2(n6963), .ZN(n4344) );
  NAND2_X1 U5838 ( .A1(n5715), .A2(n5592), .ZN(n5733) );
  NAND2_X1 U5839 ( .A1(n5954), .A2(n5955), .ZN(n4345) );
  NAND2_X1 U5840 ( .A1(n7284), .A2(n7900), .ZN(n7087) );
  INV_X1 U5841 ( .A(n7087), .ZN(n4689) );
  AND2_X1 U5842 ( .A1(n8687), .A2(n4338), .ZN(n4346) );
  INV_X1 U5843 ( .A(n9213), .ZN(n4656) );
  NAND2_X1 U5844 ( .A1(n7852), .A2(n7851), .ZN(n8576) );
  INV_X1 U5845 ( .A(n8576), .ZN(n8867) );
  AND2_X1 U5846 ( .A1(n4526), .A2(n4532), .ZN(n4347) );
  NOR2_X1 U5847 ( .A1(n6194), .A2(n4769), .ZN(n4348) );
  INV_X1 U5848 ( .A(n9498), .ZN(n9281) );
  NAND2_X1 U5849 ( .A1(n5520), .A2(n5519), .ZN(n9498) );
  AND2_X1 U5850 ( .A1(n4447), .A2(n4451), .ZN(n4349) );
  NAND2_X1 U5851 ( .A1(n5412), .A2(n5411), .ZN(n9528) );
  NOR2_X1 U5852 ( .A1(n9295), .A2(n4589), .ZN(n4350) );
  NAND2_X1 U5853 ( .A1(n5972), .A2(n5971), .ZN(n8914) );
  OR2_X1 U5854 ( .A1(n5239), .A2(n4798), .ZN(n4351) );
  NOR2_X1 U5855 ( .A1(n9599), .A2(n6511), .ZN(n4352) );
  AND2_X1 U5856 ( .A1(n7221), .A2(n7130), .ZN(n7550) );
  INV_X1 U5857 ( .A(n7550), .ZN(n4657) );
  AND2_X1 U5858 ( .A1(n5454), .A2(n5453), .ZN(n9326) );
  INV_X1 U5859 ( .A(n9326), .ZN(n9513) );
  NAND2_X1 U5860 ( .A1(n9337), .A2(n4572), .ZN(n4575) );
  AND3_X1 U5861 ( .A1(n5009), .A2(n5010), .A3(n5006), .ZN(n4353) );
  AND2_X1 U5862 ( .A1(n4487), .A2(n8162), .ZN(n4354) );
  AND2_X1 U5863 ( .A1(n9256), .A2(n7728), .ZN(n4355) );
  INV_X1 U5864 ( .A(n4834), .ZN(n4833) );
  NAND2_X1 U5865 ( .A1(n4836), .A2(n4327), .ZN(n4834) );
  INV_X1 U5866 ( .A(n4839), .ZN(n4838) );
  NAND2_X1 U5867 ( .A1(n4840), .A2(n4841), .ZN(n4839) );
  NAND2_X1 U5868 ( .A1(n9821), .A2(n6880), .ZN(n4356) );
  AND2_X1 U5869 ( .A1(n4614), .A2(n4916), .ZN(n4357) );
  INV_X1 U5870 ( .A(n5078), .ZN(n5115) );
  AND3_X1 U5871 ( .A1(n7532), .A2(n6796), .A3(n7537), .ZN(n4358) );
  AND2_X1 U5872 ( .A1(n5791), .A2(n4538), .ZN(n4359) );
  AND2_X1 U5873 ( .A1(n4746), .A2(n4747), .ZN(n4360) );
  INV_X1 U5874 ( .A(n6826), .ZN(n4778) );
  NAND2_X1 U5875 ( .A1(n4745), .A2(n4744), .ZN(n4361) );
  INV_X1 U5876 ( .A(n4791), .ZN(n4790) );
  NAND2_X1 U5877 ( .A1(n4795), .A2(n4793), .ZN(n4791) );
  AND2_X1 U5878 ( .A1(n4792), .A2(n4790), .ZN(n4362) );
  NAND2_X1 U5879 ( .A1(n5604), .A2(n5646), .ZN(n4548) );
  AND2_X1 U5880 ( .A1(n9774), .A2(n7239), .ZN(n4363) );
  INV_X1 U5881 ( .A(n4684), .ZN(n4683) );
  NOR2_X1 U5882 ( .A1(n8703), .A2(n8726), .ZN(n4684) );
  NOR2_X1 U5883 ( .A1(n9206), .A2(n9330), .ZN(n4364) );
  OR2_X1 U5884 ( .A1(n9505), .A2(n9209), .ZN(n4365) );
  NOR2_X1 U5885 ( .A1(n7498), .A2(n8207), .ZN(n4366) );
  NOR2_X1 U5886 ( .A1(n5924), .A2(n8194), .ZN(n4367) );
  NOR2_X1 U5887 ( .A1(n9519), .A2(n9202), .ZN(n4368) );
  NOR2_X1 U5888 ( .A1(n9510), .A2(n9207), .ZN(n4369) );
  AND2_X1 U5889 ( .A1(n5602), .A2(n4855), .ZN(n4370) );
  INV_X1 U5890 ( .A(n4562), .ZN(n4561) );
  NAND2_X1 U5891 ( .A1(n4563), .A2(n8719), .ZN(n4562) );
  AND2_X1 U5892 ( .A1(n8000), .A2(n8722), .ZN(n8738) );
  INV_X1 U5893 ( .A(n8738), .ZN(n4806) );
  NOR2_X1 U5894 ( .A1(n8862), .A2(n8572), .ZN(n8051) );
  NOR2_X1 U5895 ( .A1(n9281), .A2(n9295), .ZN(n4371) );
  INV_X1 U5896 ( .A(n4866), .ZN(n4865) );
  NOR2_X1 U5897 ( .A1(n4364), .A2(n9204), .ZN(n4866) );
  AND2_X1 U5898 ( .A1(n5836), .A2(n5835), .ZN(n4372) );
  AND2_X1 U5899 ( .A1(n4902), .A2(SI_4_), .ZN(n4373) );
  NAND2_X1 U5900 ( .A1(n8128), .A2(n4877), .ZN(n4374) );
  NOR2_X1 U5901 ( .A1(n9362), .A2(n9201), .ZN(n4375) );
  AND2_X1 U5902 ( .A1(n5663), .A2(n5665), .ZN(n4376) );
  AND2_X1 U5903 ( .A1(n7990), .A2(n8753), .ZN(n8764) );
  NAND2_X1 U5904 ( .A1(n5627), .A2(n4856), .ZN(n4377) );
  NAND2_X1 U5905 ( .A1(n7837), .A2(n4810), .ZN(n4378) );
  INV_X1 U5906 ( .A(n4691), .ZN(n4690) );
  NAND2_X1 U5907 ( .A1(n7876), .A2(n7280), .ZN(n4691) );
  INV_X1 U5908 ( .A(n9197), .ZN(n9634) );
  AND2_X1 U5909 ( .A1(n4442), .A2(n9030), .ZN(n4379) );
  INV_X1 U5910 ( .A(n7333), .ZN(n9642) );
  OR2_X1 U5911 ( .A1(n9484), .A2(n9773), .ZN(n4380) );
  AND2_X1 U5912 ( .A1(n4634), .A2(n4859), .ZN(n4381) );
  NOR2_X1 U5913 ( .A1(n8920), .A2(n8793), .ZN(n4382) );
  AND2_X1 U5914 ( .A1(n8649), .A2(n8023), .ZN(n8667) );
  INV_X1 U5915 ( .A(n8667), .ZN(n4679) );
  OR2_X1 U5916 ( .A1(n6374), .A2(n6210), .ZN(n4383) );
  AND2_X1 U5917 ( .A1(n7624), .A2(n7631), .ZN(n4384) );
  OR2_X1 U5918 ( .A1(n9421), .A2(n9439), .ZN(n4385) );
  AND2_X1 U5919 ( .A1(n7082), .A2(n6933), .ZN(n4386) );
  AND2_X1 U5920 ( .A1(n4443), .A2(n5444), .ZN(n4387) );
  OR2_X1 U5921 ( .A1(n4451), .A2(n5392), .ZN(n4388) );
  INV_X1 U5922 ( .A(n4879), .ZN(n4487) );
  INV_X1 U5923 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U5924 ( .A1(n5377), .A2(n5376), .ZN(n4389) );
  INV_X1 U5925 ( .A(n6542), .ZN(n4539) );
  XNOR2_X1 U5926 ( .A(n5638), .B(n5637), .ZN(n6118) );
  INV_X1 U5927 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4401) );
  AND2_X1 U5928 ( .A1(n4492), .A2(n4750), .ZN(n4390) );
  AND2_X1 U5929 ( .A1(n7495), .A2(n4559), .ZN(n4391) );
  AND2_X1 U5930 ( .A1(n4848), .A2(n7284), .ZN(n4392) );
  NAND2_X1 U5931 ( .A1(n4491), .A2(n4490), .ZN(n8130) );
  NAND2_X1 U5932 ( .A1(n5913), .A2(n5912), .ZN(n8938) );
  NAND3_X1 U5933 ( .A1(n4800), .A2(n5338), .A3(n8999), .ZN(n9104) );
  INV_X1 U5934 ( .A(n9439), .ZN(n9403) );
  AND4_X1 U5935 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n9439)
         );
  NAND2_X1 U5936 ( .A1(n8746), .A2(n4561), .ZN(n4564) );
  AND2_X1 U5937 ( .A1(n4754), .A2(n4753), .ZN(n4393) );
  AND2_X1 U5938 ( .A1(n4749), .A2(n4748), .ZN(n4394) );
  INV_X1 U5939 ( .A(n9204), .ZN(n4868) );
  NAND2_X1 U5940 ( .A1(n7121), .A2(n9315), .ZN(n7740) );
  NOR2_X1 U5941 ( .A1(n6621), .A2(n6620), .ZN(n6619) );
  XNOR2_X1 U5942 ( .A(n5007), .B(n5006), .ZN(n5539) );
  AND2_X1 U5943 ( .A1(n7862), .A2(n7909), .ZN(n4395) );
  NAND2_X1 U5944 ( .A1(n4675), .A2(n6933), .ZN(n7081) );
  INV_X1 U5945 ( .A(n9552), .ZN(n4569) );
  INV_X1 U5946 ( .A(n7424), .ZN(n4430) );
  NAND2_X1 U5947 ( .A1(n4664), .A2(n4663), .ZN(n6949) );
  AND2_X1 U5948 ( .A1(n4759), .A2(n4758), .ZN(n4396) );
  NAND2_X1 U5949 ( .A1(n4517), .A2(n4515), .ZN(n7112) );
  OR2_X1 U5950 ( .A1(n8581), .A2(n7508), .ZN(n8850) );
  INV_X1 U5951 ( .A(n8850), .ZN(n4837) );
  NAND2_X1 U5952 ( .A1(n4771), .A2(n4780), .ZN(n5165) );
  INV_X1 U5953 ( .A(n5165), .ZN(n4776) );
  NAND2_X1 U5954 ( .A1(n5014), .A2(n4998), .ZN(n4397) );
  INV_X1 U5955 ( .A(n5803), .ZN(n4518) );
  OR2_X1 U5956 ( .A1(n9561), .A2(n6743), .ZN(n9775) );
  NAND2_X1 U5957 ( .A1(n5062), .A2(n7383), .ZN(n6676) );
  OR2_X1 U5958 ( .A1(n7753), .A2(n9686), .ZN(n9438) );
  XNOR2_X1 U5959 ( .A(n5089), .B(n5508), .ZN(n6481) );
  AOI21_X1 U5960 ( .B1(n4858), .B2(n4329), .A(n4358), .ZN(n6811) );
  AND2_X1 U5961 ( .A1(n5644), .A2(n5643), .ZN(n5654) );
  INV_X1 U5962 ( .A(n5654), .ZN(n8807) );
  INV_X1 U5963 ( .A(n7383), .ZN(n9315) );
  XNOR2_X1 U5964 ( .A(n5027), .B(P1_IR_REG_19__SCAN_IN), .ZN(n7383) );
  INV_X1 U5965 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4578) );
  NAND2_X1 U5966 ( .A1(n6913), .A2(n6804), .ZN(n6898) );
  AOI21_X2 U5967 ( .B1(n9539), .B2(n9425), .A(n9544), .ZN(n9381) );
  OAI21_X2 U5968 ( .B1(n9263), .B2(n9271), .A(n4398), .ZN(n9244) );
  INV_X1 U5969 ( .A(n4629), .ZN(n4628) );
  NAND2_X1 U5970 ( .A1(n6754), .A2(n7535), .ZN(n4858) );
  NAND2_X1 U5971 ( .A1(n9416), .A2(n4385), .ZN(n4418) );
  NAND2_X1 U5972 ( .A1(n9203), .A2(n4880), .ZN(n9320) );
  OAI211_X1 U5973 ( .C1(n4576), .C2(n9775), .A(n4330), .B(n4399), .ZN(n9565)
         );
  INV_X1 U5974 ( .A(n6916), .ZN(n6803) );
  NAND2_X1 U5975 ( .A1(n4418), .A2(n4417), .ZN(n9411) );
  XNOR2_X1 U5976 ( .A(n5175), .B(n5174), .ZN(n6226) );
  OAI21_X1 U5977 ( .B1(n7242), .B2(n4869), .A(n7314), .ZN(n4629) );
  NAND2_X1 U5978 ( .A1(n4620), .A2(n4619), .ZN(n9203) );
  NAND2_X1 U5979 ( .A1(n9198), .A2(n9197), .ZN(n4626) );
  NAND2_X1 U5980 ( .A1(n4613), .A2(n4905), .ZN(n5175) );
  INV_X1 U5981 ( .A(n8051), .ZN(n4823) );
  OAI21_X2 U5982 ( .B1(n5395), .B2(n5394), .A(n4975), .ZN(n5410) );
  MUX2_X1 U5983 ( .A(n8056), .B(n8055), .S(n8054), .Z(n8057) );
  OAI21_X1 U5984 ( .B1(n6214), .B2(n4401), .A(n4400), .ZN(n4896) );
  OAI21_X2 U5985 ( .B1(n5512), .B2(n5513), .A(n5514), .ZN(n6059) );
  NAND2_X1 U5986 ( .A1(n4981), .A2(n4980), .ZN(n5425) );
  NAND2_X1 U5987 ( .A1(n6171), .A2(n6170), .ZN(n7567) );
  NAND2_X1 U5988 ( .A1(n5126), .A2(n5125), .ZN(n4522) );
  NAND2_X1 U5989 ( .A1(n7569), .A2(n7568), .ZN(n7592) );
  NAND2_X1 U5990 ( .A1(n4727), .A2(n4728), .ZN(n5464) );
  NAND2_X1 U5991 ( .A1(n5466), .A2(n5465), .ZN(n5487) );
  INV_X1 U5992 ( .A(n8571), .ZN(n8862) );
  OAI21_X1 U5993 ( .B1(n5363), .B2(n4967), .A(n4966), .ZN(n5379) );
  AOI21_X1 U5994 ( .B1(n9400), .B2(n9218), .A(n9217), .ZN(n9389) );
  NOR2_X1 U5995 ( .A1(n9328), .A2(n9329), .ZN(n9327) );
  NOR2_X1 U5996 ( .A1(n9327), .A2(n9225), .ZN(n9307) );
  OR2_X1 U5997 ( .A1(n5104), .A2(n6232), .ZN(n5106) );
  NAND2_X2 U5998 ( .A1(n7764), .A2(n6657), .ZN(n7535) );
  NAND2_X1 U5999 ( .A1(n9342), .A2(n9223), .ZN(n9328) );
  NAND2_X1 U6000 ( .A1(n7315), .A2(n7553), .ZN(n7318) );
  NAND4_X1 U6001 ( .A1(n4998), .A2(n5202), .A3(n4659), .A4(n4353), .ZN(n4408)
         );
  NAND2_X1 U6002 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U6003 ( .A1(n4696), .A2(n9315), .ZN(n4695) );
  NAND2_X1 U6004 ( .A1(n4615), .A2(n4618), .ZN(n4614) );
  NAND2_X1 U6005 ( .A1(n4971), .A2(n4970), .ZN(n5395) );
  NAND2_X1 U6006 ( .A1(n4414), .A2(n4411), .ZN(n8569) );
  NAND2_X1 U6007 ( .A1(n8566), .A2(n5654), .ZN(n4414) );
  AND2_X1 U6008 ( .A1(n7550), .A2(n7131), .ZN(n7223) );
  NAND2_X1 U6009 ( .A1(n4930), .A2(n4929), .ZN(n4631) );
  NAND2_X1 U6010 ( .A1(n4633), .A2(n4632), .ZN(n9263) );
  NAND2_X1 U6011 ( .A1(n4627), .A2(n4626), .ZN(n9431) );
  NAND2_X1 U6012 ( .A1(n5057), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U6013 ( .A1(n4419), .A2(n4357), .ZN(n5201) );
  NAND2_X1 U6014 ( .A1(n4909), .A2(n4615), .ZN(n4419) );
  INV_X1 U6015 ( .A(n6951), .ZN(n4664) );
  NAND2_X2 U6016 ( .A1(n8789), .A2(n4888), .ZN(n8790) );
  INV_X2 U6017 ( .A(n6713), .ZN(n9858) );
  NAND2_X1 U6018 ( .A1(n6713), .A2(n6696), .ZN(n7919) );
  NAND2_X1 U6019 ( .A1(n4767), .A2(n4424), .ZN(n9065) );
  NAND2_X1 U6020 ( .A1(n7301), .A2(n5281), .ZN(n4433) );
  NAND2_X1 U6021 ( .A1(n7301), .A2(n4426), .ZN(n4425) );
  INV_X1 U6022 ( .A(n5280), .ZN(n4432) );
  INV_X1 U6023 ( .A(n9091), .ZN(n4434) );
  NOR2_X2 U6024 ( .A1(n6619), .A2(n5149), .ZN(n6645) );
  NAND2_X1 U6025 ( .A1(n5445), .A2(n4387), .ZN(n9013) );
  NAND3_X1 U6026 ( .A1(n5445), .A2(n4443), .A3(n4442), .ZN(n4438) );
  NAND3_X1 U6027 ( .A1(n5445), .A2(n4443), .A3(n4379), .ZN(n4441) );
  NAND2_X1 U6028 ( .A1(n5442), .A2(n9020), .ZN(n9074) );
  INV_X1 U6029 ( .A(n5444), .ZN(n4444) );
  NOR2_X1 U6030 ( .A1(n4446), .A2(n9072), .ZN(n4445) );
  NAND3_X1 U6031 ( .A1(n5341), .A2(n4448), .A3(n9105), .ZN(n4447) );
  NAND3_X1 U6032 ( .A1(n5341), .A2(n9105), .A3(n4450), .ZN(n4449) );
  NAND2_X1 U6033 ( .A1(n5014), .A2(n4456), .ZN(n4458) );
  NAND2_X1 U6034 ( .A1(n4459), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6035 ( .A1(n5668), .A2(n4460), .ZN(n5669) );
  INV_X1 U6036 ( .A(n4464), .ZN(n4462) );
  NAND2_X1 U6037 ( .A1(n4466), .A2(n4464), .ZN(n4759) );
  NAND2_X1 U6038 ( .A1(n4471), .A2(n4470), .ZN(n4465) );
  INV_X1 U6039 ( .A(n4467), .ZN(n4466) );
  OAI21_X1 U6040 ( .B1(n4470), .B2(n4468), .A(n6588), .ZN(n4467) );
  INV_X1 U6041 ( .A(n8985), .ZN(n4476) );
  NAND3_X1 U6042 ( .A1(n4481), .A2(n4482), .A3(n4479), .ZN(n6028) );
  NAND3_X1 U6043 ( .A1(n4484), .A2(n4485), .A3(n6025), .ZN(n4482) );
  NOR2_X1 U6044 ( .A1(n8089), .A2(n4489), .ZN(n4488) );
  AND2_X1 U6045 ( .A1(n8092), .A2(n6013), .ZN(n4489) );
  NAND2_X1 U6046 ( .A1(n7435), .A2(n4493), .ZN(n4491) );
  NAND2_X1 U6047 ( .A1(n8173), .A2(n4500), .ZN(n4499) );
  NAND2_X1 U6048 ( .A1(n6973), .A2(n4508), .ZN(n4507) );
  INV_X1 U6049 ( .A(n5141), .ZN(n4521) );
  INV_X1 U6050 ( .A(n4537), .ZN(n8812) );
  INV_X2 U6051 ( .A(n4890), .ZN(n6214) );
  XNOR2_X1 U6052 ( .A(n4893), .B(SI_1_), .ZN(n5086) );
  NOR2_X1 U6053 ( .A1(n4547), .A2(n4543), .ZN(n4546) );
  AND2_X4 U6054 ( .A1(n4545), .A2(n4544), .ZN(n7859) );
  NOR2_X1 U6055 ( .A1(n8655), .A2(n8886), .ZN(n8654) );
  INV_X1 U6056 ( .A(n4564), .ZN(n8714) );
  NAND3_X1 U6057 ( .A1(n4565), .A2(n5127), .A3(n4341), .ZN(n9725) );
  INV_X1 U6058 ( .A(n4575), .ZN(n9296) );
  NAND3_X1 U6059 ( .A1(n4578), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4577) );
  NAND3_X1 U6060 ( .A1(n8570), .A2(n4581), .A3(n4580), .ZN(n4579) );
  NAND2_X1 U6061 ( .A1(n5103), .A2(n5102), .ZN(n4582) );
  NAND2_X1 U6062 ( .A1(n4891), .A2(n4892), .ZN(n4583) );
  NAND3_X1 U6063 ( .A1(n4607), .A2(n4604), .A3(n4602), .ZN(n4601) );
  MUX2_X1 U6064 ( .A(n6220), .B(n6216), .S(n6214), .Z(n5085) );
  NAND2_X1 U6065 ( .A1(n5160), .A2(n5159), .ZN(n4613) );
  NAND2_X1 U6066 ( .A1(n4873), .A2(n4621), .ZN(n4620) );
  OAI21_X1 U6067 ( .B1(n9198), .B2(n9197), .A(n9196), .ZN(n4627) );
  AOI21_X2 U6068 ( .B1(n7336), .B2(n7335), .A(n7334), .ZN(n9198) );
  NAND2_X1 U6069 ( .A1(n9320), .A2(n4322), .ZN(n4633) );
  NAND2_X1 U6070 ( .A1(n6758), .A2(n4640), .ZN(n4641) );
  NAND2_X1 U6071 ( .A1(n9452), .A2(n7539), .ZN(n6786) );
  NAND2_X1 U6072 ( .A1(n4643), .A2(n4384), .ZN(n7136) );
  NAND2_X1 U6073 ( .A1(n4644), .A2(n4649), .ZN(n4643) );
  NAND2_X1 U6074 ( .A1(n4648), .A2(n4646), .ZN(n4644) );
  NAND2_X1 U6075 ( .A1(n4652), .A2(n4651), .ZN(n9400) );
  CLKBUF_X1 U6076 ( .A(n4652), .Z(n4650) );
  AND4_X2 U6077 ( .A1(n4998), .A2(n5202), .A3(n4353), .A4(n4658), .ZN(n5030)
         );
  NAND3_X1 U6078 ( .A1(n4998), .A2(n5202), .A3(n4659), .ZN(n5004) );
  NAND3_X2 U6079 ( .A1(n5066), .A2(n5065), .A3(n4660), .ZN(n6491) );
  NAND2_X1 U6080 ( .A1(n7318), .A2(n7644), .ZN(n7358) );
  NAND2_X1 U6081 ( .A1(n9343), .A2(n9344), .ZN(n9342) );
  NAND2_X1 U6082 ( .A1(n9292), .A2(n9227), .ZN(n9283) );
  AOI21_X2 U6083 ( .B1(n9283), .B2(n9229), .A(n9228), .ZN(n9270) );
  NAND2_X1 U6084 ( .A1(n9270), .A2(n9271), .ZN(n9254) );
  AND2_X2 U6085 ( .A1(n7337), .A2(n7642), .ZN(n9214) );
  OAI21_X2 U6086 ( .B1(n9390), .B2(n9221), .A(n9220), .ZN(n9354) );
  NAND2_X1 U6087 ( .A1(n6746), .A2(n6693), .ZN(n6744) );
  NOR2_X2 U6088 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4995) );
  AND2_X2 U6089 ( .A1(n4997), .A2(n5015), .ZN(n4998) );
  NAND2_X1 U6090 ( .A1(n4665), .A2(n8080), .ZN(n7918) );
  NOR2_X1 U6091 ( .A1(n6702), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U6092 ( .A1(n7911), .A2(n4665), .ZN(n6951) );
  NAND2_X1 U6093 ( .A1(n4675), .A2(n4386), .ZN(n7086) );
  NAND2_X1 U6094 ( .A1(n7088), .A2(n4687), .ZN(n4685) );
  NAND2_X1 U6095 ( .A1(n4685), .A2(n4686), .ZN(n7405) );
  AND3_X2 U6096 ( .A1(n5627), .A2(n4856), .A3(n4370), .ZN(n6084) );
  NAND2_X1 U6097 ( .A1(n6086), .A2(n5647), .ZN(n7504) );
  NAND2_X1 U6098 ( .A1(n4695), .A2(n4694), .ZN(n7759) );
  OAI21_X1 U6099 ( .B1(n4697), .B2(n7753), .A(n7752), .ZN(n4696) );
  NAND2_X1 U6100 ( .A1(n7751), .A2(n7750), .ZN(n4699) );
  NAND2_X1 U6101 ( .A1(n4701), .A2(n4703), .ZN(n5283) );
  NAND2_X1 U6102 ( .A1(n4948), .A2(n4947), .ZN(n5304) );
  NAND2_X1 U6103 ( .A1(n5343), .A2(n5342), .ZN(n4962) );
  NAND3_X1 U6104 ( .A1(n4717), .A2(n4723), .A3(n4716), .ZN(n7720) );
  NAND2_X1 U6105 ( .A1(n7714), .A2(n7740), .ZN(n4721) );
  NAND2_X1 U6106 ( .A1(n4726), .A2(n4911), .ZN(n5193) );
  NAND2_X1 U6107 ( .A1(n5425), .A2(n4730), .ZN(n4727) );
  NAND2_X1 U6108 ( .A1(n4733), .A2(n5681), .ZN(n6555) );
  NAND2_X1 U6109 ( .A1(n6498), .A2(n6497), .ZN(n4733) );
  OAI21_X1 U6110 ( .B1(n6497), .B2(n6498), .A(n4733), .ZN(n6505) );
  INV_X1 U6111 ( .A(n5750), .ZN(n4740) );
  NAND2_X1 U6112 ( .A1(n5750), .A2(n4735), .ZN(n4734) );
  NOR2_X1 U6113 ( .A1(n5750), .A2(n4884), .ZN(n6838) );
  INV_X1 U6114 ( .A(n4884), .ZN(n4741) );
  NAND2_X2 U6115 ( .A1(n6700), .A2(n4742), .ZN(n5679) );
  INV_X1 U6116 ( .A(n6012), .ZN(n5998) );
  INV_X1 U6117 ( .A(n7444), .ZN(n4756) );
  NAND2_X1 U6118 ( .A1(n4761), .A2(n4760), .ZN(n7435) );
  OAI21_X1 U6119 ( .B1(n5928), .B2(n4765), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5642) );
  AND2_X1 U6120 ( .A1(n6044), .A2(n6043), .ZN(n8183) );
  NAND2_X1 U6121 ( .A1(n7811), .A2(n7810), .ZN(n7823) );
  NAND3_X1 U6122 ( .A1(n6044), .A2(n6081), .A3(n6043), .ZN(n7811) );
  NAND2_X1 U6123 ( .A1(n7823), .A2(n7819), .ZN(n7821) );
  NAND2_X1 U6124 ( .A1(n9023), .A2(n9021), .ZN(n5442) );
  NAND2_X1 U6125 ( .A1(n8070), .A2(n5408), .ZN(n4767) );
  NAND2_X1 U6126 ( .A1(n6207), .A2(n4768), .ZN(P1_U3218) );
  INV_X1 U6127 ( .A(n6645), .ZN(n4771) );
  OAI21_X1 U6128 ( .B1(n6645), .B2(n4779), .A(n4782), .ZN(n4781) );
  NAND2_X1 U6129 ( .A1(n6645), .A2(n4782), .ZN(n4773) );
  NAND4_X1 U6130 ( .A1(n4988), .A2(n4990), .A3(n4989), .A4(n5055), .ZN(n4783)
         );
  AND4_X2 U6131 ( .A1(n4786), .A2(n4784), .A3(n4987), .A4(n5099), .ZN(n5202)
         );
  NAND2_X1 U6132 ( .A1(n4800), .A2(n8999), .ZN(n5340) );
  NAND2_X1 U6133 ( .A1(n7919), .A2(n7021), .ZN(n7911) );
  NAND2_X1 U6134 ( .A1(n9818), .A2(n7870), .ZN(n4803) );
  OAI21_X1 U6135 ( .B1(n8790), .B2(n4809), .A(n4808), .ZN(n8739) );
  NAND2_X1 U6136 ( .A1(n8790), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U6137 ( .A1(n7848), .A2(n4813), .ZN(n4812) );
  OAI211_X1 U6138 ( .C1(n7848), .C2(n4817), .A(n4814), .B(n4812), .ZN(n8059)
         );
  NAND2_X1 U6139 ( .A1(n8720), .A2(n4826), .ZN(n4828) );
  INV_X1 U6140 ( .A(n4828), .ZN(n8704) );
  NAND2_X1 U6141 ( .A1(n7509), .A2(n4832), .ZN(n4831) );
  AND2_X1 U6142 ( .A1(n8582), .A2(n7970), .ZN(n4841) );
  NAND2_X1 U6143 ( .A1(n7091), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U6144 ( .A1(n7091), .A2(n7937), .ZN(n7092) );
  INV_X1 U6145 ( .A(n4848), .ZN(n7285) );
  INV_X1 U6146 ( .A(n7937), .ZN(n4850) );
  INV_X1 U6147 ( .A(n7876), .ZN(n4851) );
  NOR2_X1 U6148 ( .A1(n5647), .A2(n4853), .ZN(n5606) );
  NAND3_X1 U6149 ( .A1(n5646), .A2(n5648), .A3(n4854), .ZN(n4853) );
  NAND3_X1 U6150 ( .A1(n5627), .A2(n4856), .A3(n5602), .ZN(n6087) );
  NAND2_X2 U6151 ( .A1(n6210), .A2(n4409), .ZN(n5104) );
  NAND2_X4 U6152 ( .A1(n5570), .A2(n6268), .ZN(n6210) );
  XNOR2_X2 U6153 ( .A(n5001), .B(n5000), .ZN(n6268) );
  XNOR2_X2 U6154 ( .A(n4999), .B(n5029), .ZN(n5570) );
  NAND2_X1 U6155 ( .A1(n7532), .A2(n7537), .ZN(n6793) );
  NAND2_X1 U6156 ( .A1(n4858), .A2(n6675), .ZN(n6794) );
  NAND2_X1 U6157 ( .A1(n4874), .A2(n4875), .ZN(n7129) );
  NAND2_X1 U6158 ( .A1(n6902), .A2(n7043), .ZN(n4874) );
  NAND2_X2 U6159 ( .A1(n6801), .A2(n6800), .ZN(n9742) );
  AND2_X1 U6160 ( .A1(n5202), .A2(n4876), .ZN(n5014) );
  NOR2_X2 U6161 ( .A1(n9373), .A2(n9525), .ZN(n9358) );
  NAND2_X1 U6162 ( .A1(n6697), .A2(n5678), .ZN(n5666) );
  INV_X1 U6163 ( .A(n5666), .ZN(n5668) );
  AND2_X1 U6164 ( .A1(n7281), .A2(n7090), .ZN(n9904) );
  OR2_X1 U6165 ( .A1(n5704), .A2(n9600), .ZN(n5656) );
  NAND2_X1 U6166 ( .A1(n5025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6167 ( .A1(n7762), .A2(n5061), .ZN(n7753) );
  AND2_X1 U6168 ( .A1(n8991), .A2(n9678), .ZN(n5587) );
  NAND2_X1 U6169 ( .A1(n5032), .A2(n5031), .ZN(n5036) );
  BUF_X4 U6170 ( .A(n5094), .Z(n7601) );
  NAND2_X1 U6171 ( .A1(n6210), .A2(n6214), .ZN(n5143) );
  NAND2_X1 U6172 ( .A1(n5004), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5008) );
  INV_X1 U6173 ( .A(n5417), .ZN(n5077) );
  NAND2_X1 U6174 ( .A1(n6741), .A2(n9133), .ZN(n7765) );
  INV_X1 U6175 ( .A(n8392), .ZN(n6870) );
  NAND2_X1 U6176 ( .A1(n5034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5035) );
  INV_X1 U6177 ( .A(n5034), .ZN(n5032) );
  INV_X1 U6178 ( .A(n5043), .ZN(n8077) );
  NOR2_X1 U6179 ( .A1(n6566), .A2(n6565), .ZN(n6564) );
  AND2_X1 U6180 ( .A1(n5582), .A2(n5581), .ZN(n9111) );
  NAND2_X1 U6181 ( .A1(n6789), .A2(n9465), .ZN(n9460) );
  OR2_X1 U6182 ( .A1(n8769), .A2(n8588), .ZN(n4878) );
  AND2_X1 U6183 ( .A1(n6014), .A2(n8091), .ZN(n4879) );
  OR2_X1 U6184 ( .A1(n9341), .A2(n9356), .ZN(n4880) );
  XOR2_X1 U6185 ( .A(n6472), .B(n6339), .Z(n4883) );
  AND2_X1 U6186 ( .A1(n5749), .A2(n5748), .ZN(n4884) );
  OR2_X1 U6187 ( .A1(n8213), .A2(n7002), .ZN(n4885) );
  AND2_X1 U6188 ( .A1(n4929), .A2(n4928), .ZN(n4886) );
  INV_X1 U6189 ( .A(n8987), .ZN(n6366) );
  AND2_X1 U6190 ( .A1(n4923), .A2(n4922), .ZN(n4887) );
  AND2_X1 U6191 ( .A1(n8791), .A2(n8788), .ZN(n4888) );
  AND4_X1 U6192 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n9310)
         );
  INV_X1 U6193 ( .A(n6025), .ZN(n6017) );
  INV_X1 U6194 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5592) );
  NOR3_X1 U6195 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5602) );
  INV_X1 U6196 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5632) );
  INV_X1 U6197 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5367) );
  INV_X1 U6198 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4994) );
  INV_X1 U6199 ( .A(n7522), .ZN(n5906) );
  INV_X1 U6200 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5945) );
  INV_X1 U6201 ( .A(n8641), .ZN(n8595) );
  INV_X1 U6202 ( .A(n5339), .ZN(n5338) );
  NOR2_X1 U6203 ( .A1(n5385), .A2(n9084), .ZN(n5402) );
  XNOR2_X1 U6204 ( .A(n5063), .B(n5061), .ZN(n5062) );
  INV_X1 U6205 ( .A(SI_25_), .ZN(n5491) );
  INV_X1 U6206 ( .A(SI_22_), .ZN(n8314) );
  INV_X1 U6207 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4991) );
  INV_X1 U6208 ( .A(n6629), .ZN(n5731) );
  INV_X1 U6209 ( .A(n7438), .ZN(n5872) );
  OR2_X1 U6210 ( .A1(n6047), .A2(n8186), .ZN(n6071) );
  OR2_X1 U6211 ( .A1(n5973), .A2(n8156), .ZN(n5987) );
  NOR2_X1 U6212 ( .A1(n8765), .A2(n8923), .ZN(n8586) );
  OR2_X1 U6213 ( .A1(n5859), .A2(n5615), .ZN(n5878) );
  NAND2_X1 U6214 ( .A1(n6881), .A2(n4356), .ZN(n6882) );
  NOR2_X1 U6215 ( .A1(n7457), .A2(n7456), .ZN(n7477) );
  INV_X1 U6216 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6150) );
  INV_X1 U6217 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5287) );
  INV_X1 U6218 ( .A(n5110), .ZN(n5108) );
  AND2_X1 U6219 ( .A1(n5331), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5348) );
  AND2_X1 U6220 ( .A1(n5402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5413) );
  AND2_X1 U6221 ( .A1(n6195), .A2(n6180), .ZN(n9250) );
  INV_X1 U6222 ( .A(n9310), .ZN(n9209) );
  AND3_X1 U6223 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5167) );
  AND2_X1 U6224 ( .A1(n6240), .A2(n9315), .ZN(n5561) );
  INV_X1 U6225 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5305) );
  INV_X1 U6226 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8156) );
  INV_X1 U6227 ( .A(n8756), .ZN(n8725) );
  INV_X1 U6228 ( .A(n8137), .ZN(n8200) );
  OR2_X1 U6229 ( .A1(n6007), .A2(n8095), .ZN(n6019) );
  INV_X1 U6230 ( .A(n7858), .ZN(n6022) );
  INV_X1 U6231 ( .A(n6126), .ZN(n6509) );
  AND2_X1 U6232 ( .A1(n8914), .A2(n8766), .ZN(n8589) );
  INV_X1 U6233 ( .A(n8765), .ZN(n8805) );
  INV_X1 U6234 ( .A(n8209), .ZN(n7404) );
  INV_X1 U6235 ( .A(n9823), .ZN(n6886) );
  INV_X1 U6236 ( .A(n6708), .ZN(n6709) );
  INV_X1 U6237 ( .A(n8208), .ZN(n7492) );
  INV_X1 U6238 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9002) );
  XNOR2_X1 U6239 ( .A(n5146), .B(n5508), .ZN(n5151) );
  NOR2_X1 U6240 ( .A1(n5252), .A2(n6340), .ZN(n5270) );
  OR2_X1 U6241 ( .A1(n5580), .A2(n5559), .ZN(n5567) );
  OR2_X1 U6242 ( .A1(n7753), .A2(n5568), .ZN(n6490) );
  OR2_X1 U6243 ( .A1(n5404), .A2(n5133), .ZN(n5134) );
  INV_X1 U6244 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6401) );
  INV_X1 U6245 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6340) );
  INV_X1 U6246 ( .A(n9272), .ZN(n9295) );
  AND2_X1 U6247 ( .A1(n9513), .A2(n9345), .ZN(n9204) );
  INV_X1 U6248 ( .A(n9202), .ZN(n9356) );
  INV_X1 U6249 ( .A(n9533), .ZN(n9388) );
  AND2_X1 U6250 ( .A1(n7650), .A2(n9213), .ZN(n7690) );
  OR2_X1 U6251 ( .A1(n7242), .A2(n7552), .ZN(n7240) );
  AND2_X1 U6252 ( .A1(n7631), .A2(n7671), .ZN(n7547) );
  AND2_X1 U6253 ( .A1(n7541), .A2(n6799), .ZN(n9470) );
  INV_X1 U6254 ( .A(n9470), .ZN(n6800) );
  INV_X1 U6255 ( .A(n9465), .ZN(n9444) );
  AND2_X1 U6256 ( .A1(n7698), .A2(n7702), .ZN(n9410) );
  AND2_X1 U6257 ( .A1(n6660), .A2(n6659), .ZN(n9436) );
  INV_X1 U6258 ( .A(n9775), .ZN(n9749) );
  INV_X1 U6259 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5557) );
  OAI21_X1 U6260 ( .B1(n8636), .B2(n8191), .A(n6146), .ZN(n6147) );
  AOI21_X1 U6261 ( .B1(n6500), .B2(n6129), .A(P2_U3152), .ZN(n8137) );
  NAND2_X1 U6262 ( .A1(n8183), .A2(n8182), .ZN(n8181) );
  INV_X1 U6263 ( .A(n7862), .ZN(n8572) );
  AND2_X1 U6264 ( .A1(n6524), .A2(n6523), .ZN(n9804) );
  AND2_X1 U6265 ( .A1(n6545), .A2(n6142), .ZN(n9620) );
  INV_X1 U6266 ( .A(n9815), .ZN(n8824) );
  INV_X1 U6267 ( .A(n9833), .ZN(n8858) );
  INV_X1 U6268 ( .A(n6930), .ZN(n9885) );
  INV_X1 U6269 ( .A(n7076), .ZN(n7070) );
  NAND2_X1 U6270 ( .A1(n6118), .A2(n6123), .ZN(n9867) );
  INV_X1 U6271 ( .A(n9921), .ZN(n9889) );
  AND2_X1 U6272 ( .A1(n6110), .A2(n6109), .ZN(n7076) );
  AND2_X1 U6273 ( .A1(n6098), .A2(n6097), .ZN(n9838) );
  INV_X1 U6274 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6094) );
  INV_X1 U6275 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5788) );
  NOR2_X1 U6276 ( .A1(n4409), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8979) );
  INV_X1 U6277 ( .A(n9773), .ZN(n9748) );
  INV_X1 U6278 ( .A(n9683), .ZN(n9100) );
  NOR2_X2 U6279 ( .A1(n5567), .A2(n5560), .ZN(n9678) );
  AND4_X1 U6280 ( .A1(n6185), .A2(n6184), .A3(n6183), .A4(n6182), .ZN(n9235)
         );
  AND3_X1 U6281 ( .A1(n5433), .A2(n5432), .A3(n5431), .ZN(n9201) );
  INV_X1 U6282 ( .A(n9695), .ZN(n9157) );
  AND2_X1 U6283 ( .A1(n6269), .A2(n9686), .ZN(n9698) );
  OR2_X1 U6284 ( .A1(n9228), .A2(n7531), .ZN(n9284) );
  INV_X1 U6285 ( .A(n9438), .ZN(n9454) );
  INV_X1 U6286 ( .A(n9436), .ZN(n9459) );
  NOR2_X1 U6287 ( .A1(n9305), .A2(n6739), .ZN(n7372) );
  AND2_X1 U6288 ( .A1(n5543), .A2(n9581), .ZN(n7388) );
  INV_X1 U6289 ( .A(n9770), .ZN(n9655) );
  OR2_X1 U6290 ( .A1(n7740), .A2(n6743), .ZN(n9753) );
  NAND2_X1 U6291 ( .A1(n6676), .A2(n9753), .ZN(n9770) );
  INV_X1 U6292 ( .A(n9753), .ZN(n9781) );
  INV_X1 U6293 ( .A(n7388), .ZN(n7389) );
  AND2_X1 U6294 ( .A1(n5328), .A2(n5344), .ZN(n7153) );
  AND2_X1 U6295 ( .A1(n4409), .A2(P1_U3084), .ZN(n9588) );
  OAI21_X1 U6296 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9944), .ZN(n9977) );
  AND2_X1 U6297 ( .A1(n6112), .A2(n6111), .ZN(n6507) );
  INV_X1 U6298 ( .A(n8920), .ZN(n8769) );
  AND2_X1 U6299 ( .A1(n6124), .A2(n9827), .ZN(n8191) );
  NAND2_X1 U6300 ( .A1(n6140), .A2(n6119), .ZN(n8204) );
  NAND2_X1 U6301 ( .A1(n6545), .A2(n6544), .ZN(n9807) );
  OR2_X1 U6302 ( .A1(n8846), .A2(n7007), .ZN(n8781) );
  AND2_X1 U6303 ( .A1(n6710), .A2(n9827), .ZN(n9837) );
  NAND2_X1 U6304 ( .A1(n4316), .A2(n6701), .ZN(n9825) );
  OR2_X1 U6305 ( .A1(n7077), .A2(n7070), .ZN(n9937) );
  OR2_X1 U6306 ( .A1(n7077), .A2(n7076), .ZN(n9923) );
  INV_X2 U6307 ( .A(n9923), .ZN(n9924) );
  NOR2_X1 U6308 ( .A1(n9839), .A2(n9838), .ZN(n9841) );
  INV_X1 U6309 ( .A(n9841), .ZN(n9844) );
  INV_X1 U6310 ( .A(n7909), .ZN(n7895) );
  INV_X1 U6311 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6563) );
  INV_X1 U6312 ( .A(n9505), .ZN(n9208) );
  NAND2_X1 U6313 ( .A1(n9677), .A2(n9748), .ZN(n9056) );
  INV_X1 U6314 ( .A(n7530), .ZN(n9286) );
  INV_X1 U6315 ( .A(n9330), .ZN(n9207) );
  INV_X1 U6316 ( .A(n9048), .ZN(n9425) );
  INV_X1 U6317 ( .A(n7239), .ZN(n9126) );
  INV_X1 U6318 ( .A(n9698), .ZN(n7161) );
  OR2_X1 U6319 ( .A1(n9177), .A2(n9686), .ZN(n9695) );
  OR2_X1 U6320 ( .A1(P1_U3083), .A2(n6429), .ZN(n9184) );
  INV_X1 U6321 ( .A(n9429), .ZN(n9376) );
  NAND2_X1 U6322 ( .A1(n9460), .A2(n6678), .ZN(n9450) );
  AND2_X1 U6323 ( .A1(n6814), .A2(n6813), .ZN(n9737) );
  INV_X1 U6324 ( .A(n9802), .ZN(n9799) );
  AND2_X1 U6325 ( .A1(n9737), .A2(n9736), .ZN(n9790) );
  NAND2_X1 U6326 ( .A1(n6240), .A2(n6664), .ZN(n9711) );
  INV_X1 U6327 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7804) );
  INV_X1 U6328 ( .A(n7762), .ZN(n7755) );
  INV_X1 U6329 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6616) );
  AND2_X1 U6330 ( .A1(n6507), .A2(n9847), .ZN(P2_U3966) );
  NOR2_X2 U6331 ( .A1(n6286), .A2(n6241), .ZN(P1_U4006) );
  AND2_X1 U6332 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6333 ( .A1(n4890), .A2(n4889), .ZN(n5069) );
  INV_X1 U6334 ( .A(n5086), .ZN(n4892) );
  INV_X1 U6335 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6216) );
  INV_X1 U6336 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6220) );
  INV_X1 U6337 ( .A(n5085), .ZN(n4891) );
  NAND2_X1 U6338 ( .A1(n4893), .A2(SI_1_), .ZN(n4894) );
  INV_X1 U6339 ( .A(SI_2_), .ZN(n4895) );
  XNOR2_X1 U6340 ( .A(n4896), .B(n4895), .ZN(n5102) );
  NAND2_X1 U6341 ( .A1(n4896), .A2(SI_2_), .ZN(n4897) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6233) );
  INV_X1 U6343 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6215) );
  MUX2_X1 U6344 ( .A(n6233), .B(n6215), .S(n4474), .Z(n4898) );
  XNOR2_X1 U6345 ( .A(n4898), .B(SI_3_), .ZN(n5125) );
  INV_X1 U6346 ( .A(n4898), .ZN(n4899) );
  NAND2_X1 U6347 ( .A1(n4899), .A2(SI_3_), .ZN(n4900) );
  MUX2_X1 U6348 ( .A(n6230), .B(n6221), .S(n4474), .Z(n4901) );
  INV_X1 U6349 ( .A(n4901), .ZN(n4902) );
  MUX2_X1 U6350 ( .A(n6225), .B(n6218), .S(n4474), .Z(n4903) );
  XNOR2_X1 U6351 ( .A(n4903), .B(SI_5_), .ZN(n5159) );
  INV_X1 U6352 ( .A(n4903), .ZN(n4904) );
  NAND2_X1 U6353 ( .A1(n4904), .A2(SI_5_), .ZN(n4905) );
  MUX2_X1 U6354 ( .A(n6227), .B(n6222), .S(n4474), .Z(n4906) );
  XNOR2_X1 U6355 ( .A(n4906), .B(SI_6_), .ZN(n5174) );
  INV_X1 U6356 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6357 ( .A1(n4907), .A2(SI_6_), .ZN(n4908) );
  MUX2_X1 U6358 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4474), .Z(n4910) );
  INV_X1 U6359 ( .A(SI_7_), .ZN(n8381) );
  XNOR2_X1 U6360 ( .A(n4910), .B(n8381), .ZN(n5057) );
  NAND2_X1 U6361 ( .A1(n4910), .A2(SI_7_), .ZN(n4911) );
  INV_X1 U6362 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6246) );
  MUX2_X1 U6363 ( .A(n6244), .B(n6246), .S(n4474), .Z(n4913) );
  INV_X1 U6364 ( .A(SI_8_), .ZN(n4912) );
  NAND2_X1 U6365 ( .A1(n4913), .A2(n4912), .ZN(n4916) );
  INV_X1 U6366 ( .A(n4913), .ZN(n4914) );
  NAND2_X1 U6367 ( .A1(n4914), .A2(SI_8_), .ZN(n4915) );
  NAND2_X1 U6368 ( .A1(n4916), .A2(n4915), .ZN(n5192) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4918) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4917) );
  MUX2_X1 U6371 ( .A(n4918), .B(n4917), .S(n4409), .Z(n4920) );
  INV_X1 U6372 ( .A(SI_9_), .ZN(n4919) );
  NAND2_X1 U6373 ( .A1(n4920), .A2(n4919), .ZN(n4923) );
  INV_X1 U6374 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6375 ( .A1(n4921), .A2(SI_9_), .ZN(n4922) );
  NAND2_X1 U6376 ( .A1(n5201), .A2(n4887), .ZN(n4924) );
  NAND2_X1 U6377 ( .A1(n4924), .A2(n4923), .ZN(n5217) );
  INV_X1 U6378 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6291) );
  INV_X1 U6379 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6293) );
  MUX2_X1 U6380 ( .A(n6291), .B(n6293), .S(n4409), .Z(n4926) );
  INV_X1 U6381 ( .A(SI_10_), .ZN(n4925) );
  NAND2_X1 U6382 ( .A1(n4926), .A2(n4925), .ZN(n4929) );
  INV_X1 U6383 ( .A(n4926), .ZN(n4927) );
  NAND2_X1 U6384 ( .A1(n4927), .A2(SI_10_), .ZN(n4928) );
  MUX2_X1 U6385 ( .A(n6296), .B(n6295), .S(n4409), .Z(n4931) );
  XNOR2_X1 U6386 ( .A(n4931), .B(SI_11_), .ZN(n5244) );
  INV_X1 U6387 ( .A(n5244), .ZN(n4934) );
  INV_X1 U6388 ( .A(n4931), .ZN(n4932) );
  NAND2_X1 U6389 ( .A1(n4932), .A2(SI_11_), .ZN(n4933) );
  INV_X1 U6390 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n4936) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4935) );
  MUX2_X1 U6392 ( .A(n4936), .B(n4935), .S(n4409), .Z(n4938) );
  INV_X1 U6393 ( .A(SI_12_), .ZN(n4937) );
  NAND2_X1 U6394 ( .A1(n4938), .A2(n4937), .ZN(n4941) );
  INV_X1 U6395 ( .A(n4938), .ZN(n4939) );
  NAND2_X1 U6396 ( .A1(n4939), .A2(SI_12_), .ZN(n4940) );
  NAND2_X1 U6397 ( .A1(n4941), .A2(n4940), .ZN(n5265) );
  INV_X1 U6398 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4942) );
  MUX2_X1 U6399 ( .A(n6496), .B(n4942), .S(n4409), .Z(n4944) );
  INV_X1 U6400 ( .A(SI_13_), .ZN(n4943) );
  NAND2_X1 U6401 ( .A1(n4944), .A2(n4943), .ZN(n4947) );
  INV_X1 U6402 ( .A(n4944), .ZN(n4945) );
  NAND2_X1 U6403 ( .A1(n4945), .A2(SI_13_), .ZN(n4946) );
  MUX2_X1 U6404 ( .A(n6563), .B(n6561), .S(n4409), .Z(n4949) );
  XNOR2_X1 U6405 ( .A(n4949), .B(SI_14_), .ZN(n5303) );
  INV_X1 U6406 ( .A(n5303), .ZN(n4952) );
  INV_X1 U6407 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6408 ( .A1(n4950), .A2(SI_14_), .ZN(n4951) );
  MUX2_X1 U6409 ( .A(n6614), .B(n8298), .S(n4409), .Z(n4954) );
  NAND2_X1 U6410 ( .A1(n4954), .A2(n4953), .ZN(n4957) );
  INV_X1 U6411 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6412 ( .A1(n4955), .A2(SI_15_), .ZN(n4956) );
  NAND2_X1 U6413 ( .A1(n4957), .A2(n4956), .ZN(n5322) );
  MUX2_X1 U6414 ( .A(n6618), .B(n6616), .S(n4409), .Z(n4958) );
  NAND2_X1 U6415 ( .A1(n4958), .A2(n8251), .ZN(n4961) );
  INV_X1 U6416 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U6417 ( .A1(n4959), .A2(SI_16_), .ZN(n4960) );
  NAND2_X1 U6418 ( .A1(n4962), .A2(n4961), .ZN(n5363) );
  INV_X1 U6419 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4963) );
  MUX2_X1 U6420 ( .A(n6655), .B(n4963), .S(n4409), .Z(n4964) );
  XNOR2_X1 U6421 ( .A(n4964), .B(SI_17_), .ZN(n5362) );
  INV_X1 U6422 ( .A(n5362), .ZN(n4967) );
  INV_X1 U6423 ( .A(n4964), .ZN(n4965) );
  NAND2_X1 U6424 ( .A1(n4965), .A2(SI_17_), .ZN(n4966) );
  MUX2_X1 U6425 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4409), .Z(n4969) );
  XNOR2_X1 U6426 ( .A(n4969), .B(SI_18_), .ZN(n5378) );
  INV_X1 U6427 ( .A(n5378), .ZN(n4968) );
  NAND2_X1 U6428 ( .A1(n5379), .A2(n4968), .ZN(n4971) );
  NAND2_X1 U6429 ( .A1(n4969), .A2(SI_18_), .ZN(n4970) );
  MUX2_X1 U6430 ( .A(n8315), .B(n6868), .S(n4409), .Z(n4972) );
  NAND2_X1 U6431 ( .A1(n4972), .A2(n8237), .ZN(n4975) );
  INV_X1 U6432 ( .A(n4972), .ZN(n4973) );
  NAND2_X1 U6433 ( .A1(n4973), .A2(SI_19_), .ZN(n4974) );
  NAND2_X1 U6434 ( .A1(n4975), .A2(n4974), .ZN(n5394) );
  MUX2_X1 U6435 ( .A(n7063), .B(n8304), .S(n4409), .Z(n4977) );
  INV_X1 U6436 ( .A(SI_20_), .ZN(n4976) );
  NAND2_X1 U6437 ( .A1(n4977), .A2(n4976), .ZN(n4980) );
  INV_X1 U6438 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6439 ( .A1(n4978), .A2(SI_20_), .ZN(n4979) );
  NAND2_X1 U6440 ( .A1(n5410), .A2(n5409), .ZN(n4981) );
  MUX2_X1 U6441 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4409), .Z(n4982) );
  XNOR2_X1 U6442 ( .A(n4982), .B(n8297), .ZN(n5424) );
  NAND2_X1 U6443 ( .A1(n4982), .A2(SI_21_), .ZN(n4983) );
  MUX2_X1 U6444 ( .A(n7125), .B(n7122), .S(n4409), .Z(n4984) );
  NAND2_X1 U6445 ( .A1(n4984), .A2(n8314), .ZN(n5446) );
  INV_X1 U6446 ( .A(n4984), .ZN(n4985) );
  NAND2_X1 U6447 ( .A1(n4985), .A2(SI_22_), .ZN(n4986) );
  NAND2_X1 U6448 ( .A1(n5446), .A2(n4986), .ZN(n5447) );
  XNOR2_X1 U6449 ( .A(n5448), .B(n5447), .ZN(n7120) );
  INV_X2 U6450 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5055) );
  NOR2_X2 U6451 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5016) );
  NOR2_X1 U6452 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4993) );
  NOR2_X1 U6453 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4996) );
  AND4_X2 U6454 ( .A1(n4996), .A2(n4995), .A3(n5305), .A4(n4994), .ZN(n5015)
         );
  INV_X2 U6455 ( .A(n5104), .ZN(n5245) );
  NAND2_X1 U6456 ( .A1(n7120), .A2(n5245), .ZN(n5003) );
  OR2_X1 U6457 ( .A1(n7597), .A2(n7122), .ZN(n5002) );
  NAND2_X1 U6458 ( .A1(n5008), .A2(n5009), .ZN(n5005) );
  INV_X1 U6459 ( .A(n5016), .ZN(n5017) );
  NAND2_X1 U6460 ( .A1(n5017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6461 ( .A1(n5024), .A2(n5023), .ZN(n5019) );
  NAND2_X1 U6462 ( .A1(n5021), .A2(n5020), .ZN(n5025) );
  INV_X1 U6463 ( .A(n5063), .ZN(n6677) );
  INV_X1 U6464 ( .A(n5568), .ZN(n7795) );
  NOR2_X1 U6465 ( .A1(n5061), .A2(n7795), .ZN(n5028) );
  NAND2_X1 U6466 ( .A1(n5030), .A2(n5029), .ZN(n5034) );
  AND2_X2 U6467 ( .A1(n8077), .A2(n5038), .ZN(n5094) );
  NAND2_X1 U6468 ( .A1(n7601), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5047) );
  INV_X1 U6469 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6470 ( .A1(n5167), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5166) );
  INV_X1 U6471 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5048) );
  NOR2_X1 U6472 ( .A1(n5166), .A2(n5048), .ZN(n5185) );
  NAND2_X1 U6473 ( .A1(n5185), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6474 ( .A1(n5270), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6475 ( .A1(n5348), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6476 ( .A1(n5428), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6477 ( .A1(n5039), .A2(n5429), .ZN(n5041) );
  INV_X1 U6478 ( .A(n5429), .ZN(n5040) );
  NAND2_X1 U6479 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5040), .ZN(n5456) );
  AND2_X1 U6480 ( .A1(n5041), .A2(n5456), .ZN(n9339) );
  NAND2_X1 U6481 ( .A1(n6181), .A2(n9339), .ZN(n5046) );
  INV_X4 U6482 ( .A(n5404), .ZN(n7600) );
  NAND2_X1 U6483 ( .A1(n7600), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6484 ( .A1(n7587), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5044) );
  NAND4_X1 U6485 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n9202)
         );
  AOI22_X1 U6486 ( .A1(n9519), .A2(n4333), .B1(n5532), .B2(n9202), .ZN(n9072)
         );
  NAND2_X1 U6487 ( .A1(n7587), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6488 ( .A1(n7600), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5052) );
  INV_X1 U6489 ( .A(n5417), .ZN(n5473) );
  AND2_X1 U6490 ( .A1(n5166), .A2(n5048), .ZN(n5049) );
  NOR2_X1 U6491 ( .A1(n5185), .A2(n5049), .ZN(n6969) );
  NAND2_X1 U6492 ( .A1(n5473), .A2(n6969), .ZN(n5051) );
  NAND2_X1 U6493 ( .A1(n7601), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5050) );
  INV_X1 U6494 ( .A(n9095), .ZN(n9128) );
  NOR2_X1 U6495 ( .A1(n5054), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6496 ( .A1(n5157), .A2(n5055), .ZN(n5172) );
  OAI21_X1 U6497 ( .B1(n5172), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5056) );
  XNOR2_X1 U6498 ( .A(n5056), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6321) );
  INV_X1 U6499 ( .A(n6321), .ZN(n6364) );
  XNOR2_X1 U6500 ( .A(n5058), .B(n5057), .ZN(n6238) );
  OR2_X1 U6501 ( .A1(n6238), .A2(n5104), .ZN(n5060) );
  INV_X1 U6502 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6236) );
  OR2_X1 U6503 ( .A1(n7597), .A2(n6236), .ZN(n5059) );
  OAI211_X1 U6504 ( .C1(n6210), .C2(n6364), .A(n5060), .B(n5059), .ZN(n6792)
         );
  AOI22_X1 U6505 ( .A1(n9128), .A2(n5532), .B1(n5229), .B2(n6792), .ZN(n5182)
         );
  INV_X1 U6506 ( .A(n5182), .ZN(n5184) );
  INV_X2 U6507 ( .A(n6792), .ZN(n9759) );
  OAI22_X1 U6508 ( .A1(n9095), .A2(n5505), .B1(n9759), .B2(n5478), .ZN(n5064)
         );
  XNOR2_X1 U6509 ( .A(n5064), .B(n5508), .ZN(n5183) );
  NAND2_X1 U6510 ( .A1(n5077), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5066) );
  INV_X1 U6511 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U6512 ( .A1(n5094), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6513 ( .A1(n6491), .A2(n5090), .ZN(n5072) );
  NAND2_X1 U6514 ( .A1(n4409), .A2(SI_0_), .ZN(n5068) );
  INV_X1 U6515 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6516 ( .A1(n5068), .A2(n5067), .ZN(n5070) );
  AND2_X1 U6517 ( .A1(n5070), .A2(n5069), .ZN(n6212) );
  MUX2_X1 U6518 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6212), .S(n6210), .Z(n6693) );
  INV_X1 U6519 ( .A(n6286), .ZN(n5073) );
  AOI22_X1 U6520 ( .A1(n6693), .A2(n5229), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5073), .ZN(n5071) );
  AND2_X1 U6521 ( .A1(n5072), .A2(n5071), .ZN(n6425) );
  NAND2_X1 U6522 ( .A1(n6491), .A2(n4333), .ZN(n5075) );
  AOI22_X1 U6523 ( .A1(n6693), .A2(n5222), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n5073), .ZN(n5074) );
  NAND2_X1 U6524 ( .A1(n5075), .A2(n5074), .ZN(n6424) );
  NAND2_X1 U6525 ( .A1(n6425), .A2(n6424), .ZN(n6423) );
  NAND3_X1 U6526 ( .A1(n5075), .A2(n5074), .A3(n5508), .ZN(n5076) );
  AND2_X1 U6527 ( .A1(n6423), .A2(n5076), .ZN(n6482) );
  NAND2_X1 U6528 ( .A1(n5078), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6529 ( .A1(n5093), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5079) );
  NAND4_X2 U6530 ( .A1(n5082), .A2(n5081), .A3(n5080), .A4(n5079), .ZN(n9133)
         );
  INV_X1 U6531 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6532 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5083) );
  XNOR2_X1 U6533 ( .A(n5084), .B(n5083), .ZN(n6388) );
  XNOR2_X1 U6534 ( .A(n5086), .B(n5085), .ZN(n6219) );
  OR2_X1 U6535 ( .A1(n5143), .A2(n6220), .ZN(n5087) );
  OAI211_X1 U6536 ( .C1(n6210), .C2(n6388), .A(n5088), .B(n5087), .ZN(n6681)
         );
  OAI22_X1 U6537 ( .A1(n6755), .A2(n5505), .B1(n6741), .B2(n5478), .ZN(n5089)
         );
  INV_X1 U6538 ( .A(n5090), .ZN(n5319) );
  OR2_X1 U6539 ( .A1(n5319), .A2(n6755), .ZN(n5092) );
  NAND2_X1 U6540 ( .A1(n6681), .A2(n5229), .ZN(n5091) );
  NAND2_X1 U6541 ( .A1(n5092), .A2(n5091), .ZN(n6484) );
  NAND2_X1 U6542 ( .A1(n6482), .A2(n6481), .ZN(n6487) );
  NAND2_X1 U6543 ( .A1(n6483), .A2(n6487), .ZN(n6566) );
  NAND2_X1 U6544 ( .A1(n6181), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6545 ( .A1(n5078), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6546 ( .A1(n5093), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6547 ( .A1(n5094), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5095) );
  OR2_X1 U6548 ( .A1(n5099), .A2(n5247), .ZN(n5101) );
  INV_X1 U6549 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6550 ( .A1(n5101), .A2(n5100), .ZN(n5122) );
  OAI21_X1 U6551 ( .B1(n5101), .B2(n5100), .A(n5122), .ZN(n6450) );
  XNOR2_X1 U6552 ( .A(n5102), .B(n5103), .ZN(n6232) );
  OR2_X1 U6553 ( .A1(n5143), .A2(n4401), .ZN(n5105) );
  INV_X1 U6554 ( .A(n6768), .ZN(n9718) );
  OAI22_X1 U6555 ( .A1(n6674), .A2(n5505), .B1(n9718), .B2(n5478), .ZN(n5107)
         );
  XNOR2_X1 U6556 ( .A(n5107), .B(n5508), .ZN(n5109) );
  INV_X2 U6557 ( .A(n6674), .ZN(n9131) );
  AOI22_X1 U6558 ( .A1(n9131), .A2(n5532), .B1(n5229), .B2(n6768), .ZN(n5110)
         );
  NAND2_X1 U6559 ( .A1(n5109), .A2(n5108), .ZN(n5112) );
  INV_X1 U6560 ( .A(n5109), .ZN(n5111) );
  NAND2_X1 U6561 ( .A1(n5111), .A2(n5110), .ZN(n5113) );
  NAND2_X1 U6562 ( .A1(n5112), .A2(n5113), .ZN(n6565) );
  INV_X1 U6563 ( .A(n5113), .ZN(n5114) );
  NOR2_X1 U6564 ( .A1(n6564), .A2(n5114), .ZN(n6621) );
  INV_X2 U6565 ( .A(n5115), .ZN(n5571) );
  NAND2_X1 U6566 ( .A1(n5571), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5121) );
  INV_X1 U6567 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6568 ( .A1(n7601), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5119) );
  INV_X1 U6569 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6570 ( .A1(n5473), .A2(n5117), .ZN(n5118) );
  AND4_X2 U6571 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n6808)
         );
  NAND2_X1 U6572 ( .A1(n5122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5124) );
  INV_X1 U6573 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5123) );
  XNOR2_X1 U6574 ( .A(n5124), .B(n5123), .ZN(n6415) );
  OR2_X1 U6575 ( .A1(n5143), .A2(n6215), .ZN(n5127) );
  AOI22_X1 U6576 ( .A1(n9130), .A2(n5532), .B1(n5229), .B2(n9725), .ZN(n5129)
         );
  INV_X1 U6577 ( .A(n9725), .ZN(n6795) );
  OAI22_X1 U6578 ( .A1(n6808), .A2(n5505), .B1(n6795), .B2(n5478), .ZN(n5128)
         );
  XNOR2_X1 U6579 ( .A(n5128), .B(n5508), .ZN(n5131) );
  XOR2_X1 U6580 ( .A(n5129), .B(n5131), .Z(n6620) );
  INV_X1 U6581 ( .A(n5129), .ZN(n5130) );
  NOR2_X1 U6582 ( .A1(n5131), .A2(n5130), .ZN(n6644) );
  INV_X1 U6583 ( .A(n6644), .ZN(n5148) );
  INV_X2 U6584 ( .A(n5115), .ZN(n7587) );
  NAND2_X1 U6585 ( .A1(n7587), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6586 ( .A1(n7601), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5136) );
  INV_X1 U6587 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5132) );
  XNOR2_X1 U6588 ( .A(n5132), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U6589 ( .A1(n6181), .A2(n6650), .ZN(n5135) );
  INV_X1 U6590 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5133) );
  INV_X1 U6591 ( .A(n5157), .ZN(n5140) );
  NAND2_X1 U6592 ( .A1(n5054), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  MUX2_X1 U6593 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5138), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5139) );
  NAND2_X1 U6594 ( .A1(n5140), .A2(n5139), .ZN(n6431) );
  XNOR2_X1 U6595 ( .A(n5142), .B(n5141), .ZN(n6229) );
  OR2_X1 U6596 ( .A1(n5104), .A2(n6229), .ZN(n5145) );
  OR2_X1 U6597 ( .A1(n5143), .A2(n6221), .ZN(n5144) );
  OAI211_X1 U6598 ( .C1(n6210), .C2(n6431), .A(n5145), .B(n5144), .ZN(n6819)
         );
  INV_X1 U6599 ( .A(n6819), .ZN(n9732) );
  OAI22_X1 U6600 ( .A1(n6829), .A2(n5505), .B1(n9732), .B2(n5478), .ZN(n5146)
         );
  OAI22_X1 U6601 ( .A1(n6829), .A2(n5319), .B1(n9732), .B2(n5505), .ZN(n5150)
         );
  XNOR2_X1 U6602 ( .A(n5151), .B(n5150), .ZN(n6647) );
  INV_X1 U6603 ( .A(n6647), .ZN(n5147) );
  NAND2_X1 U6604 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  NAND2_X1 U6605 ( .A1(n7601), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6606 ( .A1(n7587), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5155) );
  AOI21_X1 U6607 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5152) );
  NOR2_X1 U6608 ( .A1(n5152), .A2(n5167), .ZN(n6831) );
  NAND2_X1 U6609 ( .A1(n5473), .A2(n6831), .ZN(n5154) );
  NAND2_X1 U6610 ( .A1(n7600), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5153) );
  OR2_X1 U6611 ( .A1(n5157), .A2(n5247), .ZN(n5158) );
  XNOR2_X1 U6612 ( .A(n5158), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6319) );
  INV_X1 U6613 ( .A(n6319), .ZN(n6217) );
  XNOR2_X1 U6614 ( .A(n5160), .B(n5159), .ZN(n6224) );
  OR2_X1 U6615 ( .A1(n5104), .A2(n6224), .ZN(n5162) );
  OR2_X1 U6616 ( .A1(n7597), .A2(n6218), .ZN(n5161) );
  OAI211_X1 U6617 ( .C1(n6210), .C2(n6217), .A(n5162), .B(n5161), .ZN(n9740)
         );
  OAI22_X1 U6618 ( .A1(n6918), .A2(n5505), .B1(n9466), .B2(n5478), .ZN(n5163)
         );
  XOR2_X1 U6619 ( .A(n5508), .B(n5163), .Z(n5164) );
  OAI22_X1 U6620 ( .A1(n6918), .A2(n5319), .B1(n9466), .B2(n5505), .ZN(n6826)
         );
  NAND2_X1 U6621 ( .A1(n7601), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6622 ( .A1(n7587), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5170) );
  OAI21_X1 U6623 ( .B1(n5167), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5166), .ZN(
        n6923) );
  INV_X1 U6624 ( .A(n6923), .ZN(n9099) );
  NAND2_X1 U6625 ( .A1(n6181), .A2(n9099), .ZN(n5169) );
  NAND2_X1 U6626 ( .A1(n7600), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6627 ( .A1(n5172), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5173) );
  XNOR2_X1 U6628 ( .A(n5173), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6320) );
  INV_X1 U6629 ( .A(n6320), .ZN(n6374) );
  OR2_X1 U6630 ( .A1(n7597), .A2(n6222), .ZN(n5176) );
  INV_X1 U6631 ( .A(n4315), .ZN(n6924) );
  OAI22_X1 U6632 ( .A1(n6832), .A2(n5505), .B1(n6924), .B2(n5478), .ZN(n5177)
         );
  XNOR2_X1 U6633 ( .A(n5177), .B(n5508), .ZN(n5179) );
  OAI22_X1 U6634 ( .A1(n6832), .A2(n5319), .B1(n6924), .B2(n5505), .ZN(n5178)
         );
  OR2_X1 U6635 ( .A1(n5179), .A2(n5178), .ZN(n5181) );
  NAND2_X1 U6636 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  AND2_X1 U6637 ( .A1(n5181), .A2(n5180), .ZN(n9091) );
  NAND2_X1 U6638 ( .A1(n9090), .A2(n5181), .ZN(n6962) );
  XNOR2_X1 U6639 ( .A(n5183), .B(n5182), .ZN(n6963) );
  NAND2_X1 U6640 ( .A1(n7587), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6641 ( .A1(n7600), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6642 ( .A1(n7601), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5189) );
  OR2_X1 U6643 ( .A1(n5185), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6644 ( .A1(n5207), .A2(n5186), .ZN(n9682) );
  INV_X1 U6645 ( .A(n9682), .ZN(n5187) );
  NAND2_X1 U6646 ( .A1(n6181), .A2(n5187), .ZN(n5188) );
  OR2_X1 U6647 ( .A1(n7045), .A2(n5319), .ZN(n5199) );
  XNOR2_X1 U6648 ( .A(n5193), .B(n5192), .ZN(n6243) );
  NAND2_X1 U6649 ( .A1(n6243), .A2(n5245), .ZN(n5197) );
  NAND2_X1 U6650 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5195) );
  XNOR2_X1 U6651 ( .A(n5195), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6346) );
  AOI22_X1 U6652 ( .A1(n5397), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5396), .B2(
        n6346), .ZN(n5196) );
  NAND2_X1 U6653 ( .A1(n5197), .A2(n5196), .ZN(n7042) );
  NAND2_X1 U6654 ( .A1(n7042), .A2(n5229), .ZN(n5198) );
  NAND2_X1 U6655 ( .A1(n5199), .A2(n5198), .ZN(n7197) );
  INV_X1 U6656 ( .A(n7042), .ZN(n9676) );
  OAI22_X1 U6657 ( .A1(n7045), .A2(n5505), .B1(n9676), .B2(n5478), .ZN(n5200)
         );
  XNOR2_X1 U6658 ( .A(n5200), .B(n5508), .ZN(n9674) );
  XNOR2_X1 U6659 ( .A(n5201), .B(n4887), .ZN(n6247) );
  NAND2_X1 U6660 ( .A1(n6247), .A2(n5245), .ZN(n5205) );
  OR2_X1 U6661 ( .A1(n5202), .A2(n5247), .ZN(n5203) );
  XNOR2_X1 U6662 ( .A(n5203), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9138) );
  AOI22_X1 U6663 ( .A1(n5397), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5396), .B2(
        n9138), .ZN(n5204) );
  NAND2_X1 U6664 ( .A1(n7601), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6665 ( .A1(n7587), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6666 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  AND2_X1 U6667 ( .A1(n5223), .A2(n5208), .ZN(n7208) );
  NAND2_X1 U6668 ( .A1(n6181), .A2(n7208), .ZN(n5210) );
  NAND2_X1 U6669 ( .A1(n7600), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5209) );
  OAI22_X1 U6670 ( .A1(n9774), .A2(n5478), .B1(n7239), .B2(n5505), .ZN(n5213)
         );
  XNOR2_X1 U6671 ( .A(n5213), .B(n6188), .ZN(n7200) );
  OR2_X1 U6672 ( .A1(n9774), .A2(n5505), .ZN(n5215) );
  OR2_X1 U6673 ( .A1(n7239), .A2(n5319), .ZN(n5214) );
  NAND2_X1 U6674 ( .A1(n5215), .A2(n5214), .ZN(n7199) );
  INV_X1 U6675 ( .A(n7199), .ZN(n5216) );
  NAND2_X1 U6676 ( .A1(n7200), .A2(n5216), .ZN(n7259) );
  OAI21_X1 U6677 ( .B1(n7197), .B2(n9674), .A(n7259), .ZN(n5239) );
  AOI21_X1 U6678 ( .B1(n9674), .B2(n7197), .A(n7199), .ZN(n5236) );
  NAND3_X1 U6679 ( .A1(n9674), .A2(n7199), .A3(n7197), .ZN(n5235) );
  XNOR2_X1 U6680 ( .A(n5217), .B(n4886), .ZN(n6290) );
  NAND2_X1 U6681 ( .A1(n6290), .A2(n5245), .ZN(n5221) );
  OR2_X1 U6682 ( .A1(n5218), .A2(n5247), .ZN(n5219) );
  XNOR2_X1 U6683 ( .A(n5219), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6347) );
  AOI22_X1 U6684 ( .A1(n5397), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5396), .B2(
        n6347), .ZN(n5220) );
  NAND2_X1 U6685 ( .A1(n5221), .A2(n5220), .ZN(n9556) );
  NAND2_X1 U6686 ( .A1(n9556), .A2(n5222), .ZN(n5231) );
  NAND2_X1 U6687 ( .A1(n7587), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6688 ( .A1(n7601), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6689 ( .A1(n5223), .A2(n6401), .ZN(n5224) );
  AND2_X1 U6690 ( .A1(n5252), .A2(n5224), .ZN(n7270) );
  NAND2_X1 U6691 ( .A1(n6181), .A2(n7270), .ZN(n5226) );
  NAND2_X1 U6692 ( .A1(n7600), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5225) );
  INV_X1 U6693 ( .A(n7214), .ZN(n9125) );
  NAND2_X1 U6694 ( .A1(n9125), .A2(n5229), .ZN(n5230) );
  NAND2_X1 U6695 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  XNOR2_X1 U6696 ( .A(n5232), .B(n5508), .ZN(n5240) );
  NAND2_X1 U6697 ( .A1(n9556), .A2(n5229), .ZN(n5234) );
  NAND2_X1 U6698 ( .A1(n9125), .A2(n5532), .ZN(n5233) );
  NAND2_X1 U6699 ( .A1(n5234), .A2(n5233), .ZN(n5241) );
  NAND2_X1 U6700 ( .A1(n5240), .A2(n5241), .ZN(n7262) );
  OAI211_X1 U6701 ( .C1(n5236), .C2(n7200), .A(n5235), .B(n7262), .ZN(n5237)
         );
  INV_X1 U6702 ( .A(n5237), .ZN(n5238) );
  INV_X1 U6703 ( .A(n5240), .ZN(n5243) );
  INV_X1 U6704 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6705 ( .A1(n5243), .A2(n5242), .ZN(n7261) );
  NOR2_X1 U6706 ( .A1(n5014), .A2(n5247), .ZN(n5246) );
  MUX2_X1 U6707 ( .A(n5247), .B(n5246), .S(P1_IR_REG_11__SCAN_IN), .Z(n5248)
         );
  INV_X1 U6708 ( .A(n5248), .ZN(n5250) );
  INV_X1 U6709 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6710 ( .A1(n5014), .A2(n5249), .ZN(n5284) );
  AOI22_X1 U6711 ( .A1(n5397), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5396), .B2(
        n6470), .ZN(n5251) );
  NAND2_X1 U6712 ( .A1(n9651), .A2(n5222), .ZN(n5259) );
  AND2_X1 U6713 ( .A1(n5252), .A2(n6340), .ZN(n5253) );
  NOR2_X1 U6714 ( .A1(n5270), .A2(n5253), .ZN(n7217) );
  NAND2_X1 U6715 ( .A1(n5473), .A2(n7217), .ZN(n5257) );
  NAND2_X1 U6716 ( .A1(n7600), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6717 ( .A1(n7601), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6718 ( .A1(n7587), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5254) );
  NAND4_X1 U6719 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n9124)
         );
  NAND2_X1 U6720 ( .A1(n9124), .A2(n5229), .ZN(n5258) );
  NAND2_X1 U6721 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  XNOR2_X1 U6722 ( .A(n5260), .B(n5508), .ZN(n5262) );
  AND2_X1 U6723 ( .A1(n9124), .A2(n5532), .ZN(n5261) );
  AOI21_X1 U6724 ( .B1(n9651), .B2(n4333), .A(n5261), .ZN(n5263) );
  XNOR2_X1 U6725 ( .A(n5262), .B(n5263), .ZN(n7212) );
  NAND2_X1 U6726 ( .A1(n7213), .A2(n7212), .ZN(n7211) );
  INV_X1 U6727 ( .A(n5262), .ZN(n5264) );
  NAND2_X1 U6728 ( .A1(n7211), .A2(n4882), .ZN(n7301) );
  XNOR2_X1 U6729 ( .A(n5266), .B(n5265), .ZN(n6365) );
  NAND2_X1 U6730 ( .A1(n6365), .A2(n5245), .ZN(n5269) );
  NAND2_X1 U6731 ( .A1(n5284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5267) );
  XNOR2_X1 U6732 ( .A(n5267), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6580) );
  AOI22_X1 U6733 ( .A1(n5397), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5396), .B2(
        n6580), .ZN(n5268) );
  NAND2_X1 U6734 ( .A1(n5269), .A2(n5268), .ZN(n7375) );
  NAND2_X1 U6735 ( .A1(n7375), .A2(n5222), .ZN(n5277) );
  NAND2_X1 U6736 ( .A1(n7601), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6737 ( .A1(n5571), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6738 ( .A1(n5270), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6739 ( .A1(n5271), .A2(n5288), .ZN(n7302) );
  NAND2_X1 U6740 ( .A1(n5473), .A2(n7302), .ZN(n5273) );
  NAND2_X1 U6741 ( .A1(n7600), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6742 ( .A1(n9123), .A2(n5229), .ZN(n5276) );
  NAND2_X1 U6743 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  XNOR2_X1 U6744 ( .A(n5278), .B(n6188), .ZN(n7298) );
  NOR2_X1 U6745 ( .A1(n7225), .A2(n5319), .ZN(n5279) );
  AOI21_X1 U6746 ( .B1(n7375), .B2(n4333), .A(n5279), .ZN(n7299) );
  NAND2_X1 U6747 ( .A1(n7298), .A2(n7299), .ZN(n5281) );
  NOR2_X1 U6748 ( .A1(n7298), .A2(n7299), .ZN(n5280) );
  XNOR2_X1 U6749 ( .A(n5283), .B(n5282), .ZN(n6479) );
  NAND2_X1 U6750 ( .A1(n6479), .A2(n5245), .ZN(n5286) );
  NOR2_X1 U6751 ( .A1(n5284), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5325) );
  OR2_X1 U6752 ( .A1(n5325), .A2(n5247), .ZN(n5306) );
  XNOR2_X1 U6753 ( .A(n5306), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U6754 ( .A1(n5397), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5396), .B2(
        n6856), .ZN(n5285) );
  NAND2_X1 U6755 ( .A1(n7421), .A2(n5222), .ZN(n5295) );
  NAND2_X1 U6756 ( .A1(n7600), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6757 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  AND2_X1 U6758 ( .A1(n5312), .A2(n5289), .ZN(n7432) );
  NAND2_X1 U6759 ( .A1(n5473), .A2(n7432), .ZN(n5292) );
  NAND2_X1 U6760 ( .A1(n5571), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6761 ( .A1(n7601), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5290) );
  NAND4_X1 U6762 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n9122)
         );
  NAND2_X1 U6763 ( .A1(n9122), .A2(n4333), .ZN(n5294) );
  NAND2_X1 U6764 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  XNOR2_X1 U6765 ( .A(n5296), .B(n5508), .ZN(n5299) );
  NAND2_X1 U6766 ( .A1(n7421), .A2(n4333), .ZN(n5298) );
  NAND2_X1 U6767 ( .A1(n9122), .A2(n5532), .ZN(n5297) );
  NAND2_X1 U6768 ( .A1(n5298), .A2(n5297), .ZN(n5300) );
  NAND2_X1 U6769 ( .A1(n5299), .A2(n5300), .ZN(n7425) );
  INV_X1 U6770 ( .A(n5299), .ZN(n5302) );
  INV_X1 U6771 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U6772 ( .A1(n5302), .A2(n5301), .ZN(n7424) );
  XNOR2_X1 U6773 ( .A(n5304), .B(n5303), .ZN(n6560) );
  NAND2_X1 U6774 ( .A1(n6560), .A2(n5245), .ZN(n5311) );
  NAND2_X1 U6775 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  NAND2_X1 U6776 ( .A1(n5307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5309) );
  INV_X1 U6777 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5308) );
  XNOR2_X1 U6778 ( .A(n5309), .B(n5308), .ZN(n7028) );
  INV_X1 U6779 ( .A(n7028), .ZN(n7036) );
  AOI22_X1 U6780 ( .A1(n5397), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5396), .B2(
        n7036), .ZN(n5310) );
  NAND2_X1 U6781 ( .A1(n5311), .A2(n5310), .ZN(n7333) );
  AND2_X1 U6782 ( .A1(n5312), .A2(n9002), .ZN(n5313) );
  NOR2_X1 U6783 ( .A1(n5331), .A2(n5313), .ZN(n9006) );
  NAND2_X1 U6784 ( .A1(n5077), .A2(n9006), .ZN(n5317) );
  NAND2_X1 U6785 ( .A1(n5571), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6786 ( .A1(n7600), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6787 ( .A1(n7601), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5314) );
  OAI22_X1 U6788 ( .A1(n9642), .A2(n5478), .B1(n7430), .B2(n5505), .ZN(n5318)
         );
  XOR2_X1 U6789 ( .A(n5508), .B(n5318), .Z(n5320) );
  OAI22_X1 U6790 ( .A1(n9642), .A2(n5505), .B1(n7430), .B2(n5319), .ZN(n9001)
         );
  INV_X1 U6791 ( .A(n5320), .ZN(n5321) );
  XNOR2_X1 U6792 ( .A(n5323), .B(n5322), .ZN(n6611) );
  NAND2_X1 U6793 ( .A1(n6611), .A2(n5245), .ZN(n5330) );
  NOR2_X1 U6794 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5324) );
  NAND2_X1 U6795 ( .A1(n5325), .A2(n5324), .ZN(n5327) );
  NAND2_X1 U6796 ( .A1(n5327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5326) );
  MUX2_X1 U6797 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5326), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5328) );
  AOI22_X1 U6798 ( .A1(n5397), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5396), .B2(
        n7153), .ZN(n5329) );
  NAND2_X1 U6799 ( .A1(n5330), .A2(n5329), .ZN(n9197) );
  NAND2_X1 U6800 ( .A1(n5571), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5336) );
  NOR2_X1 U6801 ( .A1(n5331), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5332) );
  OR2_X1 U6802 ( .A1(n5348), .A2(n5332), .ZN(n9113) );
  INV_X1 U6803 ( .A(n9113), .ZN(n7345) );
  NAND2_X1 U6804 ( .A1(n5473), .A2(n7345), .ZN(n5335) );
  NAND2_X1 U6805 ( .A1(n7600), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6806 ( .A1(n7601), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5333) );
  NAND4_X1 U6807 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n9196)
         );
  OAI22_X1 U6808 ( .A1(n9634), .A2(n5478), .B1(n9437), .B2(n5505), .ZN(n5337)
         );
  XNOR2_X1 U6809 ( .A(n5337), .B(n5508), .ZN(n5339) );
  OAI22_X1 U6810 ( .A1(n9634), .A2(n5505), .B1(n9437), .B2(n5319), .ZN(n9107)
         );
  NAND2_X1 U6811 ( .A1(n9104), .A2(n9107), .ZN(n5341) );
  NAND2_X1 U6812 ( .A1(n5340), .A2(n5339), .ZN(n9105) );
  XNOR2_X1 U6813 ( .A(n5343), .B(n5342), .ZN(n6615) );
  NAND2_X1 U6814 ( .A1(n6615), .A2(n5245), .ZN(n5347) );
  NAND2_X1 U6815 ( .A1(n5344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U6816 ( .A(n5345), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9148) );
  AOI22_X1 U6817 ( .A1(n5397), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5396), .B2(
        n9148), .ZN(n5346) );
  NAND2_X1 U6818 ( .A1(n7587), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6819 ( .A1(n7601), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5352) );
  OR2_X1 U6820 ( .A1(n5348), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5349) );
  AND2_X1 U6821 ( .A1(n5368), .A2(n5349), .ZN(n9445) );
  NAND2_X1 U6822 ( .A1(n5473), .A2(n9445), .ZN(n5351) );
  NAND2_X1 U6823 ( .A1(n7600), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5350) );
  NOR2_X1 U6824 ( .A1(n9108), .A2(n5319), .ZN(n5354) );
  AOI21_X1 U6825 ( .B1(n9552), .B2(n4333), .A(n5354), .ZN(n5359) );
  NAND2_X1 U6826 ( .A1(n9552), .A2(n5222), .ZN(n5356) );
  NAND2_X1 U6827 ( .A1(n9424), .A2(n4333), .ZN(n5355) );
  NAND2_X1 U6828 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  XNOR2_X1 U6829 ( .A(n5357), .B(n5508), .ZN(n5358) );
  XOR2_X1 U6830 ( .A(n5359), .B(n5358), .Z(n9036) );
  INV_X1 U6831 ( .A(n5358), .ZN(n5360) );
  NAND2_X1 U6832 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  XNOR2_X1 U6833 ( .A(n5363), .B(n5362), .ZN(n6627) );
  NAND2_X1 U6834 ( .A1(n6627), .A2(n5245), .ZN(n5366) );
  XNOR2_X1 U6835 ( .A(n5364), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9171) );
  AOI22_X1 U6836 ( .A1(n5397), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5396), .B2(
        n9171), .ZN(n5365) );
  NAND2_X1 U6837 ( .A1(n7587), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6838 ( .A1(n7600), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6839 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  AND2_X1 U6840 ( .A1(n5385), .A2(n5369), .ZN(n9419) );
  NAND2_X1 U6841 ( .A1(n6181), .A2(n9419), .ZN(n5371) );
  NAND2_X1 U6842 ( .A1(n7601), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5370) );
  OAI22_X1 U6843 ( .A1(n9421), .A2(n5478), .B1(n9439), .B2(n5505), .ZN(n5374)
         );
  XNOR2_X1 U6844 ( .A(n5374), .B(n5508), .ZN(n5375) );
  AOI22_X1 U6845 ( .A1(n9545), .A2(n4333), .B1(n5532), .B2(n9403), .ZN(n5376)
         );
  XNOR2_X1 U6846 ( .A(n5375), .B(n5376), .ZN(n9045) );
  INV_X1 U6847 ( .A(n5375), .ZN(n5377) );
  XNOR2_X1 U6848 ( .A(n5379), .B(n5378), .ZN(n6823) );
  NAND2_X1 U6849 ( .A1(n6823), .A2(n5245), .ZN(n5384) );
  INV_X1 U6850 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6851 ( .A1(n5364), .A2(n5380), .ZN(n5381) );
  NAND2_X1 U6852 ( .A1(n5381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5382) );
  XNOR2_X1 U6853 ( .A(n5382), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U6854 ( .A1(n5397), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5396), .B2(
        n9699), .ZN(n5383) );
  NAND2_X1 U6855 ( .A1(n7601), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6856 ( .A1(n7587), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5389) );
  AND2_X1 U6857 ( .A1(n5385), .A2(n9084), .ZN(n5386) );
  NOR2_X1 U6858 ( .A1(n5402), .A2(n5386), .ZN(n9406) );
  NAND2_X1 U6859 ( .A1(n6181), .A2(n9406), .ZN(n5388) );
  NAND2_X1 U6860 ( .A1(n7600), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5387) );
  AOI22_X1 U6861 ( .A1(n9539), .A2(n5222), .B1(n4333), .B2(n9425), .ZN(n5391)
         );
  XOR2_X1 U6862 ( .A(n5508), .B(n5391), .Z(n5392) );
  INV_X1 U6863 ( .A(n9539), .ZN(n9408) );
  OAI22_X1 U6864 ( .A1(n9408), .A2(n5505), .B1(n9048), .B2(n5319), .ZN(n9083)
         );
  NAND2_X1 U6865 ( .A1(n9081), .A2(n9083), .ZN(n5393) );
  NAND2_X1 U6866 ( .A1(n4349), .A2(n5392), .ZN(n9080) );
  XNOR2_X1 U6867 ( .A(n5395), .B(n5394), .ZN(n6865) );
  NAND2_X1 U6868 ( .A1(n6865), .A2(n5245), .ZN(n5399) );
  AOI22_X1 U6869 ( .A1(n5397), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5396), .B2(
        n9315), .ZN(n5398) );
  NAND2_X1 U6870 ( .A1(n7587), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6871 ( .A1(n7601), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6872 ( .A1(n5401), .A2(n5400), .ZN(n5406) );
  NOR2_X1 U6873 ( .A1(n5402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5403) );
  OR2_X1 U6874 ( .A1(n5413), .A2(n5403), .ZN(n9385) );
  INV_X1 U6875 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8325) );
  OAI22_X1 U6876 ( .A1(n9385), .A2(n5417), .B1(n5404), .B2(n8325), .ZN(n5405)
         );
  OAI22_X1 U6877 ( .A1(n9388), .A2(n5478), .B1(n9199), .B2(n5505), .ZN(n5407)
         );
  XNOR2_X1 U6878 ( .A(n5407), .B(n5508), .ZN(n5408) );
  INV_X1 U6879 ( .A(n5408), .ZN(n8068) );
  OAI22_X1 U6880 ( .A1(n9388), .A2(n5505), .B1(n9199), .B2(n5319), .ZN(n8067)
         );
  XNOR2_X1 U6881 ( .A(n5410), .B(n5409), .ZN(n6991) );
  NAND2_X1 U6882 ( .A1(n6991), .A2(n5245), .ZN(n5412) );
  OR2_X1 U6883 ( .A1(n7597), .A2(n8304), .ZN(n5411) );
  NAND2_X1 U6884 ( .A1(n9528), .A2(n5222), .ZN(n5419) );
  NOR2_X1 U6885 ( .A1(n5413), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5414) );
  OR2_X1 U6886 ( .A1(n5428), .A2(n5414), .ZN(n9371) );
  AOI22_X1 U6887 ( .A1(n7587), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n7600), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6888 ( .A1(n7601), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U6889 ( .C1(n9371), .C2(n5417), .A(n5416), .B(n5415), .ZN(n9394)
         );
  NAND2_X1 U6890 ( .A1(n9394), .A2(n4333), .ZN(n5418) );
  NAND2_X1 U6891 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  XNOR2_X1 U6892 ( .A(n5420), .B(n6188), .ZN(n5423) );
  AND2_X1 U6893 ( .A1(n9394), .A2(n5532), .ZN(n5421) );
  AOI21_X1 U6894 ( .B1(n9528), .B2(n4333), .A(n5421), .ZN(n5422) );
  NAND2_X1 U6895 ( .A1(n5423), .A2(n5422), .ZN(n9061) );
  NOR2_X1 U6896 ( .A1(n5423), .A2(n5422), .ZN(n9063) );
  XNOR2_X1 U6897 ( .A(n5425), .B(n5424), .ZN(n7058) );
  NAND2_X1 U6898 ( .A1(n7058), .A2(n5245), .ZN(n5427) );
  INV_X1 U6899 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7059) );
  OR2_X1 U6900 ( .A1(n7597), .A2(n7059), .ZN(n5426) );
  NAND2_X1 U6901 ( .A1(n9525), .A2(n5222), .ZN(n5435) );
  OR2_X1 U6902 ( .A1(n5428), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5430) );
  AND2_X1 U6903 ( .A1(n5430), .A2(n5429), .ZN(n9359) );
  NAND2_X1 U6904 ( .A1(n9359), .A2(n5473), .ZN(n5433) );
  AOI22_X1 U6905 ( .A1(n7587), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n7601), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6906 ( .A1(n7600), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6907 ( .A1(n9201), .A2(n5505), .ZN(n5434) );
  NAND2_X1 U6908 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  XNOR2_X1 U6909 ( .A(n5436), .B(n6188), .ZN(n5439) );
  NOR2_X1 U6910 ( .A1(n9201), .A2(n5319), .ZN(n5437) );
  AOI21_X1 U6911 ( .B1(n9525), .B2(n4333), .A(n5437), .ZN(n5438) );
  OR2_X1 U6912 ( .A1(n5439), .A2(n5438), .ZN(n9021) );
  NAND2_X1 U6913 ( .A1(n5439), .A2(n5438), .ZN(n9020) );
  OAI22_X1 U6914 ( .A1(n9341), .A2(n5478), .B1(n9356), .B2(n5505), .ZN(n5440)
         );
  XNOR2_X1 U6915 ( .A(n5440), .B(n5508), .ZN(n9071) );
  AND2_X1 U6916 ( .A1(n9020), .A2(n9071), .ZN(n5441) );
  NAND2_X1 U6917 ( .A1(n5442), .A2(n5441), .ZN(n5445) );
  INV_X1 U6918 ( .A(n9071), .ZN(n5443) );
  OR2_X1 U6919 ( .A1(n5443), .A2(n9072), .ZN(n5444) );
  MUX2_X1 U6920 ( .A(n7258), .B(n7255), .S(n4409), .Z(n5450) );
  INV_X1 U6921 ( .A(SI_23_), .ZN(n5449) );
  NAND2_X1 U6922 ( .A1(n5450), .A2(n5449), .ZN(n5465) );
  INV_X1 U6923 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6924 ( .A1(n5451), .A2(SI_23_), .ZN(n5452) );
  XNOR2_X1 U6925 ( .A(n5464), .B(n5463), .ZN(n7256) );
  NAND2_X1 U6926 ( .A1(n7256), .A2(n5245), .ZN(n5454) );
  OR2_X1 U6927 ( .A1(n7597), .A2(n7255), .ZN(n5453) );
  NAND2_X1 U6928 ( .A1(n7587), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6929 ( .A1(n7601), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5460) );
  INV_X1 U6930 ( .A(n5456), .ZN(n5455) );
  NAND2_X1 U6931 ( .A1(n5455), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5471) );
  INV_X1 U6932 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U6933 ( .A1(n5456), .A2(n9014), .ZN(n5457) );
  AND2_X1 U6934 ( .A1(n5471), .A2(n5457), .ZN(n9324) );
  NAND2_X1 U6935 ( .A1(n5473), .A2(n9324), .ZN(n5459) );
  NAND2_X1 U6936 ( .A1(n7600), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5458) );
  OAI22_X1 U6937 ( .A1(n9326), .A2(n5478), .B1(n9309), .B2(n5505), .ZN(n5462)
         );
  XNOR2_X1 U6938 ( .A(n5462), .B(n5508), .ZN(n9009) );
  OAI22_X1 U6939 ( .A1(n9326), .A2(n5505), .B1(n9309), .B2(n5319), .ZN(n9010)
         );
  NAND2_X1 U6940 ( .A1(n5464), .A2(n5463), .ZN(n5466) );
  INV_X1 U6941 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7353) );
  INV_X1 U6942 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7351) );
  MUX2_X1 U6943 ( .A(n7353), .B(n7351), .S(n4409), .Z(n5488) );
  XNOR2_X1 U6944 ( .A(n5488), .B(SI_24_), .ZN(n5485) );
  XNOR2_X1 U6945 ( .A(n5487), .B(n5485), .ZN(n7350) );
  NAND2_X1 U6946 ( .A1(n7350), .A2(n5245), .ZN(n5468) );
  OR2_X1 U6947 ( .A1(n7597), .A2(n7351), .ZN(n5467) );
  NAND2_X1 U6948 ( .A1(n5571), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6949 ( .A1(n7601), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5476) );
  INV_X1 U6950 ( .A(n5471), .ZN(n5469) );
  NAND2_X1 U6951 ( .A1(n5469), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5499) );
  INV_X1 U6952 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6953 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  AND2_X1 U6954 ( .A1(n5499), .A2(n5472), .ZN(n9313) );
  NAND2_X1 U6955 ( .A1(n5473), .A2(n9313), .ZN(n5475) );
  NAND2_X1 U6956 ( .A1(n7600), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5474) );
  OAI22_X1 U6957 ( .A1(n9206), .A2(n5478), .B1(n9330), .B2(n5505), .ZN(n5479)
         );
  XNOR2_X1 U6958 ( .A(n5479), .B(n6188), .ZN(n5483) );
  OR2_X1 U6959 ( .A1(n9206), .A2(n5505), .ZN(n5481) );
  NAND2_X1 U6960 ( .A1(n9207), .A2(n5532), .ZN(n5480) );
  NAND2_X1 U6961 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  OAI21_X1 U6962 ( .B1(n5483), .B2(n5482), .A(n5484), .ZN(n9053) );
  INV_X1 U6963 ( .A(n5485), .ZN(n5486) );
  INV_X1 U6964 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U6965 ( .A1(n5489), .A2(SI_24_), .ZN(n5490) );
  INV_X1 U6966 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7452) );
  INV_X1 U6967 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7455) );
  MUX2_X1 U6968 ( .A(n7452), .B(n7455), .S(n4409), .Z(n5492) );
  NAND2_X1 U6969 ( .A1(n5492), .A2(n5491), .ZN(n5514) );
  INV_X1 U6970 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U6971 ( .A1(n5493), .A2(SI_25_), .ZN(n5494) );
  NAND2_X1 U6972 ( .A1(n5514), .A2(n5494), .ZN(n5513) );
  NAND2_X1 U6973 ( .A1(n7450), .A2(n5245), .ZN(n5496) );
  OR2_X1 U6974 ( .A1(n7597), .A2(n7455), .ZN(n5495) );
  NAND2_X1 U6975 ( .A1(n7601), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U6976 ( .A1(n7587), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5503) );
  INV_X1 U6977 ( .A(n5499), .ZN(n5497) );
  NAND2_X1 U6978 ( .A1(n5497), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5523) );
  INV_X1 U6979 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6980 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AND2_X1 U6981 ( .A1(n5523), .A2(n5500), .ZN(n9297) );
  NAND2_X1 U6982 ( .A1(n6181), .A2(n9297), .ZN(n5502) );
  NAND2_X1 U6983 ( .A1(n7600), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5501) );
  OAI22_X1 U6984 ( .A1(n9208), .A2(n5505), .B1(n9310), .B2(n5319), .ZN(n5510)
         );
  NAND2_X1 U6985 ( .A1(n9505), .A2(n5222), .ZN(n5507) );
  OR2_X1 U6986 ( .A1(n9310), .A2(n5505), .ZN(n5506) );
  NAND2_X1 U6987 ( .A1(n5507), .A2(n5506), .ZN(n5509) );
  XNOR2_X1 U6988 ( .A(n5509), .B(n5508), .ZN(n5511) );
  XOR2_X1 U6989 ( .A(n5510), .B(n5511), .Z(n9030) );
  INV_X1 U6990 ( .A(n5538), .ZN(n5534) );
  NOR2_X1 U6991 ( .A1(n5511), .A2(n5510), .ZN(n5535) );
  INV_X1 U6992 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7503) );
  MUX2_X1 U6993 ( .A(n7503), .B(n7804), .S(n4409), .Z(n5516) );
  INV_X1 U6994 ( .A(SI_26_), .ZN(n5515) );
  NAND2_X1 U6995 ( .A1(n5516), .A2(n5515), .ZN(n6060) );
  INV_X1 U6996 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U6997 ( .A1(n5517), .A2(SI_26_), .ZN(n5518) );
  XNOR2_X1 U6998 ( .A(n6059), .B(n6058), .ZN(n7502) );
  NAND2_X1 U6999 ( .A1(n7502), .A2(n5245), .ZN(n5520) );
  OR2_X1 U7000 ( .A1(n7597), .A2(n7804), .ZN(n5519) );
  NAND2_X1 U7001 ( .A1(n9498), .A2(n5222), .ZN(n5530) );
  INV_X1 U7002 ( .A(n5523), .ZN(n5521) );
  NAND2_X1 U7003 ( .A1(n5521), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5574) );
  INV_X1 U7004 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7005 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  AND2_X1 U7006 ( .A1(n5574), .A2(n5524), .ZN(n9279) );
  NAND2_X1 U7007 ( .A1(n6181), .A2(n9279), .ZN(n5528) );
  NAND2_X1 U7008 ( .A1(n7600), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7009 ( .A1(n5571), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7010 ( .A1(n7601), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5525) );
  NAND4_X1 U7011 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n9272)
         );
  NAND2_X1 U7012 ( .A1(n9272), .A2(n4333), .ZN(n5529) );
  NAND2_X1 U7013 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  XNOR2_X1 U7014 ( .A(n5531), .B(n6188), .ZN(n6161) );
  AND2_X1 U7015 ( .A1(n9272), .A2(n5532), .ZN(n5533) );
  AOI21_X1 U7016 ( .B1(n9498), .B2(n4333), .A(n5533), .ZN(n6162) );
  XNOR2_X1 U7017 ( .A(n6161), .B(n6162), .ZN(n5536) );
  OAI21_X1 U7018 ( .B1(n5534), .B2(n5535), .A(n5536), .ZN(n5588) );
  NOR2_X1 U7019 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  NAND3_X1 U7020 ( .A1(n7453), .A2(P1_B_REG_SCAN_IN), .A3(n7352), .ZN(n5540)
         );
  OAI21_X1 U7021 ( .B1(P1_B_REG_SCAN_IN), .B2(n7352), .A(n5540), .ZN(n5541) );
  INV_X1 U7022 ( .A(n6664), .ZN(n6667) );
  INV_X1 U7023 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7024 ( .A1(n6667), .A2(n5542), .ZN(n5543) );
  NAND2_X1 U7025 ( .A1(n5539), .A2(n7352), .ZN(n9581) );
  NOR4_X1 U7026 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5547) );
  NOR4_X1 U7027 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5546) );
  NOR4_X1 U7028 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n5545) );
  NOR4_X1 U7029 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5544) );
  NAND4_X1 U7030 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n5553)
         );
  NOR2_X1 U7031 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .ZN(
        n5551) );
  NOR4_X1 U7032 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5550) );
  NOR4_X1 U7033 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5549) );
  NOR4_X1 U7034 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5548) );
  NAND4_X1 U7035 ( .A1(n5551), .A2(n5550), .A3(n5549), .A4(n5548), .ZN(n5552)
         );
  NOR2_X1 U7036 ( .A1(n5553), .A2(n5552), .ZN(n6663) );
  AND2_X1 U7037 ( .A1(n6663), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7038 ( .A1(n5539), .A2(n7453), .ZN(n6668) );
  OAI21_X1 U7039 ( .B1(n6664), .B2(n5554), .A(n6668), .ZN(n5555) );
  INV_X1 U7040 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7041 ( .A1(n7388), .A2(n5556), .ZN(n5580) );
  NAND2_X1 U7042 ( .A1(n4397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5558) );
  INV_X1 U7043 ( .A(n6240), .ZN(n5559) );
  NAND2_X1 U7044 ( .A1(n9773), .A2(n7753), .ZN(n5560) );
  NAND2_X1 U7045 ( .A1(n5567), .A2(n9465), .ZN(n9677) );
  NAND2_X1 U7046 ( .A1(n5580), .A2(n9773), .ZN(n5562) );
  NAND3_X1 U7047 ( .A1(n5562), .A2(n6490), .A3(n6286), .ZN(n5563) );
  NAND2_X1 U7048 ( .A1(n5563), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5566) );
  NOR2_X1 U7049 ( .A1(n9561), .A2(n7792), .ZN(n6679) );
  AND2_X1 U7050 ( .A1(n6679), .A2(n6240), .ZN(n5564) );
  OR2_X1 U7051 ( .A1(n6284), .A2(P1_U3084), .ZN(n7798) );
  INV_X1 U7052 ( .A(n7798), .ZN(n7793) );
  AOI21_X1 U7053 ( .B1(n5580), .B2(n5564), .A(n7793), .ZN(n5565) );
  INV_X1 U7054 ( .A(n5567), .ZN(n5569) );
  NAND2_X1 U7055 ( .A1(n5569), .A2(n5568), .ZN(n9667) );
  INV_X1 U7056 ( .A(n7753), .ZN(n6688) );
  NAND2_X1 U7057 ( .A1(n5571), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7058 ( .A1(n7600), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5578) );
  INV_X1 U7059 ( .A(n5574), .ZN(n5572) );
  NAND2_X1 U7060 ( .A1(n5572), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6179) );
  INV_X1 U7061 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7062 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  NAND2_X1 U7063 ( .A1(n5473), .A2(n9267), .ZN(n5577) );
  NAND2_X1 U7064 ( .A1(n7601), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5576) );
  INV_X1 U7065 ( .A(n5580), .ZN(n5582) );
  NAND2_X1 U7066 ( .A1(n6240), .A2(n6490), .ZN(n7797) );
  NOR2_X1 U7067 ( .A1(n7797), .A2(n9438), .ZN(n5581) );
  AOI22_X1 U7068 ( .A1(n9209), .A2(n9111), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n5583) );
  OAI21_X1 U7069 ( .B1(n9096), .B2(n7530), .A(n5583), .ZN(n5584) );
  AOI21_X1 U7070 ( .B1(n9279), .B2(n9100), .A(n5584), .ZN(n5585) );
  INV_X1 U7071 ( .A(n5589), .ZN(P1_U3238) );
  AND2_X2 U7072 ( .A1(n5768), .A2(n5593), .ZN(n5627) );
  NOR2_X1 U7073 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5597) );
  NOR2_X1 U7074 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5596) );
  NOR2_X1 U7075 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5595) );
  NOR2_X1 U7076 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5594) );
  NAND4_X1 U7077 ( .A1(n5597), .A2(n5596), .A3(n5595), .A4(n5594), .ZN(n5600)
         );
  NAND4_X1 U7078 ( .A1(n5598), .A2(n5888), .A3(n5837), .A4(n5822), .ZN(n5599)
         );
  NAND2_X1 U7079 ( .A1(n6084), .A2(n5603), .ZN(n5647) );
  INV_X1 U7080 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5604) );
  INV_X1 U7081 ( .A(n5606), .ZN(n8977) );
  NAND2_X1 U7082 ( .A1(n5607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5608) );
  MUX2_X1 U7083 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5608), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5609) );
  NAND2_X1 U7084 ( .A1(n6021), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7085 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5740) );
  INV_X1 U7086 ( .A(n5740), .ZN(n5610) );
  NAND2_X1 U7087 ( .A1(n5610), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5775) );
  INV_X1 U7088 ( .A(n5775), .ZN(n5612) );
  AND2_X1 U7089 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5611) );
  NAND2_X1 U7090 ( .A1(n5612), .A2(n5611), .ZN(n5793) );
  INV_X1 U7091 ( .A(n5793), .ZN(n5613) );
  NAND2_X1 U7092 ( .A1(n5613), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5808) );
  INV_X1 U7093 ( .A(n5827), .ZN(n5614) );
  NAND2_X1 U7094 ( .A1(n5614), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7095 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5615) );
  INV_X1 U7096 ( .A(n5878), .ZN(n5616) );
  NAND2_X1 U7097 ( .A1(n5616), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5894) );
  INV_X1 U7098 ( .A(n5917), .ZN(n5617) );
  NAND2_X1 U7099 ( .A1(n5617), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5933) );
  INV_X1 U7100 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7101 ( .A1(n5917), .A2(n5618), .ZN(n5619) );
  NAND2_X1 U7102 ( .A1(n5933), .A2(n5619), .ZN(n8133) );
  OR2_X1 U7103 ( .A1(n7824), .A2(n8133), .ZN(n5625) );
  INV_X1 U7104 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8508) );
  OR2_X1 U7105 ( .A1(n7854), .A2(n8508), .ZN(n5624) );
  INV_X1 U7106 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5622) );
  OR2_X1 U7107 ( .A1(n7858), .A2(n5622), .ZN(n5623) );
  NAND4_X1 U7108 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .ZN(n8584)
         );
  INV_X1 U7109 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7110 ( .A1(n5804), .A2(n5629), .ZN(n5853) );
  NAND3_X1 U7111 ( .A1(n5888), .A2(n5908), .A3(n5632), .ZN(n5633) );
  NAND2_X1 U7112 ( .A1(n5650), .A2(n5634), .ZN(n5928) );
  INV_X1 U7113 ( .A(n8063), .ZN(n7123) );
  NAND2_X1 U7114 ( .A1(n5639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7115 ( .A1(n5642), .A2(n5641), .ZN(n5644) );
  NAND2_X1 U7116 ( .A1(n8584), .A2(n5678), .ZN(n5923) );
  INV_X1 U7117 ( .A(n5923), .ZN(n5927) );
  INV_X2 U7118 ( .A(n5767), .ZN(n5790) );
  NAND2_X1 U7119 ( .A1(n6615), .A2(n5790), .ZN(n5653) );
  OR2_X1 U7120 ( .A1(n5650), .A2(n5604), .ZN(n5651) );
  XNOR2_X1 U7121 ( .A(n5651), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8532) );
  AOI22_X1 U7122 ( .A1(n5964), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6252), .B2(
        n8532), .ZN(n5652) );
  NAND2_X1 U7123 ( .A1(n5654), .A2(n8063), .ZN(n7891) );
  XNOR2_X1 U7124 ( .A(n8933), .B(n5679), .ZN(n5926) );
  INV_X1 U7125 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U7126 ( .A1(n5703), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5655) );
  INV_X1 U7127 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6511) );
  OR2_X1 U7128 ( .A1(n7854), .A2(n6511), .ZN(n5658) );
  INV_X1 U7129 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6707) );
  OR2_X1 U7130 ( .A1(n5721), .A2(n6707), .ZN(n5657) );
  NAND3_X2 U7131 ( .A1(n5659), .A2(n5658), .A3(n5657), .ZN(n6697) );
  OR2_X1 U7132 ( .A1(n5767), .A2(n6219), .ZN(n5664) );
  INV_X1 U7133 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7134 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5660) );
  OR2_X1 U7135 ( .A1(n5662), .A2(n9599), .ZN(n5663) );
  NAND2_X1 U7136 ( .A1(n5666), .A2(n5667), .ZN(n5681) );
  INV_X1 U7137 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5670) );
  OR2_X1 U7138 ( .A1(n5704), .A2(n5670), .ZN(n5676) );
  INV_X1 U7139 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5671) );
  INV_X1 U7140 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9925) );
  INV_X1 U7141 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U7142 ( .A1(n6214), .A2(SI_0_), .ZN(n5677) );
  XNOR2_X1 U7143 ( .A(n5677), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8988) );
  MUX2_X1 U7144 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8988), .S(n5662), .Z(n8082) );
  NOR2_X1 U7145 ( .A1(n5679), .A2(n8082), .ZN(n5680) );
  AOI21_X1 U7146 ( .B1(n6871), .B2(n5678), .A(n5680), .ZN(n6497) );
  INV_X1 U7147 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6231) );
  OR2_X1 U7148 ( .A1(n7859), .A2(n6231), .ZN(n5689) );
  OR2_X1 U7149 ( .A1(n5767), .A2(n6232), .ZN(n5688) );
  NOR2_X1 U7150 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5684) );
  INV_X1 U7151 ( .A(n5684), .ZN(n5682) );
  NAND2_X1 U7152 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5682), .ZN(n5683) );
  INV_X1 U7153 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5685) );
  MUX2_X1 U7154 ( .A(n5683), .B(P2_IR_REG_31__SCAN_IN), .S(n5685), .Z(n5686)
         );
  NAND2_X1 U7155 ( .A1(n5685), .A2(n5684), .ZN(n5699) );
  NAND2_X1 U7156 ( .A1(n5686), .A2(n5699), .ZN(n6535) );
  OR2_X1 U7157 ( .A1(n5662), .A2(n6535), .ZN(n5687) );
  AND3_X2 U7158 ( .A1(n5689), .A2(n5688), .A3(n5687), .ZN(n9862) );
  XNOR2_X1 U7159 ( .A(n5679), .B(n9862), .ZN(n5698) );
  INV_X1 U7160 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6512) );
  OR2_X1 U7161 ( .A1(n7854), .A2(n6512), .ZN(n5696) );
  INV_X1 U7162 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5690) );
  OR2_X1 U7163 ( .A1(n5704), .A2(n5690), .ZN(n5695) );
  INV_X1 U7164 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5691) );
  INV_X1 U7165 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6534) );
  OR2_X1 U7166 ( .A1(n5721), .A2(n6534), .ZN(n5692) );
  NAND2_X1 U7167 ( .A1(n8394), .A2(n5678), .ZN(n5697) );
  XNOR2_X1 U7168 ( .A(n5698), .B(n5697), .ZN(n6554) );
  NAND2_X1 U7169 ( .A1(n5699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5700) );
  XNOR2_X1 U7170 ( .A(n5700), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8401) );
  INV_X1 U7171 ( .A(n8401), .ZN(n6235) );
  OR2_X1 U7172 ( .A1(n7859), .A2(n6233), .ZN(n5702) );
  OR2_X1 U7173 ( .A1(n5767), .A2(n6234), .ZN(n5701) );
  OAI211_X1 U7174 ( .C1(n5662), .C2(n6235), .A(n5702), .B(n5701), .ZN(n6869)
         );
  XNOR2_X1 U7175 ( .A(n5679), .B(n6869), .ZN(n5712) );
  NAND2_X1 U7176 ( .A1(n5703), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5710) );
  OR2_X1 U7177 ( .A1(n5704), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5709) );
  INV_X1 U7178 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5705) );
  OR2_X1 U7179 ( .A1(n7854), .A2(n5705), .ZN(n5708) );
  INV_X1 U7180 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5706) );
  OR2_X1 U7181 ( .A1(n5721), .A2(n5706), .ZN(n5707) );
  NAND2_X1 U7182 ( .A1(n8393), .A2(n5678), .ZN(n5711) );
  XNOR2_X1 U7183 ( .A(n5712), .B(n5711), .ZN(n6588) );
  INV_X1 U7184 ( .A(n5711), .ZN(n5713) );
  NAND2_X1 U7185 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  OR2_X1 U7186 ( .A1(n5767), .A2(n6229), .ZN(n5719) );
  OR2_X1 U7187 ( .A1(n7859), .A2(n6230), .ZN(n5718) );
  OR2_X1 U7188 ( .A1(n5715), .A2(n5604), .ZN(n5716) );
  XNOR2_X1 U7189 ( .A(n5716), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8414) );
  INV_X1 U7190 ( .A(n8414), .ZN(n6228) );
  OR2_X1 U7191 ( .A1(n5662), .A2(n6228), .ZN(n5717) );
  XNOR2_X1 U7192 ( .A(n5679), .B(n9876), .ZN(n5727) );
  OAI21_X1 U7193 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5740), .ZN(n9828) );
  OR2_X1 U7194 ( .A1(n7824), .A2(n9828), .ZN(n5725) );
  NAND2_X1 U7195 ( .A1(n6021), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5724) );
  INV_X1 U7196 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5720) );
  OR2_X1 U7197 ( .A1(n7854), .A2(n5720), .ZN(n5723) );
  INV_X1 U7198 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6532) );
  OR2_X1 U7199 ( .A1(n5721), .A2(n6532), .ZN(n5722) );
  NAND4_X2 U7200 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n8392)
         );
  NAND2_X1 U7201 ( .A1(n8392), .A2(n5678), .ZN(n5726) );
  NAND2_X1 U7202 ( .A1(n5727), .A2(n5726), .ZN(n5732) );
  INV_X1 U7203 ( .A(n5726), .ZN(n5729) );
  INV_X1 U7204 ( .A(n5727), .ZN(n5728) );
  NAND2_X1 U7205 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  NAND2_X1 U7206 ( .A1(n5732), .A2(n5730), .ZN(n6629) );
  OR2_X1 U7207 ( .A1(n5767), .A2(n6224), .ZN(n5739) );
  OR2_X1 U7208 ( .A1(n7859), .A2(n6225), .ZN(n5738) );
  NAND2_X1 U7209 ( .A1(n5733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  MUX2_X1 U7210 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5734), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5736) );
  AND2_X1 U7211 ( .A1(n5736), .A2(n5735), .ZN(n8428) );
  INV_X1 U7212 ( .A(n8428), .ZN(n6223) );
  OR2_X1 U7213 ( .A1(n5662), .A2(n6223), .ZN(n5737) );
  XNOR2_X1 U7214 ( .A(n5679), .B(n6930), .ZN(n5747) );
  NAND2_X1 U7215 ( .A1(n7825), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7216 ( .A1(n6021), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5744) );
  INV_X1 U7217 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U7218 ( .A1(n5740), .A2(n8426), .ZN(n5741) );
  NAND2_X1 U7219 ( .A1(n5775), .A2(n5741), .ZN(n6640) );
  OR2_X1 U7220 ( .A1(n7824), .A2(n6640), .ZN(n5743) );
  INV_X1 U7221 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6892) );
  OR2_X1 U7222 ( .A1(n7858), .A2(n6892), .ZN(n5742) );
  NAND4_X1 U7223 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n8391)
         );
  NAND2_X1 U7224 ( .A1(n8391), .A2(n5678), .ZN(n5746) );
  XNOR2_X1 U7225 ( .A(n5747), .B(n5746), .ZN(n6635) );
  NOR2_X1 U7226 ( .A1(n6636), .A2(n6635), .ZN(n5750) );
  INV_X1 U7227 ( .A(n5746), .ZN(n5749) );
  INV_X1 U7228 ( .A(n5747), .ZN(n5748) );
  OR2_X1 U7229 ( .A1(n5767), .A2(n6226), .ZN(n5755) );
  OR2_X1 U7230 ( .A1(n7859), .A2(n6227), .ZN(n5754) );
  NAND2_X1 U7231 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5752) );
  INV_X1 U7232 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5751) );
  XNOR2_X1 U7233 ( .A(n5752), .B(n5751), .ZN(n6539) );
  OR2_X1 U7234 ( .A1(n5662), .A2(n6539), .ZN(n5753) );
  XNOR2_X1 U7235 ( .A(n5679), .B(n9894), .ZN(n5762) );
  NAND2_X1 U7236 ( .A1(n6021), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5760) );
  INV_X1 U7237 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U7238 ( .A(n5775), .B(n5774), .ZN(n7003) );
  OR2_X1 U7239 ( .A1(n7824), .A2(n7003), .ZN(n5759) );
  INV_X1 U7240 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5756) );
  OR2_X1 U7241 ( .A1(n7854), .A2(n5756), .ZN(n5758) );
  INV_X1 U7242 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6540) );
  OR2_X1 U7243 ( .A1(n7858), .A2(n6540), .ZN(n5757) );
  NAND4_X1 U7244 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n8213)
         );
  NAND2_X1 U7245 ( .A1(n8213), .A2(n5678), .ZN(n5761) );
  NAND2_X1 U7246 ( .A1(n5762), .A2(n5761), .ZN(n5766) );
  INV_X1 U7247 ( .A(n5761), .ZN(n5764) );
  INV_X1 U7248 ( .A(n5762), .ZN(n5763) );
  NAND2_X1 U7249 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  AND2_X1 U7250 ( .A1(n5766), .A2(n5765), .ZN(n6839) );
  OR2_X1 U7251 ( .A1(n5767), .A2(n6238), .ZN(n5772) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7253 ( .A1(n7859), .A2(n6239), .ZN(n5771) );
  OR2_X1 U7254 ( .A1(n5768), .A2(n5604), .ZN(n5769) );
  XNOR2_X1 U7255 ( .A(n5769), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8454) );
  INV_X1 U7256 ( .A(n8454), .ZN(n6237) );
  OR2_X1 U7257 ( .A1(n5662), .A2(n6237), .ZN(n5770) );
  XNOR2_X1 U7258 ( .A(n5679), .B(n7083), .ZN(n5784) );
  NAND2_X1 U7259 ( .A1(n6021), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5782) );
  INV_X1 U7260 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5773) );
  OAI21_X1 U7261 ( .B1(n5775), .B2(n5774), .A(n5773), .ZN(n5776) );
  NAND2_X1 U7262 ( .A1(n5776), .A2(n5793), .ZN(n6940) );
  OR2_X1 U7263 ( .A1(n7824), .A2(n6940), .ZN(n5781) );
  INV_X1 U7264 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5777) );
  OR2_X1 U7265 ( .A1(n7854), .A2(n5777), .ZN(n5780) );
  INV_X1 U7266 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5778) );
  OR2_X1 U7267 ( .A1(n7858), .A2(n5778), .ZN(n5779) );
  NAND4_X1 U7268 ( .A1(n5782), .A2(n5781), .A3(n5780), .A4(n5779), .ZN(n8212)
         );
  NAND2_X1 U7269 ( .A1(n8212), .A2(n5678), .ZN(n5783) );
  XNOR2_X1 U7270 ( .A(n5784), .B(n5783), .ZN(n6845) );
  INV_X1 U7271 ( .A(n5783), .ZN(n5786) );
  INV_X1 U7272 ( .A(n5784), .ZN(n5785) );
  NAND2_X1 U7273 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  XNOR2_X1 U7274 ( .A(n5789), .B(n5788), .ZN(n6542) );
  NAND2_X1 U7275 ( .A1(n6243), .A2(n5790), .ZN(n5792) );
  OR2_X1 U7276 ( .A1(n7859), .A2(n6244), .ZN(n5791) );
  XNOR2_X1 U7277 ( .A(n7279), .B(n5679), .ZN(n5801) );
  NAND2_X1 U7278 ( .A1(n6021), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5799) );
  INV_X1 U7279 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U7280 ( .A1(n5793), .A2(n8466), .ZN(n5794) );
  NAND2_X1 U7281 ( .A1(n5808), .A2(n5794), .ZN(n7096) );
  OR2_X1 U7282 ( .A1(n7824), .A2(n7096), .ZN(n5798) );
  INV_X1 U7283 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5795) );
  OR2_X1 U7284 ( .A1(n7854), .A2(n5795), .ZN(n5797) );
  INV_X1 U7285 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7097) );
  OR2_X1 U7286 ( .A1(n7858), .A2(n7097), .ZN(n5796) );
  NAND4_X1 U7287 ( .A1(n5799), .A2(n5798), .A3(n5797), .A4(n5796), .ZN(n8211)
         );
  NAND2_X1 U7288 ( .A1(n8211), .A2(n5678), .ZN(n5800) );
  XNOR2_X1 U7289 ( .A(n5801), .B(n5800), .ZN(n6972) );
  INV_X1 U7290 ( .A(n5800), .ZN(n5802) );
  AND2_X1 U7291 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  NAND2_X1 U7292 ( .A1(n6247), .A2(n5790), .ZN(n5806) );
  OR2_X1 U7293 ( .A1(n5804), .A2(n5604), .ZN(n5823) );
  XNOR2_X1 U7294 ( .A(n5823), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8479) );
  AOI22_X1 U7295 ( .A1(n5964), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6252), .B2(
        n8479), .ZN(n5805) );
  NAND2_X1 U7296 ( .A1(n5806), .A2(n5805), .ZN(n7394) );
  XNOR2_X1 U7297 ( .A(n7394), .B(n6068), .ZN(n5816) );
  NAND2_X1 U7298 ( .A1(n6021), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7299 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  NAND2_X1 U7300 ( .A1(n5827), .A2(n5809), .ZN(n7116) );
  OR2_X1 U7301 ( .A1(n7824), .A2(n7116), .ZN(n5814) );
  INV_X1 U7302 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7303 ( .A1(n7854), .A2(n5810), .ZN(n5813) );
  INV_X1 U7304 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7305 ( .A1(n7858), .A2(n5811), .ZN(n5812) );
  NAND4_X1 U7306 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n8210)
         );
  NAND2_X1 U7307 ( .A1(n8210), .A2(n5678), .ZN(n5817) );
  NAND2_X1 U7308 ( .A1(n5816), .A2(n5817), .ZN(n5821) );
  INV_X1 U7309 ( .A(n5816), .ZN(n5819) );
  INV_X1 U7310 ( .A(n5817), .ZN(n5818) );
  NAND2_X1 U7311 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  AND2_X1 U7312 ( .A1(n5821), .A2(n5820), .ZN(n7113) );
  NAND2_X1 U7313 ( .A1(n6290), .A2(n5790), .ZN(n5826) );
  NAND2_X1 U7314 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  NAND2_X1 U7315 ( .A1(n5824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  XNOR2_X1 U7316 ( .A(n5838), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7317 ( .A1(n5964), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6252), .B2(
        n6602), .ZN(n5825) );
  XNOR2_X1 U7318 ( .A(n9907), .B(n6068), .ZN(n5833) );
  NAND2_X1 U7319 ( .A1(n6021), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5832) );
  INV_X1 U7320 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U7321 ( .A1(n5827), .A2(n7107), .ZN(n5828) );
  NAND2_X1 U7322 ( .A1(n5859), .A2(n5828), .ZN(n7411) );
  OR2_X1 U7323 ( .A1(n7824), .A2(n7411), .ZN(n5831) );
  OR2_X1 U7324 ( .A1(n7854), .A2(n9935), .ZN(n5830) );
  INV_X1 U7325 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7412) );
  OR2_X1 U7326 ( .A1(n7858), .A2(n7412), .ZN(n5829) );
  NAND4_X1 U7327 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n8209)
         );
  NAND2_X1 U7328 ( .A1(n8209), .A2(n5678), .ZN(n5834) );
  XNOR2_X1 U7329 ( .A(n5833), .B(n5834), .ZN(n7105) );
  INV_X1 U7330 ( .A(n5833), .ZN(n5836) );
  INV_X1 U7331 ( .A(n5834), .ZN(n5835) );
  NAND2_X1 U7332 ( .A1(n6294), .A2(n5790), .ZN(n5842) );
  NAND2_X1 U7333 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  NAND2_X1 U7334 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7335 ( .A(n5840), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U7336 ( .A1(n5964), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6252), .B2(
        n6724), .ZN(n5841) );
  XNOR2_X1 U7337 ( .A(n8948), .B(n5679), .ZN(n5851) );
  NAND2_X1 U7338 ( .A1(n7825), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5848) );
  INV_X1 U7339 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5844) );
  OR2_X1 U7340 ( .A1(n5843), .A2(n5844), .ZN(n5847) );
  INV_X1 U7341 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5858) );
  XNOR2_X1 U7342 ( .A(n5859), .B(n5858), .ZN(n7482) );
  OR2_X1 U7343 ( .A1(n7824), .A2(n7482), .ZN(n5846) );
  INV_X1 U7344 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6598) );
  OR2_X1 U7345 ( .A1(n7858), .A2(n6598), .ZN(n5845) );
  NAND4_X1 U7346 ( .A1(n5848), .A2(n5847), .A3(n5846), .A4(n5845), .ZN(n8208)
         );
  NAND2_X1 U7347 ( .A1(n8208), .A2(n5678), .ZN(n5849) );
  XNOR2_X1 U7348 ( .A(n5851), .B(n5849), .ZN(n7273) );
  INV_X1 U7349 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U7350 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  NAND2_X1 U7351 ( .A1(n6365), .A2(n5790), .ZN(n5856) );
  NAND2_X1 U7352 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U7353 ( .A(n5854), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8494) );
  AOI22_X1 U7354 ( .A1(n5964), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6252), .B2(
        n8494), .ZN(n5855) );
  NAND2_X1 U7355 ( .A1(n5856), .A2(n5855), .ZN(n7498) );
  XNOR2_X1 U7356 ( .A(n7498), .B(n6068), .ZN(n5867) );
  NAND2_X1 U7357 ( .A1(n6022), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5866) );
  INV_X1 U7358 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5857) );
  OAI21_X1 U7359 ( .B1(n5859), .B2(n5858), .A(n5857), .ZN(n5860) );
  NAND2_X1 U7360 ( .A1(n5860), .A2(n5878), .ZN(n7493) );
  OR2_X1 U7361 ( .A1(n7824), .A2(n7493), .ZN(n5865) );
  INV_X1 U7362 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5861) );
  OR2_X1 U7363 ( .A1(n7854), .A2(n5861), .ZN(n5864) );
  INV_X1 U7364 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5862) );
  OR2_X1 U7365 ( .A1(n5843), .A2(n5862), .ZN(n5863) );
  NAND4_X1 U7366 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n8207)
         );
  NAND2_X1 U7367 ( .A1(n8207), .A2(n5678), .ZN(n5868) );
  NAND2_X1 U7368 ( .A1(n5867), .A2(n5868), .ZN(n5873) );
  INV_X1 U7369 ( .A(n5867), .ZN(n5870) );
  INV_X1 U7370 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U7371 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7372 ( .A1(n5873), .A2(n5871), .ZN(n7438) );
  NAND2_X1 U7373 ( .A1(n6479), .A2(n5790), .ZN(n5876) );
  NAND2_X1 U7374 ( .A1(n5874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7375 ( .A(n5889), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6782) );
  AOI22_X1 U7376 ( .A1(n5964), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6252), .B2(
        n6782), .ZN(n5875) );
  XNOR2_X1 U7377 ( .A(n8943), .B(n6068), .ZN(n5887) );
  NAND2_X1 U7378 ( .A1(n6021), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5885) );
  INV_X1 U7379 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7380 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  NAND2_X1 U7381 ( .A1(n5894), .A2(n5879), .ZN(n7470) );
  OR2_X1 U7382 ( .A1(n7824), .A2(n7470), .ZN(n5884) );
  INV_X1 U7383 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7384 ( .A1(n7854), .A2(n5880), .ZN(n5883) );
  INV_X1 U7385 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5881) );
  OR2_X1 U7386 ( .A1(n7858), .A2(n5881), .ZN(n5882) );
  NAND4_X1 U7387 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n8206)
         );
  NAND2_X1 U7388 ( .A1(n8206), .A2(n5678), .ZN(n5886) );
  XNOR2_X1 U7389 ( .A(n5887), .B(n5886), .ZN(n7443) );
  NAND2_X1 U7390 ( .A1(n6560), .A2(n5790), .ZN(n5892) );
  NAND2_X1 U7391 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NAND2_X1 U7392 ( .A1(n5890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7393 ( .A(n5909), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U7394 ( .A1(n5964), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6252), .B2(
        n6982), .ZN(n5891) );
  XNOR2_X1 U7395 ( .A(n8581), .B(n6068), .ZN(n5901) );
  NAND2_X1 U7396 ( .A1(n6021), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7397 ( .A1(n5894), .A2(n5893), .ZN(n5895) );
  NAND2_X1 U7398 ( .A1(n5915), .A2(n5895), .ZN(n7526) );
  OR2_X1 U7399 ( .A1(n7824), .A2(n7526), .ZN(n5899) );
  INV_X1 U7400 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5896) );
  OR2_X1 U7401 ( .A1(n7854), .A2(n5896), .ZN(n5898) );
  INV_X1 U7402 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7515) );
  OR2_X1 U7403 ( .A1(n7858), .A2(n7515), .ZN(n5897) );
  NAND4_X1 U7404 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n8580)
         );
  NAND2_X1 U7405 ( .A1(n8580), .A2(n5678), .ZN(n5902) );
  NAND2_X1 U7406 ( .A1(n5901), .A2(n5902), .ZN(n5907) );
  INV_X1 U7407 ( .A(n5901), .ZN(n5904) );
  INV_X1 U7408 ( .A(n5902), .ZN(n5903) );
  NAND2_X1 U7409 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  NAND2_X1 U7410 ( .A1(n5907), .A2(n5905), .ZN(n7522) );
  NAND2_X1 U7411 ( .A1(n6611), .A2(n5790), .ZN(n5913) );
  NAND2_X1 U7412 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  NAND2_X1 U7413 ( .A1(n5910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  XNOR2_X1 U7414 ( .A(n5911), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8514) );
  AOI22_X1 U7415 ( .A1(n5964), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6252), .B2(
        n8514), .ZN(n5912) );
  XNOR2_X1 U7416 ( .A(n8938), .B(n5679), .ZN(n5924) );
  NAND2_X1 U7417 ( .A1(n6021), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7418 ( .A1(n5915), .A2(n5914), .ZN(n5916) );
  NAND2_X1 U7419 ( .A1(n5917), .A2(n5916), .ZN(n8843) );
  OR2_X1 U7420 ( .A1(n7824), .A2(n8843), .ZN(n5921) );
  INV_X1 U7421 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8227) );
  OR2_X1 U7422 ( .A1(n7854), .A2(n8227), .ZN(n5920) );
  INV_X1 U7423 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7424 ( .A1(n7858), .A2(n5918), .ZN(n5919) );
  NAND4_X1 U7425 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n8820)
         );
  AND2_X1 U7426 ( .A1(n8820), .A2(n5678), .ZN(n8194) );
  XNOR2_X1 U7427 ( .A(n5926), .B(n5923), .ZN(n8128) );
  INV_X1 U7428 ( .A(n5924), .ZN(n8126) );
  INV_X1 U7429 ( .A(n8194), .ZN(n5925) );
  OAI21_X1 U7430 ( .B1(n5927), .B2(n5926), .A(n8130), .ZN(n8141) );
  NAND2_X1 U7431 ( .A1(n6627), .A2(n5790), .ZN(n5931) );
  NAND2_X1 U7432 ( .A1(n5928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  XNOR2_X1 U7433 ( .A(n5929), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8546) );
  AOI22_X1 U7434 ( .A1(n5964), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6252), .B2(
        n8546), .ZN(n5930) );
  XNOR2_X1 U7435 ( .A(n8930), .B(n6068), .ZN(n5941) );
  NAND2_X1 U7436 ( .A1(n6021), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5939) );
  INV_X1 U7437 ( .A(n5933), .ZN(n5932) );
  NAND2_X1 U7438 ( .A1(n5932), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5946) );
  INV_X1 U7439 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U7440 ( .A1(n5933), .A2(n8530), .ZN(n5934) );
  NAND2_X1 U7441 ( .A1(n5946), .A2(n5934), .ZN(n8808) );
  OR2_X1 U7442 ( .A1(n7824), .A2(n8808), .ZN(n5938) );
  INV_X1 U7443 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5935) );
  OR2_X1 U7444 ( .A1(n7854), .A2(n5935), .ZN(n5937) );
  INV_X1 U7445 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8809) );
  OR2_X1 U7446 ( .A1(n7858), .A2(n8809), .ZN(n5936) );
  NAND4_X1 U7447 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n8822)
         );
  NAND2_X1 U7448 ( .A1(n8822), .A2(n5678), .ZN(n5940) );
  XNOR2_X1 U7449 ( .A(n5941), .B(n5940), .ZN(n8140) );
  NAND2_X1 U7450 ( .A1(n6823), .A2(n5790), .ZN(n5944) );
  XNOR2_X1 U7451 ( .A(n5942), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8551) );
  AOI22_X1 U7452 ( .A1(n5964), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6252), .B2(
        n8551), .ZN(n5943) );
  XNOR2_X1 U7453 ( .A(n8923), .B(n5679), .ZN(n5954) );
  NAND2_X1 U7454 ( .A1(n5703), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5952) );
  INV_X1 U7455 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8557) );
  OR2_X1 U7456 ( .A1(n7854), .A2(n8557), .ZN(n5951) );
  NAND2_X1 U7457 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  NAND2_X1 U7458 ( .A1(n5957), .A2(n5947), .ZN(n8784) );
  OR2_X1 U7459 ( .A1(n7824), .A2(n8784), .ZN(n5950) );
  INV_X1 U7460 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7461 ( .A1(n7858), .A2(n5948), .ZN(n5949) );
  NAND4_X1 U7462 ( .A1(n5952), .A2(n5951), .A3(n5950), .A4(n5949), .ZN(n8765)
         );
  NAND2_X1 U7463 ( .A1(n8765), .A2(n5678), .ZN(n5953) );
  XNOR2_X1 U7464 ( .A(n5954), .B(n5953), .ZN(n8172) );
  INV_X1 U7465 ( .A(n5953), .ZN(n5955) );
  NAND2_X1 U7466 ( .A1(n6021), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5963) );
  INV_X1 U7467 ( .A(n5957), .ZN(n5956) );
  NAND2_X1 U7468 ( .A1(n5956), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5973) );
  INV_X1 U7469 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U7470 ( .A1(n5957), .A2(n8312), .ZN(n5958) );
  NAND2_X1 U7471 ( .A1(n5973), .A2(n5958), .ZN(n8776) );
  OR2_X1 U7472 ( .A1(n7824), .A2(n8776), .ZN(n5962) );
  INV_X1 U7473 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7474 ( .A1(n7854), .A2(n5959), .ZN(n5961) );
  INV_X1 U7475 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8777) );
  OR2_X1 U7476 ( .A1(n7858), .A2(n8777), .ZN(n5960) );
  NAND4_X1 U7477 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n8793)
         );
  AND2_X1 U7478 ( .A1(n8793), .A2(n5678), .ZN(n5968) );
  NAND2_X1 U7479 ( .A1(n6865), .A2(n5790), .ZN(n5966) );
  AOI22_X1 U7480 ( .A1(n5964), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5654), .B2(
        n6252), .ZN(n5965) );
  XNOR2_X1 U7481 ( .A(n8920), .B(n5679), .ZN(n5967) );
  NOR2_X1 U7482 ( .A1(n5967), .A2(n5968), .ZN(n5969) );
  AOI21_X1 U7483 ( .B1(n5968), .B2(n5967), .A(n5969), .ZN(n8102) );
  INV_X1 U7484 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U7485 ( .A1(n6991), .A2(n5790), .ZN(n5972) );
  OR2_X1 U7486 ( .A1(n7859), .A2(n7063), .ZN(n5971) );
  XNOR2_X1 U7487 ( .A(n8914), .B(n5679), .ZN(n5982) );
  NAND2_X1 U7488 ( .A1(n5973), .A2(n8156), .ZN(n5974) );
  NAND2_X1 U7489 ( .A1(n5987), .A2(n5974), .ZN(n8749) );
  OR2_X1 U7490 ( .A1(n7824), .A2(n8749), .ZN(n5980) );
  INV_X1 U7491 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8300) );
  OR2_X1 U7492 ( .A1(n5843), .A2(n8300), .ZN(n5979) );
  INV_X1 U7493 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7494 ( .A1(n7854), .A2(n5975), .ZN(n5978) );
  INV_X1 U7495 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5976) );
  OR2_X1 U7496 ( .A1(n7858), .A2(n5976), .ZN(n5977) );
  NAND4_X1 U7497 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n8766)
         );
  NAND2_X1 U7498 ( .A1(n8766), .A2(n5678), .ZN(n5981) );
  XNOR2_X1 U7499 ( .A(n5982), .B(n5981), .ZN(n8155) );
  INV_X1 U7500 ( .A(n5981), .ZN(n5983) );
  NAND2_X1 U7501 ( .A1(n7058), .A2(n5790), .ZN(n5985) );
  INV_X1 U7502 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7061) );
  OR2_X1 U7503 ( .A1(n7859), .A2(n7061), .ZN(n5984) );
  XNOR2_X1 U7504 ( .A(n8909), .B(n6068), .ZN(n5995) );
  INV_X1 U7505 ( .A(n5987), .ZN(n5986) );
  NAND2_X1 U7506 ( .A1(n5986), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5999) );
  INV_X1 U7507 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U7508 ( .A1(n5987), .A2(n8110), .ZN(n5988) );
  NAND2_X1 U7509 ( .A1(n5999), .A2(n5988), .ZN(n8733) );
  OR2_X1 U7510 ( .A1(n8733), .A2(n7824), .ZN(n5993) );
  NAND2_X1 U7511 ( .A1(n6021), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7512 ( .A1(n7825), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5991) );
  INV_X1 U7513 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7514 ( .A1(n7858), .A2(n5989), .ZN(n5990) );
  NAND4_X1 U7515 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n8756)
         );
  NAND2_X1 U7516 ( .A1(n8756), .A2(n5678), .ZN(n5994) );
  XNOR2_X1 U7517 ( .A(n5995), .B(n5994), .ZN(n8109) );
  NAND2_X1 U7518 ( .A1(n7120), .A2(n5790), .ZN(n5997) );
  OR2_X1 U7519 ( .A1(n7859), .A2(n7125), .ZN(n5996) );
  XNOR2_X1 U7520 ( .A(n8904), .B(n5679), .ZN(n6011) );
  INV_X1 U7521 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U7522 ( .A1(n5999), .A2(n8165), .ZN(n6000) );
  NAND2_X1 U7523 ( .A1(n6007), .A2(n6000), .ZN(n8716) );
  NAND2_X1 U7524 ( .A1(n7825), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7525 ( .A1(n6021), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6001) );
  AND2_X1 U7526 ( .A1(n6002), .A2(n6001), .ZN(n6004) );
  NAND2_X1 U7527 ( .A1(n6022), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6003) );
  OAI211_X1 U7528 ( .C1(n8716), .C2(n7824), .A(n6004), .B(n6003), .ZN(n8740)
         );
  NAND2_X1 U7529 ( .A1(n8740), .A2(n5678), .ZN(n8162) );
  NAND2_X1 U7530 ( .A1(n7256), .A2(n5790), .ZN(n6006) );
  OR2_X1 U7531 ( .A1(n7859), .A2(n7258), .ZN(n6005) );
  XNOR2_X1 U7532 ( .A(n8899), .B(n6068), .ZN(n8092) );
  INV_X1 U7533 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U7534 ( .A1(n6007), .A2(n8095), .ZN(n6008) );
  NAND2_X1 U7535 ( .A1(n6019), .A2(n6008), .ZN(n8700) );
  AOI22_X1 U7536 ( .A1(n6022), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5703), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7537 ( .A1(n7825), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U7538 ( .C1(n8700), .C2(n7824), .A(n6010), .B(n6009), .ZN(n8689)
         );
  NAND2_X1 U7539 ( .A1(n8689), .A2(n5678), .ZN(n6013) );
  NOR2_X1 U7540 ( .A1(n6012), .A2(n6011), .ZN(n8089) );
  INV_X1 U7541 ( .A(n8092), .ZN(n6014) );
  INV_X1 U7542 ( .A(n6013), .ZN(n8091) );
  NAND2_X1 U7543 ( .A1(n7350), .A2(n5790), .ZN(n6016) );
  OR2_X1 U7544 ( .A1(n7859), .A2(n7353), .ZN(n6015) );
  XNOR2_X1 U7545 ( .A(n8894), .B(n5679), .ZN(n6025) );
  INV_X1 U7546 ( .A(n6019), .ZN(n6018) );
  NAND2_X1 U7547 ( .A1(n6018), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6033) );
  INV_X1 U7548 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U7549 ( .A1(n6019), .A2(n8148), .ZN(n6020) );
  NAND2_X1 U7550 ( .A1(n6033), .A2(n6020), .ZN(n8682) );
  AOI22_X1 U7551 ( .A1(n6022), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n6021), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7552 ( .A1(n7825), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7553 ( .A1(n8708), .A2(n5678), .ZN(n8146) );
  OR2_X1 U7554 ( .A1(n6026), .A2(n6017), .ZN(n6027) );
  NAND2_X1 U7555 ( .A1(n7450), .A2(n5790), .ZN(n6030) );
  OR2_X1 U7556 ( .A1(n7859), .A2(n7452), .ZN(n6029) );
  XNOR2_X1 U7557 ( .A(n8891), .B(n5679), .ZN(n8117) );
  NAND2_X1 U7558 ( .A1(n8119), .A2(n8117), .ZN(n6040) );
  INV_X1 U7559 ( .A(n6033), .ZN(n6031) );
  NAND2_X1 U7560 ( .A1(n6031), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6047) );
  INV_X1 U7561 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7562 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7563 ( .A1(n6047), .A2(n6034), .ZN(n8664) );
  OR2_X1 U7564 ( .A1(n8664), .A2(n7824), .ZN(n6039) );
  INV_X1 U7565 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U7566 ( .A1(n7825), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7567 ( .A1(n6021), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7568 ( .C1(n8665), .C2(n7858), .A(n6036), .B(n6035), .ZN(n6037)
         );
  INV_X1 U7569 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7570 ( .A1(n6039), .A2(n6038), .ZN(n8690) );
  NAND2_X1 U7571 ( .A1(n8690), .A2(n5678), .ZN(n8116) );
  NAND2_X1 U7572 ( .A1(n6040), .A2(n8116), .ZN(n6044) );
  INV_X1 U7573 ( .A(n8119), .ZN(n6042) );
  INV_X1 U7574 ( .A(n8117), .ZN(n6041) );
  NAND2_X1 U7575 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  NAND2_X1 U7576 ( .A1(n7502), .A2(n5790), .ZN(n6046) );
  OR2_X1 U7577 ( .A1(n7859), .A2(n7503), .ZN(n6045) );
  XNOR2_X1 U7578 ( .A(n8886), .B(n6068), .ZN(n6056) );
  INV_X1 U7579 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U7580 ( .A1(n6047), .A2(n8186), .ZN(n6048) );
  NAND2_X1 U7581 ( .A1(n8656), .A2(n6049), .ZN(n6054) );
  INV_X1 U7582 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U7583 ( .A1(n7825), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7584 ( .A1(n6021), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6050) );
  OAI211_X1 U7585 ( .C1(n8658), .C2(n7858), .A(n6051), .B(n6050), .ZN(n6052)
         );
  INV_X1 U7586 ( .A(n6052), .ZN(n6053) );
  NAND2_X1 U7587 ( .A1(n6054), .A2(n6053), .ZN(n8640) );
  NAND2_X1 U7588 ( .A1(n8640), .A2(n5678), .ZN(n6055) );
  NOR2_X1 U7589 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  AOI21_X1 U7590 ( .B1(n6056), .B2(n6055), .A(n6057), .ZN(n8182) );
  INV_X1 U7591 ( .A(n6057), .ZN(n6082) );
  NAND2_X1 U7592 ( .A1(n8181), .A2(n6082), .ZN(n6122) );
  NAND2_X1 U7593 ( .A1(n6059), .A2(n6058), .ZN(n6061) );
  INV_X1 U7594 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8986) );
  MUX2_X1 U7595 ( .A(n8986), .B(n6150), .S(n4409), .Z(n6063) );
  INV_X1 U7596 ( .A(SI_27_), .ZN(n6062) );
  NAND2_X1 U7597 ( .A1(n6063), .A2(n6062), .ZN(n6170) );
  INV_X1 U7598 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7599 ( .A1(n6064), .A2(SI_27_), .ZN(n6065) );
  NAND2_X1 U7600 ( .A1(n8984), .A2(n5790), .ZN(n6067) );
  OR2_X1 U7601 ( .A1(n7859), .A2(n8986), .ZN(n6066) );
  XNOR2_X1 U7602 ( .A(n8880), .B(n6068), .ZN(n6080) );
  INV_X1 U7603 ( .A(n6071), .ZN(n6069) );
  NAND2_X1 U7604 ( .A1(n6069), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6132) );
  INV_X1 U7605 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7606 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  NAND2_X1 U7607 ( .A1(n6132), .A2(n6072), .ZN(n8633) );
  OR2_X1 U7608 ( .A1(n8633), .A2(n7824), .ZN(n6078) );
  INV_X1 U7609 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7610 ( .A1(n6021), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7611 ( .A1(n7825), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6073) );
  OAI211_X1 U7612 ( .C1(n6075), .C2(n7858), .A(n6074), .B(n6073), .ZN(n6076)
         );
  INV_X1 U7613 ( .A(n6076), .ZN(n6077) );
  NAND2_X1 U7614 ( .A1(n8619), .A2(n5678), .ZN(n6079) );
  NOR2_X1 U7615 ( .A1(n6080), .A2(n6079), .ZN(n7807) );
  AOI21_X1 U7616 ( .B1(n6080), .B2(n6079), .A(n7807), .ZN(n6121) );
  AND2_X1 U7617 ( .A1(n8182), .A2(n6121), .ZN(n6081) );
  INV_X1 U7618 ( .A(n6121), .ZN(n6083) );
  OR2_X1 U7619 ( .A1(n6083), .A2(n6082), .ZN(n7809) );
  AND2_X1 U7620 ( .A1(n7811), .A2(n7809), .ZN(n6120) );
  NAND2_X1 U7621 ( .A1(n6089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6085) );
  MUX2_X1 U7622 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6085), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6086) );
  INV_X1 U7623 ( .A(n7504), .ZN(n6098) );
  NAND2_X1 U7624 ( .A1(n6087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6088) );
  MUX2_X1 U7625 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6088), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6090) );
  NAND2_X1 U7626 ( .A1(n6090), .A2(n6089), .ZN(n7451) );
  NAND2_X1 U7627 ( .A1(n6092), .A2(n6091), .ZN(n6093) );
  XNOR2_X1 U7628 ( .A(n7355), .B(P2_B_REG_SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7629 ( .A1(n7451), .A2(n6096), .ZN(n6097) );
  INV_X1 U7630 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9845) );
  AND2_X1 U7631 ( .A1(n7451), .A2(n7504), .ZN(n9846) );
  AOI21_X1 U7632 ( .B1(n9838), .B2(n9845), .A(n9846), .ZN(n7064) );
  NOR4_X1 U7633 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6102) );
  NOR4_X1 U7634 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6101) );
  NOR4_X1 U7635 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6100) );
  NOR4_X1 U7636 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6099) );
  NAND4_X1 U7637 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n6108)
         );
  NOR2_X1 U7638 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .ZN(
        n6106) );
  NOR4_X1 U7639 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6105) );
  NOR4_X1 U7640 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6104) );
  NOR4_X1 U7641 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6103) );
  NAND4_X1 U7642 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n6107)
         );
  OAI21_X1 U7643 ( .B1(n6108), .B2(n6107), .A(n9838), .ZN(n7065) );
  AND2_X1 U7644 ( .A1(n7064), .A2(n7065), .ZN(n6699) );
  INV_X1 U7645 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U7646 ( .A1(n9838), .A2(n9842), .ZN(n6110) );
  AND2_X1 U7647 ( .A1(n7355), .A2(n7504), .ZN(n9843) );
  INV_X1 U7648 ( .A(n9843), .ZN(n6109) );
  NAND2_X1 U7649 ( .A1(n6699), .A2(n7076), .ZN(n6125) );
  INV_X1 U7650 ( .A(n7355), .ZN(n6112) );
  NOR2_X1 U7651 ( .A1(n7504), .A2(n7451), .ZN(n6111) );
  NAND2_X1 U7652 ( .A1(n6116), .A2(n6115), .ZN(n6127) );
  INV_X1 U7653 ( .A(n9847), .ZN(n6117) );
  NAND2_X1 U7654 ( .A1(n8063), .A2(n7909), .ZN(n6126) );
  AND2_X1 U7655 ( .A1(n9915), .A2(n6126), .ZN(n6119) );
  OAI211_X1 U7656 ( .C1(n6122), .C2(n6121), .A(n6120), .B(n8180), .ZN(n6149)
         );
  INV_X1 U7657 ( .A(n6118), .ZN(n7892) );
  AND2_X1 U7658 ( .A1(n7892), .A2(n7865), .ZN(n6708) );
  NAND2_X1 U7659 ( .A1(n6140), .A2(n6708), .ZN(n6124) );
  NOR2_X1 U7660 ( .A1(n8807), .A2(n8063), .ZN(n6123) );
  NAND2_X1 U7661 ( .A1(n6125), .A2(n7067), .ZN(n6500) );
  INV_X1 U7662 ( .A(n6127), .ZN(n6251) );
  NOR2_X1 U7663 ( .A1(n6507), .A2(n6251), .ZN(n6128) );
  AND2_X1 U7664 ( .A1(n7066), .A2(n6128), .ZN(n6129) );
  NOR2_X1 U7665 ( .A1(n8633), .A2(n8200), .ZN(n6145) );
  INV_X1 U7666 ( .A(n6132), .ZN(n6130) );
  NAND2_X1 U7667 ( .A1(n6130), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8607) );
  INV_X1 U7668 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7669 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  NAND2_X1 U7670 ( .A1(n8607), .A2(n6133), .ZN(n8623) );
  OR2_X1 U7671 ( .A1(n8623), .A2(n7824), .ZN(n6138) );
  INV_X1 U7672 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U7673 ( .A1(n7825), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7674 ( .A1(n6021), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6134) );
  OAI211_X1 U7675 ( .C1(n8622), .C2(n7858), .A(n6135), .B(n6134), .ZN(n6136)
         );
  INV_X1 U7676 ( .A(n6136), .ZN(n6137) );
  NAND2_X1 U7677 ( .A1(n6138), .A2(n6137), .ZN(n8641) );
  INV_X1 U7678 ( .A(n6139), .ZN(n8061) );
  NAND2_X1 U7679 ( .A1(n6140), .A2(n8061), .ZN(n6590) );
  INV_X1 U7680 ( .A(n6142), .ZN(n6143) );
  NOR2_X1 U7681 ( .A1(n6590), .A2(n8806), .ZN(n8174) );
  NOR2_X1 U7682 ( .A1(n6590), .A2(n8804), .ZN(n8175) );
  OAI22_X1 U7683 ( .A1(n8595), .A2(n8166), .B1(n8594), .B2(n8167), .ZN(n6144)
         );
  AOI211_X1 U7684 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n6145), 
        .B(n6144), .ZN(n6146) );
  INV_X1 U7685 ( .A(n6147), .ZN(n6148) );
  NAND2_X1 U7686 ( .A1(n6149), .A2(n6148), .ZN(P2_U3216) );
  NAND2_X1 U7687 ( .A1(n8984), .A2(n5245), .ZN(n6152) );
  OR2_X1 U7688 ( .A1(n7597), .A2(n6150), .ZN(n6151) );
  NAND2_X1 U7689 ( .A1(n9493), .A2(n5222), .ZN(n6154) );
  OR2_X1 U7690 ( .A1(n7530), .A2(n5505), .ZN(n6153) );
  NAND2_X1 U7691 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  XNOR2_X1 U7692 ( .A(n6155), .B(n6188), .ZN(n6158) );
  INV_X1 U7693 ( .A(n6158), .ZN(n6160) );
  NOR2_X1 U7694 ( .A1(n7530), .A2(n5319), .ZN(n6156) );
  AOI21_X1 U7695 ( .B1(n9493), .B2(n4333), .A(n6156), .ZN(n6157) );
  INV_X1 U7696 ( .A(n6157), .ZN(n6159) );
  AOI21_X1 U7697 ( .B1(n6160), .B2(n6159), .A(n6193), .ZN(n8989) );
  INV_X1 U7698 ( .A(n8989), .ZN(n6166) );
  INV_X1 U7699 ( .A(n6161), .ZN(n6164) );
  INV_X1 U7700 ( .A(n6162), .ZN(n6163) );
  NAND2_X1 U7701 ( .A1(n6164), .A2(n6163), .ZN(n8990) );
  INV_X1 U7702 ( .A(n8990), .ZN(n6165) );
  NOR2_X1 U7703 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  NAND2_X1 U7704 ( .A1(n6169), .A2(n6168), .ZN(n6171) );
  INV_X1 U7705 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8088) );
  INV_X1 U7706 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U7707 ( .A(n8088), .B(n9592), .S(n4409), .Z(n6172) );
  INV_X1 U7708 ( .A(SI_28_), .ZN(n8238) );
  NAND2_X1 U7709 ( .A1(n6172), .A2(n8238), .ZN(n7568) );
  INV_X1 U7710 ( .A(n6172), .ZN(n6173) );
  NAND2_X1 U7711 ( .A1(n6173), .A2(SI_28_), .ZN(n6174) );
  NAND2_X1 U7712 ( .A1(n9589), .A2(n5245), .ZN(n6176) );
  OR2_X1 U7713 ( .A1(n7597), .A2(n9592), .ZN(n6175) );
  NAND2_X1 U7714 ( .A1(n9488), .A2(n5222), .ZN(n6187) );
  NAND2_X1 U7715 ( .A1(n7587), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7716 ( .A1(n7601), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6184) );
  INV_X1 U7717 ( .A(n6179), .ZN(n6177) );
  NAND2_X1 U7718 ( .A1(n6177), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6195) );
  INV_X1 U7719 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7720 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  NAND2_X1 U7721 ( .A1(n6181), .A2(n9250), .ZN(n6183) );
  NAND2_X1 U7722 ( .A1(n7600), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6182) );
  OR2_X1 U7723 ( .A1(n9235), .A2(n5505), .ZN(n6186) );
  NAND2_X1 U7724 ( .A1(n6187), .A2(n6186), .ZN(n6189) );
  XNOR2_X1 U7725 ( .A(n6189), .B(n6188), .ZN(n6192) );
  NAND2_X1 U7726 ( .A1(n9488), .A2(n4333), .ZN(n6190) );
  OAI21_X1 U7727 ( .B1(n9235), .B2(n5319), .A(n6190), .ZN(n6191) );
  XNOR2_X1 U7728 ( .A(n6192), .B(n6191), .ZN(n6194) );
  AND2_X1 U7729 ( .A1(n6194), .A2(n9678), .ZN(n6206) );
  NAND3_X1 U7730 ( .A1(n6194), .A2(n9678), .A3(n6193), .ZN(n6204) );
  NAND2_X1 U7731 ( .A1(n7600), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6199) );
  INV_X1 U7732 ( .A(n6195), .ZN(n9238) );
  NAND2_X1 U7733 ( .A1(n6181), .A2(n9238), .ZN(n6198) );
  NAND2_X1 U7734 ( .A1(n7587), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7735 ( .A1(n7601), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6196) );
  NAND4_X1 U7736 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n9258)
         );
  INV_X1 U7737 ( .A(n9258), .ZN(n7741) );
  AOI22_X1 U7738 ( .A1(n9286), .A2(n9111), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6200) );
  OAI21_X1 U7739 ( .B1(n9096), .B2(n7741), .A(n6200), .ZN(n6202) );
  INV_X1 U7740 ( .A(n9488), .ZN(n9252) );
  NOR2_X1 U7741 ( .A1(n9252), .A2(n9056), .ZN(n6201) );
  AOI211_X1 U7742 ( .C1(n9250), .C2(n9100), .A(n6202), .B(n6201), .ZN(n6203)
         );
  NAND2_X1 U7743 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  AOI21_X1 U7744 ( .B1(n8992), .B2(n6206), .A(n6205), .ZN(n6207) );
  NAND2_X1 U7745 ( .A1(n7753), .A2(n6286), .ZN(n6209) );
  NAND2_X1 U7746 ( .A1(n6209), .A2(n6284), .ZN(n6280) );
  NAND2_X1 U7747 ( .A1(n6280), .A2(n6210), .ZN(n6211) );
  NAND2_X1 U7748 ( .A1(n6211), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7749 ( .A(n6212), .ZN(n6213) );
  NAND2_X1 U7750 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), .ZN(
        n6427) );
  OAI21_X1 U7751 ( .B1(n6213), .B2(P1_STATE_REG_SCAN_IN), .A(n6427), .ZN(
        P1_U3353) );
  NAND2_X2 U7752 ( .A1(n6214), .A2(P1_U3084), .ZN(n9593) );
  OAI222_X1 U7753 ( .A1(n9593), .A2(n6215), .B1(n9597), .B2(n6234), .C1(
        P1_U3084), .C2(n6415), .ZN(P1_U3350) );
  INV_X2 U7754 ( .A(n8979), .ZN(n6866) );
  NAND2_X2 U7755 ( .A1(n4409), .A2(P2_U3152), .ZN(n8987) );
  OAI222_X1 U7756 ( .A1(P2_U3152), .A2(n9599), .B1(n6866), .B2(n6219), .C1(
        n6216), .C2(n8987), .ZN(P2_U3357) );
  OAI222_X1 U7757 ( .A1(n9593), .A2(n6218), .B1(n9597), .B2(n6224), .C1(
        P1_U3084), .C2(n6217), .ZN(P1_U3348) );
  OAI222_X1 U7758 ( .A1(n9593), .A2(n6220), .B1(n9597), .B2(n6219), .C1(
        P1_U3084), .C2(n6388), .ZN(P1_U3352) );
  OAI222_X1 U7759 ( .A1(n9593), .A2(n6221), .B1(n9597), .B2(n6229), .C1(
        P1_U3084), .C2(n6431), .ZN(P1_U3349) );
  OAI222_X1 U7760 ( .A1(n9593), .A2(n6222), .B1(n9597), .B2(n6226), .C1(
        P1_U3084), .C2(n6374), .ZN(P1_U3347) );
  OAI222_X1 U7761 ( .A1(n9593), .A2(n4401), .B1(n9597), .B2(n6232), .C1(
        P1_U3084), .C2(n6450), .ZN(P1_U3351) );
  OAI222_X1 U7762 ( .A1(n8987), .A2(n6225), .B1(n6866), .B2(n6224), .C1(
        P2_U3152), .C2(n6223), .ZN(P2_U3353) );
  OAI222_X1 U7763 ( .A1(n8987), .A2(n6227), .B1(n6866), .B2(n6226), .C1(
        P2_U3152), .C2(n6539), .ZN(P2_U3352) );
  OAI222_X1 U7764 ( .A1(n8987), .A2(n6230), .B1(n6866), .B2(n6229), .C1(
        P2_U3152), .C2(n6228), .ZN(P2_U3354) );
  OAI222_X1 U7765 ( .A1(P2_U3152), .A2(n6535), .B1(n6866), .B2(n6232), .C1(
        n6231), .C2(n8987), .ZN(P2_U3356) );
  OAI222_X1 U7766 ( .A1(P2_U3152), .A2(n6235), .B1(n6866), .B2(n6234), .C1(
        n6233), .C2(n8987), .ZN(P2_U3355) );
  OAI222_X1 U7767 ( .A1(n9593), .A2(n6236), .B1(n9597), .B2(n6238), .C1(
        P1_U3084), .C2(n6364), .ZN(P1_U3346) );
  OAI222_X1 U7768 ( .A1(n8987), .A2(n6239), .B1(n6866), .B2(n6238), .C1(
        P2_U3152), .C2(n6237), .ZN(P2_U3351) );
  INV_X1 U7769 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6666) );
  NOR2_X1 U7770 ( .A1(n6668), .A2(n6241), .ZN(n6242) );
  AOI21_X1 U7771 ( .B1(n9711), .B2(n6666), .A(n6242), .ZN(P1_U3441) );
  INV_X1 U7772 ( .A(n6243), .ZN(n6245) );
  OAI222_X1 U7773 ( .A1(n8987), .A2(n6244), .B1(n6866), .B2(n6245), .C1(
        P2_U3152), .C2(n6542), .ZN(P2_U3350) );
  INV_X1 U7774 ( .A(n6346), .ZN(n6325) );
  OAI222_X1 U7775 ( .A1(n9593), .A2(n6246), .B1(n9597), .B2(n6245), .C1(
        P1_U3084), .C2(n6325), .ZN(P1_U3345) );
  INV_X1 U7776 ( .A(n6247), .ZN(n6250) );
  AOI22_X1 U7777 ( .A1(n8479), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n6366), .ZN(n6248) );
  OAI21_X1 U7778 ( .B1(n6250), .B2(n6866), .A(n6248), .ZN(P2_U3349) );
  INV_X1 U7779 ( .A(n9593), .ZN(n9595) );
  AOI22_X1 U7780 ( .A1(n9138), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9595), .ZN(n6249) );
  OAI21_X1 U7781 ( .B1(n6250), .B2(n9597), .A(n6249), .ZN(P1_U3344) );
  INV_X1 U7782 ( .A(n9839), .ZN(n8060) );
  NAND2_X1 U7783 ( .A1(n8060), .A2(n6509), .ZN(n6255) );
  NAND2_X1 U7784 ( .A1(n6251), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8065) );
  NAND2_X1 U7785 ( .A1(n9839), .A2(n8065), .ZN(n6253) );
  NAND2_X1 U7786 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  AND2_X1 U7787 ( .A1(n6255), .A2(n6254), .ZN(n9602) );
  INV_X1 U7788 ( .A(n9602), .ZN(n9809) );
  NOR2_X1 U7789 ( .A1(n9809), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7790 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6256) );
  MUX2_X1 U7791 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6256), .S(n6319), .Z(n6257)
         );
  INV_X1 U7792 ( .A(n6257), .ZN(n6267) );
  INV_X1 U7793 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6265) );
  INV_X1 U7794 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6761) );
  MUX2_X1 U7795 ( .A(n6761), .B(P1_REG2_REG_2__SCAN_IN), .S(n6450), .Z(n6260)
         );
  INV_X1 U7796 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6752) );
  MUX2_X1 U7797 ( .A(n6752), .B(P1_REG2_REG_1__SCAN_IN), .S(n6388), .Z(n6391)
         );
  AND2_X1 U7798 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6258) );
  OR2_X1 U7799 ( .A1(n6388), .A2(n6752), .ZN(n6451) );
  NAND2_X1 U7800 ( .A1(n6452), .A2(n6451), .ZN(n6259) );
  NAND2_X1 U7801 ( .A1(n6260), .A2(n6259), .ZN(n6455) );
  OR2_X1 U7802 ( .A1(n6450), .A2(n6761), .ZN(n6261) );
  NAND2_X1 U7803 ( .A1(n6455), .A2(n6261), .ZN(n6414) );
  INV_X1 U7804 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6262) );
  MUX2_X1 U7805 ( .A(n6262), .B(P1_REG2_REG_3__SCAN_IN), .S(n6415), .Z(n6263)
         );
  NAND2_X1 U7806 ( .A1(n6414), .A2(n6263), .ZN(n6416) );
  INV_X1 U7807 ( .A(n6415), .ZN(n6274) );
  NAND2_X1 U7808 ( .A1(n6274), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7809 ( .A1(n6416), .A2(n6264), .ZN(n6439) );
  MUX2_X1 U7810 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6265), .S(n6431), .Z(n6438)
         );
  AOI21_X1 U7811 ( .B1(n6431), .B2(n6265), .A(n6437), .ZN(n6266) );
  AOI21_X1 U7812 ( .B1(n6267), .B2(n6266), .A(n6306), .ZN(n6289) );
  NOR2_X1 U7813 ( .A1(n6268), .A2(P1_U3084), .ZN(n9594) );
  NAND2_X1 U7814 ( .A1(n6280), .A2(n9594), .ZN(n9177) );
  INV_X1 U7815 ( .A(n9177), .ZN(n6269) );
  AND2_X1 U7816 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6827) );
  INV_X1 U7817 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9787) );
  MUX2_X1 U7818 ( .A(n9787), .B(P1_REG1_REG_2__SCAN_IN), .S(n6450), .Z(n6448)
         );
  INV_X1 U7819 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9785) );
  MUX2_X1 U7820 ( .A(n9785), .B(P1_REG1_REG_1__SCAN_IN), .S(n6388), .Z(n6383)
         );
  NAND2_X1 U7821 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6387) );
  INV_X1 U7822 ( .A(n6387), .ZN(n6270) );
  NAND2_X1 U7823 ( .A1(n6383), .A2(n6270), .ZN(n6384) );
  INV_X1 U7824 ( .A(n6388), .ZN(n6271) );
  NAND2_X1 U7825 ( .A1(n6271), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7826 ( .A1(n6384), .A2(n6272), .ZN(n6447) );
  NAND2_X1 U7827 ( .A1(n6448), .A2(n6447), .ZN(n6446) );
  INV_X1 U7828 ( .A(n6450), .ZN(n6460) );
  NAND2_X1 U7829 ( .A1(n6460), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7830 ( .A1(n6446), .A2(n6273), .ZN(n6411) );
  XNOR2_X1 U7831 ( .A(n6415), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U7832 ( .A1(n6411), .A2(n6412), .ZN(n6410) );
  NAND2_X1 U7833 ( .A1(n6274), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7834 ( .A1(n6410), .A2(n6275), .ZN(n6433) );
  XNOR2_X1 U7835 ( .A(n6431), .B(n5133), .ZN(n6434) );
  NOR2_X1 U7836 ( .A1(n6433), .A2(n6434), .ZN(n6432) );
  AND2_X1 U7837 ( .A1(n6431), .A2(n5133), .ZN(n6276) );
  OR2_X1 U7838 ( .A1(n6432), .A2(n6276), .ZN(n6282) );
  OR2_X1 U7839 ( .A1(n6319), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7840 ( .A1(n6319), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7841 ( .A1(n6278), .A2(n6277), .ZN(n6281) );
  NOR2_X1 U7842 ( .A1(n6282), .A2(n6281), .ZN(n6318) );
  OR2_X1 U7843 ( .A1(n9686), .A2(P1_U3084), .ZN(n9590) );
  INV_X1 U7844 ( .A(n6268), .ZN(n9186) );
  NOR2_X1 U7845 ( .A1(n9590), .A2(n9186), .ZN(n6279) );
  NAND2_X1 U7846 ( .A1(n6280), .A2(n6279), .ZN(n9173) );
  AOI211_X1 U7847 ( .C1(n6282), .C2(n6281), .A(n6318), .B(n9173), .ZN(n6283)
         );
  AOI211_X1 U7848 ( .C1(n9698), .C2(n6319), .A(n6827), .B(n6283), .ZN(n6288)
         );
  INV_X1 U7849 ( .A(n6284), .ZN(n6285) );
  NOR2_X1 U7850 ( .A1(n6286), .A2(n6285), .ZN(n6429) );
  INV_X1 U7851 ( .A(n9184), .ZN(n9703) );
  NAND2_X1 U7852 ( .A1(n9703), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6287) );
  OAI211_X1 U7853 ( .C1(n6289), .C2(n9695), .A(n6288), .B(n6287), .ZN(P1_U3246) );
  INV_X1 U7854 ( .A(n6290), .ZN(n6292) );
  INV_X1 U7855 ( .A(n6602), .ZN(n6550) );
  OAI222_X1 U7856 ( .A1(n8987), .A2(n6291), .B1(n6866), .B2(n6292), .C1(n6550), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7857 ( .A(n6347), .ZN(n6402) );
  OAI222_X1 U7858 ( .A1(n9593), .A2(n6293), .B1(n9597), .B2(n6292), .C1(n6402), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7859 ( .A(n6294), .ZN(n6297) );
  INV_X1 U7860 ( .A(n6470), .ZN(n6342) );
  OAI222_X1 U7861 ( .A1(n9593), .A2(n6295), .B1(n9597), .B2(n6297), .C1(n6342), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7862 ( .A(n6724), .ZN(n6717) );
  OAI222_X1 U7863 ( .A1(P2_U3152), .A2(n6717), .B1(n6866), .B2(n6297), .C1(
        n6296), .C2(n8987), .ZN(P2_U3347) );
  INV_X1 U7864 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7865 ( .A1(n6021), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6302) );
  INV_X1 U7866 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6298) );
  OR2_X1 U7867 ( .A1(n7854), .A2(n6298), .ZN(n6301) );
  INV_X1 U7868 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6299) );
  OR2_X1 U7869 ( .A1(n7858), .A2(n6299), .ZN(n6300) );
  AND3_X1 U7870 ( .A1(n6302), .A2(n6301), .A3(n6300), .ZN(n7862) );
  NAND2_X1 U7871 ( .A1(n8572), .A2(P2_U3966), .ZN(n6303) );
  OAI21_X1 U7872 ( .B1(n6304), .B2(P2_U3966), .A(n6303), .ZN(P2_U3583) );
  NOR2_X1 U7873 ( .A1(n6321), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6311) );
  INV_X1 U7874 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6305) );
  MUX2_X1 U7875 ( .A(n6305), .B(P1_REG2_REG_7__SCAN_IN), .S(n6321), .Z(n6354)
         );
  NAND2_X1 U7876 ( .A1(n6320), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6310) );
  NOR2_X1 U7877 ( .A1(n6319), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6307) );
  NOR2_X1 U7878 ( .A1(n6307), .A2(n6306), .ZN(n6379) );
  INV_X1 U7879 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6308) );
  MUX2_X1 U7880 ( .A(n6308), .B(P1_REG2_REG_6__SCAN_IN), .S(n6320), .Z(n6309)
         );
  INV_X1 U7881 ( .A(n6309), .ZN(n6378) );
  NAND2_X1 U7882 ( .A1(n6379), .A2(n6378), .ZN(n6377) );
  NAND2_X1 U7883 ( .A1(n6310), .A2(n6377), .ZN(n6355) );
  NOR2_X1 U7884 ( .A1(n6311), .A2(n6353), .ZN(n6314) );
  INV_X1 U7885 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6312) );
  AOI22_X1 U7886 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6325), .B1(n6346), .B2(
        n6312), .ZN(n6313) );
  AOI21_X1 U7887 ( .B1(n6314), .B2(n6313), .A(n6334), .ZN(n6329) );
  INV_X1 U7888 ( .A(n9173), .ZN(n9704) );
  NOR2_X1 U7889 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6346), .ZN(n6315) );
  AOI21_X1 U7890 ( .B1(n6346), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6315), .ZN(
        n6323) );
  NOR2_X1 U7891 ( .A1(n6321), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6316) );
  AOI21_X1 U7892 ( .B1(n6321), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6316), .ZN(
        n6360) );
  NOR2_X1 U7893 ( .A1(n6320), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6317) );
  AOI21_X1 U7894 ( .B1(n6320), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6317), .ZN(
        n6371) );
  AOI21_X1 U7895 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6319), .A(n6318), .ZN(
        n6372) );
  NAND2_X1 U7896 ( .A1(n6371), .A2(n6372), .ZN(n6370) );
  OAI21_X1 U7897 ( .B1(n6320), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6370), .ZN(
        n6359) );
  NAND2_X1 U7898 ( .A1(n6360), .A2(n6359), .ZN(n6358) );
  OAI21_X1 U7899 ( .B1(n6321), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6358), .ZN(
        n6322) );
  NAND2_X1 U7900 ( .A1(n6323), .A2(n6322), .ZN(n6345) );
  OAI21_X1 U7901 ( .B1(n6323), .B2(n6322), .A(n6345), .ZN(n6327) );
  NAND2_X1 U7902 ( .A1(n9703), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7903 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9668) );
  OAI211_X1 U7904 ( .C1(n7161), .C2(n6325), .A(n6324), .B(n9668), .ZN(n6326)
         );
  AOI21_X1 U7905 ( .B1(n9704), .B2(n6327), .A(n6326), .ZN(n6328) );
  OAI21_X1 U7906 ( .B1(n6329), .B2(n9695), .A(n6328), .ZN(P1_U3249) );
  NAND2_X1 U7907 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6347), .ZN(n6337) );
  INV_X1 U7908 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6330) );
  MUX2_X1 U7909 ( .A(n6330), .B(P1_REG2_REG_10__SCAN_IN), .S(n6347), .Z(n6331)
         );
  INV_X1 U7910 ( .A(n6331), .ZN(n6396) );
  NAND2_X1 U7911 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9138), .ZN(n6336) );
  INV_X1 U7912 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6332) );
  MUX2_X1 U7913 ( .A(n6332), .B(P1_REG2_REG_9__SCAN_IN), .S(n9138), .Z(n6333)
         );
  INV_X1 U7914 ( .A(n6333), .ZN(n9135) );
  NOR2_X1 U7915 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6346), .ZN(n6335) );
  NOR2_X1 U7916 ( .A1(n6335), .A2(n6334), .ZN(n9136) );
  NAND2_X1 U7917 ( .A1(n9135), .A2(n9136), .ZN(n9134) );
  NAND2_X1 U7918 ( .A1(n6336), .A2(n9134), .ZN(n6397) );
  NAND2_X1 U7919 ( .A1(n6396), .A2(n6397), .ZN(n6395) );
  NAND2_X1 U7920 ( .A1(n6337), .A2(n6395), .ZN(n6472) );
  INV_X1 U7921 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7922 ( .A1(n6338), .A2(n6342), .ZN(n6471) );
  OAI21_X1 U7923 ( .B1(n6342), .B2(n6338), .A(n6471), .ZN(n6339) );
  OAI22_X1 U7924 ( .A1(n7161), .A2(n6342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6340), .ZN(n6341) );
  AOI21_X1 U7925 ( .B1(n9703), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6341), .ZN(
        n6352) );
  INV_X1 U7926 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9658) );
  AOI22_X1 U7927 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6470), .B1(n6342), .B2(
        n9658), .ZN(n6349) );
  INV_X1 U7928 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6343) );
  MUX2_X1 U7929 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6343), .S(n6347), .Z(n6400)
         );
  NOR2_X1 U7930 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9138), .ZN(n6344) );
  AOI21_X1 U7931 ( .B1(n9138), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6344), .ZN(
        n9140) );
  OAI21_X1 U7932 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6346), .A(n6345), .ZN(
        n9141) );
  NAND2_X1 U7933 ( .A1(n9140), .A2(n9141), .ZN(n9139) );
  OAI21_X1 U7934 ( .B1(n9138), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9139), .ZN(
        n6399) );
  NAND2_X1 U7935 ( .A1(n6400), .A2(n6399), .ZN(n6398) );
  OAI21_X1 U7936 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6347), .A(n6398), .ZN(
        n6348) );
  NAND2_X1 U7937 ( .A1(n6349), .A2(n6348), .ZN(n6463) );
  OAI21_X1 U7938 ( .B1(n6349), .B2(n6348), .A(n6463), .ZN(n6350) );
  NAND2_X1 U7939 ( .A1(n6350), .A2(n9704), .ZN(n6351) );
  OAI211_X1 U7940 ( .C1(n4883), .C2(n9695), .A(n6352), .B(n6351), .ZN(P1_U3252) );
  AOI21_X1 U7941 ( .B1(n6355), .B2(n6354), .A(n6353), .ZN(n6356) );
  NOR2_X1 U7942 ( .A1(n9695), .A2(n6356), .ZN(n6357) );
  AOI21_X1 U7943 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(n9703), .A(n6357), .ZN(
        n6363) );
  OAI21_X1 U7944 ( .B1(n6360), .B2(n6359), .A(n6358), .ZN(n6361) );
  AND2_X1 U7945 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6965) );
  AOI21_X1 U7946 ( .B1(n9704), .B2(n6361), .A(n6965), .ZN(n6362) );
  OAI211_X1 U7947 ( .C1(n6364), .C2(n7161), .A(n6363), .B(n6362), .ZN(P1_U3248) );
  INV_X1 U7948 ( .A(n6365), .ZN(n6369) );
  AOI22_X1 U7949 ( .A1(n8494), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n6366), .ZN(n6367) );
  OAI21_X1 U7950 ( .B1(n6369), .B2(n6866), .A(n6367), .ZN(P2_U3346) );
  AOI22_X1 U7951 ( .A1(n6580), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9595), .ZN(n6368) );
  OAI21_X1 U7952 ( .B1(n6369), .B2(n9597), .A(n6368), .ZN(P1_U3341) );
  INV_X1 U7953 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6382) );
  OAI21_X1 U7954 ( .B1(n6372), .B2(n6371), .A(n6370), .ZN(n6376) );
  INV_X1 U7955 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6373) );
  NOR2_X1 U7956 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6373), .ZN(n9098) );
  NOR2_X1 U7957 ( .A1(n7161), .A2(n6374), .ZN(n6375) );
  AOI211_X1 U7958 ( .C1(n9704), .C2(n6376), .A(n9098), .B(n6375), .ZN(n6381)
         );
  OAI211_X1 U7959 ( .C1(n6379), .C2(n6378), .A(n9157), .B(n6377), .ZN(n6380)
         );
  OAI211_X1 U7960 ( .C1(n9184), .C2(n6382), .A(n6381), .B(n6380), .ZN(P1_U3247) );
  INV_X1 U7961 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6394) );
  INV_X1 U7962 ( .A(n6383), .ZN(n6386) );
  INV_X1 U7963 ( .A(n6384), .ZN(n6385) );
  AOI211_X1 U7964 ( .C1(n6387), .C2(n6386), .A(n6385), .B(n9173), .ZN(n6390)
         );
  NOR2_X1 U7965 ( .A1(n7161), .A2(n6388), .ZN(n6389) );
  AOI211_X1 U7966 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n6390), .B(
        n6389), .ZN(n6393) );
  NAND2_X1 U7967 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6426) );
  OAI211_X1 U7968 ( .C1(n6258), .C2(n6391), .A(n9157), .B(n6452), .ZN(n6392)
         );
  OAI211_X1 U7969 ( .C1(n9184), .C2(n6394), .A(n6393), .B(n6392), .ZN(P1_U3242) );
  INV_X1 U7970 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6407) );
  OAI211_X1 U7971 ( .C1(n6397), .C2(n6396), .A(n9157), .B(n6395), .ZN(n6406)
         );
  OAI21_X1 U7972 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6404) );
  NOR2_X1 U7973 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6401), .ZN(n7265) );
  NOR2_X1 U7974 ( .A1(n7161), .A2(n6402), .ZN(n6403) );
  AOI211_X1 U7975 ( .C1(n9704), .C2(n6404), .A(n7265), .B(n6403), .ZN(n6405)
         );
  OAI211_X1 U7976 ( .C1(n9184), .C2(n6407), .A(n6406), .B(n6405), .ZN(P1_U3251) );
  INV_X1 U7977 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U7978 ( .A1(n6491), .A2(n9132), .ZN(n6408) );
  OAI21_X1 U7979 ( .B1(n9132), .B2(n6409), .A(n6408), .ZN(P1_U3555) );
  NAND2_X1 U7980 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6622) );
  OAI211_X1 U7981 ( .C1(n6412), .C2(n6411), .A(n9704), .B(n6410), .ZN(n6413)
         );
  OAI211_X1 U7982 ( .C1(n7161), .C2(n6415), .A(n6622), .B(n6413), .ZN(n6421)
         );
  INV_X1 U7983 ( .A(n6414), .ZN(n6419) );
  MUX2_X1 U7984 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6262), .S(n6415), .Z(n6418)
         );
  INV_X1 U7985 ( .A(n6416), .ZN(n6417) );
  AOI211_X1 U7986 ( .C1(n6419), .C2(n6418), .A(n6417), .B(n9695), .ZN(n6420)
         );
  AOI211_X1 U7987 ( .C1(n9703), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n6421), .B(
        n6420), .ZN(n6422) );
  INV_X1 U7988 ( .A(n6422), .ZN(P1_U3244) );
  OAI21_X1 U7989 ( .B1(n6425), .B2(n6424), .A(n6423), .ZN(n6551) );
  MUX2_X1 U7990 ( .A(n6426), .B(n6551), .S(n6268), .Z(n6430) );
  INV_X1 U7991 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6691) );
  AND2_X1 U7992 ( .A1(n9186), .A2(n6691), .ZN(n6428) );
  OAI21_X1 U7993 ( .B1(n9590), .B2(n6428), .A(n6427), .ZN(n9684) );
  OAI211_X1 U7994 ( .C1(n6430), .C2(n9686), .A(n6429), .B(n9684), .ZN(n6462)
         );
  INV_X1 U7995 ( .A(n6431), .ZN(n6444) );
  AOI21_X1 U7996 ( .B1(n6434), .B2(n6433), .A(n6432), .ZN(n6436) );
  AND2_X1 U7997 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6648) );
  INV_X1 U7998 ( .A(n6648), .ZN(n6435) );
  OAI21_X1 U7999 ( .B1(n9173), .B2(n6436), .A(n6435), .ZN(n6443) );
  INV_X1 U8000 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6441) );
  AOI21_X1 U8001 ( .B1(n6439), .B2(n6438), .A(n6437), .ZN(n6440) );
  OAI22_X1 U8002 ( .A1(n9184), .A2(n6441), .B1(n9695), .B2(n6440), .ZN(n6442)
         );
  AOI211_X1 U8003 ( .C1(n6444), .C2(n9698), .A(n6443), .B(n6442), .ZN(n6445)
         );
  NAND2_X1 U8004 ( .A1(n6462), .A2(n6445), .ZN(P1_U3245) );
  INV_X1 U8005 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6766) );
  OAI211_X1 U8006 ( .C1(n6448), .C2(n6447), .A(n9704), .B(n6446), .ZN(n6449)
         );
  OAI21_X1 U8007 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6766), .A(n6449), .ZN(n6459) );
  INV_X1 U8008 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6457) );
  MUX2_X1 U8009 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6761), .S(n6450), .Z(n6453)
         );
  NAND3_X1 U8010 ( .A1(n6453), .A2(n6452), .A3(n6451), .ZN(n6454) );
  NAND2_X1 U8011 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  OAI22_X1 U8012 ( .A1(n9184), .A2(n6457), .B1(n9695), .B2(n6456), .ZN(n6458)
         );
  AOI211_X1 U8013 ( .C1(n6460), .C2(n9698), .A(n6459), .B(n6458), .ZN(n6461)
         );
  NAND2_X1 U8014 ( .A1(n6462), .A2(n6461), .ZN(P1_U3243) );
  OAI21_X1 U8015 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6470), .A(n6463), .ZN(
        n6466) );
  INV_X1 U8016 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6464) );
  MUX2_X1 U8017 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6464), .S(n6580), .Z(n6465)
         );
  NAND2_X1 U8018 ( .A1(n6466), .A2(n6465), .ZN(n6573) );
  OAI21_X1 U8019 ( .B1(n6466), .B2(n6465), .A(n6573), .ZN(n6477) );
  INV_X1 U8020 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6469) );
  INV_X1 U8021 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6467) );
  NOR2_X1 U8022 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6467), .ZN(n7303) );
  AOI21_X1 U8023 ( .B1(n9698), .B2(n6580), .A(n7303), .ZN(n6468) );
  OAI21_X1 U8024 ( .B1(n9184), .B2(n6469), .A(n6468), .ZN(n6476) );
  XNOR2_X1 U8025 ( .A(n6580), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U8026 ( .A1(n6474), .A2(n6473), .ZN(n6579) );
  AOI211_X1 U8027 ( .C1(n6474), .C2(n6473), .A(n9695), .B(n6579), .ZN(n6475)
         );
  AOI211_X1 U8028 ( .C1(n9704), .C2(n6477), .A(n6476), .B(n6475), .ZN(n6478)
         );
  INV_X1 U8029 ( .A(n6478), .ZN(P1_U3253) );
  INV_X1 U8030 ( .A(n6479), .ZN(n6495) );
  AOI22_X1 U8031 ( .A1(n6856), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9595), .ZN(n6480) );
  OAI21_X1 U8032 ( .B1(n6495), .B2(n9597), .A(n6480), .ZN(P1_U3340) );
  INV_X1 U8033 ( .A(n6484), .ZN(n6488) );
  XOR2_X1 U8034 ( .A(n6482), .B(n6481), .Z(n6485) );
  OAI21_X1 U8035 ( .B1(n6485), .B2(n6484), .A(n6483), .ZN(n6486) );
  OAI21_X1 U8036 ( .B1(n6488), .B2(n6487), .A(n6486), .ZN(n6489) );
  NAND2_X1 U8037 ( .A1(n6489), .A2(n9678), .ZN(n6494) );
  NAND2_X1 U8038 ( .A1(n9677), .A2(n6490), .ZN(n6567) );
  NAND2_X1 U8039 ( .A1(n9131), .A2(n9456), .ZN(n6745) );
  INV_X1 U8040 ( .A(n9111), .ZN(n6830) );
  OAI22_X1 U8041 ( .A1(n6745), .A2(n9667), .B1(n6830), .B2(n6746), .ZN(n6492)
         );
  AOI21_X1 U8042 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6567), .A(n6492), .ZN(
        n6493) );
  OAI211_X1 U8043 ( .C1(n6741), .C2(n9056), .A(n6494), .B(n6493), .ZN(P1_U3220) );
  INV_X1 U8044 ( .A(n6782), .ZN(n6723) );
  OAI222_X1 U8045 ( .A1(n8987), .A2(n6496), .B1(n6866), .B2(n6495), .C1(n6723), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  AND2_X1 U8046 ( .A1(n7066), .A2(n8060), .ZN(n6499) );
  NAND2_X1 U8047 ( .A1(n6500), .A2(n6499), .ZN(n8079) );
  INV_X1 U8048 ( .A(n8079), .ZN(n6501) );
  OAI22_X1 U8049 ( .A1(n8191), .A2(n9858), .B1(n6501), .B2(n9600), .ZN(n6504)
         );
  OAI22_X1 U8050 ( .A1(n6704), .A2(n8167), .B1(n8166), .B2(n6876), .ZN(n6503)
         );
  AOI211_X1 U8051 ( .C1(n8180), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6506)
         );
  INV_X1 U8052 ( .A(n6506), .ZN(P2_U3224) );
  NAND2_X1 U8053 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6507), .ZN(n6508) );
  OAI211_X1 U8054 ( .C1(n9839), .C2(n6509), .A(n8065), .B(n6508), .ZN(n6524)
         );
  NAND2_X1 U8055 ( .A1(n6524), .A2(n5662), .ZN(n6510) );
  NAND2_X1 U8056 ( .A1(n6510), .A2(n8395), .ZN(n6545) );
  INV_X1 U8057 ( .A(n9620), .ZN(n9806) );
  NOR2_X1 U8058 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7107), .ZN(n6528) );
  XNOR2_X1 U8059 ( .A(n6539), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U8060 ( .A1(n8428), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6517) );
  INV_X1 U8061 ( .A(n6535), .ZN(n9619) );
  INV_X1 U8062 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9812) );
  MUX2_X1 U8063 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6511), .S(n9599), .Z(n9604)
         );
  MUX2_X1 U8064 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6512), .S(n6535), .Z(n9616)
         );
  NOR2_X1 U8065 ( .A1(n9617), .A2(n9616), .ZN(n9615) );
  AOI21_X1 U8066 ( .B1(n9619), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9615), .ZN(
        n8404) );
  OR2_X1 U8067 ( .A1(n8401), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8068 ( .A1(n8401), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8069 ( .A1(n6514), .A2(n6513), .ZN(n8403) );
  AOI21_X1 U8070 ( .B1(n8401), .B2(P2_REG1_REG_3__SCAN_IN), .A(n8402), .ZN(
        n8416) );
  NAND2_X1 U8071 ( .A1(n8414), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U8072 ( .B1(n8414), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6515), .ZN(
        n8417) );
  NOR2_X1 U8073 ( .A1(n8416), .A2(n8417), .ZN(n8415) );
  AOI21_X1 U8074 ( .B1(n8414), .B2(P2_REG1_REG_4__SCAN_IN), .A(n8415), .ZN(
        n8430) );
  OAI21_X1 U8075 ( .B1(n8428), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6517), .ZN(
        n8431) );
  INV_X1 U8076 ( .A(n8429), .ZN(n6516) );
  NAND2_X1 U8077 ( .A1(n6517), .A2(n6516), .ZN(n8444) );
  NAND2_X1 U8078 ( .A1(n8445), .A2(n8444), .ZN(n8443) );
  INV_X1 U8079 ( .A(n6539), .ZN(n8442) );
  NAND2_X1 U8080 ( .A1(n8442), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6518) );
  AND2_X1 U8081 ( .A1(n8443), .A2(n6518), .ZN(n8456) );
  NAND2_X1 U8082 ( .A1(n8454), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6519) );
  OAI21_X1 U8083 ( .B1(n8454), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6519), .ZN(
        n8455) );
  XNOR2_X1 U8084 ( .A(n6542), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U8085 ( .A1(n8469), .A2(n8470), .ZN(n8468) );
  NAND2_X1 U8086 ( .A1(n4539), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8087 ( .A1(n8468), .A2(n6520), .ZN(n8482) );
  NAND2_X1 U8088 ( .A1(n8479), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6521) );
  OAI21_X1 U8089 ( .B1(n8479), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6521), .ZN(
        n6522) );
  INV_X1 U8090 ( .A(n6522), .ZN(n8483) );
  AOI21_X1 U8091 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n8479), .A(n8480), .ZN(
        n6526) );
  MUX2_X1 U8092 ( .A(n9935), .B(P2_REG1_REG_10__SCAN_IN), .S(n6602), .Z(n6525)
         );
  AND2_X1 U8093 ( .A1(n5662), .A2(n8985), .ZN(n6523) );
  INV_X1 U8094 ( .A(n9804), .ZN(n9614) );
  AOI211_X1 U8095 ( .C1(n6526), .C2(n6525), .A(n6601), .B(n9614), .ZN(n6527)
         );
  AOI211_X1 U8096 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9809), .A(n6528), .B(
        n6527), .ZN(n6549) );
  NAND2_X1 U8097 ( .A1(n8479), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6543) );
  MUX2_X1 U8098 ( .A(n5811), .B(P2_REG2_REG_9__SCAN_IN), .S(n8479), .Z(n6529)
         );
  INV_X1 U8099 ( .A(n6529), .ZN(n8477) );
  NAND2_X1 U8100 ( .A1(n8454), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6541) );
  MUX2_X1 U8101 ( .A(n5778), .B(P2_REG2_REG_7__SCAN_IN), .S(n8454), .Z(n6530)
         );
  INV_X1 U8102 ( .A(n6530), .ZN(n8451) );
  NAND2_X1 U8103 ( .A1(n8428), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6538) );
  MUX2_X1 U8104 ( .A(n6892), .B(P2_REG2_REG_5__SCAN_IN), .S(n8428), .Z(n6531)
         );
  INV_X1 U8105 ( .A(n6531), .ZN(n8424) );
  NAND2_X1 U8106 ( .A1(n8414), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U8107 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6532), .S(n8414), .Z(n8411)
         );
  NAND2_X1 U8108 ( .A1(n8401), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6536) );
  MUX2_X1 U8109 ( .A(n5706), .B(P2_REG2_REG_3__SCAN_IN), .S(n8401), .Z(n6533)
         );
  INV_X1 U8110 ( .A(n6533), .ZN(n8397) );
  XNOR2_X1 U8111 ( .A(n6535), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9623) );
  MUX2_X1 U8112 ( .A(n6707), .B(P2_REG2_REG_1__SCAN_IN), .S(n9599), .Z(n9610)
         );
  NAND3_X1 U8113 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9610), .ZN(n9609) );
  OAI21_X1 U8114 ( .B1(n9599), .B2(n6707), .A(n9609), .ZN(n9622) );
  NAND2_X1 U8115 ( .A1(n9623), .A2(n9622), .ZN(n9621) );
  OAI21_X1 U8116 ( .B1(n6535), .B2(n6534), .A(n9621), .ZN(n8398) );
  NAND2_X1 U8117 ( .A1(n8397), .A2(n8398), .ZN(n8396) );
  NAND2_X1 U8118 ( .A1(n6536), .A2(n8396), .ZN(n8412) );
  NAND2_X1 U8119 ( .A1(n8411), .A2(n8412), .ZN(n8410) );
  NAND2_X1 U8120 ( .A1(n6537), .A2(n8410), .ZN(n8425) );
  NAND2_X1 U8121 ( .A1(n8424), .A2(n8425), .ZN(n8423) );
  NAND2_X1 U8122 ( .A1(n6538), .A2(n8423), .ZN(n8439) );
  MUX2_X1 U8123 ( .A(n6540), .B(P2_REG2_REG_6__SCAN_IN), .S(n6539), .Z(n8438)
         );
  NAND2_X1 U8124 ( .A1(n8439), .A2(n8438), .ZN(n8437) );
  OAI21_X1 U8125 ( .B1(n6540), .B2(n6539), .A(n8437), .ZN(n8452) );
  NAND2_X1 U8126 ( .A1(n8451), .A2(n8452), .ZN(n8450) );
  NAND2_X1 U8127 ( .A1(n6541), .A2(n8450), .ZN(n8465) );
  MUX2_X1 U8128 ( .A(n7097), .B(P2_REG2_REG_8__SCAN_IN), .S(n6542), .Z(n8464)
         );
  NAND2_X1 U8129 ( .A1(n8465), .A2(n8464), .ZN(n8463) );
  OAI21_X1 U8130 ( .B1(n7097), .B2(n6542), .A(n8463), .ZN(n8476) );
  NAND2_X1 U8131 ( .A1(n8477), .A2(n8476), .ZN(n8475) );
  NAND2_X1 U8132 ( .A1(n6543), .A2(n8475), .ZN(n6547) );
  MUX2_X1 U8133 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7412), .S(n6602), .Z(n6546)
         );
  NOR2_X1 U8134 ( .A1(n6142), .A2(n8985), .ZN(n6544) );
  INV_X1 U8135 ( .A(n9807), .ZN(n9803) );
  NAND2_X1 U8136 ( .A1(n6546), .A2(n6547), .ZN(n6596) );
  OAI211_X1 U8137 ( .C1(n6547), .C2(n6546), .A(n9803), .B(n6596), .ZN(n6548)
         );
  OAI211_X1 U8138 ( .C1(n9806), .C2(n6550), .A(n6549), .B(n6548), .ZN(P2_U3255) );
  INV_X1 U8139 ( .A(n9096), .ZN(n6568) );
  AOI22_X1 U8140 ( .A1(n6551), .A2(n9678), .B1(n6568), .B2(n9133), .ZN(n6553)
         );
  AOI22_X1 U8141 ( .A1(n9115), .A2(n6693), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6567), .ZN(n6552) );
  NAND2_X1 U8142 ( .A1(n6553), .A2(n6552), .ZN(P1_U3230) );
  XNOR2_X1 U8143 ( .A(n6555), .B(n6554), .ZN(n6559) );
  NOR2_X1 U8144 ( .A1(n8191), .A2(n9862), .ZN(n6557) );
  INV_X2 U8145 ( .A(n6697), .ZN(n6696) );
  OAI22_X1 U8146 ( .A1(n6696), .A2(n8167), .B1(n8166), .B2(n6953), .ZN(n6556)
         );
  AOI211_X1 U8147 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n8079), .A(n6557), .B(
        n6556), .ZN(n6558) );
  OAI21_X1 U8148 ( .B1(n6559), .B2(n8204), .A(n6558), .ZN(P2_U3239) );
  INV_X1 U8149 ( .A(n6560), .ZN(n6562) );
  OAI222_X1 U8150 ( .A1(n9593), .A2(n6561), .B1(n9597), .B2(n6562), .C1(n7028), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8151 ( .A(n6982), .ZN(n6722) );
  OAI222_X1 U8152 ( .A1(n8987), .A2(n6563), .B1(n6866), .B2(n6562), .C1(n6722), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  AOI21_X1 U8153 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6571) );
  AOI22_X1 U8154 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n6567), .B1(n9133), .B2(
        n9111), .ZN(n6570) );
  AOI22_X1 U8155 ( .A1(n6568), .A2(n9130), .B1(n9115), .B2(n6768), .ZN(n6569)
         );
  OAI211_X1 U8156 ( .C1(n6571), .C2(n9117), .A(n6570), .B(n6569), .ZN(P1_U3235) );
  INV_X1 U8157 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6572) );
  MUX2_X1 U8158 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6572), .S(n6856), .Z(n6575)
         );
  OAI21_X1 U8159 ( .B1(n6580), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6573), .ZN(
        n6574) );
  NAND2_X1 U8160 ( .A1(n6574), .A2(n6575), .ZN(n6851) );
  OAI21_X1 U8161 ( .B1(n6575), .B2(n6574), .A(n6851), .ZN(n6586) );
  INV_X1 U8162 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U8163 ( .A1(n9698), .A2(n6856), .ZN(n6577) );
  NOR2_X1 U8164 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5287), .ZN(n7428) );
  INV_X1 U8165 ( .A(n7428), .ZN(n6576) );
  OAI211_X1 U8166 ( .C1(n9184), .C2(n6578), .A(n6577), .B(n6576), .ZN(n6585)
         );
  AOI21_X1 U8167 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6580), .A(n6579), .ZN(
        n6583) );
  NAND2_X1 U8168 ( .A1(n6856), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6581) );
  OAI21_X1 U8169 ( .B1(n6856), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6581), .ZN(
        n6582) );
  NOR2_X1 U8170 ( .A1(n6583), .A2(n6582), .ZN(n6855) );
  AOI211_X1 U8171 ( .C1(n6583), .C2(n6582), .A(n9695), .B(n6855), .ZN(n6584)
         );
  AOI211_X1 U8172 ( .C1(n9704), .C2(n6586), .A(n6585), .B(n6584), .ZN(n6587)
         );
  INV_X1 U8173 ( .A(n6587), .ZN(P1_U3254) );
  XNOR2_X1 U8174 ( .A(n6589), .B(n6588), .ZN(n6595) );
  INV_X1 U8175 ( .A(n6590), .ZN(n8197) );
  NAND2_X1 U8176 ( .A1(n8394), .A2(n8819), .ZN(n6592) );
  NAND2_X1 U8177 ( .A1(n8392), .A2(n8821), .ZN(n6591) );
  NAND2_X1 U8178 ( .A1(n6592), .A2(n6591), .ZN(n7013) );
  AOI22_X1 U8179 ( .A1(n8197), .A2(n7013), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6594) );
  INV_X1 U8180 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8399) );
  AOI22_X1 U8181 ( .A1(n8202), .A2(n6869), .B1(n8399), .B2(n8137), .ZN(n6593)
         );
  OAI211_X1 U8182 ( .C1(n6595), .C2(n8204), .A(n6594), .B(n6593), .ZN(P2_U3220) );
  NAND2_X1 U8183 ( .A1(n6602), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8184 ( .A1(n6597), .A2(n6596), .ZN(n6600) );
  MUX2_X1 U8185 ( .A(n6598), .B(P2_REG2_REG_11__SCAN_IN), .S(n6724), .Z(n6599)
         );
  NOR2_X1 U8186 ( .A1(n6600), .A2(n6599), .ZN(n6716) );
  AOI21_X1 U8187 ( .B1(n6600), .B2(n6599), .A(n6716), .ZN(n6610) );
  NOR2_X1 U8188 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5858), .ZN(n6607) );
  AOI21_X1 U8189 ( .B1(n6602), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6601), .ZN(
        n6605) );
  INV_X1 U8190 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U8191 ( .A(n6603), .B(P2_REG1_REG_11__SCAN_IN), .S(n6724), .Z(n6604)
         );
  NOR2_X1 U8192 ( .A1(n6605), .A2(n6604), .ZN(n6725) );
  AOI211_X1 U8193 ( .C1(n6605), .C2(n6604), .A(n6725), .B(n9614), .ZN(n6606)
         );
  AOI211_X1 U8194 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9809), .A(n6607), .B(
        n6606), .ZN(n6609) );
  NAND2_X1 U8195 ( .A1(n9620), .A2(n6724), .ZN(n6608) );
  OAI211_X1 U8196 ( .C1(n6610), .C2(n9807), .A(n6609), .B(n6608), .ZN(P2_U3256) );
  INV_X1 U8197 ( .A(n6611), .ZN(n6613) );
  INV_X1 U8198 ( .A(n7153), .ZN(n6612) );
  OAI222_X1 U8199 ( .A1(n9593), .A2(n8298), .B1(n9597), .B2(n6613), .C1(
        P1_U3084), .C2(n6612), .ZN(P1_U3338) );
  INV_X1 U8200 ( .A(n8514), .ZN(n8505) );
  OAI222_X1 U8201 ( .A1(n8987), .A2(n6614), .B1(n6866), .B2(n6613), .C1(
        P2_U3152), .C2(n8505), .ZN(P2_U3343) );
  INV_X1 U8202 ( .A(n6615), .ZN(n6617) );
  INV_X1 U8203 ( .A(n9148), .ZN(n7162) );
  OAI222_X1 U8204 ( .A1(n9593), .A2(n6616), .B1(n9597), .B2(n6617), .C1(n7162), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8205 ( .A(n8532), .ZN(n8518) );
  OAI222_X1 U8206 ( .A1(n8987), .A2(n6618), .B1(n6866), .B2(n6617), .C1(n8518), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  AOI21_X1 U8207 ( .B1(n6621), .B2(n6620), .A(n6619), .ZN(n6626) );
  OAI21_X1 U8208 ( .B1(n6830), .B2(n6674), .A(n6622), .ZN(n6624) );
  OAI22_X1 U8209 ( .A1(n9096), .A2(n6829), .B1(n9683), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n6623) );
  AOI211_X1 U8210 ( .C1(n9115), .C2(n9725), .A(n6624), .B(n6623), .ZN(n6625)
         );
  OAI21_X1 U8211 ( .B1(n6626), .B2(n9117), .A(n6625), .ZN(P1_U3216) );
  INV_X1 U8212 ( .A(n6627), .ZN(n6654) );
  AOI22_X1 U8213 ( .A1(n9171), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9595), .ZN(n6628) );
  OAI21_X1 U8214 ( .B1(n6654), .B2(n9597), .A(n6628), .ZN(P1_U3336) );
  AOI21_X1 U8215 ( .B1(n6630), .B2(n6629), .A(n4396), .ZN(n6634) );
  INV_X1 U8216 ( .A(n8391), .ZN(n6931) );
  OAI22_X1 U8217 ( .A1(n6931), .A2(n8806), .B1(n6953), .B2(n8804), .ZN(n9817)
         );
  AOI22_X1 U8218 ( .A1(n8197), .A2(n9817), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6633) );
  INV_X1 U8219 ( .A(n9828), .ZN(n6631) );
  AOI22_X1 U8220 ( .A1(n8202), .A2(n9830), .B1(n8137), .B2(n6631), .ZN(n6632)
         );
  OAI211_X1 U8221 ( .C1(n6634), .C2(n8204), .A(n6633), .B(n6632), .ZN(P2_U3232) );
  XNOR2_X1 U8222 ( .A(n6636), .B(n6635), .ZN(n6643) );
  NAND2_X1 U8223 ( .A1(n8392), .A2(n8819), .ZN(n6638) );
  NAND2_X1 U8224 ( .A1(n8213), .A2(n8821), .ZN(n6637) );
  AND2_X1 U8225 ( .A1(n6638), .A2(n6637), .ZN(n6890) );
  INV_X1 U8226 ( .A(n6890), .ZN(n6639) );
  AOI22_X1 U8227 ( .A1(n8197), .A2(n6639), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6642) );
  INV_X1 U8228 ( .A(n6640), .ZN(n6894) );
  AOI22_X1 U8229 ( .A1(n8202), .A2(n9885), .B1(n8137), .B2(n6894), .ZN(n6641)
         );
  OAI211_X1 U8230 ( .C1(n6643), .C2(n8204), .A(n6642), .B(n6641), .ZN(P2_U3229) );
  OR2_X1 U8231 ( .A1(n6619), .A2(n6644), .ZN(n6646) );
  AOI211_X1 U8232 ( .C1(n6647), .C2(n6646), .A(n9117), .B(n6645), .ZN(n6653)
         );
  AOI21_X1 U8233 ( .B1(n9130), .B2(n9111), .A(n6648), .ZN(n6649) );
  OAI21_X1 U8234 ( .B1(n9732), .B2(n9056), .A(n6649), .ZN(n6652) );
  INV_X1 U8235 ( .A(n6650), .ZN(n6817) );
  OAI22_X1 U8236 ( .A1(n9096), .A2(n6918), .B1(n9683), .B2(n6817), .ZN(n6651)
         );
  OR3_X1 U8237 ( .A1(n6653), .A2(n6652), .A3(n6651), .ZN(P1_U3228) );
  INV_X1 U8238 ( .A(n8546), .ZN(n8539) );
  OAI222_X1 U8239 ( .A1(n8987), .A2(n6655), .B1(n6866), .B2(n6654), .C1(n8539), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U8240 ( .A1(n6755), .A2(n6681), .ZN(n6671) );
  NAND2_X1 U8241 ( .A1(n6744), .A2(n6671), .ZN(n6656) );
  NAND2_X1 U8242 ( .A1(n6656), .A2(n7765), .ZN(n6756) );
  NAND2_X1 U8243 ( .A1(n6674), .A2(n6768), .ZN(n6657) );
  NAND2_X1 U8244 ( .A1(n6808), .A2(n9725), .ZN(n7537) );
  INV_X1 U8245 ( .A(n6793), .ZN(n6658) );
  XNOR2_X1 U8246 ( .A(n7636), .B(n6658), .ZN(n6662) );
  NAND2_X1 U8247 ( .A1(n5061), .A2(n9315), .ZN(n6660) );
  NAND2_X1 U8248 ( .A1(n7762), .A2(n6743), .ZN(n6659) );
  OAI22_X1 U8249 ( .A1(n6674), .A2(n9438), .B1(n6829), .B2(n9440), .ZN(n6661)
         );
  AOI21_X1 U8250 ( .B1(n6662), .B2(n9459), .A(n6661), .ZN(n9730) );
  NOR2_X1 U8251 ( .A1(n6664), .A2(n6663), .ZN(n6665) );
  NAND2_X1 U8252 ( .A1(n6667), .A2(n6666), .ZN(n6669) );
  NAND2_X1 U8253 ( .A1(n6669), .A2(n6668), .ZN(n7382) );
  NOR2_X1 U8254 ( .A1(n7388), .A2(n7382), .ZN(n6670) );
  NAND2_X1 U8255 ( .A1(n7386), .A2(n6670), .ZN(n6789) );
  NAND2_X1 U8256 ( .A1(n6491), .A2(n6693), .ZN(n6738) );
  NAND2_X1 U8257 ( .A1(n6737), .A2(n6738), .ZN(n6673) );
  NAND2_X1 U8258 ( .A1(n6755), .A2(n6741), .ZN(n6672) );
  NAND2_X1 U8259 ( .A1(n6673), .A2(n6672), .ZN(n6754) );
  NAND2_X1 U8260 ( .A1(n6674), .A2(n9718), .ZN(n6675) );
  XNOR2_X1 U8261 ( .A(n6794), .B(n6793), .ZN(n9727) );
  NAND2_X1 U8262 ( .A1(n6677), .A2(n9315), .ZN(n6739) );
  NAND2_X1 U8263 ( .A1(n6676), .A2(n6739), .ZN(n6678) );
  INV_X1 U8264 ( .A(n9450), .ZN(n9472) );
  NOR2_X1 U8265 ( .A1(n9561), .A2(n7795), .ZN(n6680) );
  NAND2_X1 U8266 ( .A1(n6763), .A2(n6795), .ZN(n6815) );
  OR2_X1 U8267 ( .A1(n6763), .A2(n6795), .ZN(n6682) );
  AND2_X1 U8268 ( .A1(n6815), .A2(n6682), .ZN(n9726) );
  OAI22_X1 U8269 ( .A1(n9460), .A2(n6262), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9465), .ZN(n6683) );
  AOI21_X1 U8270 ( .B1(n9429), .B2(n9726), .A(n6683), .ZN(n6684) );
  OAI21_X1 U8271 ( .B1(n6795), .B2(n9467), .A(n6684), .ZN(n6685) );
  AOI21_X1 U8272 ( .B1(n9727), .B2(n9472), .A(n6685), .ZN(n6686) );
  OAI21_X1 U8273 ( .B1(n9730), .B2(n9305), .A(n6686), .ZN(P1_U3288) );
  INV_X1 U8274 ( .A(n6693), .ZN(n9562) );
  NAND2_X1 U8275 ( .A1(n6491), .A2(n9562), .ZN(n7763) );
  NAND2_X1 U8276 ( .A1(n6744), .A2(n7763), .ZN(n7534) );
  INV_X1 U8277 ( .A(n9561), .ZN(n6687) );
  NOR2_X1 U8278 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  AOI22_X1 U8279 ( .A1(n7534), .A2(n6689), .B1(n9456), .B2(n9133), .ZN(n9560)
         );
  INV_X1 U8280 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6690) );
  OAI22_X1 U8281 ( .A1(n9460), .A2(n6691), .B1(n6690), .B2(n9465), .ZN(n6692)
         );
  INV_X1 U8282 ( .A(n6692), .ZN(n6695) );
  OAI21_X1 U8283 ( .B1(n9374), .B2(n9429), .A(n6693), .ZN(n6694) );
  OAI211_X1 U8284 ( .C1(n9560), .C2(n9305), .A(n6695), .B(n6694), .ZN(P1_U3291) );
  XNOR2_X1 U8285 ( .A(n6873), .B(n6871), .ZN(n9853) );
  NOR2_X1 U8286 ( .A1(n7076), .A2(n9839), .ZN(n6698) );
  NAND3_X1 U8287 ( .A1(n6699), .A2(n6698), .A3(n7066), .ZN(n6710) );
  XNOR2_X1 U8288 ( .A(n6700), .B(n8063), .ZN(n8772) );
  NAND2_X1 U8289 ( .A1(n8772), .A2(n8807), .ZN(n7465) );
  OR2_X1 U8290 ( .A1(n6700), .A2(n8807), .ZN(n7007) );
  NAND2_X1 U8291 ( .A1(n7465), .A2(n7007), .ZN(n6701) );
  INV_X1 U8292 ( .A(n7021), .ZN(n8083) );
  OR2_X1 U8293 ( .A1(n6118), .A2(n7895), .ZN(n7864) );
  OAI21_X1 U8294 ( .B1(n7911), .B2(n6702), .A(n8824), .ZN(n6703) );
  AOI21_X1 U8295 ( .B1(n8083), .B2(n6873), .A(n6703), .ZN(n6706) );
  OAI22_X1 U8296 ( .A1(n6704), .A2(n8804), .B1(n6876), .B2(n8806), .ZN(n6705)
         );
  NOR2_X1 U8297 ( .A1(n6706), .A2(n6705), .ZN(n9857) );
  MUX2_X1 U8298 ( .A(n6707), .B(n9857), .S(n4316), .Z(n6715) );
  NOR2_X2 U8299 ( .A1(n8846), .A2(n6709), .ZN(n9831) );
  INV_X1 U8300 ( .A(n8082), .ZN(n9849) );
  NAND2_X1 U8301 ( .A1(n9849), .A2(n9858), .ZN(n9854) );
  OR2_X1 U8302 ( .A1(n9858), .A2(n9849), .ZN(n9855) );
  NAND3_X1 U8303 ( .A1(n8858), .A2(n9854), .A3(n9855), .ZN(n6711) );
  OAI21_X1 U8304 ( .B1(n9827), .B2(n9600), .A(n6711), .ZN(n6712) );
  AOI21_X1 U8305 ( .B1(n9831), .B2(n6713), .A(n6712), .ZN(n6714) );
  OAI211_X1 U8306 ( .C1(n9853), .C2(n9825), .A(n6715), .B(n6714), .ZN(P2_U3295) );
  NOR2_X1 U8307 ( .A1(n6782), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U8308 ( .A1(n8494), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6718) );
  INV_X1 U8309 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8488) );
  AOI21_X1 U8310 ( .B1(n6717), .B2(n6598), .A(n6716), .ZN(n8491) );
  OAI211_X1 U8311 ( .C1(n8494), .C2(P2_REG2_REG_12__SCAN_IN), .A(n8491), .B(
        n6718), .ZN(n8489) );
  NAND2_X1 U8312 ( .A1(n6718), .A2(n8489), .ZN(n6774) );
  AOI22_X1 U8313 ( .A1(n6782), .A2(n5881), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6723), .ZN(n6773) );
  NOR2_X1 U8314 ( .A1(n6774), .A2(n6773), .ZN(n6772) );
  NOR2_X1 U8315 ( .A1(n6719), .A2(n6772), .ZN(n6721) );
  AOI22_X1 U8316 ( .A1(n6982), .A2(n7515), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n6722), .ZN(n6720) );
  NOR2_X1 U8317 ( .A1(n6721), .A2(n6720), .ZN(n6978) );
  AOI21_X1 U8318 ( .B1(n6721), .B2(n6720), .A(n6978), .ZN(n6736) );
  AOI22_X1 U8319 ( .A1(n6982), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n5896), .B2(
        n6722), .ZN(n6730) );
  AOI22_X1 U8320 ( .A1(n6782), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5880), .B2(
        n6723), .ZN(n6776) );
  NAND2_X1 U8321 ( .A1(n6724), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6727) );
  INV_X1 U8322 ( .A(n6725), .ZN(n6726) );
  NAND2_X1 U8323 ( .A1(n6727), .A2(n6726), .ZN(n8496) );
  MUX2_X1 U8324 ( .A(n5861), .B(P2_REG1_REG_12__SCAN_IN), .S(n8494), .Z(n8495)
         );
  OR2_X1 U8325 ( .A1(n8494), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8326 ( .A1(n8498), .A2(n6728), .ZN(n6777) );
  NAND2_X1 U8327 ( .A1(n6776), .A2(n6777), .ZN(n6775) );
  OAI21_X1 U8328 ( .B1(n6782), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6775), .ZN(
        n6729) );
  OAI21_X1 U8329 ( .B1(n6730), .B2(n6729), .A(n6981), .ZN(n6731) );
  NAND2_X1 U8330 ( .A1(n6731), .A2(n9804), .ZN(n6735) );
  INV_X1 U8331 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U8332 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7525) );
  OAI21_X1 U8333 ( .B1(n9602), .B2(n6732), .A(n7525), .ZN(n6733) );
  AOI21_X1 U8334 ( .B1(n9620), .B2(n6982), .A(n6733), .ZN(n6734) );
  OAI211_X1 U8335 ( .C1(n6736), .C2(n9807), .A(n6735), .B(n6734), .ZN(P2_U3259) );
  XOR2_X1 U8336 ( .A(n6737), .B(n6738), .Z(n9712) );
  INV_X1 U8337 ( .A(n7372), .ZN(n7250) );
  OAI21_X1 U8338 ( .B1(n6741), .B2(n9562), .A(n9749), .ZN(n6740) );
  OAI21_X1 U8339 ( .B1(n6741), .B2(n9773), .A(n6740), .ZN(n6742) );
  NAND2_X1 U8340 ( .A1(n6742), .A2(n6762), .ZN(n9713) );
  NOR2_X1 U8341 ( .A1(n9713), .A2(n9770), .ZN(n6750) );
  XNOR2_X1 U8342 ( .A(n6737), .B(n6744), .ZN(n6748) );
  OAI21_X1 U8343 ( .B1(n6746), .B2(n9438), .A(n6745), .ZN(n6747) );
  AOI21_X1 U8344 ( .B1(n6748), .B2(n9459), .A(n6747), .ZN(n6749) );
  OAI21_X1 U8345 ( .B1(n9712), .B2(n6676), .A(n6749), .ZN(n9714) );
  AOI211_X1 U8346 ( .C1(n9444), .C2(P1_REG3_REG_1__SCAN_IN), .A(n6750), .B(
        n9714), .ZN(n6751) );
  MUX2_X1 U8347 ( .A(n6752), .B(n6751), .S(n9460), .Z(n6753) );
  OAI21_X1 U8348 ( .B1(n9712), .B2(n7250), .A(n6753), .ZN(P1_U3290) );
  XNOR2_X1 U8349 ( .A(n6754), .B(n7535), .ZN(n9723) );
  INV_X1 U8350 ( .A(n9723), .ZN(n6771) );
  INV_X1 U8351 ( .A(n6676), .ZN(n7362) );
  OAI22_X1 U8352 ( .A1(n6808), .A2(n9440), .B1(n6755), .B2(n9438), .ZN(n6760)
         );
  NAND2_X1 U8353 ( .A1(n6756), .A2(n7535), .ZN(n6757) );
  AOI21_X1 U8354 ( .B1(n6758), .B2(n6757), .A(n9436), .ZN(n6759) );
  AOI211_X1 U8355 ( .C1(n7362), .C2(n9723), .A(n6760), .B(n6759), .ZN(n9720)
         );
  MUX2_X1 U8356 ( .A(n6761), .B(n9720), .S(n9460), .Z(n6770) );
  INV_X1 U8357 ( .A(n6762), .ZN(n6765) );
  INV_X1 U8358 ( .A(n6763), .ZN(n6764) );
  OAI21_X1 U8359 ( .B1(n9718), .B2(n6765), .A(n6764), .ZN(n9719) );
  OAI22_X1 U8360 ( .A1(n9376), .A2(n9719), .B1(n6766), .B2(n9465), .ZN(n6767)
         );
  AOI21_X1 U8361 ( .B1(n9374), .B2(n6768), .A(n6767), .ZN(n6769) );
  OAI211_X1 U8362 ( .C1(n6771), .C2(n7250), .A(n6770), .B(n6769), .ZN(P1_U3289) );
  AOI21_X1 U8363 ( .B1(n6774), .B2(n6773), .A(n6772), .ZN(n6784) );
  INV_X1 U8364 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6780) );
  OAI21_X1 U8365 ( .B1(n6777), .B2(n6776), .A(n6775), .ZN(n6778) );
  NAND2_X1 U8366 ( .A1(n9804), .A2(n6778), .ZN(n6779) );
  NAND2_X1 U8367 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7445) );
  OAI211_X1 U8368 ( .C1(n9602), .C2(n6780), .A(n6779), .B(n7445), .ZN(n6781)
         );
  AOI21_X1 U8369 ( .B1(n6782), .B2(n9620), .A(n6781), .ZN(n6783) );
  OAI21_X1 U8370 ( .B1(n6784), .B2(n9807), .A(n6783), .ZN(P2_U3258) );
  INV_X1 U8371 ( .A(n7537), .ZN(n6785) );
  NAND2_X1 U8372 ( .A1(n6829), .A2(n6819), .ZN(n7538) );
  INV_X1 U8373 ( .A(n6829), .ZN(n9455) );
  NAND2_X1 U8374 ( .A1(n9455), .A2(n9732), .ZN(n9451) );
  NAND2_X1 U8375 ( .A1(n9129), .A2(n9466), .ZN(n6799) );
  AND2_X1 U8376 ( .A1(n9451), .A2(n6799), .ZN(n7539) );
  NAND2_X1 U8377 ( .A1(n6918), .A2(n9740), .ZN(n7541) );
  NAND2_X1 U8378 ( .A1(n6832), .A2(n4315), .ZN(n7542) );
  NAND2_X1 U8379 ( .A1(n9457), .A2(n6924), .ZN(n7637) );
  NAND2_X1 U8380 ( .A1(n9095), .A2(n6792), .ZN(n7630) );
  NAND2_X1 U8381 ( .A1(n9128), .A2(n9759), .ZN(n7768) );
  NAND2_X1 U8382 ( .A1(n7630), .A2(n7768), .ZN(n6897) );
  INV_X1 U8383 ( .A(n6897), .ZN(n7546) );
  XNOR2_X1 U8384 ( .A(n7770), .B(n7546), .ZN(n6787) );
  AOI222_X1 U8385 ( .A1(n9459), .A2(n6787), .B1(n9127), .B2(n9456), .C1(n9457), 
        .C2(n9454), .ZN(n9758) );
  INV_X1 U8386 ( .A(n6969), .ZN(n6788) );
  OAI22_X1 U8387 ( .A1(n9460), .A2(n6305), .B1(n6788), .B2(n9465), .ZN(n6791)
         );
  OR2_X1 U8388 ( .A1(n9463), .A2(n9740), .ZN(n9461) );
  NAND2_X1 U8389 ( .A1(n6922), .A2(n9759), .ZN(n6907) );
  OAI211_X1 U8390 ( .C1(n6922), .C2(n9759), .A(n6907), .B(n9749), .ZN(n9757)
         );
  NOR2_X1 U8391 ( .A1(n6789), .A2(n9315), .ZN(n9469) );
  INV_X1 U8392 ( .A(n9469), .ZN(n7329) );
  NOR2_X1 U8393 ( .A1(n9757), .A2(n7329), .ZN(n6790) );
  AOI211_X1 U8394 ( .C1(n9374), .C2(n6792), .A(n6791), .B(n6790), .ZN(n6806)
         );
  NAND2_X1 U8395 ( .A1(n6808), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U8396 ( .A1(n7538), .A2(n9451), .ZN(n6812) );
  NAND2_X1 U8397 ( .A1(n6811), .A2(n6812), .ZN(n6798) );
  NAND2_X1 U8398 ( .A1(n6829), .A2(n9732), .ZN(n6797) );
  INV_X1 U8399 ( .A(n9471), .ZN(n6801) );
  NAND2_X1 U8400 ( .A1(n9129), .A2(n9740), .ZN(n6802) );
  NAND2_X1 U8401 ( .A1(n6832), .A2(n6924), .ZN(n6804) );
  XNOR2_X1 U8402 ( .A(n6898), .B(n6897), .ZN(n9761) );
  NAND2_X1 U8403 ( .A1(n9761), .A2(n9472), .ZN(n6805) );
  OAI211_X1 U8404 ( .C1(n9758), .C2(n9305), .A(n6806), .B(n6805), .ZN(P1_U3284) );
  XNOR2_X1 U8405 ( .A(n6807), .B(n6812), .ZN(n6810) );
  OAI22_X1 U8406 ( .A1(n6808), .A2(n9438), .B1(n6918), .B2(n9440), .ZN(n6809)
         );
  AOI21_X1 U8407 ( .B1(n6810), .B2(n9459), .A(n6809), .ZN(n6814) );
  XNOR2_X1 U8408 ( .A(n6811), .B(n6812), .ZN(n9735) );
  NAND2_X1 U8409 ( .A1(n9735), .A2(n7362), .ZN(n6813) );
  NAND2_X1 U8410 ( .A1(n6815), .A2(n6819), .ZN(n6816) );
  NAND2_X1 U8411 ( .A1(n9463), .A2(n6816), .ZN(n9733) );
  OAI22_X1 U8412 ( .A1(n9460), .A2(n6265), .B1(n6817), .B2(n9465), .ZN(n6818)
         );
  AOI21_X1 U8413 ( .B1(n9374), .B2(n6819), .A(n6818), .ZN(n6820) );
  OAI21_X1 U8414 ( .B1(n9376), .B2(n9733), .A(n6820), .ZN(n6821) );
  AOI21_X1 U8415 ( .B1(n9735), .B2(n7372), .A(n6821), .ZN(n6822) );
  OAI21_X1 U8416 ( .B1(n9737), .B2(n9305), .A(n6822), .ZN(P1_U3287) );
  INV_X1 U8417 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8215) );
  INV_X1 U8418 ( .A(n6823), .ZN(n6824) );
  INV_X1 U8419 ( .A(n9699), .ZN(n9169) );
  OAI222_X1 U8420 ( .A1(n9593), .A2(n8215), .B1(n9597), .B2(n6824), .C1(
        P1_U3084), .C2(n9169), .ZN(P1_U3335) );
  INV_X1 U8421 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8382) );
  INV_X1 U8422 ( .A(n8551), .ZN(n8558) );
  OAI222_X1 U8423 ( .A1(n8987), .A2(n8382), .B1(n6866), .B2(n6824), .C1(
        P2_U3152), .C2(n8558), .ZN(P2_U3340) );
  AOI21_X1 U8424 ( .B1(n6826), .B2(n6825), .A(n9092), .ZN(n6836) );
  INV_X1 U8425 ( .A(n6827), .ZN(n6828) );
  OAI21_X1 U8426 ( .B1(n6830), .B2(n6829), .A(n6828), .ZN(n6834) );
  INV_X1 U8427 ( .A(n6831), .ZN(n9464) );
  OAI22_X1 U8428 ( .A1(n9096), .A2(n6832), .B1(n9683), .B2(n9464), .ZN(n6833)
         );
  AOI211_X1 U8429 ( .C1(n9115), .C2(n9740), .A(n6834), .B(n6833), .ZN(n6835)
         );
  OAI21_X1 U8430 ( .B1(n6836), .B2(n9117), .A(n6835), .ZN(P1_U3225) );
  OAI21_X1 U8431 ( .B1(n6839), .B2(n6838), .A(n6837), .ZN(n6843) );
  INV_X1 U8432 ( .A(n8212), .ZN(n7084) );
  OAI22_X1 U8433 ( .A1(n8166), .A2(n7084), .B1(n9894), .B2(n8191), .ZN(n6842)
         );
  NAND2_X1 U8434 ( .A1(n8175), .A2(n8391), .ZN(n6840) );
  NAND2_X1 U8435 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8440) );
  OAI211_X1 U8436 ( .C1(n8200), .C2(n7003), .A(n6840), .B(n8440), .ZN(n6841)
         );
  AOI211_X1 U8437 ( .C1(n6843), .C2(n8180), .A(n6842), .B(n6841), .ZN(n6844)
         );
  INV_X1 U8438 ( .A(n6844), .ZN(P2_U3241) );
  XNOR2_X1 U8439 ( .A(n6846), .B(n6845), .ZN(n6850) );
  INV_X1 U8440 ( .A(n7083), .ZN(n6942) );
  AOI22_X1 U8441 ( .A1(n6942), .A2(n8202), .B1(n8174), .B2(n8211), .ZN(n6849)
         );
  AND2_X1 U8442 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8453) );
  NOR2_X1 U8443 ( .A1(n8200), .A2(n6940), .ZN(n6847) );
  AOI211_X1 U8444 ( .C1(n8175), .C2(n8213), .A(n8453), .B(n6847), .ZN(n6848)
         );
  OAI211_X1 U8445 ( .C1(n6850), .C2(n8204), .A(n6849), .B(n6848), .ZN(P2_U3215) );
  OAI21_X1 U8446 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6856), .A(n6851), .ZN(
        n6854) );
  INV_X1 U8447 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6852) );
  MUX2_X1 U8448 ( .A(n6852), .B(P1_REG1_REG_14__SCAN_IN), .S(n7028), .Z(n6853)
         );
  NAND2_X1 U8449 ( .A1(n6853), .A2(n6854), .ZN(n7035) );
  OAI21_X1 U8450 ( .B1(n6854), .B2(n6853), .A(n7035), .ZN(n6863) );
  XNOR2_X1 U8451 ( .A(n7028), .B(n7029), .ZN(n6858) );
  INV_X1 U8452 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6857) );
  NOR2_X1 U8453 ( .A1(n6857), .A2(n6858), .ZN(n7030) );
  AOI211_X1 U8454 ( .C1(n6858), .C2(n6857), .A(n7030), .B(n9695), .ZN(n6859)
         );
  AOI21_X1 U8455 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9703), .A(n6859), .ZN(
        n6861) );
  NAND2_X1 U8456 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n6860) );
  OAI211_X1 U8457 ( .C1(n7028), .C2(n7161), .A(n6861), .B(n6860), .ZN(n6862)
         );
  AOI21_X1 U8458 ( .B1(n6863), .B2(n9704), .A(n6862), .ZN(n6864) );
  INV_X1 U8459 ( .A(n6864), .ZN(P1_U3255) );
  INV_X1 U8460 ( .A(n6865), .ZN(n6867) );
  OAI222_X1 U8461 ( .A1(n8987), .A2(n8315), .B1(n6866), .B2(n6867), .C1(n8807), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8462 ( .A1(n6868), .A2(n9593), .B1(P1_U3084), .B2(n7383), .C1(
        n9597), .C2(n6867), .ZN(P1_U3334) );
  NAND2_X1 U8463 ( .A1(n6953), .A2(n6869), .ZN(n7903) );
  INV_X1 U8464 ( .A(n6869), .ZN(n9871) );
  NAND2_X1 U8465 ( .A1(n8393), .A2(n9871), .ZN(n7869) );
  NAND2_X1 U8466 ( .A1(n6870), .A2(n9876), .ZN(n6880) );
  NAND3_X1 U8467 ( .A1(n7904), .A2(n6880), .A3(n7868), .ZN(n6881) );
  AND2_X1 U8468 ( .A1(n9820), .A2(n6881), .ZN(n6879) );
  INV_X1 U8469 ( .A(n6871), .ZN(n6872) );
  NAND2_X1 U8470 ( .A1(n6873), .A2(n6872), .ZN(n6875) );
  NAND2_X1 U8471 ( .A1(n6696), .A2(n9858), .ZN(n6874) );
  NAND2_X1 U8472 ( .A1(n6875), .A2(n6874), .ZN(n6948) );
  INV_X1 U8473 ( .A(n9862), .ZN(n6954) );
  NAND2_X1 U8474 ( .A1(n8394), .A2(n9862), .ZN(n7921) );
  NAND2_X1 U8475 ( .A1(n6948), .A2(n6947), .ZN(n6878) );
  NAND2_X1 U8476 ( .A1(n6876), .A2(n9862), .ZN(n6877) );
  NAND2_X1 U8477 ( .A1(n6878), .A2(n6877), .ZN(n7008) );
  NAND2_X1 U8478 ( .A1(n6879), .A2(n7008), .ZN(n6883) );
  NAND2_X1 U8479 ( .A1(n6953), .A2(n9871), .ZN(n9821) );
  NAND2_X1 U8480 ( .A1(n6883), .A2(n6882), .ZN(n6929) );
  NAND2_X1 U8481 ( .A1(n6931), .A2(n9885), .ZN(n7906) );
  NAND2_X1 U8482 ( .A1(n8391), .A2(n6930), .ZN(n7926) );
  NAND2_X1 U8483 ( .A1(n7906), .A2(n7926), .ZN(n6928) );
  INV_X1 U8484 ( .A(n6928), .ZN(n6888) );
  XNOR2_X1 U8485 ( .A(n6929), .B(n6888), .ZN(n9888) );
  NAND2_X1 U8486 ( .A1(n7009), .A2(n9871), .ZN(n9826) );
  OAI21_X1 U8487 ( .B1(n9826), .B2(n9830), .A(n9885), .ZN(n6884) );
  AND3_X1 U8488 ( .A1(n6884), .A2(n9868), .A3(n7001), .ZN(n9884) );
  NAND2_X1 U8489 ( .A1(n6949), .A2(n7920), .ZN(n7012) );
  INV_X1 U8490 ( .A(n9820), .ZN(n7914) );
  NAND2_X1 U8491 ( .A1(n7012), .A2(n7914), .ZN(n6885) );
  NAND2_X1 U8492 ( .A1(n6885), .A2(n7903), .ZN(n9816) );
  INV_X1 U8493 ( .A(n9816), .ZN(n6887) );
  NAND2_X1 U8494 ( .A1(n7904), .A2(n7868), .ZN(n9823) );
  NAND3_X1 U8495 ( .A1(n9818), .A2(n6928), .A3(n7868), .ZN(n6889) );
  NAND3_X1 U8496 ( .A1(n6934), .A2(n8824), .A3(n6889), .ZN(n6891) );
  NAND2_X1 U8497 ( .A1(n6891), .A2(n6890), .ZN(n9883) );
  AOI21_X1 U8498 ( .B1(n9884), .B2(n8807), .A(n9883), .ZN(n6893) );
  MUX2_X1 U8499 ( .A(n6893), .B(n6892), .S(n8846), .Z(n6896) );
  INV_X1 U8500 ( .A(n9827), .ZN(n8844) );
  AOI22_X1 U8501 ( .A1(n9831), .A2(n9885), .B1(n8844), .B2(n6894), .ZN(n6895)
         );
  OAI211_X1 U8502 ( .C1(n9888), .C2(n9825), .A(n6896), .B(n6895), .ZN(P2_U3291) );
  NAND2_X1 U8503 ( .A1(n6898), .A2(n6897), .ZN(n6900) );
  NAND2_X1 U8504 ( .A1(n9095), .A2(n9759), .ZN(n6899) );
  NAND2_X1 U8505 ( .A1(n6900), .A2(n6899), .ZN(n6902) );
  NAND2_X1 U8506 ( .A1(n7045), .A2(n7042), .ZN(n7631) );
  NAND2_X1 U8507 ( .A1(n9127), .A2(n9676), .ZN(n7671) );
  NAND2_X1 U8508 ( .A1(n6902), .A2(n7547), .ZN(n6903) );
  NAND2_X1 U8509 ( .A1(n7044), .A2(n6903), .ZN(n9763) );
  NAND2_X1 U8510 ( .A1(n7770), .A2(n7768), .ZN(n6904) );
  NAND2_X1 U8511 ( .A1(n6904), .A2(n7630), .ZN(n7674) );
  XNOR2_X1 U8512 ( .A(n7674), .B(n7547), .ZN(n6905) );
  OAI22_X1 U8513 ( .A1(n7239), .A2(n9440), .B1(n9095), .B2(n9438), .ZN(n9671)
         );
  AOI21_X1 U8514 ( .B1(n6905), .B2(n9459), .A(n9671), .ZN(n9767) );
  OAI21_X1 U8515 ( .B1(n9763), .B2(n6676), .A(n9767), .ZN(n6906) );
  NAND2_X1 U8516 ( .A1(n6906), .A2(n9460), .ZN(n6912) );
  OAI22_X1 U8517 ( .A1(n9460), .A2(n6312), .B1(n9682), .B2(n9465), .ZN(n6910)
         );
  OR2_X1 U8518 ( .A1(n6907), .A2(n7042), .ZN(n7052) );
  NAND2_X1 U8519 ( .A1(n6907), .A2(n7042), .ZN(n6908) );
  NAND2_X1 U8520 ( .A1(n7052), .A2(n6908), .ZN(n9766) );
  NOR2_X1 U8521 ( .A1(n9766), .A2(n9376), .ZN(n6909) );
  AOI211_X1 U8522 ( .C1(n9374), .C2(n7042), .A(n6910), .B(n6909), .ZN(n6911)
         );
  OAI211_X1 U8523 ( .C1(n9763), .C2(n7250), .A(n6912), .B(n6911), .ZN(P1_U3283) );
  INV_X1 U8524 ( .A(n6913), .ZN(n6914) );
  AOI21_X1 U8525 ( .B1(n6916), .B2(n6915), .A(n6914), .ZN(n9754) );
  XNOR2_X1 U8526 ( .A(n6917), .B(n6916), .ZN(n6921) );
  OAI22_X1 U8527 ( .A1(n6918), .A2(n9438), .B1(n9095), .B2(n9440), .ZN(n6920)
         );
  NOR2_X1 U8528 ( .A1(n9754), .A2(n6676), .ZN(n6919) );
  AOI211_X1 U8529 ( .C1(n6921), .C2(n9459), .A(n6920), .B(n6919), .ZN(n9752)
         );
  MUX2_X1 U8530 ( .A(n6308), .B(n9752), .S(n9460), .Z(n6927) );
  AOI21_X1 U8531 ( .B1(n4315), .B2(n9461), .A(n6922), .ZN(n9750) );
  OAI22_X1 U8532 ( .A1(n9467), .A2(n6924), .B1(n9465), .B2(n6923), .ZN(n6925)
         );
  AOI21_X1 U8533 ( .B1(n9750), .B2(n9429), .A(n6925), .ZN(n6926) );
  OAI211_X1 U8534 ( .C1(n9754), .C2(n7250), .A(n6927), .B(n6926), .ZN(P1_U3285) );
  NAND2_X1 U8535 ( .A1(n6929), .A2(n6928), .ZN(n6993) );
  NAND2_X1 U8536 ( .A1(n6931), .A2(n6930), .ZN(n6992) );
  AND2_X1 U8537 ( .A1(n6992), .A2(n4885), .ZN(n6932) );
  NAND2_X1 U8538 ( .A1(n8213), .A2(n7002), .ZN(n6933) );
  NAND2_X1 U8539 ( .A1(n7084), .A2(n6942), .ZN(n7951) );
  NAND2_X1 U8540 ( .A1(n8212), .A2(n7083), .ZN(n7937) );
  XNOR2_X1 U8541 ( .A(n7081), .B(n7931), .ZN(n7074) );
  INV_X1 U8542 ( .A(n7074), .ZN(n6946) );
  XNOR2_X1 U8543 ( .A(n8213), .B(n7002), .ZN(n7874) );
  NOR2_X1 U8544 ( .A1(n8213), .A2(n9894), .ZN(n7933) );
  NAND2_X1 U8545 ( .A1(n6935), .A2(n7931), .ZN(n7091) );
  OAI211_X1 U8546 ( .C1(n6935), .C2(n7931), .A(n7091), .B(n8824), .ZN(n6937)
         );
  AOI22_X1 U8547 ( .A1(n8819), .A2(n8213), .B1(n8211), .B2(n8821), .ZN(n6936)
         );
  NAND2_X1 U8548 ( .A1(n6937), .A2(n6936), .ZN(n7072) );
  NOR2_X1 U8549 ( .A1(n7000), .A2(n7083), .ZN(n6938) );
  OR2_X1 U8550 ( .A1(n7098), .A2(n6938), .ZN(n7071) );
  NAND2_X1 U8551 ( .A1(n8846), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6939) );
  OAI21_X1 U8552 ( .B1(n9827), .B2(n6940), .A(n6939), .ZN(n6941) );
  AOI21_X1 U8553 ( .B1(n9831), .B2(n6942), .A(n6941), .ZN(n6943) );
  OAI21_X1 U8554 ( .B1(n7071), .B2(n9833), .A(n6943), .ZN(n6944) );
  AOI21_X1 U8555 ( .B1(n7072), .B2(n4316), .A(n6944), .ZN(n6945) );
  OAI21_X1 U8556 ( .B1(n9825), .B2(n6946), .A(n6945), .ZN(P2_U3289) );
  XNOR2_X1 U8557 ( .A(n6947), .B(n6948), .ZN(n9866) );
  INV_X1 U8558 ( .A(n9866), .ZN(n6960) );
  INV_X1 U8559 ( .A(n6949), .ZN(n6950) );
  AOI21_X1 U8560 ( .B1(n6947), .B2(n6951), .A(n6950), .ZN(n6952) );
  OAI222_X1 U8561 ( .A1(n8806), .A2(n6953), .B1(n8804), .B2(n6696), .C1(n9815), 
        .C2(n6952), .ZN(n9864) );
  AND2_X1 U8562 ( .A1(n9854), .A2(n6954), .ZN(n6955) );
  OR2_X1 U8563 ( .A1(n7009), .A2(n6955), .ZN(n9863) );
  OAI22_X1 U8564 ( .A1(n9863), .A2(n9833), .B1(n5690), .B2(n9827), .ZN(n6956)
         );
  AOI21_X1 U8565 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n8846), .A(n6956), .ZN(
        n6957) );
  OAI21_X1 U8566 ( .B1(n9862), .B2(n8848), .A(n6957), .ZN(n6958) );
  AOI21_X1 U8567 ( .B1(n9864), .B2(n4316), .A(n6958), .ZN(n6959) );
  OAI21_X1 U8568 ( .B1(n6960), .B2(n9825), .A(n6959), .ZN(P2_U3294) );
  OAI21_X1 U8569 ( .B1(n6963), .B2(n6962), .A(n6961), .ZN(n6964) );
  NAND2_X1 U8570 ( .A1(n6964), .A2(n9678), .ZN(n6971) );
  NOR2_X1 U8571 ( .A1(n9056), .A2(n9759), .ZN(n6968) );
  AOI21_X1 U8572 ( .B1(n9457), .B2(n9111), .A(n6965), .ZN(n6966) );
  OAI21_X1 U8573 ( .B1(n9096), .B2(n7045), .A(n6966), .ZN(n6967) );
  AOI211_X1 U8574 ( .C1(n6969), .C2(n9100), .A(n6968), .B(n6967), .ZN(n6970)
         );
  NAND2_X1 U8575 ( .A1(n6971), .A2(n6970), .ZN(P1_U3211) );
  XNOR2_X1 U8576 ( .A(n6973), .B(n6972), .ZN(n6977) );
  OAI22_X1 U8577 ( .A1(n8200), .A2(n7096), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8466), .ZN(n6975) );
  OAI22_X1 U8578 ( .A1(n7084), .A2(n8167), .B1(n8166), .B2(n7407), .ZN(n6974)
         );
  AOI211_X1 U8579 ( .C1(n7279), .C2(n8202), .A(n6975), .B(n6974), .ZN(n6976)
         );
  OAI21_X1 U8580 ( .B1(n6977), .B2(n8204), .A(n6976), .ZN(P2_U3223) );
  NOR2_X1 U8581 ( .A1(n6982), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6979) );
  NOR2_X1 U8582 ( .A1(n6979), .A2(n6978), .ZN(n8513) );
  XNOR2_X1 U8583 ( .A(n8513), .B(n8514), .ZN(n6980) );
  NOR2_X1 U8584 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n6980), .ZN(n8515) );
  AOI21_X1 U8585 ( .B1(n6980), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8515), .ZN(
        n6990) );
  XNOR2_X1 U8586 ( .A(n8504), .B(n8505), .ZN(n6983) );
  INV_X1 U8587 ( .A(n6983), .ZN(n6985) );
  NOR2_X1 U8588 ( .A1(n8227), .A2(n6983), .ZN(n8506) );
  INV_X1 U8589 ( .A(n8506), .ZN(n6984) );
  OAI211_X1 U8590 ( .C1(n6985), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9804), .B(
        n6984), .ZN(n6989) );
  INV_X1 U8591 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U8592 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8199) );
  OAI21_X1 U8593 ( .B1(n9602), .B2(n6986), .A(n8199), .ZN(n6987) );
  AOI21_X1 U8594 ( .B1(n9620), .B2(n8514), .A(n6987), .ZN(n6988) );
  OAI211_X1 U8595 ( .C1(n6990), .C2(n9807), .A(n6989), .B(n6988), .ZN(P2_U3260) );
  INV_X1 U8596 ( .A(n6991), .ZN(n7062) );
  OAI222_X1 U8597 ( .A1(n9593), .A2(n8304), .B1(n9597), .B2(n7062), .C1(n7792), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  NAND2_X1 U8598 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  XNOR2_X1 U8599 ( .A(n6994), .B(n7874), .ZN(n9892) );
  XNOR2_X1 U8600 ( .A(n6995), .B(n7874), .ZN(n6996) );
  NAND2_X1 U8601 ( .A1(n6996), .A2(n8824), .ZN(n6998) );
  AOI22_X1 U8602 ( .A1(n8819), .A2(n8391), .B1(n8212), .B2(n8821), .ZN(n6997)
         );
  NAND2_X1 U8603 ( .A1(n6998), .A2(n6997), .ZN(n9896) );
  MUX2_X1 U8604 ( .A(n9896), .B(P2_REG2_REG_6__SCAN_IN), .S(n8846), .Z(n6999)
         );
  INV_X1 U8605 ( .A(n6999), .ZN(n7006) );
  AOI21_X1 U8606 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n9893) );
  OAI22_X1 U8607 ( .A1(n8848), .A2(n9894), .B1(n9827), .B2(n7003), .ZN(n7004)
         );
  AOI21_X1 U8608 ( .B1(n9893), .B2(n8858), .A(n7004), .ZN(n7005) );
  OAI211_X1 U8609 ( .C1(n9825), .C2(n9892), .A(n7006), .B(n7005), .ZN(P2_U3290) );
  INV_X1 U8610 ( .A(n8781), .ZN(n7019) );
  XNOR2_X1 U8611 ( .A(n9820), .B(n7008), .ZN(n9874) );
  OR2_X1 U8612 ( .A1(n7009), .A2(n9871), .ZN(n7010) );
  AND2_X1 U8613 ( .A1(n9826), .A2(n7010), .ZN(n9869) );
  AOI22_X1 U8614 ( .A1(n9869), .A2(n8858), .B1(n8844), .B2(n8399), .ZN(n7011)
         );
  OAI21_X1 U8615 ( .B1(n8848), .B2(n9871), .A(n7011), .ZN(n7018) );
  XNOR2_X1 U8616 ( .A(n7012), .B(n7914), .ZN(n7014) );
  AOI21_X1 U8617 ( .B1(n7014), .B2(n8824), .A(n7013), .ZN(n7016) );
  INV_X1 U8618 ( .A(n7465), .ZN(n7289) );
  NAND2_X1 U8619 ( .A1(n9874), .A2(n7289), .ZN(n7015) );
  NAND2_X1 U8620 ( .A1(n7016), .A2(n7015), .ZN(n9872) );
  MUX2_X1 U8621 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9872), .S(n4316), .Z(n7017)
         );
  AOI211_X1 U8622 ( .C1(n7019), .C2(n9874), .A(n7018), .B(n7017), .ZN(n7020)
         );
  INV_X1 U8623 ( .A(n7020), .ZN(P2_U3293) );
  NAND2_X1 U8624 ( .A1(n6502), .A2(n9849), .ZN(n8080) );
  NAND2_X1 U8625 ( .A1(n7021), .A2(n8080), .ZN(n9852) );
  INV_X1 U8626 ( .A(n9852), .ZN(n7027) );
  AND2_X1 U8627 ( .A1(n6697), .A2(n8821), .ZN(n7022) );
  AOI21_X1 U8628 ( .B1(n9852), .B2(n8824), .A(n7022), .ZN(n9848) );
  INV_X1 U8629 ( .A(n9848), .ZN(n7025) );
  OAI22_X1 U8630 ( .A1(n4316), .A2(n5672), .B1(n5670), .B2(n9827), .ZN(n7024)
         );
  AOI21_X1 U8631 ( .B1(n8848), .B2(n9833), .A(n9849), .ZN(n7023) );
  AOI211_X1 U8632 ( .C1(n4316), .C2(n7025), .A(n7024), .B(n7023), .ZN(n7026)
         );
  OAI21_X1 U8633 ( .B1(n7027), .B2(n9825), .A(n7026), .ZN(P2_U3296) );
  INV_X1 U8634 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7041) );
  INV_X1 U8635 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7033) );
  NOR2_X1 U8636 ( .A1(n7029), .A2(n7028), .ZN(n7031) );
  XOR2_X1 U8637 ( .A(n7153), .B(n7146), .Z(n7032) );
  NOR2_X1 U8638 ( .A1(n7032), .A2(n7033), .ZN(n7147) );
  AOI211_X1 U8639 ( .C1(n7033), .C2(n7032), .A(n9695), .B(n7147), .ZN(n7034)
         );
  INV_X1 U8640 ( .A(n7034), .ZN(n7040) );
  AND2_X1 U8641 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9110) );
  INV_X1 U8642 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9640) );
  OAI21_X1 U8643 ( .B1(n7036), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7035), .ZN(
        n7151) );
  XOR2_X1 U8644 ( .A(n7153), .B(n7151), .Z(n7037) );
  NOR2_X1 U8645 ( .A1(n7037), .A2(n9640), .ZN(n7152) );
  AOI211_X1 U8646 ( .C1(n9640), .C2(n7037), .A(n9173), .B(n7152), .ZN(n7038)
         );
  AOI211_X1 U8647 ( .C1(n9698), .C2(n7153), .A(n9110), .B(n7038), .ZN(n7039)
         );
  OAI211_X1 U8648 ( .C1(n9184), .C2(n7041), .A(n7040), .B(n7039), .ZN(P1_U3256) );
  NAND2_X1 U8649 ( .A1(n9774), .A2(n9126), .ZN(n7672) );
  NAND2_X1 U8650 ( .A1(n7239), .A2(n7127), .ZN(n7624) );
  NAND2_X1 U8651 ( .A1(n7672), .A2(n7624), .ZN(n7548) );
  NAND2_X1 U8652 ( .A1(n9127), .A2(n7042), .ZN(n7043) );
  XOR2_X1 U8653 ( .A(n7548), .B(n7126), .Z(n9780) );
  OAI22_X1 U8654 ( .A1(n7045), .A2(n9438), .B1(n7214), .B2(n9440), .ZN(n7051)
         );
  INV_X1 U8655 ( .A(n7630), .ZN(n7046) );
  NAND2_X1 U8656 ( .A1(n7134), .A2(n7631), .ZN(n7049) );
  INV_X1 U8657 ( .A(n7631), .ZN(n7673) );
  NOR2_X1 U8658 ( .A1(n7548), .A2(n7673), .ZN(n7047) );
  NAND2_X1 U8659 ( .A1(n7134), .A2(n7047), .ZN(n7237) );
  INV_X1 U8660 ( .A(n7237), .ZN(n7048) );
  AOI211_X1 U8661 ( .C1(n7548), .C2(n7049), .A(n9436), .B(n7048), .ZN(n7050)
         );
  AOI211_X1 U8662 ( .C1(n9780), .C2(n7362), .A(n7051), .B(n7050), .ZN(n9777)
         );
  AND2_X1 U8663 ( .A1(n7052), .A2(n7127), .ZN(n7053) );
  OR2_X1 U8664 ( .A1(n7053), .A2(n7246), .ZN(n9776) );
  AOI22_X1 U8665 ( .A1(n9305), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7208), .B2(
        n9444), .ZN(n7055) );
  NAND2_X1 U8666 ( .A1(n9374), .A2(n7127), .ZN(n7054) );
  OAI211_X1 U8667 ( .C1(n9776), .C2(n9376), .A(n7055), .B(n7054), .ZN(n7056)
         );
  AOI21_X1 U8668 ( .B1(n9780), .B2(n7372), .A(n7056), .ZN(n7057) );
  OAI21_X1 U8669 ( .B1(n9777), .B2(n9305), .A(n7057), .ZN(P1_U3282) );
  INV_X1 U8670 ( .A(n7058), .ZN(n7060) );
  OAI222_X1 U8671 ( .A1(n9593), .A2(n7059), .B1(n9597), .B2(n7060), .C1(n7755), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI222_X1 U8672 ( .A1(n8987), .A2(n7061), .B1(P2_U3152), .B2(n7895), .C1(
        n6866), .C2(n7060), .ZN(P2_U3337) );
  OAI222_X1 U8673 ( .A1(n8987), .A2(n7063), .B1(P2_U3152), .B2(n6118), .C1(
        n6866), .C2(n7062), .ZN(P2_U3338) );
  INV_X1 U8674 ( .A(n7064), .ZN(n7069) );
  AND2_X1 U8675 ( .A1(n7065), .A2(n8060), .ZN(n7068) );
  NAND4_X1 U8676 ( .A1(n7069), .A2(n7068), .A3(n7067), .A4(n7066), .ZN(n7077)
         );
  OAI22_X1 U8677 ( .A1(n7071), .A2(n9917), .B1(n7083), .B2(n9915), .ZN(n7073)
         );
  AOI211_X1 U8678 ( .C1(n7074), .C2(n9921), .A(n7073), .B(n7072), .ZN(n7078)
         );
  OR2_X1 U8679 ( .A1(n7078), .A2(n9937), .ZN(n7075) );
  OAI21_X1 U8680 ( .B1(n9939), .B2(n5777), .A(n7075), .ZN(P2_U3527) );
  INV_X1 U8681 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7080) );
  OR2_X1 U8682 ( .A1(n7078), .A2(n9923), .ZN(n7079) );
  OAI21_X1 U8683 ( .B1(n9924), .B2(n7080), .A(n7079), .ZN(P2_U3472) );
  INV_X1 U8684 ( .A(n7931), .ZN(n7082) );
  NAND2_X1 U8685 ( .A1(n7084), .A2(n7083), .ZN(n7085) );
  NAND2_X1 U8686 ( .A1(n7086), .A2(n7085), .ZN(n7089) );
  INV_X1 U8687 ( .A(n7089), .ZN(n7088) );
  INV_X1 U8688 ( .A(n8211), .ZN(n7283) );
  NAND2_X1 U8689 ( .A1(n7089), .A2(n4689), .ZN(n7090) );
  INV_X1 U8690 ( .A(n9904), .ZN(n7104) );
  AOI21_X1 U8691 ( .B1(n7087), .B2(n7092), .A(n7285), .ZN(n7095) );
  AOI22_X1 U8692 ( .A1(n8819), .A2(n8212), .B1(n8210), .B2(n8821), .ZN(n7094)
         );
  NAND2_X1 U8693 ( .A1(n9904), .A2(n7289), .ZN(n7093) );
  OAI211_X1 U8694 ( .C1(n7095), .C2(n9815), .A(n7094), .B(n7093), .ZN(n9902)
         );
  NAND2_X1 U8695 ( .A1(n9902), .A2(n4316), .ZN(n7103) );
  OAI22_X1 U8696 ( .A1(n4316), .A2(n7097), .B1(n7096), .B2(n9827), .ZN(n7101)
         );
  OR2_X1 U8697 ( .A1(n7098), .A2(n9900), .ZN(n7099) );
  NAND2_X1 U8698 ( .A1(n7291), .A2(n7099), .ZN(n9901) );
  NOR2_X1 U8699 ( .A1(n9901), .A2(n9833), .ZN(n7100) );
  AOI211_X1 U8700 ( .C1(n9831), .C2(n7279), .A(n7101), .B(n7100), .ZN(n7102)
         );
  OAI211_X1 U8701 ( .C1(n7104), .C2(n8781), .A(n7103), .B(n7102), .ZN(P2_U3288) );
  XNOR2_X1 U8702 ( .A(n7106), .B(n7105), .ZN(n7111) );
  OAI22_X1 U8703 ( .A1(n8200), .A2(n7411), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7107), .ZN(n7109) );
  OAI22_X1 U8704 ( .A1(n7407), .A2(n8167), .B1(n8166), .B2(n7492), .ZN(n7108)
         );
  AOI211_X1 U8705 ( .C1(n9907), .C2(n8202), .A(n7109), .B(n7108), .ZN(n7110)
         );
  OAI21_X1 U8706 ( .B1(n7111), .B2(n8204), .A(n7110), .ZN(P2_U3219) );
  INV_X1 U8707 ( .A(n7394), .ZN(n7401) );
  OAI21_X1 U8708 ( .B1(n7114), .B2(n7113), .A(n7112), .ZN(n7115) );
  NAND2_X1 U8709 ( .A1(n7115), .A2(n8180), .ZN(n7119) );
  INV_X1 U8710 ( .A(n7116), .ZN(n7292) );
  AND2_X1 U8711 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8478) );
  OAI22_X1 U8712 ( .A1(n7283), .A2(n8167), .B1(n8166), .B2(n7404), .ZN(n7117)
         );
  AOI211_X1 U8713 ( .C1(n7292), .C2(n8137), .A(n8478), .B(n7117), .ZN(n7118)
         );
  OAI211_X1 U8714 ( .C1(n7401), .C2(n8191), .A(n7119), .B(n7118), .ZN(P2_U3233) );
  INV_X1 U8715 ( .A(n7120), .ZN(n7124) );
  OAI222_X1 U8716 ( .A1(n9593), .A2(n7122), .B1(n9597), .B2(n7124), .C1(
        P1_U3084), .C2(n7121), .ZN(P1_U3331) );
  OAI222_X1 U8717 ( .A1(n8987), .A2(n7125), .B1(n6866), .B2(n7124), .C1(n7123), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U8718 ( .A1(n7127), .A2(n9126), .ZN(n7128) );
  NAND2_X1 U8719 ( .A1(n7129), .A2(n7128), .ZN(n7242) );
  OR2_X1 U8720 ( .A1(n9556), .A2(n7214), .ZN(n7675) );
  NAND2_X1 U8721 ( .A1(n9556), .A2(n7214), .ZN(n7625) );
  OR2_X1 U8722 ( .A1(n9556), .A2(n9125), .ZN(n7131) );
  AND2_X1 U8723 ( .A1(n7240), .A2(n7131), .ZN(n7133) );
  NAND2_X1 U8724 ( .A1(n9651), .A2(n9124), .ZN(n7221) );
  OR2_X1 U8725 ( .A1(n9651), .A2(n9124), .ZN(n7130) );
  NAND2_X1 U8726 ( .A1(n7240), .A2(n7223), .ZN(n7132) );
  OAI21_X1 U8727 ( .B1(n7133), .B2(n7550), .A(n7132), .ZN(n9656) );
  AND2_X1 U8728 ( .A1(n7675), .A2(n7672), .ZN(n7646) );
  INV_X1 U8729 ( .A(n7625), .ZN(n7135) );
  AOI21_X1 U8730 ( .B1(n7137), .B2(n7550), .A(n9436), .ZN(n7139) );
  OAI22_X1 U8731 ( .A1(n7214), .A2(n9438), .B1(n7225), .B2(n9440), .ZN(n7138)
         );
  AOI21_X1 U8732 ( .B1(n7139), .B2(n7227), .A(n7138), .ZN(n9654) );
  INV_X1 U8733 ( .A(n9654), .ZN(n7144) );
  INV_X1 U8734 ( .A(n9651), .ZN(n7220) );
  INV_X1 U8735 ( .A(n9556), .ZN(n7267) );
  AND2_X1 U8736 ( .A1(n7246), .A2(n7267), .ZN(n7247) );
  NAND2_X1 U8737 ( .A1(n7247), .A2(n7220), .ZN(n7231) );
  OR2_X1 U8738 ( .A1(n7247), .A2(n7220), .ZN(n7140) );
  AND2_X1 U8739 ( .A1(n7231), .A2(n7140), .ZN(n9652) );
  NAND2_X1 U8740 ( .A1(n9652), .A2(n9429), .ZN(n7142) );
  AOI22_X1 U8741 ( .A1(n9305), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7217), .B2(
        n9444), .ZN(n7141) );
  OAI211_X1 U8742 ( .C1(n7220), .C2(n9467), .A(n7142), .B(n7141), .ZN(n7143)
         );
  AOI21_X1 U8743 ( .B1(n7144), .B2(n9460), .A(n7143), .ZN(n7145) );
  OAI21_X1 U8744 ( .B1(n9656), .B2(n9450), .A(n7145), .ZN(P1_U3280) );
  INV_X1 U8745 ( .A(n7146), .ZN(n7148) );
  NAND2_X1 U8746 ( .A1(n9148), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9156) );
  OAI21_X1 U8747 ( .B1(n9148), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9156), .ZN(
        n7149) );
  NOR2_X1 U8748 ( .A1(n7150), .A2(n7149), .ZN(n9154) );
  AOI211_X1 U8749 ( .C1(n7150), .C2(n7149), .A(n9154), .B(n9695), .ZN(n7164)
         );
  INV_X1 U8750 ( .A(n7151), .ZN(n7154) );
  AOI21_X1 U8751 ( .B1(n7154), .B2(n7153), .A(n7152), .ZN(n7157) );
  INV_X1 U8752 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7155) );
  MUX2_X1 U8753 ( .A(n7155), .B(P1_REG1_REG_16__SCAN_IN), .S(n9148), .Z(n7156)
         );
  NOR2_X1 U8754 ( .A1(n7157), .A2(n7156), .ZN(n9147) );
  AOI211_X1 U8755 ( .C1(n7157), .C2(n7156), .A(n9147), .B(n9173), .ZN(n7158)
         );
  AOI21_X1 U8756 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n9703), .A(n7158), .ZN(
        n7160) );
  NAND2_X1 U8757 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7159) );
  OAI211_X1 U8758 ( .C1(n7162), .C2(n7161), .A(n7160), .B(n7159), .ZN(n7163)
         );
  OR2_X1 U8759 ( .A1(n7164), .A2(n7163), .ZN(P1_U3257) );
  INV_X1 U8760 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9978) );
  NOR2_X1 U8761 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7165) );
  AOI21_X1 U8762 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7165), .ZN(n9946) );
  NOR2_X1 U8763 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7166) );
  AOI21_X1 U8764 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7166), .ZN(n9949) );
  NOR2_X1 U8765 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7167) );
  AOI21_X1 U8766 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7167), .ZN(n9952) );
  NOR2_X1 U8767 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7168) );
  AOI21_X1 U8768 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7168), .ZN(n9955) );
  NOR2_X1 U8769 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7169) );
  AOI21_X1 U8770 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7169), .ZN(n9958) );
  NOR2_X1 U8771 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7175) );
  XNOR2_X1 U8772 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9986) );
  NAND2_X1 U8773 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7173) );
  XOR2_X1 U8774 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9984) );
  NAND2_X1 U8775 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7171) );
  XOR2_X1 U8776 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9981) );
  AOI21_X1 U8777 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9940) );
  INV_X1 U8778 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9601) );
  NAND3_X1 U8779 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9942) );
  OAI21_X1 U8780 ( .B1(n9940), .B2(n9601), .A(n9942), .ZN(n9980) );
  NAND2_X1 U8781 ( .A1(n9981), .A2(n9980), .ZN(n7170) );
  NAND2_X1 U8782 ( .A1(n7171), .A2(n7170), .ZN(n9983) );
  NAND2_X1 U8783 ( .A1(n9984), .A2(n9983), .ZN(n7172) );
  NAND2_X1 U8784 ( .A1(n7173), .A2(n7172), .ZN(n9985) );
  NOR2_X1 U8785 ( .A1(n9986), .A2(n9985), .ZN(n7174) );
  NOR2_X1 U8786 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  NOR2_X1 U8787 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7176), .ZN(n9974) );
  AND2_X1 U8788 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7176), .ZN(n9973) );
  NOR2_X1 U8789 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9973), .ZN(n7177) );
  NOR2_X1 U8790 ( .A1(n9974), .A2(n7177), .ZN(n7178) );
  NAND2_X1 U8791 ( .A1(n7178), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7180) );
  XOR2_X1 U8792 ( .A(n7178), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9972) );
  NAND2_X1 U8793 ( .A1(n9972), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8794 ( .A1(n7180), .A2(n7179), .ZN(n7181) );
  NAND2_X1 U8795 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7181), .ZN(n7183) );
  XOR2_X1 U8796 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7181), .Z(n9968) );
  NAND2_X1 U8797 ( .A1(n9968), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7182) );
  NAND2_X1 U8798 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  NAND2_X1 U8799 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7184), .ZN(n7186) );
  XOR2_X1 U8800 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7184), .Z(n9982) );
  NAND2_X1 U8801 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9982), .ZN(n7185) );
  NAND2_X1 U8802 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  AND2_X1 U8803 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7187), .ZN(n7188) );
  XNOR2_X1 U8804 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7187), .ZN(n9971) );
  INV_X1 U8805 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U8806 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  NOR2_X1 U8807 ( .A1(n7188), .A2(n9969), .ZN(n9967) );
  NAND2_X1 U8808 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7189) );
  OAI21_X1 U8809 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7189), .ZN(n9966) );
  NOR2_X1 U8810 ( .A1(n9967), .A2(n9966), .ZN(n9965) );
  AOI21_X1 U8811 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9965), .ZN(n9964) );
  NAND2_X1 U8812 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7190) );
  OAI21_X1 U8813 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7190), .ZN(n9963) );
  NOR2_X1 U8814 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  AOI21_X1 U8815 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9962), .ZN(n9961) );
  NOR2_X1 U8816 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7191) );
  AOI21_X1 U8817 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7191), .ZN(n9960) );
  NAND2_X1 U8818 ( .A1(n9961), .A2(n9960), .ZN(n9959) );
  OAI21_X1 U8819 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9959), .ZN(n9957) );
  NAND2_X1 U8820 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  OAI21_X1 U8821 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9956), .ZN(n9954) );
  NAND2_X1 U8822 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  OAI21_X1 U8823 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9953), .ZN(n9951) );
  NAND2_X1 U8824 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  OAI21_X1 U8825 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9950), .ZN(n9948) );
  NAND2_X1 U8826 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  OAI21_X1 U8827 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9947), .ZN(n9945) );
  NAND2_X1 U8828 ( .A1(n9946), .A2(n9945), .ZN(n9944) );
  NOR2_X1 U8829 ( .A1(n9978), .A2(n9977), .ZN(n7192) );
  NAND2_X1 U8830 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  OAI21_X1 U8831 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7192), .A(n9976), .ZN(
        n7194) );
  XNOR2_X1 U8832 ( .A(n4581), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7193) );
  XNOR2_X1 U8833 ( .A(n7194), .B(n7193), .ZN(ADD_1071_U4) );
  INV_X1 U8834 ( .A(n7197), .ZN(n7195) );
  NAND2_X1 U8835 ( .A1(n7196), .A2(n7195), .ZN(n9672) );
  NAND2_X1 U8836 ( .A1(n9672), .A2(n9674), .ZN(n7202) );
  INV_X1 U8837 ( .A(n7196), .ZN(n7198) );
  NAND2_X1 U8838 ( .A1(n7198), .A2(n7197), .ZN(n9673) );
  XNOR2_X1 U8839 ( .A(n7200), .B(n7199), .ZN(n7201) );
  NAND3_X1 U8840 ( .A1(n7202), .A2(n9673), .A3(n7201), .ZN(n7260) );
  INV_X1 U8841 ( .A(n7260), .ZN(n7204) );
  AOI21_X1 U8842 ( .B1(n7202), .B2(n9673), .A(n7201), .ZN(n7203) );
  OAI21_X1 U8843 ( .B1(n7204), .B2(n7203), .A(n9678), .ZN(n7210) );
  NOR2_X1 U8844 ( .A1(n9056), .A2(n9774), .ZN(n7207) );
  AND2_X1 U8845 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9137) );
  AOI21_X1 U8846 ( .B1(n9127), .B2(n9111), .A(n9137), .ZN(n7205) );
  OAI21_X1 U8847 ( .B1(n9096), .B2(n7214), .A(n7205), .ZN(n7206) );
  AOI211_X1 U8848 ( .C1(n7208), .C2(n9100), .A(n7207), .B(n7206), .ZN(n7209)
         );
  NAND2_X1 U8849 ( .A1(n7210), .A2(n7209), .ZN(P1_U3229) );
  OAI211_X1 U8850 ( .C1(n7213), .C2(n7212), .A(n7211), .B(n9678), .ZN(n7219)
         );
  NOR2_X1 U8851 ( .A1(n9096), .A2(n7225), .ZN(n7216) );
  OAI22_X1 U8852 ( .A1(n6830), .A2(n7214), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6340), .ZN(n7215) );
  AOI211_X1 U8853 ( .C1(n7217), .C2(n9100), .A(n7216), .B(n7215), .ZN(n7218)
         );
  OAI211_X1 U8854 ( .C1(n7220), .C2(n9056), .A(n7219), .B(n7218), .ZN(P1_U3234) );
  INV_X1 U8855 ( .A(n7221), .ZN(n7224) );
  OR2_X1 U8856 ( .A1(n7552), .A2(n7224), .ZN(n7222) );
  OR2_X1 U8857 ( .A1(n7224), .A2(n7223), .ZN(n7309) );
  AND2_X1 U8858 ( .A1(n7312), .A2(n7309), .ZN(n7226) );
  OR2_X1 U8859 ( .A1(n7375), .A2(n7225), .ZN(n7679) );
  NAND2_X1 U8860 ( .A1(n7375), .A2(n7225), .ZN(n7683) );
  NAND2_X1 U8861 ( .A1(n7679), .A2(n7683), .ZN(n7310) );
  XNOR2_X1 U8862 ( .A(n7226), .B(n7553), .ZN(n7379) );
  INV_X1 U8863 ( .A(n9124), .ZN(n7627) );
  OR2_X1 U8864 ( .A1(n9651), .A2(n7627), .ZN(n7316) );
  XNOR2_X1 U8865 ( .A(n7315), .B(n7553), .ZN(n7229) );
  AOI22_X1 U8866 ( .A1(n9454), .A2(n9124), .B1(n9122), .B2(n9456), .ZN(n7228)
         );
  OAI21_X1 U8867 ( .B1(n7229), .B2(n9436), .A(n7228), .ZN(n7230) );
  AOI21_X1 U8868 ( .B1(n7379), .B2(n7362), .A(n7230), .ZN(n7381) );
  AOI21_X1 U8869 ( .B1(n7231), .B2(n7375), .A(n9775), .ZN(n7232) );
  OR2_X1 U8870 ( .A1(n7231), .A2(n7375), .ZN(n7366) );
  NAND2_X1 U8871 ( .A1(n7232), .A2(n7366), .ZN(n7376) );
  AOI22_X1 U8872 ( .A1(n9305), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7302), .B2(
        n9444), .ZN(n7234) );
  NAND2_X1 U8873 ( .A1(n7375), .A2(n9374), .ZN(n7233) );
  OAI211_X1 U8874 ( .C1(n7376), .C2(n7329), .A(n7234), .B(n7233), .ZN(n7235)
         );
  AOI21_X1 U8875 ( .B1(n7379), .B2(n7372), .A(n7235), .ZN(n7236) );
  OAI21_X1 U8876 ( .B1(n7381), .B2(n9305), .A(n7236), .ZN(P1_U3279) );
  NAND2_X1 U8877 ( .A1(n7237), .A2(n7672), .ZN(n7238) );
  XOR2_X1 U8878 ( .A(n7552), .B(n7238), .Z(n7245) );
  OAI22_X1 U8879 ( .A1(n7627), .A2(n9440), .B1(n7239), .B2(n9438), .ZN(n7244)
         );
  INV_X1 U8880 ( .A(n7240), .ZN(n7241) );
  AOI21_X1 U8881 ( .B1(n7552), .B2(n7242), .A(n7241), .ZN(n9559) );
  NOR2_X1 U8882 ( .A1(n9559), .A2(n6676), .ZN(n7243) );
  AOI211_X1 U8883 ( .C1(n9459), .C2(n7245), .A(n7244), .B(n7243), .ZN(n9558)
         );
  INV_X1 U8884 ( .A(n7246), .ZN(n7248) );
  AOI211_X1 U8885 ( .C1(n9556), .C2(n7248), .A(n9775), .B(n7247), .ZN(n9555)
         );
  AOI22_X1 U8886 ( .A1(n9305), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7270), .B2(
        n9444), .ZN(n7249) );
  OAI21_X1 U8887 ( .B1(n7267), .B2(n9467), .A(n7249), .ZN(n7252) );
  NOR2_X1 U8888 ( .A1(n9559), .A2(n7250), .ZN(n7251) );
  AOI211_X1 U8889 ( .C1(n9555), .C2(n9469), .A(n7252), .B(n7251), .ZN(n7253)
         );
  OAI21_X1 U8890 ( .B1(n9558), .B2(n9305), .A(n7253), .ZN(P1_U3281) );
  NAND2_X1 U8891 ( .A1(n7256), .A2(n9588), .ZN(n7254) );
  OAI211_X1 U8892 ( .C1(n7255), .C2(n9593), .A(n7254), .B(n7798), .ZN(P1_U3330) );
  NAND2_X1 U8893 ( .A1(n7256), .A2(n8979), .ZN(n7257) );
  OAI211_X1 U8894 ( .C1(n7258), .C2(n8987), .A(n7257), .B(n8065), .ZN(P2_U3335) );
  NAND2_X1 U8895 ( .A1(n7260), .A2(n7259), .ZN(n7264) );
  NAND2_X1 U8896 ( .A1(n7262), .A2(n7261), .ZN(n7263) );
  XNOR2_X1 U8897 ( .A(n7264), .B(n7263), .ZN(n7272) );
  AOI21_X1 U8898 ( .B1(n9126), .B2(n9111), .A(n7265), .ZN(n7266) );
  OAI21_X1 U8899 ( .B1(n9096), .B2(n7627), .A(n7266), .ZN(n7269) );
  NOR2_X1 U8900 ( .A1(n7267), .A2(n9056), .ZN(n7268) );
  AOI211_X1 U8901 ( .C1(n7270), .C2(n9100), .A(n7269), .B(n7268), .ZN(n7271)
         );
  OAI21_X1 U8902 ( .B1(n7272), .B2(n9117), .A(n7271), .ZN(P1_U3215) );
  XNOR2_X1 U8903 ( .A(n7274), .B(n7273), .ZN(n7278) );
  OAI22_X1 U8904 ( .A1(n8200), .A2(n7482), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5858), .ZN(n7276) );
  INV_X1 U8905 ( .A(n8207), .ZN(n7466) );
  OAI22_X1 U8906 ( .A1(n7404), .A2(n8167), .B1(n8166), .B2(n7466), .ZN(n7275)
         );
  AOI211_X1 U8907 ( .C1(n8948), .C2(n8202), .A(n7276), .B(n7275), .ZN(n7277)
         );
  OAI21_X1 U8908 ( .B1(n7278), .B2(n8204), .A(n7277), .ZN(P2_U3238) );
  NAND2_X1 U8909 ( .A1(n8211), .A2(n7279), .ZN(n7280) );
  NAND2_X1 U8910 ( .A1(n7401), .A2(n8210), .ZN(n7941) );
  NAND2_X1 U8911 ( .A1(n7407), .A2(n7394), .ZN(n7946) );
  NAND2_X1 U8912 ( .A1(n7941), .A2(n7946), .ZN(n7876) );
  OAI21_X1 U8913 ( .B1(n7282), .B2(n7876), .A(n7403), .ZN(n7294) );
  OAI22_X1 U8914 ( .A1(n7283), .A2(n8804), .B1(n7404), .B2(n8806), .ZN(n7288)
         );
  XOR2_X1 U8915 ( .A(n7876), .B(n4392), .Z(n7286) );
  NOR2_X1 U8916 ( .A1(n7286), .A2(n9815), .ZN(n7287) );
  AOI211_X1 U8917 ( .C1(n7289), .C2(n7294), .A(n7288), .B(n7287), .ZN(n7397)
         );
  INV_X1 U8918 ( .A(n7413), .ZN(n7290) );
  AOI21_X1 U8919 ( .B1(n7394), .B2(n7291), .A(n7290), .ZN(n7395) );
  AOI22_X1 U8920 ( .A1(n8846), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7292), .B2(
        n8844), .ZN(n7293) );
  OAI21_X1 U8921 ( .B1(n8848), .B2(n7401), .A(n7293), .ZN(n7296) );
  INV_X1 U8922 ( .A(n7294), .ZN(n7398) );
  NOR2_X1 U8923 ( .A1(n7398), .A2(n8781), .ZN(n7295) );
  AOI211_X1 U8924 ( .C1(n7395), .C2(n8858), .A(n7296), .B(n7295), .ZN(n7297)
         );
  OAI21_X1 U8925 ( .B1(n7397), .B2(n9837), .A(n7297), .ZN(P2_U3287) );
  XOR2_X1 U8926 ( .A(n7299), .B(n7298), .Z(n7300) );
  XNOR2_X1 U8927 ( .A(n7301), .B(n7300), .ZN(n7308) );
  INV_X1 U8928 ( .A(n9122), .ZN(n7319) );
  NAND2_X1 U8929 ( .A1(n9100), .A2(n7302), .ZN(n7305) );
  AOI21_X1 U8930 ( .B1(n9111), .B2(n9124), .A(n7303), .ZN(n7304) );
  OAI211_X1 U8931 ( .C1(n7319), .C2(n9096), .A(n7305), .B(n7304), .ZN(n7306)
         );
  AOI21_X1 U8932 ( .B1(n9115), .B2(n7375), .A(n7306), .ZN(n7307) );
  OAI21_X1 U8933 ( .B1(n7308), .B2(n9117), .A(n7307), .ZN(P1_U3222) );
  AND2_X1 U8934 ( .A1(n7310), .A2(n7309), .ZN(n7311) );
  NAND2_X1 U8935 ( .A1(n7421), .A2(n9122), .ZN(n7313) );
  NAND2_X1 U8936 ( .A1(n7375), .A2(n9123), .ZN(n7359) );
  OR2_X1 U8937 ( .A1(n7421), .A2(n9122), .ZN(n7314) );
  OR2_X1 U8938 ( .A1(n7333), .A2(n7430), .ZN(n7642) );
  NAND2_X1 U8939 ( .A1(n7333), .A2(n7430), .ZN(n7623) );
  NAND2_X1 U8940 ( .A1(n7642), .A2(n7623), .ZN(n7335) );
  XNOR2_X1 U8941 ( .A(n7336), .B(n7335), .ZN(n9645) );
  INV_X1 U8942 ( .A(n9645), .ZN(n7332) );
  NAND2_X1 U8943 ( .A1(n7679), .A2(n7316), .ZN(n7317) );
  NAND2_X1 U8944 ( .A1(n7317), .A2(n7683), .ZN(n7644) );
  OR2_X1 U8945 ( .A1(n7421), .A2(n7319), .ZN(n7641) );
  NAND2_X1 U8946 ( .A1(n7421), .A2(n7319), .ZN(n7622) );
  NAND2_X1 U8947 ( .A1(n7641), .A2(n7622), .ZN(n7554) );
  OR2_X2 U8948 ( .A1(n7358), .A2(n7554), .ZN(n7356) );
  INV_X1 U8949 ( .A(n7622), .ZN(n7320) );
  NOR2_X1 U8950 ( .A1(n7335), .A2(n7320), .ZN(n7321) );
  NAND2_X1 U8951 ( .A1(n7337), .A2(n9459), .ZN(n7325) );
  INV_X1 U8952 ( .A(n7335), .ZN(n7557) );
  AOI21_X1 U8953 ( .B1(n7356), .B2(n7622), .A(n7557), .ZN(n7324) );
  NAND2_X1 U8954 ( .A1(n9196), .A2(n9456), .ZN(n7323) );
  NAND2_X1 U8955 ( .A1(n9122), .A2(n9454), .ZN(n7322) );
  AND2_X1 U8956 ( .A1(n7323), .A2(n7322), .ZN(n9003) );
  OAI21_X1 U8957 ( .B1(n7325), .B2(n7324), .A(n9003), .ZN(n9644) );
  INV_X1 U8958 ( .A(n7343), .ZN(n7326) );
  OAI211_X1 U8959 ( .C1(n9642), .C2(n7367), .A(n7326), .B(n9749), .ZN(n9641)
         );
  AOI22_X1 U8960 ( .A1(n9305), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9006), .B2(
        n9444), .ZN(n7328) );
  NAND2_X1 U8961 ( .A1(n7333), .A2(n9374), .ZN(n7327) );
  OAI211_X1 U8962 ( .C1(n9641), .C2(n7329), .A(n7328), .B(n7327), .ZN(n7330)
         );
  AOI21_X1 U8963 ( .B1(n9644), .B2(n9460), .A(n7330), .ZN(n7331) );
  OAI21_X1 U8964 ( .B1(n7332), .B2(n9450), .A(n7331), .ZN(P1_U3277) );
  INV_X1 U8965 ( .A(n7430), .ZN(n9121) );
  NOR2_X1 U8966 ( .A1(n7333), .A2(n9121), .ZN(n7334) );
  AND2_X1 U8967 ( .A1(n9197), .A2(n9437), .ZN(n9212) );
  INV_X1 U8968 ( .A(n9212), .ZN(n7650) );
  OR2_X1 U8969 ( .A1(n9197), .A2(n9437), .ZN(n9213) );
  XNOR2_X1 U8970 ( .A(n9198), .B(n7690), .ZN(n9637) );
  XNOR2_X1 U8971 ( .A(n9214), .B(n7690), .ZN(n7338) );
  NAND2_X1 U8972 ( .A1(n7338), .A2(n9459), .ZN(n7341) );
  OAI22_X1 U8973 ( .A1(n7430), .A2(n9438), .B1(n9108), .B2(n9440), .ZN(n7339)
         );
  INV_X1 U8974 ( .A(n7339), .ZN(n7340) );
  NAND2_X1 U8975 ( .A1(n7341), .A2(n7340), .ZN(n7342) );
  AOI21_X1 U8976 ( .B1(n9637), .B2(n7362), .A(n7342), .ZN(n9639) );
  OR2_X1 U8977 ( .A1(n7343), .A2(n9634), .ZN(n7344) );
  NAND2_X1 U8978 ( .A1(n9443), .A2(n7344), .ZN(n9635) );
  AOI22_X1 U8979 ( .A1(n9305), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7345), .B2(
        n9444), .ZN(n7347) );
  NAND2_X1 U8980 ( .A1(n9197), .A2(n9374), .ZN(n7346) );
  OAI211_X1 U8981 ( .C1(n9635), .C2(n9376), .A(n7347), .B(n7346), .ZN(n7348)
         );
  AOI21_X1 U8982 ( .B1(n9637), .B2(n7372), .A(n7348), .ZN(n7349) );
  OAI21_X1 U8983 ( .B1(n9639), .B2(n9305), .A(n7349), .ZN(P1_U3276) );
  INV_X1 U8984 ( .A(n7350), .ZN(n7354) );
  OAI222_X1 U8985 ( .A1(P1_U3084), .A2(n7352), .B1(n9597), .B2(n7354), .C1(
        n7351), .C2(n9593), .ZN(P1_U3329) );
  OAI222_X1 U8986 ( .A1(P2_U3152), .A2(n7355), .B1(n6866), .B2(n7354), .C1(
        n7353), .C2(n8987), .ZN(P2_U3334) );
  INV_X1 U8987 ( .A(n7356), .ZN(n7357) );
  AOI21_X1 U8988 ( .B1(n7358), .B2(n7554), .A(n7357), .ZN(n7365) );
  NAND2_X1 U8989 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  XOR2_X1 U8990 ( .A(n7554), .B(n7361), .Z(n9650) );
  NAND2_X1 U8991 ( .A1(n9650), .A2(n7362), .ZN(n7364) );
  AOI22_X1 U8992 ( .A1(n9454), .A2(n9123), .B1(n9121), .B2(n9456), .ZN(n7363)
         );
  OAI211_X1 U8993 ( .C1(n9436), .C2(n7365), .A(n7364), .B(n7363), .ZN(n9648)
         );
  INV_X1 U8994 ( .A(n9648), .ZN(n7374) );
  AND2_X1 U8995 ( .A1(n7366), .A2(n7421), .ZN(n7368) );
  OR2_X1 U8996 ( .A1(n7368), .A2(n7367), .ZN(n9647) );
  AOI22_X1 U8997 ( .A1(n9305), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7432), .B2(
        n9444), .ZN(n7370) );
  NAND2_X1 U8998 ( .A1(n7421), .A2(n9374), .ZN(n7369) );
  OAI211_X1 U8999 ( .C1(n9647), .C2(n9376), .A(n7370), .B(n7369), .ZN(n7371)
         );
  AOI21_X1 U9000 ( .B1(n9650), .B2(n7372), .A(n7371), .ZN(n7373) );
  OAI21_X1 U9001 ( .B1(n7374), .B2(n9305), .A(n7373), .ZN(P1_U3278) );
  INV_X1 U9002 ( .A(n7375), .ZN(n7377) );
  OAI21_X1 U9003 ( .B1(n7377), .B2(n9773), .A(n7376), .ZN(n7378) );
  AOI21_X1 U9004 ( .B1(n7379), .B2(n9781), .A(n7378), .ZN(n7380) );
  AND2_X1 U9005 ( .A1(n7381), .A2(n7380), .ZN(n7391) );
  OAI21_X1 U9006 ( .B1(n9775), .B2(n7383), .A(n7382), .ZN(n7384) );
  INV_X1 U9007 ( .A(n7384), .ZN(n7385) );
  MUX2_X1 U9008 ( .A(n6464), .B(n7391), .S(n9802), .Z(n7387) );
  INV_X1 U9009 ( .A(n7387), .ZN(P1_U3535) );
  INV_X1 U9010 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7392) );
  MUX2_X1 U9011 ( .A(n7392), .B(n7391), .S(n9784), .Z(n7393) );
  INV_X1 U9012 ( .A(n7393), .ZN(P1_U3490) );
  INV_X1 U9013 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7400) );
  AOI22_X1 U9014 ( .A1(n7395), .A2(n9868), .B1(n9886), .B2(n7394), .ZN(n7396)
         );
  OAI211_X1 U9015 ( .C1(n7398), .C2(n9867), .A(n7397), .B(n7396), .ZN(n7419)
         );
  NAND2_X1 U9016 ( .A1(n7419), .A2(n9924), .ZN(n7399) );
  OAI21_X1 U9017 ( .B1(n9924), .B2(n7400), .A(n7399), .ZN(P2_U3478) );
  NAND2_X1 U9018 ( .A1(n7401), .A2(n7407), .ZN(n7402) );
  NAND2_X1 U9019 ( .A1(n9907), .A2(n7404), .ZN(n7948) );
  NAND2_X1 U9020 ( .A1(n7954), .A2(n7948), .ZN(n7942) );
  NAND2_X1 U9021 ( .A1(n7405), .A2(n7942), .ZN(n7461) );
  OAI21_X1 U9022 ( .B1(n7405), .B2(n7942), .A(n7461), .ZN(n9906) );
  AOI211_X1 U9023 ( .C1(n7942), .C2(n7406), .A(n9815), .B(n7457), .ZN(n7409)
         );
  OAI22_X1 U9024 ( .A1(n7407), .A2(n8804), .B1(n7492), .B2(n8806), .ZN(n7408)
         );
  NOR2_X1 U9025 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  OAI21_X1 U9026 ( .B1(n7465), .B2(n9906), .A(n7410), .ZN(n9910) );
  NAND2_X1 U9027 ( .A1(n9910), .A2(n4316), .ZN(n7418) );
  OAI22_X1 U9028 ( .A1(n4316), .A2(n7412), .B1(n7411), .B2(n9827), .ZN(n7416)
         );
  NAND2_X1 U9029 ( .A1(n7413), .A2(n9907), .ZN(n7414) );
  NAND2_X1 U9030 ( .A1(n7479), .A2(n7414), .ZN(n9909) );
  NOR2_X1 U9031 ( .A1(n9909), .A2(n9833), .ZN(n7415) );
  AOI211_X1 U9032 ( .C1(n9831), .C2(n9907), .A(n7416), .B(n7415), .ZN(n7417)
         );
  OAI211_X1 U9033 ( .C1(n9906), .C2(n8781), .A(n7418), .B(n7417), .ZN(P2_U3286) );
  NAND2_X1 U9034 ( .A1(n7419), .A2(n9939), .ZN(n7420) );
  OAI21_X1 U9035 ( .B1(n9939), .B2(n5810), .A(n7420), .ZN(P2_U3529) );
  INV_X1 U9036 ( .A(n7421), .ZN(n9646) );
  NOR2_X1 U9037 ( .A1(n7422), .A2(n4430), .ZN(n7427) );
  AOI21_X1 U9038 ( .B1(n7425), .B2(n7424), .A(n7423), .ZN(n7426) );
  OAI21_X1 U9039 ( .B1(n7427), .B2(n7426), .A(n9678), .ZN(n7434) );
  AOI21_X1 U9040 ( .B1(n9123), .B2(n9111), .A(n7428), .ZN(n7429) );
  OAI21_X1 U9041 ( .B1(n9096), .B2(n7430), .A(n7429), .ZN(n7431) );
  AOI21_X1 U9042 ( .B1(n7432), .B2(n9100), .A(n7431), .ZN(n7433) );
  OAI211_X1 U9043 ( .C1(n9646), .C2(n9056), .A(n7434), .B(n7433), .ZN(P1_U3232) );
  INV_X1 U9044 ( .A(n7435), .ZN(n7436) );
  AOI21_X1 U9045 ( .B1(n7438), .B2(n7437), .A(n7436), .ZN(n7442) );
  AOI22_X1 U9046 ( .A1(n8175), .A2(n8208), .B1(n8174), .B2(n8206), .ZN(n7439)
         );
  NAND2_X1 U9047 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8492) );
  OAI211_X1 U9048 ( .C1(n7493), .C2(n8200), .A(n7439), .B(n8492), .ZN(n7440)
         );
  AOI21_X1 U9049 ( .B1(n7498), .B2(n8202), .A(n7440), .ZN(n7441) );
  OAI21_X1 U9050 ( .B1(n7442), .B2(n8204), .A(n7441), .ZN(P2_U3226) );
  XNOR2_X1 U9051 ( .A(n7444), .B(n7443), .ZN(n7449) );
  AOI22_X1 U9052 ( .A1(n8175), .A2(n8207), .B1(n8174), .B2(n8580), .ZN(n7446)
         );
  OAI211_X1 U9053 ( .C1(n8200), .C2(n7470), .A(n7446), .B(n7445), .ZN(n7447)
         );
  AOI21_X1 U9054 ( .B1(n8943), .B2(n8202), .A(n7447), .ZN(n7448) );
  OAI21_X1 U9055 ( .B1(n7449), .B2(n8204), .A(n7448), .ZN(P2_U3236) );
  INV_X1 U9056 ( .A(n7450), .ZN(n7454) );
  OAI222_X1 U9057 ( .A1(n8987), .A2(n7452), .B1(n6866), .B2(n7454), .C1(
        P2_U3152), .C2(n7451), .ZN(P2_U3333) );
  OAI222_X1 U9058 ( .A1(n9593), .A2(n7455), .B1(n9597), .B2(n7454), .C1(
        P1_U3084), .C2(n7453), .ZN(P1_U3328) );
  OR2_X1 U9059 ( .A1(n8943), .A2(n7506), .ZN(n7971) );
  NAND2_X1 U9060 ( .A1(n8943), .A2(n7506), .ZN(n7970) );
  INV_X1 U9061 ( .A(n7954), .ZN(n7456) );
  OR2_X1 U9062 ( .A1(n8948), .A2(n7492), .ZN(n7958) );
  NAND2_X1 U9063 ( .A1(n8948), .A2(n7492), .ZN(n7949) );
  NAND2_X1 U9064 ( .A1(n7958), .A2(n7949), .ZN(n7877) );
  NAND2_X1 U9065 ( .A1(n7477), .A2(n4527), .ZN(n7489) );
  NAND2_X1 U9066 ( .A1(n7498), .A2(n7466), .ZN(n7965) );
  AND2_X1 U9067 ( .A1(n7965), .A2(n7949), .ZN(n7959) );
  OR2_X1 U9068 ( .A1(n7498), .A2(n7466), .ZN(n7964) );
  INV_X1 U9069 ( .A(n7964), .ZN(n7458) );
  AOI21_X1 U9070 ( .B1(n7489), .B2(n7959), .A(n7458), .ZN(n7459) );
  OAI21_X1 U9071 ( .B1(n7968), .B2(n7459), .A(n7509), .ZN(n7469) );
  NAND2_X1 U9072 ( .A1(n9907), .A2(n8209), .ZN(n7460) );
  NAND2_X1 U9073 ( .A1(n7461), .A2(n7460), .ZN(n7476) );
  NAND2_X1 U9074 ( .A1(n8948), .A2(n8208), .ZN(n7462) );
  NAND2_X1 U9075 ( .A1(n7463), .A2(n7968), .ZN(n7464) );
  NAND2_X1 U9076 ( .A1(n7505), .A2(n7464), .ZN(n8947) );
  NOR2_X1 U9077 ( .A1(n8947), .A2(n7465), .ZN(n7468) );
  INV_X1 U9078 ( .A(n8580), .ZN(n7508) );
  OAI22_X1 U9079 ( .A1(n7466), .A2(n8804), .B1(n7508), .B2(n8806), .ZN(n7467)
         );
  AOI211_X1 U9080 ( .C1(n7469), .C2(n8824), .A(n7468), .B(n7467), .ZN(n8946)
         );
  INV_X1 U9081 ( .A(n7498), .ZN(n9916) );
  AOI21_X1 U9082 ( .B1(n8943), .B2(n7494), .A(n4391), .ZN(n8944) );
  INV_X1 U9083 ( .A(n8943), .ZN(n7507) );
  INV_X1 U9084 ( .A(n7470), .ZN(n7471) );
  AOI22_X1 U9085 ( .A1(n8846), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7471), .B2(
        n8844), .ZN(n7472) );
  OAI21_X1 U9086 ( .B1(n7507), .B2(n8848), .A(n7472), .ZN(n7474) );
  NOR2_X1 U9087 ( .A1(n8947), .A2(n8781), .ZN(n7473) );
  AOI211_X1 U9088 ( .C1(n8944), .C2(n8858), .A(n7474), .B(n7473), .ZN(n7475)
         );
  OAI21_X1 U9089 ( .B1(n8946), .B2(n9837), .A(n7475), .ZN(P2_U3283) );
  XNOR2_X1 U9090 ( .A(n7476), .B(n7877), .ZN(n8954) );
  OAI21_X1 U9091 ( .B1(n4527), .B2(n7477), .A(n7489), .ZN(n7478) );
  AOI222_X1 U9092 ( .A1(n8824), .A2(n7478), .B1(n8207), .B2(n8821), .C1(n8209), 
        .C2(n8819), .ZN(n8953) );
  INV_X1 U9093 ( .A(n8953), .ZN(n7486) );
  AND2_X1 U9094 ( .A1(n7479), .A2(n8948), .ZN(n7480) );
  OR2_X1 U9095 ( .A1(n7480), .A2(n7495), .ZN(n8950) );
  NAND2_X1 U9096 ( .A1(n8846), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7481) );
  OAI21_X1 U9097 ( .B1(n9827), .B2(n7482), .A(n7481), .ZN(n7483) );
  AOI21_X1 U9098 ( .B1(n9831), .B2(n8948), .A(n7483), .ZN(n7484) );
  OAI21_X1 U9099 ( .B1(n8950), .B2(n9833), .A(n7484), .ZN(n7485) );
  AOI21_X1 U9100 ( .B1(n7486), .B2(n4316), .A(n7485), .ZN(n7487) );
  OAI21_X1 U9101 ( .B1(n9825), .B2(n8954), .A(n7487), .ZN(P2_U3285) );
  XNOR2_X1 U9102 ( .A(n7488), .B(n7880), .ZN(n9922) );
  INV_X1 U9103 ( .A(n9922), .ZN(n7501) );
  NAND2_X1 U9104 ( .A1(n7489), .A2(n7949), .ZN(n7490) );
  XOR2_X1 U9105 ( .A(n7880), .B(n7490), .Z(n7491) );
  OAI222_X1 U9106 ( .A1(n8806), .A2(n7506), .B1(n8804), .B2(n7492), .C1(n7491), 
        .C2(n9815), .ZN(n9919) );
  NAND2_X1 U9107 ( .A1(n9919), .A2(n4316), .ZN(n7500) );
  OAI22_X1 U9108 ( .A1(n4316), .A2(n8488), .B1(n7493), .B2(n9827), .ZN(n7497)
         );
  OAI21_X1 U9109 ( .B1(n7495), .B2(n9916), .A(n7494), .ZN(n9918) );
  NOR2_X1 U9110 ( .A1(n9918), .A2(n9833), .ZN(n7496) );
  AOI211_X1 U9111 ( .C1(n9831), .C2(n7498), .A(n7497), .B(n7496), .ZN(n7499)
         );
  OAI211_X1 U9112 ( .C1(n7501), .C2(n9825), .A(n7500), .B(n7499), .ZN(P2_U3284) );
  INV_X1 U9113 ( .A(n7502), .ZN(n7805) );
  OAI222_X1 U9114 ( .A1(P2_U3152), .A2(n7504), .B1(n6866), .B2(n7805), .C1(
        n7503), .C2(n8987), .ZN(P2_U3332) );
  NAND2_X1 U9115 ( .A1(n8581), .A2(n7508), .ZN(n7974) );
  XNOR2_X1 U9116 ( .A(n8583), .B(n8582), .ZN(n9631) );
  INV_X1 U9117 ( .A(n9631), .ZN(n7520) );
  NAND2_X1 U9118 ( .A1(n8852), .A2(n8824), .ZN(n7514) );
  AOI21_X1 U9119 ( .B1(n7509), .B2(n7970), .A(n8582), .ZN(n7513) );
  NAND2_X1 U9120 ( .A1(n8206), .A2(n8819), .ZN(n7511) );
  NAND2_X1 U9121 ( .A1(n8820), .A2(n8821), .ZN(n7510) );
  NAND2_X1 U9122 ( .A1(n7511), .A2(n7510), .ZN(n7523) );
  INV_X1 U9123 ( .A(n7523), .ZN(n7512) );
  OAI21_X1 U9124 ( .B1(n7514), .B2(n7513), .A(n7512), .ZN(n9629) );
  INV_X1 U9125 ( .A(n8581), .ZN(n9627) );
  OAI21_X1 U9126 ( .B1(n9627), .B2(n4391), .A(n4331), .ZN(n9628) );
  OAI22_X1 U9127 ( .A1(n4316), .A2(n7515), .B1(n7526), .B2(n9827), .ZN(n7516)
         );
  AOI21_X1 U9128 ( .B1(n8581), .B2(n9831), .A(n7516), .ZN(n7517) );
  OAI21_X1 U9129 ( .B1(n9628), .B2(n9833), .A(n7517), .ZN(n7518) );
  AOI21_X1 U9130 ( .B1(n9629), .B2(n4316), .A(n7518), .ZN(n7519) );
  OAI21_X1 U9131 ( .B1(n9825), .B2(n7520), .A(n7519), .ZN(P2_U3282) );
  AOI21_X1 U9132 ( .B1(n7522), .B2(n7521), .A(n4393), .ZN(n7529) );
  NAND2_X1 U9133 ( .A1(n8197), .A2(n7523), .ZN(n7524) );
  OAI211_X1 U9134 ( .C1(n8200), .C2(n7526), .A(n7525), .B(n7524), .ZN(n7527)
         );
  AOI21_X1 U9135 ( .B1(n8581), .B2(n8202), .A(n7527), .ZN(n7528) );
  OAI21_X1 U9136 ( .B1(n7529), .B2(n8204), .A(n7528), .ZN(P2_U3217) );
  OR2_X1 U9137 ( .A1(n9488), .A2(n9235), .ZN(n7730) );
  NAND2_X1 U9138 ( .A1(n9488), .A2(n9235), .ZN(n9230) );
  INV_X1 U9139 ( .A(n9256), .ZN(n9246) );
  NAND2_X1 U9140 ( .A1(n9493), .A2(n7530), .ZN(n7727) );
  INV_X1 U9141 ( .A(n9271), .ZN(n7565) );
  AND2_X1 U9142 ( .A1(n9498), .A2(n9295), .ZN(n9228) );
  NOR2_X1 U9143 ( .A1(n9498), .A2(n9295), .ZN(n7531) );
  NAND2_X1 U9144 ( .A1(n9505), .A2(n9310), .ZN(n9227) );
  OR2_X1 U9145 ( .A1(n9513), .A2(n9309), .ZN(n9224) );
  NAND2_X1 U9146 ( .A1(n9513), .A2(n9309), .ZN(n7714) );
  NAND2_X1 U9147 ( .A1(n9224), .A2(n7714), .ZN(n9329) );
  OR2_X1 U9148 ( .A1(n9519), .A2(n9356), .ZN(n7712) );
  NAND2_X1 U9149 ( .A1(n9519), .A2(n9356), .ZN(n9223) );
  NAND2_X1 U9150 ( .A1(n9525), .A2(n9201), .ZN(n7704) );
  NAND2_X1 U9151 ( .A1(n7709), .A2(n7704), .ZN(n9351) );
  INV_X1 U9152 ( .A(n9394), .ZN(n9357) );
  OR2_X1 U9153 ( .A1(n9528), .A2(n9357), .ZN(n9220) );
  NAND2_X1 U9154 ( .A1(n9528), .A2(n9357), .ZN(n7701) );
  OR2_X1 U9155 ( .A1(n9539), .A2(n9048), .ZN(n7698) );
  NAND2_X1 U9156 ( .A1(n9539), .A2(n9048), .ZN(n7702) );
  OR2_X1 U9157 ( .A1(n9533), .A2(n9199), .ZN(n7699) );
  NAND2_X1 U9158 ( .A1(n9533), .A2(n9199), .ZN(n7700) );
  NAND2_X1 U9159 ( .A1(n7699), .A2(n7700), .ZN(n9219) );
  INV_X1 U9160 ( .A(n9219), .ZN(n9393) );
  OR2_X1 U9161 ( .A1(n9552), .A2(n9108), .ZN(n7691) );
  NAND2_X1 U9162 ( .A1(n9552), .A2(n9108), .ZN(n9215) );
  NAND2_X1 U9163 ( .A1(n7691), .A2(n9215), .ZN(n9433) );
  NAND2_X1 U9164 ( .A1(n7539), .A2(n7532), .ZN(n7634) );
  INV_X1 U9165 ( .A(n7637), .ZN(n7533) );
  NOR2_X1 U9166 ( .A1(n7634), .A2(n7533), .ZN(n7761) );
  OR2_X1 U9167 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NOR2_X1 U9168 ( .A1(n7536), .A2(n6737), .ZN(n7545) );
  NAND2_X1 U9169 ( .A1(n7538), .A2(n7537), .ZN(n7540) );
  NAND2_X1 U9170 ( .A1(n7540), .A2(n7539), .ZN(n7544) );
  AND2_X1 U9171 ( .A1(n7542), .A2(n7541), .ZN(n7543) );
  AND2_X1 U9172 ( .A1(n7544), .A2(n7543), .ZN(n7639) );
  NAND4_X1 U9173 ( .A1(n7761), .A2(n7546), .A3(n7545), .A4(n7639), .ZN(n7549)
         );
  NOR3_X1 U9174 ( .A1(n7549), .A2(n6901), .A3(n7548), .ZN(n7551) );
  NAND4_X1 U9175 ( .A1(n7553), .A2(n7552), .A3(n7551), .A4(n4657), .ZN(n7555)
         );
  NOR2_X1 U9176 ( .A1(n7555), .A2(n7554), .ZN(n7556) );
  NAND4_X1 U9177 ( .A1(n4654), .A2(n7557), .A3(n7690), .A4(n7556), .ZN(n7558)
         );
  OR2_X1 U9178 ( .A1(n9545), .A2(n9439), .ZN(n9399) );
  NAND2_X1 U9179 ( .A1(n9545), .A2(n9439), .ZN(n9216) );
  INV_X1 U9180 ( .A(n9415), .ZN(n9422) );
  NOR2_X1 U9181 ( .A1(n7558), .A2(n9422), .ZN(n7559) );
  NAND4_X1 U9182 ( .A1(n9368), .A2(n9410), .A3(n9393), .A4(n7559), .ZN(n7560)
         );
  NOR2_X1 U9183 ( .A1(n9351), .A2(n7560), .ZN(n7561) );
  NAND2_X1 U9184 ( .A1(n9344), .A2(n7561), .ZN(n7562) );
  NOR2_X1 U9185 ( .A1(n9329), .A2(n7562), .ZN(n7563) );
  XNOR2_X1 U9186 ( .A(n9510), .B(n9330), .ZN(n9306) );
  INV_X1 U9187 ( .A(n9306), .ZN(n9303) );
  NAND3_X1 U9188 ( .A1(n4861), .A2(n7563), .A3(n9303), .ZN(n7564) );
  NOR4_X1 U9189 ( .A1(n9246), .A2(n7565), .A3(n9284), .A4(n7564), .ZN(n7605)
         );
  NAND2_X1 U9190 ( .A1(n7567), .A2(n7566), .ZN(n7569) );
  INV_X1 U9191 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8981) );
  INV_X1 U9192 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7806) );
  MUX2_X1 U9193 ( .A(n8981), .B(n7806), .S(n4409), .Z(n7571) );
  INV_X1 U9194 ( .A(SI_29_), .ZN(n7570) );
  NAND2_X1 U9195 ( .A1(n7571), .A2(n7570), .ZN(n7574) );
  INV_X1 U9196 ( .A(n7571), .ZN(n7572) );
  NAND2_X1 U9197 ( .A1(n7572), .A2(SI_29_), .ZN(n7573) );
  NAND2_X1 U9198 ( .A1(n7592), .A2(n7591), .ZN(n7575) );
  NAND2_X1 U9199 ( .A1(n7575), .A2(n7574), .ZN(n7596) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7850) );
  INV_X1 U9201 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8076) );
  MUX2_X1 U9202 ( .A(n7850), .B(n8076), .S(n4409), .Z(n7577) );
  INV_X1 U9203 ( .A(SI_30_), .ZN(n7576) );
  NAND2_X1 U9204 ( .A1(n7577), .A2(n7576), .ZN(n7580) );
  INV_X1 U9205 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U9206 ( .A1(n7578), .A2(SI_30_), .ZN(n7579) );
  NAND2_X1 U9207 ( .A1(n7596), .A2(n7595), .ZN(n7581) );
  NAND2_X1 U9208 ( .A1(n7581), .A2(n7580), .ZN(n7584) );
  INV_X1 U9209 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8975) );
  MUX2_X1 U9210 ( .A(n8975), .B(n6304), .S(n4409), .Z(n7582) );
  XNOR2_X1 U9211 ( .A(n7582), .B(SI_31_), .ZN(n7583) );
  NAND2_X1 U9212 ( .A1(n9586), .A2(n5245), .ZN(n7586) );
  OR2_X1 U9213 ( .A1(n7597), .A2(n6304), .ZN(n7585) );
  NAND2_X2 U9214 ( .A1(n7586), .A2(n7585), .ZN(n9476) );
  NAND2_X1 U9215 ( .A1(n7601), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9216 ( .A1(n7587), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U9217 ( .A1(n7600), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7588) );
  AND3_X1 U9218 ( .A1(n7590), .A2(n7589), .A3(n7588), .ZN(n9188) );
  XNOR2_X1 U9219 ( .A(n7592), .B(n7591), .ZN(n7845) );
  NAND2_X1 U9220 ( .A1(n7845), .A2(n5245), .ZN(n7594) );
  OR2_X1 U9221 ( .A1(n7597), .A2(n7806), .ZN(n7593) );
  XNOR2_X1 U9222 ( .A(n9237), .B(n9258), .ZN(n9231) );
  XNOR2_X1 U9223 ( .A(n7596), .B(n7595), .ZN(n7849) );
  NAND2_X1 U9224 ( .A1(n7849), .A2(n5245), .ZN(n7599) );
  OR2_X1 U9225 ( .A1(n7597), .A2(n8076), .ZN(n7598) );
  NAND2_X1 U9226 ( .A1(n7600), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9227 ( .A1(n7587), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9228 ( .A1(n7601), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9229 ( .A1(n9480), .A2(n9233), .ZN(n7784) );
  NAND4_X1 U9230 ( .A1(n7605), .A2(n7790), .A3(n9231), .A4(n7784), .ZN(n7607)
         );
  NAND2_X1 U9231 ( .A1(n9476), .A2(n9188), .ZN(n7735) );
  NOR2_X1 U9232 ( .A1(n9480), .A2(n9233), .ZN(n7608) );
  INV_X1 U9233 ( .A(n7608), .ZN(n7606) );
  NAND2_X1 U9234 ( .A1(n7735), .A2(n7606), .ZN(n7760) );
  OAI21_X1 U9235 ( .B1(n7607), .B2(n7760), .A(n7755), .ZN(n7752) );
  INV_X1 U9236 ( .A(n7752), .ZN(n7670) );
  NAND2_X1 U9237 ( .A1(n7608), .A2(n9476), .ZN(n7737) );
  NAND2_X1 U9238 ( .A1(n7737), .A2(n7735), .ZN(n7746) );
  INV_X1 U9239 ( .A(n7746), .ZN(n7668) );
  OR2_X1 U9240 ( .A1(n9237), .A2(n7741), .ZN(n7609) );
  AND2_X1 U9241 ( .A1(n7609), .A2(n7730), .ZN(n7664) );
  INV_X1 U9242 ( .A(n7664), .ZN(n7612) );
  NAND2_X1 U9243 ( .A1(n9498), .A2(n9282), .ZN(n7610) );
  NAND2_X1 U9244 ( .A1(n9282), .A2(n9295), .ZN(n7721) );
  NAND2_X1 U9245 ( .A1(n7610), .A2(n7721), .ZN(n9229) );
  INV_X1 U9246 ( .A(n9229), .ZN(n7611) );
  OR2_X1 U9247 ( .A1(n7612), .A2(n7611), .ZN(n7787) );
  INV_X1 U9248 ( .A(n7701), .ZN(n7613) );
  NAND2_X1 U9249 ( .A1(n7709), .A2(n7613), .ZN(n7614) );
  AND2_X1 U9250 ( .A1(n7614), .A2(n7704), .ZN(n7615) );
  AND2_X1 U9251 ( .A1(n9223), .A2(n7615), .ZN(n7710) );
  NAND2_X1 U9252 ( .A1(n9220), .A2(n7699), .ZN(n7703) );
  INV_X1 U9253 ( .A(n7703), .ZN(n7617) );
  AND2_X1 U9254 ( .A1(n7698), .A2(n9399), .ZN(n9218) );
  INV_X1 U9255 ( .A(n9218), .ZN(n7694) );
  NAND3_X1 U9256 ( .A1(n7694), .A2(n7702), .A3(n7700), .ZN(n7616) );
  NAND3_X1 U9257 ( .A1(n7709), .A2(n7617), .A3(n7616), .ZN(n7618) );
  NAND2_X1 U9258 ( .A1(n7710), .A2(n7618), .ZN(n7619) );
  AND2_X1 U9259 ( .A1(n7619), .A2(n7712), .ZN(n7778) );
  INV_X1 U9260 ( .A(n7710), .ZN(n7620) );
  INV_X1 U9261 ( .A(n7700), .ZN(n9366) );
  NOR2_X1 U9262 ( .A1(n7620), .A2(n9366), .ZN(n7776) );
  AND2_X1 U9263 ( .A1(n9216), .A2(n9215), .ZN(n7621) );
  NAND2_X1 U9264 ( .A1(n7702), .A2(n7621), .ZN(n7655) );
  NAND2_X1 U9265 ( .A1(n7623), .A2(n7622), .ZN(n7682) );
  AND2_X1 U9266 ( .A1(n7625), .A2(n7624), .ZN(n7676) );
  INV_X1 U9267 ( .A(n7676), .ZN(n7626) );
  NAND2_X1 U9268 ( .A1(n7626), .A2(n7675), .ZN(n7628) );
  NAND2_X1 U9269 ( .A1(n9651), .A2(n7627), .ZN(n7678) );
  AND2_X1 U9270 ( .A1(n7628), .A2(n7678), .ZN(n7629) );
  NAND2_X1 U9271 ( .A1(n7683), .A2(n7629), .ZN(n7647) );
  NAND2_X1 U9272 ( .A1(n7631), .A2(n7630), .ZN(n7632) );
  OR3_X1 U9273 ( .A1(n7682), .A2(n7647), .A3(n7632), .ZN(n7633) );
  OR3_X1 U9274 ( .A1(n7655), .A2(n9212), .A3(n7633), .ZN(n7774) );
  INV_X1 U9275 ( .A(n7634), .ZN(n7635) );
  NAND2_X1 U9276 ( .A1(n7636), .A2(n7635), .ZN(n7640) );
  NAND2_X1 U9277 ( .A1(n7768), .A2(n7637), .ZN(n7638) );
  AOI21_X1 U9278 ( .B1(n7640), .B2(n7639), .A(n7638), .ZN(n7656) );
  OR2_X1 U9279 ( .A1(n7682), .A2(n7641), .ZN(n7643) );
  NAND2_X1 U9280 ( .A1(n7643), .A2(n7642), .ZN(n7681) );
  NOR2_X1 U9281 ( .A1(n7682), .A2(n7644), .ZN(n7645) );
  NOR2_X1 U9282 ( .A1(n7681), .A2(n7645), .ZN(n7685) );
  INV_X1 U9283 ( .A(n7685), .ZN(n7652) );
  AND2_X1 U9284 ( .A1(n7646), .A2(n7671), .ZN(n7648) );
  OR3_X1 U9285 ( .A1(n7682), .A2(n7648), .A3(n7647), .ZN(n7649) );
  NAND2_X1 U9286 ( .A1(n9213), .A2(n7649), .ZN(n7651) );
  OAI21_X1 U9287 ( .B1(n7652), .B2(n7651), .A(n7650), .ZN(n7653) );
  AND2_X1 U9288 ( .A1(n7653), .A2(n7691), .ZN(n7654) );
  OR2_X1 U9289 ( .A1(n7655), .A2(n7654), .ZN(n7772) );
  OAI21_X1 U9290 ( .B1(n7774), .B2(n7656), .A(n7772), .ZN(n7657) );
  NAND2_X1 U9291 ( .A1(n7776), .A2(n7657), .ZN(n7658) );
  INV_X1 U9292 ( .A(n7714), .ZN(n7777) );
  AOI21_X1 U9293 ( .B1(n7778), .B2(n7658), .A(n7777), .ZN(n7659) );
  OR2_X1 U9294 ( .A1(n9510), .A2(n9330), .ZN(n7716) );
  NAND2_X1 U9295 ( .A1(n7716), .A2(n9224), .ZN(n7781) );
  NAND2_X1 U9296 ( .A1(n9510), .A2(n9330), .ZN(n7713) );
  AND2_X1 U9297 ( .A1(n9227), .A2(n7713), .ZN(n7780) );
  OAI21_X1 U9298 ( .B1(n7659), .B2(n7781), .A(n7780), .ZN(n7660) );
  NAND2_X1 U9299 ( .A1(n9253), .A2(n7660), .ZN(n7666) );
  NAND2_X1 U9300 ( .A1(n9253), .A2(n9228), .ZN(n7661) );
  NAND3_X1 U9301 ( .A1(n9230), .A2(n7727), .A3(n7661), .ZN(n7663) );
  AND2_X1 U9302 ( .A1(n9237), .A2(n7741), .ZN(n7662) );
  AOI21_X1 U9303 ( .B1(n7664), .B2(n7663), .A(n7662), .ZN(n7785) );
  INV_X1 U9304 ( .A(n9233), .ZN(n9120) );
  INV_X1 U9305 ( .A(n9188), .ZN(n9119) );
  NAND2_X1 U9306 ( .A1(n9120), .A2(n9119), .ZN(n7665) );
  NAND2_X1 U9307 ( .A1(n9480), .A2(n7665), .ZN(n7743) );
  OAI211_X1 U9308 ( .C1(n7787), .C2(n7666), .A(n7785), .B(n7743), .ZN(n7667)
         );
  INV_X1 U9309 ( .A(n7790), .ZN(n7756) );
  AOI211_X1 U9310 ( .C1(n7668), .C2(n7667), .A(n7755), .B(n7756), .ZN(n7669)
         );
  NOR2_X1 U9311 ( .A1(n7670), .A2(n7669), .ZN(n7754) );
  NAND3_X1 U9312 ( .A1(n7687), .A2(n7683), .A3(n7678), .ZN(n7680) );
  INV_X1 U9313 ( .A(n7682), .ZN(n7684) );
  NAND2_X1 U9314 ( .A1(n7684), .A2(n7683), .ZN(n7686) );
  OAI21_X1 U9315 ( .B1(n7687), .B2(n7686), .A(n7685), .ZN(n7688) );
  MUX2_X1 U9316 ( .A(n9212), .B(n4656), .S(n7740), .Z(n7689) );
  MUX2_X1 U9317 ( .A(n9215), .B(n7691), .S(n7740), .Z(n7692) );
  OAI21_X1 U9318 ( .B1(n7693), .B2(n9433), .A(n7692), .ZN(n7697) );
  NAND2_X1 U9319 ( .A1(n7702), .A2(n9216), .ZN(n7695) );
  MUX2_X1 U9320 ( .A(n7695), .B(n7694), .S(n7740), .Z(n7696) );
  NAND2_X1 U9321 ( .A1(n7701), .A2(n7700), .ZN(n9221) );
  INV_X1 U9322 ( .A(n7702), .ZN(n9217) );
  INV_X1 U9323 ( .A(n9220), .ZN(n7705) );
  OAI21_X1 U9324 ( .B1(n7708), .B2(n7705), .A(n7704), .ZN(n7706) );
  NAND3_X1 U9325 ( .A1(n7706), .A2(n7709), .A3(n7712), .ZN(n7707) );
  AOI211_X1 U9326 ( .C1(n7707), .C2(n9223), .A(n7781), .B(n7740), .ZN(n7719)
         );
  INV_X1 U9327 ( .A(n7708), .ZN(n7711) );
  INV_X1 U9328 ( .A(n7709), .ZN(n9222) );
  NOR2_X1 U9329 ( .A1(n7714), .A2(n7740), .ZN(n7715) );
  AOI22_X1 U9330 ( .A1(n4722), .A2(n4589), .B1(n7716), .B2(n7715), .ZN(n7717)
         );
  OAI21_X1 U9331 ( .B1(n7740), .B2(n9227), .A(n7717), .ZN(n7718) );
  NAND2_X1 U9332 ( .A1(n7720), .A2(n9282), .ZN(n7724) );
  INV_X1 U9333 ( .A(n7721), .ZN(n7722) );
  NOR2_X1 U9334 ( .A1(n9228), .A2(n7722), .ZN(n7723) );
  MUX2_X1 U9335 ( .A(n9498), .B(n7723), .S(n4589), .Z(n7725) );
  OAI21_X1 U9336 ( .B1(n7726), .B2(n7725), .A(n9271), .ZN(n7729) );
  MUX2_X1 U9337 ( .A(n9253), .B(n7727), .S(n7740), .Z(n7728) );
  NAND4_X1 U9338 ( .A1(n7737), .A2(n7740), .A3(n9237), .A4(n7730), .ZN(n7733)
         );
  INV_X1 U9339 ( .A(n7735), .ZN(n7732) );
  NAND4_X1 U9340 ( .A1(n7743), .A2(n4589), .A3(n9230), .A4(n9258), .ZN(n7731)
         );
  OAI21_X1 U9341 ( .B1(n7733), .B2(n7732), .A(n7731), .ZN(n7750) );
  OAI21_X1 U9342 ( .B1(n4589), .B2(n7743), .A(n7735), .ZN(n7734) );
  OAI21_X1 U9343 ( .B1(n4589), .B2(n7735), .A(n7734), .ZN(n7736) );
  OAI211_X1 U9344 ( .C1(n7740), .C2(n7737), .A(n7736), .B(n7790), .ZN(n7749)
         );
  INV_X1 U9345 ( .A(n9235), .ZN(n9273) );
  NAND3_X1 U9346 ( .A1(n9252), .A2(n7740), .A3(n9273), .ZN(n7738) );
  INV_X1 U9347 ( .A(n9237), .ZN(n9484) );
  INV_X1 U9348 ( .A(n9230), .ZN(n7739) );
  AOI21_X1 U9349 ( .B1(n7741), .B2(n7739), .A(n9237), .ZN(n7742) );
  MUX2_X1 U9350 ( .A(n7742), .B(n7741), .S(n7740), .Z(n7744) );
  NAND2_X1 U9351 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  AOI211_X1 U9352 ( .C1(n7747), .C2(n9484), .A(n7746), .B(n7745), .ZN(n7748)
         );
  NOR4_X1 U9353 ( .A1(n7757), .A2(n5061), .A3(n7756), .A4(n7755), .ZN(n7758)
         );
  NOR3_X1 U9354 ( .A1(n7759), .A2(n7758), .A3(n7792), .ZN(n7802) );
  INV_X1 U9355 ( .A(n7760), .ZN(n7789) );
  INV_X1 U9356 ( .A(n7761), .ZN(n7767) );
  NAND4_X1 U9357 ( .A1(n7765), .A2(n7764), .A3(n7763), .A4(n7762), .ZN(n7766)
         );
  NOR2_X1 U9358 ( .A1(n7767), .A2(n7766), .ZN(n7769) );
  OAI21_X1 U9359 ( .B1(n7770), .B2(n7769), .A(n7768), .ZN(n7771) );
  INV_X1 U9360 ( .A(n7771), .ZN(n7773) );
  OAI21_X1 U9361 ( .B1(n7774), .B2(n7773), .A(n7772), .ZN(n7775) );
  NAND2_X1 U9362 ( .A1(n7776), .A2(n7775), .ZN(n7779) );
  AOI21_X1 U9363 ( .B1(n7779), .B2(n7778), .A(n7777), .ZN(n7782) );
  OAI21_X1 U9364 ( .B1(n7782), .B2(n7781), .A(n7780), .ZN(n7783) );
  NAND2_X1 U9365 ( .A1(n9253), .A2(n7783), .ZN(n7786) );
  OAI211_X1 U9366 ( .C1(n7787), .C2(n7786), .A(n7785), .B(n7784), .ZN(n7788)
         );
  NAND2_X1 U9367 ( .A1(n7789), .A2(n7788), .ZN(n7791) );
  NAND2_X1 U9368 ( .A1(n7791), .A2(n7790), .ZN(n7796) );
  NAND3_X1 U9369 ( .A1(n7796), .A2(n9315), .A3(n7792), .ZN(n7794) );
  OAI211_X1 U9370 ( .C1(n7796), .C2(n7795), .A(n7794), .B(n7793), .ZN(n7801)
         );
  NOR3_X1 U9371 ( .A1(n7797), .A2(n6268), .A3(n9438), .ZN(n7800) );
  OAI21_X1 U9372 ( .B1(n5061), .B2(n7798), .A(P1_B_REG_SCAN_IN), .ZN(n7799) );
  OAI22_X1 U9373 ( .A1(n7802), .A2(n7801), .B1(n7800), .B2(n7799), .ZN(
        P1_U3240) );
  INV_X1 U9374 ( .A(n7849), .ZN(n8078) );
  OAI222_X1 U9375 ( .A1(P1_U3084), .A2(n5539), .B1(n9597), .B2(n7805), .C1(
        n7804), .C2(n9593), .ZN(P1_U3327) );
  INV_X1 U9376 ( .A(n7845), .ZN(n8983) );
  OAI222_X1 U9377 ( .A1(n9593), .A2(n7806), .B1(n9597), .B2(n8983), .C1(n5038), 
        .C2(P1_U3084), .ZN(P1_U3324) );
  INV_X1 U9378 ( .A(n7807), .ZN(n7808) );
  AND2_X1 U9379 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  NAND2_X1 U9380 ( .A1(n9589), .A2(n5790), .ZN(n7813) );
  OR2_X1 U9381 ( .A1(n7859), .A2(n8088), .ZN(n7812) );
  NAND2_X1 U9382 ( .A1(n8641), .A2(n5678), .ZN(n7815) );
  XNOR2_X1 U9383 ( .A(n7815), .B(n5679), .ZN(n7818) );
  NOR3_X1 U9384 ( .A1(n8621), .A2(n8202), .A3(n7818), .ZN(n7816) );
  AOI21_X1 U9385 ( .B1(n8621), .B2(n7818), .A(n7816), .ZN(n7822) );
  NAND3_X1 U9386 ( .A1(n8875), .A2(n8191), .A3(n7818), .ZN(n7817) );
  OAI21_X1 U9387 ( .B1(n8875), .B2(n7818), .A(n7817), .ZN(n7819) );
  OAI21_X1 U9388 ( .B1(n8621), .B2(n8191), .A(n8204), .ZN(n7820) );
  OAI211_X1 U9389 ( .C1(n7823), .C2(n7822), .A(n7821), .B(n7820), .ZN(n7835)
         );
  OR2_X1 U9390 ( .A1(n8607), .A2(n7824), .ZN(n7830) );
  INV_X1 U9391 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8606) );
  NAND2_X1 U9392 ( .A1(n6021), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U9393 ( .A1(n7825), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7826) );
  OAI211_X1 U9394 ( .C1(n8606), .C2(n7858), .A(n7827), .B(n7826), .ZN(n7828)
         );
  INV_X1 U9395 ( .A(n7828), .ZN(n7829) );
  NAND2_X1 U9396 ( .A1(n7830), .A2(n7829), .ZN(n8618) );
  AOI22_X1 U9397 ( .A1(n8174), .A2(n8618), .B1(n8619), .B2(n8175), .ZN(n7833)
         );
  INV_X1 U9398 ( .A(n8623), .ZN(n7831) );
  AOI22_X1 U9399 ( .A1(n7831), .A2(n8137), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7832) );
  AND2_X1 U9400 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  NAND2_X1 U9401 ( .A1(n7835), .A2(n7834), .ZN(P2_U3222) );
  INV_X1 U9402 ( .A(n8938), .ZN(n8849) );
  INV_X1 U9403 ( .A(n8820), .ZN(n8135) );
  XNOR2_X1 U9404 ( .A(n8938), .B(n8135), .ZN(n8839) );
  INV_X1 U9405 ( .A(n8584), .ZN(n8803) );
  NAND2_X1 U9406 ( .A1(n8933), .A2(n8803), .ZN(n7981) );
  INV_X1 U9407 ( .A(n7981), .ZN(n7836) );
  INV_X1 U9408 ( .A(n8822), .ZN(n8134) );
  OR2_X1 U9409 ( .A1(n8930), .A2(n8134), .ZN(n8788) );
  NAND2_X1 U9410 ( .A1(n8930), .A2(n8134), .ZN(n7985) );
  NAND2_X1 U9411 ( .A1(n8788), .A2(n7985), .ZN(n8811) );
  INV_X1 U9412 ( .A(n8811), .ZN(n8800) );
  NAND2_X1 U9413 ( .A1(n8801), .A2(n8800), .ZN(n8789) );
  OR2_X1 U9414 ( .A1(n8923), .A2(n8805), .ZN(n7989) );
  NAND2_X1 U9415 ( .A1(n8923), .A2(n8805), .ZN(n7997) );
  INV_X1 U9416 ( .A(n8793), .ZN(n8588) );
  OR2_X1 U9417 ( .A1(n8920), .A2(n8588), .ZN(n7990) );
  NAND2_X1 U9418 ( .A1(n8920), .A2(n8588), .ZN(n8753) );
  INV_X1 U9419 ( .A(n8766), .ZN(n8111) );
  NAND2_X1 U9420 ( .A1(n8914), .A2(n8111), .ZN(n7999) );
  NAND2_X1 U9421 ( .A1(n8001), .A2(n7999), .ZN(n8755) );
  INV_X1 U9422 ( .A(n8753), .ZN(n7991) );
  NOR2_X1 U9423 ( .A1(n8755), .A2(n7991), .ZN(n7837) );
  INV_X1 U9424 ( .A(n8001), .ZN(n7993) );
  OR2_X1 U9425 ( .A1(n8909), .A2(n8725), .ZN(n8000) );
  NAND2_X1 U9426 ( .A1(n8909), .A2(n8725), .ZN(n8722) );
  INV_X1 U9427 ( .A(n8740), .ZN(n8591) );
  NAND2_X1 U9428 ( .A1(n8904), .A2(n8591), .ZN(n8011) );
  NAND2_X1 U9429 ( .A1(n8005), .A2(n8011), .ZN(n8592) );
  NAND3_X1 U9430 ( .A1(n8737), .A2(n8721), .A3(n8722), .ZN(n8720) );
  XNOR2_X1 U9431 ( .A(n8899), .B(n8726), .ZN(n8706) );
  NAND2_X1 U9432 ( .A1(n8894), .A2(n8708), .ZN(n7838) );
  NAND2_X1 U9433 ( .A1(n8593), .A2(n7838), .ZN(n8687) );
  INV_X1 U9434 ( .A(n8894), .ZN(n8685) );
  NAND2_X1 U9435 ( .A1(n8685), .A2(n8708), .ZN(n7897) );
  NAND2_X1 U9436 ( .A1(n8686), .A2(n7897), .ZN(n7839) );
  INV_X1 U9437 ( .A(n8690), .ZN(n8149) );
  NAND2_X1 U9438 ( .A1(n8891), .A2(n8149), .ZN(n8023) );
  NAND2_X1 U9439 ( .A1(n7839), .A2(n8667), .ZN(n8671) );
  INV_X1 U9440 ( .A(n8020), .ZN(n7841) );
  INV_X1 U9441 ( .A(n8649), .ZN(n7840) );
  NOR2_X1 U9442 ( .A1(n7841), .A2(n7840), .ZN(n7894) );
  NAND2_X1 U9443 ( .A1(n8886), .A2(n8594), .ZN(n8021) );
  INV_X1 U9444 ( .A(n8021), .ZN(n7842) );
  AOI21_X1 U9445 ( .B1(n8671), .B2(n7894), .A(n7842), .ZN(n8639) );
  NAND2_X1 U9446 ( .A1(n8639), .A2(n8638), .ZN(n8637) );
  NAND2_X1 U9447 ( .A1(n8636), .A2(n8619), .ZN(n8028) );
  NAND2_X1 U9448 ( .A1(n8637), .A2(n8028), .ZN(n8617) );
  NAND2_X1 U9449 ( .A1(n8875), .A2(n8595), .ZN(n8033) );
  NAND2_X1 U9450 ( .A1(n8032), .A2(n8033), .ZN(n8616) );
  INV_X1 U9451 ( .A(n8616), .ZN(n8614) );
  INV_X1 U9452 ( .A(n8032), .ZN(n7843) );
  NOR2_X1 U9453 ( .A1(n7859), .A2(n8981), .ZN(n7844) );
  AOI21_X1 U9454 ( .B1(n7845), .B2(n5790), .A(n7844), .ZN(n8869) );
  NOR2_X1 U9455 ( .A1(n8869), .A2(n8618), .ZN(n8036) );
  INV_X1 U9456 ( .A(n8869), .ZN(n8609) );
  INV_X1 U9457 ( .A(n8618), .ZN(n7846) );
  NOR2_X1 U9458 ( .A1(n8609), .A2(n7846), .ZN(n8037) );
  NAND2_X1 U9459 ( .A1(n8601), .A2(n8600), .ZN(n7848) );
  INV_X1 U9460 ( .A(n8036), .ZN(n7847) );
  NAND2_X1 U9461 ( .A1(n7849), .A2(n5790), .ZN(n7852) );
  OR2_X1 U9462 ( .A1(n7859), .A2(n7850), .ZN(n7851) );
  INV_X1 U9463 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U9464 ( .A1(n5703), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7856) );
  INV_X1 U9465 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7853) );
  OR2_X1 U9466 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  OAI211_X1 U9467 ( .C1(n7858), .C2(n7857), .A(n7856), .B(n7855), .ZN(n8602)
         );
  NAND2_X1 U9468 ( .A1(n8867), .A2(n8602), .ZN(n8038) );
  NAND2_X1 U9469 ( .A1(n9586), .A2(n5790), .ZN(n7861) );
  OR2_X1 U9470 ( .A1(n7859), .A2(n8975), .ZN(n7860) );
  NAND2_X1 U9471 ( .A1(n7861), .A2(n7860), .ZN(n8571) );
  OR2_X1 U9472 ( .A1(n8571), .A2(n7862), .ZN(n8048) );
  INV_X1 U9473 ( .A(n8602), .ZN(n7863) );
  NAND2_X1 U9474 ( .A1(n8576), .A2(n7863), .ZN(n8039) );
  NAND2_X1 U9475 ( .A1(n8048), .A2(n8039), .ZN(n8044) );
  NAND2_X1 U9476 ( .A1(n5678), .A2(n7864), .ZN(n8058) );
  INV_X1 U9477 ( .A(n7891), .ZN(n7866) );
  NOR2_X1 U9478 ( .A1(n7866), .A2(n7865), .ZN(n8056) );
  NAND2_X1 U9479 ( .A1(n4823), .A2(n8038), .ZN(n8043) );
  INV_X1 U9480 ( .A(n8043), .ZN(n7889) );
  INV_X1 U9481 ( .A(n8044), .ZN(n7888) );
  INV_X1 U9482 ( .A(n8638), .ZN(n8628) );
  NAND2_X1 U9483 ( .A1(n8020), .A2(n8021), .ZN(n8650) );
  INV_X1 U9484 ( .A(n8833), .ZN(n7882) );
  NOR2_X1 U9485 ( .A1(n9852), .A2(n6873), .ZN(n7873) );
  NAND2_X1 U9486 ( .A1(n7903), .A2(n7892), .ZN(n7867) );
  NOR2_X1 U9487 ( .A1(n6947), .A2(n7867), .ZN(n7872) );
  NAND2_X1 U9488 ( .A1(n7926), .A2(n7868), .ZN(n7901) );
  INV_X1 U9489 ( .A(n7901), .ZN(n7870) );
  AND2_X1 U9490 ( .A1(n7870), .A2(n7869), .ZN(n7925) );
  NAND2_X1 U9491 ( .A1(n7906), .A2(n7904), .ZN(n7902) );
  INV_X1 U9492 ( .A(n7902), .ZN(n7871) );
  AND4_X1 U9493 ( .A1(n7873), .A2(n7872), .A3(n7925), .A4(n7871), .ZN(n7875)
         );
  NAND4_X1 U9494 ( .A1(n7875), .A2(n7931), .A3(n4689), .A4(n7874), .ZN(n7878)
         );
  NOR4_X1 U9495 ( .A1(n7878), .A2(n7877), .A3(n7942), .A4(n7876), .ZN(n7879)
         );
  NAND4_X1 U9496 ( .A1(n8582), .A2(n7968), .A3(n7880), .A4(n7879), .ZN(n7881)
         );
  NOR4_X1 U9497 ( .A1(n8811), .A2(n7882), .A3(n8839), .A4(n7881), .ZN(n7883)
         );
  NAND3_X1 U9498 ( .A1(n8764), .A2(n8791), .A3(n7883), .ZN(n7884) );
  NOR4_X1 U9499 ( .A1(n8592), .A2(n4806), .A3(n8755), .A4(n7884), .ZN(n7885)
         );
  INV_X1 U9500 ( .A(n8706), .ZN(n8009) );
  NAND4_X1 U9501 ( .A1(n8667), .A2(n7885), .A3(n8009), .A4(n8687), .ZN(n7886)
         );
  NOR4_X1 U9502 ( .A1(n8616), .A2(n8628), .A3(n8650), .A4(n7886), .ZN(n7887)
         );
  NAND4_X1 U9503 ( .A1(n7889), .A2(n8600), .A3(n7888), .A4(n7887), .ZN(n7890)
         );
  XNOR2_X1 U9504 ( .A(n7890), .B(n8807), .ZN(n7893) );
  OAI22_X1 U9505 ( .A1(n7893), .A2(n7909), .B1(n7892), .B2(n7891), .ZN(n8055)
         );
  INV_X1 U9506 ( .A(n7894), .ZN(n8019) );
  NOR2_X1 U9507 ( .A1(n8063), .A2(n7895), .ZN(n7896) );
  NAND2_X1 U9508 ( .A1(n5654), .A2(n7896), .ZN(n8049) );
  INV_X1 U9509 ( .A(n8049), .ZN(n8018) );
  NOR2_X1 U9510 ( .A1(n8685), .A2(n8708), .ZN(n7898) );
  INV_X1 U9511 ( .A(n7897), .ZN(n8666) );
  MUX2_X1 U9512 ( .A(n7898), .B(n8666), .S(n8049), .Z(n7899) );
  NOR2_X1 U9513 ( .A1(n4679), .A2(n7899), .ZN(n8017) );
  AND2_X1 U9514 ( .A1(n7941), .A2(n7900), .ZN(n7940) );
  MUX2_X1 U9515 ( .A(n7902), .B(n7901), .S(n8049), .Z(n7927) );
  AND2_X1 U9516 ( .A1(n7904), .A2(n7903), .ZN(n7907) );
  INV_X1 U9517 ( .A(n7933), .ZN(n7905) );
  OAI211_X1 U9518 ( .C1(n7927), .C2(n7907), .A(n7906), .B(n7905), .ZN(n7908)
         );
  NAND2_X1 U9519 ( .A1(n7908), .A2(n8049), .ZN(n7917) );
  INV_X1 U9520 ( .A(n7927), .ZN(n7915) );
  AND2_X1 U9521 ( .A1(n8080), .A2(n7909), .ZN(n7910) );
  NAND3_X1 U9522 ( .A1(n7912), .A2(n7920), .A3(n8049), .ZN(n7913) );
  NAND3_X1 U9523 ( .A1(n7915), .A2(n7914), .A3(n7913), .ZN(n7916) );
  NAND2_X1 U9524 ( .A1(n7917), .A2(n7916), .ZN(n7924) );
  NAND3_X1 U9525 ( .A1(n7920), .A2(n7919), .A3(n7918), .ZN(n7922) );
  NAND3_X1 U9526 ( .A1(n7922), .A2(n8018), .A3(n7921), .ZN(n7923) );
  NAND2_X1 U9527 ( .A1(n7924), .A2(n7923), .ZN(n7930) );
  AOI21_X1 U9528 ( .B1(n7927), .B2(n7926), .A(n7925), .ZN(n7928) );
  AND2_X1 U9529 ( .A1(n8213), .A2(n9894), .ZN(n7932) );
  OAI21_X1 U9530 ( .B1(n7928), .B2(n7932), .A(n8018), .ZN(n7929) );
  NAND2_X1 U9531 ( .A1(n7930), .A2(n7929), .ZN(n7936) );
  MUX2_X1 U9532 ( .A(n7933), .B(n7932), .S(n8049), .Z(n7934) );
  NOR2_X1 U9533 ( .A1(n7082), .A2(n7934), .ZN(n7935) );
  NAND2_X1 U9534 ( .A1(n7936), .A2(n7935), .ZN(n7953) );
  AND2_X1 U9535 ( .A1(n4689), .A2(n7937), .ZN(n7938) );
  AOI21_X1 U9536 ( .B1(n7953), .B2(n7938), .A(n4847), .ZN(n7939) );
  MUX2_X1 U9537 ( .A(n7940), .B(n7939), .S(n8018), .Z(n7947) );
  NAND2_X1 U9538 ( .A1(n7954), .A2(n7941), .ZN(n7945) );
  INV_X1 U9539 ( .A(n7942), .ZN(n7943) );
  NAND2_X1 U9540 ( .A1(n7943), .A2(n7946), .ZN(n7944) );
  MUX2_X1 U9541 ( .A(n7945), .B(n7944), .S(n8049), .Z(n7950) );
  AOI21_X1 U9542 ( .B1(n7947), .B2(n7946), .A(n7950), .ZN(n7963) );
  NAND2_X1 U9543 ( .A1(n7949), .A2(n7948), .ZN(n7957) );
  INV_X1 U9544 ( .A(n7950), .ZN(n7952) );
  NAND4_X1 U9545 ( .A1(n7953), .A2(n4689), .A3(n7952), .A4(n7951), .ZN(n7955)
         );
  NAND3_X1 U9546 ( .A1(n7955), .A2(n7958), .A3(n7954), .ZN(n7956) );
  MUX2_X1 U9547 ( .A(n7957), .B(n7956), .S(n8049), .Z(n7962) );
  AND2_X1 U9548 ( .A1(n7964), .A2(n7958), .ZN(n7960) );
  MUX2_X1 U9549 ( .A(n7960), .B(n7959), .S(n8049), .Z(n7961) );
  OAI21_X1 U9550 ( .B1(n7963), .B2(n7962), .A(n7961), .ZN(n7967) );
  MUX2_X1 U9551 ( .A(n7965), .B(n7964), .S(n8049), .Z(n7966) );
  NAND2_X1 U9552 ( .A1(n7967), .A2(n7966), .ZN(n7969) );
  NAND2_X1 U9553 ( .A1(n7969), .A2(n7968), .ZN(n7973) );
  MUX2_X1 U9554 ( .A(n7971), .B(n7970), .S(n8018), .Z(n7972) );
  NAND3_X1 U9555 ( .A1(n7973), .A2(n8582), .A3(n7972), .ZN(n7976) );
  MUX2_X1 U9556 ( .A(n8850), .B(n7974), .S(n8049), .Z(n7975) );
  NAND3_X1 U9557 ( .A1(n7976), .A2(n4840), .A3(n7975), .ZN(n7980) );
  NAND2_X1 U9558 ( .A1(n8820), .A2(n8049), .ZN(n7978) );
  NAND2_X1 U9559 ( .A1(n8135), .A2(n8018), .ZN(n7977) );
  MUX2_X1 U9560 ( .A(n7978), .B(n7977), .S(n8938), .Z(n7979) );
  NAND3_X1 U9561 ( .A1(n7980), .A2(n8833), .A3(n7979), .ZN(n7984) );
  MUX2_X1 U9562 ( .A(n7982), .B(n7981), .S(n8049), .Z(n7983) );
  NAND3_X1 U9563 ( .A1(n7984), .A2(n8800), .A3(n7983), .ZN(n7988) );
  AND2_X1 U9564 ( .A1(n7997), .A2(n7985), .ZN(n7986) );
  MUX2_X1 U9565 ( .A(n8788), .B(n7986), .S(n8018), .Z(n7987) );
  NAND2_X1 U9566 ( .A1(n7988), .A2(n7987), .ZN(n7998) );
  NAND2_X1 U9567 ( .A1(n7990), .A2(n7989), .ZN(n7996) );
  INV_X1 U9568 ( .A(n7996), .ZN(n7992) );
  AOI21_X1 U9569 ( .B1(n7998), .B2(n7992), .A(n7991), .ZN(n7994) );
  OAI211_X1 U9570 ( .C1(n7994), .C2(n7993), .A(n8722), .B(n7999), .ZN(n7995)
         );
  NAND3_X1 U9571 ( .A1(n7995), .A2(n8005), .A3(n8000), .ZN(n8008) );
  AOI21_X1 U9572 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n8003) );
  NAND2_X1 U9573 ( .A1(n7999), .A2(n8753), .ZN(n8002) );
  OAI211_X1 U9574 ( .C1(n8003), .C2(n8002), .A(n8001), .B(n8000), .ZN(n8004)
         );
  NAND3_X1 U9575 ( .A1(n8004), .A2(n8011), .A3(n8722), .ZN(n8006) );
  AND2_X1 U9576 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  MUX2_X1 U9577 ( .A(n8008), .B(n8007), .S(n8049), .Z(n8010) );
  OAI211_X1 U9578 ( .C1(n8011), .C2(n8049), .A(n8010), .B(n8009), .ZN(n8015)
         );
  NAND2_X1 U9579 ( .A1(n8689), .A2(n8018), .ZN(n8013) );
  NAND2_X1 U9580 ( .A1(n8726), .A2(n8049), .ZN(n8012) );
  MUX2_X1 U9581 ( .A(n8013), .B(n8012), .S(n8899), .Z(n8014) );
  NAND3_X1 U9582 ( .A1(n8015), .A2(n8687), .A3(n8014), .ZN(n8016) );
  AOI22_X1 U9583 ( .A1(n8019), .A2(n8018), .B1(n8017), .B2(n8016), .ZN(n8031)
         );
  MUX2_X1 U9584 ( .A(n8021), .B(n8020), .S(n8049), .Z(n8022) );
  NAND2_X1 U9585 ( .A1(n8638), .A2(n8022), .ZN(n8030) );
  INV_X1 U9586 ( .A(n8619), .ZN(n8026) );
  INV_X1 U9587 ( .A(n8033), .ZN(n8025) );
  INV_X1 U9588 ( .A(n8650), .ZN(n8647) );
  AOI21_X1 U9589 ( .B1(n8647), .B2(n8023), .A(n8030), .ZN(n8024) );
  AOI211_X1 U9590 ( .C1(n8026), .C2(n8880), .A(n8025), .B(n8024), .ZN(n8027)
         );
  MUX2_X1 U9591 ( .A(n8028), .B(n8027), .S(n8049), .Z(n8029) );
  OAI211_X1 U9592 ( .C1(n8031), .C2(n8030), .A(n8029), .B(n8032), .ZN(n8035)
         );
  MUX2_X1 U9593 ( .A(n8033), .B(n8032), .S(n8049), .Z(n8034) );
  NAND3_X1 U9594 ( .A1(n8035), .A2(n8600), .A3(n8034), .ZN(n8047) );
  MUX2_X1 U9595 ( .A(n8037), .B(n8036), .S(n8049), .Z(n8042) );
  INV_X1 U9596 ( .A(n8038), .ZN(n8041) );
  INV_X1 U9597 ( .A(n8039), .ZN(n8040) );
  NOR3_X1 U9598 ( .A1(n8042), .A2(n8041), .A3(n8040), .ZN(n8046) );
  MUX2_X1 U9599 ( .A(n8044), .B(n8043), .S(n8049), .Z(n8045) );
  AOI21_X1 U9600 ( .B1(n8047), .B2(n8046), .A(n8045), .ZN(n8053) );
  INV_X1 U9601 ( .A(n8048), .ZN(n8050) );
  MUX2_X1 U9602 ( .A(n8051), .B(n8050), .S(n8049), .Z(n8052) );
  OAI21_X1 U9603 ( .B1(n8053), .B2(n8052), .A(n6118), .ZN(n8054) );
  NAND4_X1 U9604 ( .A1(n8061), .A2(n4476), .A3(n8060), .A4(n8819), .ZN(n8062)
         );
  OAI211_X1 U9605 ( .C1(n8063), .C2(n8065), .A(n8062), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8064) );
  OAI21_X1 U9606 ( .B1(n8066), .B2(n8065), .A(n8064), .ZN(P2_U3244) );
  XNOR2_X1 U9607 ( .A(n8068), .B(n8067), .ZN(n8069) );
  XNOR2_X1 U9608 ( .A(n8070), .B(n8069), .ZN(n8075) );
  NOR2_X1 U9609 ( .A1(n9683), .A2(n9385), .ZN(n8073) );
  NAND2_X1 U9610 ( .A1(n9425), .A2(n9111), .ZN(n8071) );
  NAND2_X1 U9611 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9182) );
  OAI211_X1 U9612 ( .C1(n9096), .C2(n9357), .A(n8071), .B(n9182), .ZN(n8072)
         );
  AOI211_X1 U9613 ( .C1(n9533), .C2(n9115), .A(n8073), .B(n8072), .ZN(n8074)
         );
  OAI21_X1 U9614 ( .B1(n8075), .B2(n9117), .A(n8074), .ZN(P1_U3217) );
  OAI222_X1 U9615 ( .A1(n9597), .A2(n8078), .B1(P1_U3084), .B2(n8077), .C1(
        n8076), .C2(n9593), .ZN(P1_U3323) );
  AOI22_X1 U9616 ( .A1(n8202), .A2(n8082), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8079), .ZN(n8086) );
  INV_X1 U9617 ( .A(n8080), .ZN(n8081) );
  MUX2_X1 U9618 ( .A(n8082), .B(n8081), .S(n5678), .Z(n8084) );
  OAI21_X1 U9619 ( .B1(n8084), .B2(n8083), .A(n8180), .ZN(n8085) );
  OAI211_X1 U9620 ( .C1(n8166), .C2(n6696), .A(n8086), .B(n8085), .ZN(P2_U3234) );
  INV_X1 U9621 ( .A(n9589), .ZN(n8087) );
  OAI222_X1 U9622 ( .A1(n8987), .A2(n8088), .B1(P2_U3152), .B2(n6142), .C1(
        n6866), .C2(n8087), .ZN(P2_U3330) );
  INV_X1 U9623 ( .A(n8161), .ZN(n8090) );
  NOR2_X1 U9624 ( .A1(n8090), .A2(n8089), .ZN(n8094) );
  XNOR2_X1 U9625 ( .A(n8092), .B(n8091), .ZN(n8093) );
  XNOR2_X1 U9626 ( .A(n8094), .B(n8093), .ZN(n8100) );
  OAI22_X1 U9627 ( .A1(n8200), .A2(n8700), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8095), .ZN(n8098) );
  INV_X1 U9628 ( .A(n8708), .ZN(n8096) );
  OAI22_X1 U9629 ( .A1(n8096), .A2(n8166), .B1(n8167), .B2(n8591), .ZN(n8097)
         );
  AOI211_X1 U9630 ( .C1(n8899), .C2(n8202), .A(n8098), .B(n8097), .ZN(n8099)
         );
  OAI21_X1 U9631 ( .B1(n8100), .B2(n8204), .A(n8099), .ZN(P2_U3218) );
  OAI21_X1 U9632 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8104) );
  NAND2_X1 U9633 ( .A1(n8104), .A2(n8180), .ZN(n8108) );
  INV_X1 U9634 ( .A(n8776), .ZN(n8106) );
  NOR2_X1 U9635 ( .A1(n8312), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8567) );
  OAI22_X1 U9636 ( .A1(n8805), .A2(n8167), .B1(n8166), .B2(n8111), .ZN(n8105)
         );
  AOI211_X1 U9637 ( .C1(n8137), .C2(n8106), .A(n8567), .B(n8105), .ZN(n8107)
         );
  OAI211_X1 U9638 ( .C1(n8769), .C2(n8191), .A(n8108), .B(n8107), .ZN(P2_U3221) );
  XNOR2_X1 U9639 ( .A(n4394), .B(n8109), .ZN(n8115) );
  OAI22_X1 U9640 ( .A1(n8200), .A2(n8733), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8110), .ZN(n8113) );
  OAI22_X1 U9641 ( .A1(n8111), .A2(n8167), .B1(n8166), .B2(n8591), .ZN(n8112)
         );
  AOI211_X1 U9642 ( .C1(n8909), .C2(n8202), .A(n8113), .B(n8112), .ZN(n8114)
         );
  OAI21_X1 U9643 ( .B1(n8115), .B2(n8204), .A(n8114), .ZN(P2_U3225) );
  XNOR2_X1 U9644 ( .A(n8117), .B(n8116), .ZN(n8118) );
  XNOR2_X1 U9645 ( .A(n8119), .B(n8118), .ZN(n8125) );
  NAND2_X1 U9646 ( .A1(n8640), .A2(n8821), .ZN(n8121) );
  NAND2_X1 U9647 ( .A1(n8708), .A2(n8819), .ZN(n8120) );
  NAND2_X1 U9648 ( .A1(n8121), .A2(n8120), .ZN(n8669) );
  AOI22_X1 U9649 ( .A1(n8669), .A2(n8197), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8122) );
  OAI21_X1 U9650 ( .B1(n8664), .B2(n8200), .A(n8122), .ZN(n8123) );
  AOI21_X1 U9651 ( .B1(n8891), .B2(n8202), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9652 ( .B1(n8125), .B2(n8204), .A(n8124), .ZN(P2_U3227) );
  INV_X1 U9653 ( .A(n8933), .ZN(n8830) );
  NAND2_X1 U9654 ( .A1(n4390), .A2(n8126), .ZN(n8127) );
  OAI21_X1 U9655 ( .B1(n4390), .B2(n8126), .A(n8127), .ZN(n8193) );
  NOR2_X1 U9656 ( .A1(n8193), .A2(n8194), .ZN(n8192) );
  INV_X1 U9657 ( .A(n8127), .ZN(n8129) );
  NOR3_X1 U9658 ( .A1(n8192), .A2(n8129), .A3(n8128), .ZN(n8132) );
  INV_X1 U9659 ( .A(n8130), .ZN(n8131) );
  OAI21_X1 U9660 ( .B1(n8132), .B2(n8131), .A(n8180), .ZN(n8139) );
  INV_X1 U9661 ( .A(n8133), .ZN(n8828) );
  AND2_X1 U9662 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8512) );
  OAI22_X1 U9663 ( .A1(n8135), .A2(n8167), .B1(n8166), .B2(n8134), .ZN(n8136)
         );
  AOI211_X1 U9664 ( .C1(n8137), .C2(n8828), .A(n8512), .B(n8136), .ZN(n8138)
         );
  OAI211_X1 U9665 ( .C1(n8830), .C2(n8191), .A(n8139), .B(n8138), .ZN(P2_U3228) );
  XNOR2_X1 U9666 ( .A(n8141), .B(n8140), .ZN(n8145) );
  OAI22_X1 U9667 ( .A1(n8200), .A2(n8808), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8530), .ZN(n8143) );
  OAI22_X1 U9668 ( .A1(n8803), .A2(n8167), .B1(n8166), .B2(n8805), .ZN(n8142)
         );
  AOI211_X1 U9669 ( .C1(n8930), .C2(n8202), .A(n8143), .B(n8142), .ZN(n8144)
         );
  OAI21_X1 U9670 ( .B1(n8145), .B2(n8204), .A(n8144), .ZN(P2_U3230) );
  XNOR2_X1 U9671 ( .A(n8147), .B(n8146), .ZN(n8153) );
  OAI22_X1 U9672 ( .A1(n8200), .A2(n8682), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8148), .ZN(n8151) );
  OAI22_X1 U9673 ( .A1(n8726), .A2(n8167), .B1(n8166), .B2(n8149), .ZN(n8150)
         );
  AOI211_X1 U9674 ( .C1(n8894), .C2(n8202), .A(n8151), .B(n8150), .ZN(n8152)
         );
  OAI21_X1 U9675 ( .B1(n8153), .B2(n8204), .A(n8152), .ZN(P2_U3231) );
  XNOR2_X1 U9676 ( .A(n8154), .B(n8155), .ZN(n8160) );
  OAI22_X1 U9677 ( .A1(n8200), .A2(n8749), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8156), .ZN(n8158) );
  OAI22_X1 U9678 ( .A1(n8588), .A2(n8167), .B1(n8166), .B2(n8725), .ZN(n8157)
         );
  AOI211_X1 U9679 ( .C1(n8914), .C2(n8202), .A(n8158), .B(n8157), .ZN(n8159)
         );
  OAI21_X1 U9680 ( .B1(n8160), .B2(n8204), .A(n8159), .ZN(P2_U3235) );
  OAI21_X1 U9681 ( .B1(n8163), .B2(n8162), .A(n8161), .ZN(n8164) );
  NAND2_X1 U9682 ( .A1(n8164), .A2(n8180), .ZN(n8171) );
  OAI22_X1 U9683 ( .A1(n8200), .A2(n8716), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8165), .ZN(n8169) );
  OAI22_X1 U9684 ( .A1(n8725), .A2(n8167), .B1(n8166), .B2(n8726), .ZN(n8168)
         );
  AOI211_X1 U9685 ( .C1(n8904), .C2(n8202), .A(n8169), .B(n8168), .ZN(n8170)
         );
  NAND2_X1 U9686 ( .A1(n8171), .A2(n8170), .ZN(P2_U3237) );
  XNOR2_X1 U9687 ( .A(n8173), .B(n8172), .ZN(n8179) );
  AOI22_X1 U9688 ( .A1(n8175), .A2(n8822), .B1(n8174), .B2(n8793), .ZN(n8176)
         );
  NAND2_X1 U9689 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8548) );
  OAI211_X1 U9690 ( .C1(n8200), .C2(n8784), .A(n8176), .B(n8548), .ZN(n8177)
         );
  AOI21_X1 U9691 ( .B1(n8923), .B2(n8202), .A(n8177), .ZN(n8178) );
  OAI21_X1 U9692 ( .B1(n8179), .B2(n8204), .A(n8178), .ZN(P2_U3240) );
  OAI211_X1 U9693 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8190)
         );
  NAND2_X1 U9694 ( .A1(n8619), .A2(n8821), .ZN(n8185) );
  NAND2_X1 U9695 ( .A1(n8690), .A2(n8819), .ZN(n8184) );
  NAND2_X1 U9696 ( .A1(n8185), .A2(n8184), .ZN(n8652) );
  INV_X1 U9697 ( .A(n8656), .ZN(n8187) );
  OAI22_X1 U9698 ( .A1(n8187), .A2(n8200), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8186), .ZN(n8188) );
  AOI21_X1 U9699 ( .B1(n8652), .B2(n8197), .A(n8188), .ZN(n8189) );
  OAI211_X1 U9700 ( .C1(n8659), .C2(n8191), .A(n8190), .B(n8189), .ZN(P2_U3242) );
  AOI21_X1 U9701 ( .B1(n8194), .B2(n8193), .A(n8192), .ZN(n8205) );
  NAND2_X1 U9702 ( .A1(n8584), .A2(n8821), .ZN(n8196) );
  NAND2_X1 U9703 ( .A1(n8580), .A2(n8819), .ZN(n8195) );
  NAND2_X1 U9704 ( .A1(n8196), .A2(n8195), .ZN(n8854) );
  NAND2_X1 U9705 ( .A1(n8197), .A2(n8854), .ZN(n8198) );
  OAI211_X1 U9706 ( .C1(n8200), .C2(n8843), .A(n8199), .B(n8198), .ZN(n8201)
         );
  AOI21_X1 U9707 ( .B1(n8938), .B2(n8202), .A(n8201), .ZN(n8203) );
  OAI21_X1 U9708 ( .B1(n8205), .B2(n8204), .A(n8203), .ZN(P2_U3243) );
  MUX2_X1 U9709 ( .A(n8602), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8395), .Z(
        P2_U3582) );
  MUX2_X1 U9710 ( .A(n8618), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8395), .Z(
        P2_U3581) );
  MUX2_X1 U9711 ( .A(n8641), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8395), .Z(
        P2_U3580) );
  MUX2_X1 U9712 ( .A(n8619), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8395), .Z(
        P2_U3579) );
  MUX2_X1 U9713 ( .A(n8640), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8395), .Z(
        P2_U3578) );
  MUX2_X1 U9714 ( .A(n8690), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8395), .Z(
        P2_U3577) );
  MUX2_X1 U9715 ( .A(n8708), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8395), .Z(
        P2_U3576) );
  MUX2_X1 U9716 ( .A(n8689), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8395), .Z(
        P2_U3575) );
  MUX2_X1 U9717 ( .A(n8740), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8395), .Z(
        P2_U3574) );
  MUX2_X1 U9718 ( .A(n8756), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8395), .Z(
        P2_U3573) );
  MUX2_X1 U9719 ( .A(n8766), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8395), .Z(
        P2_U3572) );
  MUX2_X1 U9720 ( .A(n8793), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8395), .Z(
        P2_U3571) );
  MUX2_X1 U9721 ( .A(n8765), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8395), .Z(
        P2_U3570) );
  MUX2_X1 U9722 ( .A(n8822), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8395), .Z(
        P2_U3569) );
  MUX2_X1 U9723 ( .A(n8584), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8395), .Z(
        P2_U3568) );
  MUX2_X1 U9724 ( .A(n8820), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8395), .Z(
        P2_U3567) );
  MUX2_X1 U9725 ( .A(n8580), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8395), .Z(
        P2_U3566) );
  MUX2_X1 U9726 ( .A(n8206), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8395), .Z(
        P2_U3565) );
  MUX2_X1 U9727 ( .A(n8207), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8395), .Z(
        P2_U3564) );
  MUX2_X1 U9728 ( .A(n8208), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8395), .Z(
        P2_U3563) );
  MUX2_X1 U9729 ( .A(n8209), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8395), .Z(
        P2_U3562) );
  MUX2_X1 U9730 ( .A(n8210), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8395), .Z(
        P2_U3561) );
  MUX2_X1 U9731 ( .A(n8211), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8395), .Z(
        P2_U3560) );
  MUX2_X1 U9732 ( .A(n8212), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8395), .Z(
        P2_U3559) );
  MUX2_X1 U9733 ( .A(n8213), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8395), .Z(n8390)
         );
  AOI22_X1 U9734 ( .A1(n7412), .A2(keyinput101), .B1(n8215), .B2(keyinput79), 
        .ZN(n8214) );
  OAI221_X1 U9735 ( .B1(n7412), .B2(keyinput101), .C1(n8215), .C2(keyinput79), 
        .A(n8214), .ZN(n8223) );
  XNOR2_X1 U9736 ( .A(keyinput97), .B(n5287), .ZN(n8222) );
  INV_X1 U9737 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9731) );
  XNOR2_X1 U9738 ( .A(keyinput112), .B(n9731), .ZN(n8221) );
  XNOR2_X1 U9739 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput83), .ZN(n8219) );
  XNOR2_X1 U9740 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput75), .ZN(n8218) );
  XNOR2_X1 U9741 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput90), .ZN(n8217) );
  XNOR2_X1 U9742 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput120), .ZN(n8216) );
  NAND4_X1 U9743 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n8220)
         );
  NOR4_X1 U9744 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n8259)
         );
  AOI22_X1 U9745 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput99), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput74), .ZN(n8224) );
  OAI221_X1 U9746 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput99), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput74), .A(n8224), .ZN(n8232) );
  AOI22_X1 U9747 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(keyinput69), .B1(SI_21_), 
        .B2(keyinput68), .ZN(n8225) );
  OAI221_X1 U9748 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(keyinput69), .C1(SI_21_), 
        .C2(keyinput68), .A(n8225), .ZN(n8231) );
  INV_X1 U9749 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9038) );
  AOI22_X1 U9750 ( .A1(n9038), .A2(keyinput103), .B1(keyinput108), .B2(n8227), 
        .ZN(n8226) );
  OAI221_X1 U9751 ( .B1(n9038), .B2(keyinput103), .C1(n8227), .C2(keyinput108), 
        .A(n8226), .ZN(n8230) );
  AOI22_X1 U9752 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput115), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(keyinput104), .ZN(n8228) );
  OAI221_X1 U9753 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput115), .C1(
        P1_DATAO_REG_18__SCAN_IN), .C2(keyinput104), .A(n8228), .ZN(n8229) );
  NOR4_X1 U9754 ( .A1(n8232), .A2(n8231), .A3(n8230), .A4(n8229), .ZN(n8258)
         );
  INV_X1 U9755 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9709) );
  AOI22_X1 U9756 ( .A1(n9709), .A2(keyinput72), .B1(keyinput119), .B2(n5705), 
        .ZN(n8233) );
  OAI221_X1 U9757 ( .B1(n9709), .B2(keyinput72), .C1(n5705), .C2(keyinput119), 
        .A(n8233), .ZN(n8244) );
  INV_X1 U9758 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8235) );
  AOI22_X1 U9759 ( .A1(n8314), .A2(keyinput93), .B1(n8235), .B2(keyinput80), 
        .ZN(n8234) );
  OAI221_X1 U9760 ( .B1(n8314), .B2(keyinput93), .C1(n8235), .C2(keyinput80), 
        .A(n8234), .ZN(n8243) );
  AOI22_X1 U9761 ( .A1(n8238), .A2(keyinput107), .B1(n8237), .B2(keyinput77), 
        .ZN(n8236) );
  OAI221_X1 U9762 ( .B1(n8238), .B2(keyinput107), .C1(n8237), .C2(keyinput77), 
        .A(n8236), .ZN(n8242) );
  XNOR2_X1 U9763 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput95), .ZN(n8240) );
  XNOR2_X1 U9764 ( .A(SI_2_), .B(keyinput121), .ZN(n8239) );
  NAND2_X1 U9765 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NOR4_X1 U9766 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8257)
         );
  INV_X1 U9767 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9738) );
  AOI22_X1 U9768 ( .A1(n5116), .A2(keyinput110), .B1(n9738), .B2(keyinput124), 
        .ZN(n8245) );
  OAI221_X1 U9769 ( .B1(n5116), .B2(keyinput110), .C1(n9738), .C2(keyinput124), 
        .A(n8245), .ZN(n8255) );
  INV_X1 U9770 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U9771 ( .A1(n5862), .A2(keyinput88), .B1(n9708), .B2(keyinput76), 
        .ZN(n8246) );
  OAI221_X1 U9772 ( .B1(n5862), .B2(keyinput88), .C1(n9708), .C2(keyinput76), 
        .A(n8246), .ZN(n8254) );
  INV_X1 U9773 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8249) );
  INV_X1 U9774 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8248) );
  AOI22_X1 U9775 ( .A1(n8249), .A2(keyinput122), .B1(keyinput71), .B2(n8248), 
        .ZN(n8247) );
  OAI221_X1 U9776 ( .B1(n8249), .B2(keyinput122), .C1(n8248), .C2(keyinput71), 
        .A(n8247), .ZN(n8253) );
  AOI22_X1 U9777 ( .A1(n8557), .A2(keyinput116), .B1(n8251), .B2(keyinput100), 
        .ZN(n8250) );
  OAI221_X1 U9778 ( .B1(n8557), .B2(keyinput116), .C1(n8251), .C2(keyinput100), 
        .A(n8250), .ZN(n8252) );
  NOR4_X1 U9779 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n8256)
         );
  NAND4_X1 U9780 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n8323)
         );
  AOI22_X1 U9781 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(keyinput73), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput117), .ZN(n8260) );
  OAI221_X1 U9782 ( .B1(P1_DATAO_REG_6__SCAN_IN), .B2(keyinput73), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput117), .A(n8260), .ZN(n8267) );
  AOI22_X1 U9783 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput113), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput114), .ZN(n8261) );
  OAI221_X1 U9784 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput113), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput114), .A(n8261), .ZN(n8266) );
  AOI22_X1 U9785 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput89), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput82), .ZN(n8262) );
  OAI221_X1 U9786 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput89), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput82), .A(n8262), .ZN(n8265) );
  AOI22_X1 U9787 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(keyinput70), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput127), .ZN(n8263) );
  OAI221_X1 U9788 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(keyinput70), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput127), .A(n8263), .ZN(n8264) );
  NOR4_X1 U9789 ( .A1(n8267), .A2(n8266), .A3(n8265), .A4(n8264), .ZN(n8295)
         );
  AOI22_X1 U9790 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(keyinput67), .B1(
        P2_IR_REG_12__SCAN_IN), .B2(keyinput102), .ZN(n8268) );
  OAI221_X1 U9791 ( .B1(P2_IR_REG_5__SCAN_IN), .B2(keyinput67), .C1(
        P2_IR_REG_12__SCAN_IN), .C2(keyinput102), .A(n8268), .ZN(n8275) );
  AOI22_X1 U9792 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput118), .B1(
        P1_REG1_REG_11__SCAN_IN), .B2(keyinput125), .ZN(n8269) );
  OAI221_X1 U9793 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput118), .C1(
        P1_REG1_REG_11__SCAN_IN), .C2(keyinput125), .A(n8269), .ZN(n8274) );
  AOI22_X1 U9794 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(keyinput96), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput78), .ZN(n8270) );
  OAI221_X1 U9795 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(keyinput96), .C1(
        P1_D_REG_28__SCAN_IN), .C2(keyinput78), .A(n8270), .ZN(n8273) );
  AOI22_X1 U9796 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(keyinput66), .B1(SI_7_), 
        .B2(keyinput87), .ZN(n8271) );
  OAI221_X1 U9797 ( .B1(P2_REG0_REG_20__SCAN_IN), .B2(keyinput66), .C1(SI_7_), 
        .C2(keyinput87), .A(n8271), .ZN(n8272) );
  NOR4_X1 U9798 ( .A1(n8275), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n8294)
         );
  AOI22_X1 U9799 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput106), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput111), .ZN(n8276) );
  OAI221_X1 U9800 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput106), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput111), .A(n8276), .ZN(n8283) );
  AOI22_X1 U9801 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput94), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput86), .ZN(n8277) );
  OAI221_X1 U9802 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput94), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput86), .A(n8277), .ZN(n8282) );
  AOI22_X1 U9803 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(keyinput98), .B1(
        P1_REG1_REG_27__SCAN_IN), .B2(keyinput65), .ZN(n8278) );
  OAI221_X1 U9804 ( .B1(P1_REG0_REG_20__SCAN_IN), .B2(keyinput98), .C1(
        P1_REG1_REG_27__SCAN_IN), .C2(keyinput65), .A(n8278), .ZN(n8281) );
  AOI22_X1 U9805 ( .A1(P1_REG1_REG_19__SCAN_IN), .A2(keyinput109), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput81), .ZN(n8279) );
  OAI221_X1 U9806 ( .B1(P1_REG1_REG_19__SCAN_IN), .B2(keyinput109), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput81), .A(n8279), .ZN(n8280) );
  NOR4_X1 U9807 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n8293)
         );
  AOI22_X1 U9808 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput85), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput84), .ZN(n8284) );
  OAI221_X1 U9809 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput85), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput84), .A(n8284), .ZN(n8291) );
  AOI22_X1 U9810 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(keyinput64), .B1(
        P1_REG0_REG_21__SCAN_IN), .B2(keyinput126), .ZN(n8285) );
  OAI221_X1 U9811 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(keyinput64), .C1(
        P1_REG0_REG_21__SCAN_IN), .C2(keyinput126), .A(n8285), .ZN(n8290) );
  AOI22_X1 U9812 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(keyinput105), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput123), .ZN(n8286) );
  OAI221_X1 U9813 ( .B1(P1_DATAO_REG_1__SCAN_IN), .B2(keyinput105), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput123), .A(n8286), .ZN(n8289) );
  AOI22_X1 U9814 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(keyinput91), .B1(
        P2_REG0_REG_0__SCAN_IN), .B2(keyinput92), .ZN(n8287) );
  OAI221_X1 U9815 ( .B1(P1_REG1_REG_31__SCAN_IN), .B2(keyinput91), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput92), .A(n8287), .ZN(n8288) );
  NOR4_X1 U9816 ( .A1(n8291), .A2(n8290), .A3(n8289), .A4(n8288), .ZN(n8292)
         );
  NAND4_X1 U9817 ( .A1(n8295), .A2(n8294), .A3(n8293), .A4(n8292), .ZN(n8322)
         );
  AOI22_X1 U9818 ( .A1(n8298), .A2(keyinput10), .B1(n8297), .B2(keyinput4), 
        .ZN(n8296) );
  OAI221_X1 U9819 ( .B1(n8298), .B2(keyinput10), .C1(n8297), .C2(keyinput4), 
        .A(n8296), .ZN(n8308) );
  AOI22_X1 U9820 ( .A1(n4578), .A2(keyinput17), .B1(keyinput2), .B2(n8300), 
        .ZN(n8299) );
  OAI221_X1 U9821 ( .B1(n4578), .B2(keyinput17), .C1(n8300), .C2(keyinput2), 
        .A(n8299), .ZN(n8307) );
  INV_X1 U9822 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8302) );
  INV_X1 U9823 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U9824 ( .A1(n8302), .A2(keyinput32), .B1(n9840), .B2(keyinput54), 
        .ZN(n8301) );
  OAI221_X1 U9825 ( .B1(n8302), .B2(keyinput32), .C1(n9840), .C2(keyinput54), 
        .A(n8301), .ZN(n8306) );
  AOI22_X1 U9826 ( .A1(n8304), .A2(keyinput22), .B1(keyinput37), .B2(n7412), 
        .ZN(n8303) );
  OAI221_X1 U9827 ( .B1(n8304), .B2(keyinput22), .C1(n7412), .C2(keyinput37), 
        .A(n8303), .ZN(n8305) );
  NOR4_X1 U9828 ( .A1(n8308), .A2(n8307), .A3(n8306), .A4(n8305), .ZN(n8321)
         );
  AOI22_X1 U9829 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput31), .B1(n5116), 
        .B2(keyinput46), .ZN(n8309) );
  OAI221_X1 U9830 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput31), .C1(n5116), 
        .C2(keyinput46), .A(n8309), .ZN(n8319) );
  AOI22_X1 U9831 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(keyinput24), .B1(
        P2_REG1_REG_18__SCAN_IN), .B2(keyinput52), .ZN(n8310) );
  OAI221_X1 U9832 ( .B1(P2_REG0_REG_12__SCAN_IN), .B2(keyinput24), .C1(
        P2_REG1_REG_18__SCAN_IN), .C2(keyinput52), .A(n8310), .ZN(n8318) );
  AOI22_X1 U9833 ( .A1(n8312), .A2(keyinput56), .B1(keyinput55), .B2(n5705), 
        .ZN(n8311) );
  OAI221_X1 U9834 ( .B1(n8312), .B2(keyinput56), .C1(n5705), .C2(keyinput55), 
        .A(n8311), .ZN(n8317) );
  AOI22_X1 U9835 ( .A1(n8315), .A2(keyinput53), .B1(n8314), .B2(keyinput29), 
        .ZN(n8313) );
  OAI221_X1 U9836 ( .B1(n8315), .B2(keyinput53), .C1(n8314), .C2(keyinput29), 
        .A(n8313), .ZN(n8316) );
  NOR4_X1 U9837 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(n8320)
         );
  OAI211_X1 U9838 ( .C1(n8323), .C2(n8322), .A(n8321), .B(n8320), .ZN(n8388)
         );
  INV_X1 U9839 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8326) );
  OAI22_X1 U9840 ( .A1(n8326), .A2(keyinput1), .B1(n8325), .B2(keyinput45), 
        .ZN(n8324) );
  AOI221_X1 U9841 ( .B1(n8326), .B2(keyinput1), .C1(keyinput45), .C2(n8325), 
        .A(n8324), .ZN(n8332) );
  XNOR2_X1 U9842 ( .A(P2_REG1_REG_15__SCAN_IN), .B(keyinput44), .ZN(n8328) );
  XNOR2_X1 U9843 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput59), .ZN(n8327) );
  AND2_X1 U9844 ( .A1(n8328), .A2(n8327), .ZN(n8331) );
  XNOR2_X1 U9845 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput11), .ZN(n8330) );
  XNOR2_X1 U9846 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput58), .ZN(n8329) );
  AND4_X1 U9847 ( .A1(n8332), .A2(n8331), .A3(n8330), .A4(n8329), .ZN(n8376)
         );
  INV_X1 U9848 ( .A(P2_WR_REG_SCAN_IN), .ZN(n8334) );
  OAI22_X1 U9849 ( .A1(n9708), .A2(keyinput12), .B1(n8334), .B2(keyinput25), 
        .ZN(n8333) );
  AOI221_X1 U9850 ( .B1(n9708), .B2(keyinput12), .C1(keyinput25), .C2(n8334), 
        .A(n8333), .ZN(n8375) );
  INV_X1 U9851 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8336) );
  OAI22_X1 U9852 ( .A1(n8336), .A2(keyinput62), .B1(n5720), .B2(keyinput21), 
        .ZN(n8335) );
  AOI221_X1 U9853 ( .B1(n8336), .B2(keyinput62), .C1(keyinput21), .C2(n5720), 
        .A(n8335), .ZN(n8374) );
  AOI22_X1 U9854 ( .A1(SI_2_), .A2(keyinput57), .B1(SI_19_), .B2(keyinput13), 
        .ZN(n8337) );
  OAI221_X1 U9855 ( .B1(SI_2_), .B2(keyinput57), .C1(SI_19_), .C2(keyinput13), 
        .A(n8337), .ZN(n8344) );
  AOI22_X1 U9856 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(keyinput0), .B1(
        P2_ADDR_REG_13__SCAN_IN), .B2(keyinput6), .ZN(n8338) );
  OAI221_X1 U9857 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(keyinput0), .C1(
        P2_ADDR_REG_13__SCAN_IN), .C2(keyinput6), .A(n8338), .ZN(n8343) );
  AOI22_X1 U9858 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput35), .B1(
        P1_REG2_REG_19__SCAN_IN), .B2(keyinput30), .ZN(n8339) );
  OAI221_X1 U9859 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput35), .C1(
        P1_REG2_REG_19__SCAN_IN), .C2(keyinput30), .A(n8339), .ZN(n8342) );
  AOI22_X1 U9860 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput19), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput50), .ZN(n8340) );
  OAI221_X1 U9861 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput19), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput50), .A(n8340), .ZN(n8341) );
  NOR4_X1 U9862 ( .A1(n8344), .A2(n8343), .A3(n8342), .A4(n8341), .ZN(n8372)
         );
  AOI22_X1 U9863 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput7), .B1(
        P2_REG0_REG_0__SCAN_IN), .B2(keyinput28), .ZN(n8345) );
  OAI221_X1 U9864 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput7), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput28), .A(n8345), .ZN(n8352) );
  AOI22_X1 U9865 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput51), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(keyinput9), .ZN(n8346) );
  OAI221_X1 U9866 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput51), .C1(
        P1_DATAO_REG_6__SCAN_IN), .C2(keyinput9), .A(n8346), .ZN(n8351) );
  AOI22_X1 U9867 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput49), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput14), .ZN(n8347) );
  OAI221_X1 U9868 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput49), .C1(
        P1_D_REG_28__SCAN_IN), .C2(keyinput14), .A(n8347), .ZN(n8350) );
  AOI22_X1 U9869 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(keyinput38), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput26), .ZN(n8348) );
  OAI221_X1 U9870 ( .B1(P2_IR_REG_12__SCAN_IN), .B2(keyinput38), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput26), .A(n8348), .ZN(n8349) );
  NOR4_X1 U9871 ( .A1(n8352), .A2(n8351), .A3(n8350), .A4(n8349), .ZN(n8371)
         );
  AOI22_X1 U9872 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput42), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput16), .ZN(n8353) );
  OAI221_X1 U9873 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput42), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput16), .A(n8353), .ZN(n8360) );
  AOI22_X1 U9874 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(keyinput27), .B1(SI_28_), 
        .B2(keyinput43), .ZN(n8354) );
  OAI221_X1 U9875 ( .B1(P1_REG1_REG_31__SCAN_IN), .B2(keyinput27), .C1(SI_28_), 
        .C2(keyinput43), .A(n8354), .ZN(n8359) );
  AOI22_X1 U9876 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput61), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput47), .ZN(n8355) );
  OAI221_X1 U9877 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput61), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput47), .A(n8355), .ZN(n8358) );
  AOI22_X1 U9878 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(keyinput34), .B1(
        P1_REG3_REG_16__SCAN_IN), .B2(keyinput39), .ZN(n8356) );
  OAI221_X1 U9879 ( .B1(P1_REG0_REG_20__SCAN_IN), .B2(keyinput34), .C1(
        P1_REG3_REG_16__SCAN_IN), .C2(keyinput39), .A(n8356), .ZN(n8357) );
  NOR4_X1 U9880 ( .A1(n8360), .A2(n8359), .A3(n8358), .A4(n8357), .ZN(n8370)
         );
  AOI22_X1 U9881 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput20), .B1(SI_16_), 
        .B2(keyinput36), .ZN(n8361) );
  OAI221_X1 U9882 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput20), .C1(SI_16_), 
        .C2(keyinput36), .A(n8361), .ZN(n8368) );
  AOI22_X1 U9883 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput60), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput15), .ZN(n8362) );
  OAI221_X1 U9884 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput60), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput15), .A(n8362), .ZN(n8367) );
  AOI22_X1 U9885 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput18), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(keyinput41), .ZN(n8363) );
  OAI221_X1 U9886 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput18), .C1(
        P1_DATAO_REG_1__SCAN_IN), .C2(keyinput41), .A(n8363), .ZN(n8366) );
  AOI22_X1 U9887 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(keyinput5), .B1(
        P1_REG0_REG_3__SCAN_IN), .B2(keyinput48), .ZN(n8364) );
  OAI221_X1 U9888 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(keyinput5), .C1(
        P1_REG0_REG_3__SCAN_IN), .C2(keyinput48), .A(n8364), .ZN(n8365) );
  NOR4_X1 U9889 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8369)
         );
  AND4_X1 U9890 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n8373)
         );
  NAND4_X1 U9891 ( .A1(n8376), .A2(n8375), .A3(n8374), .A4(n8373), .ZN(n8387)
         );
  OAI22_X1 U9892 ( .A1(n9709), .A2(keyinput8), .B1(n5287), .B2(keyinput33), 
        .ZN(n8377) );
  AOI221_X1 U9893 ( .B1(n9709), .B2(keyinput8), .C1(keyinput33), .C2(n5287), 
        .A(n8377), .ZN(n8385) );
  INV_X1 U9894 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8379) );
  OAI22_X1 U9895 ( .A1(n8379), .A2(keyinput3), .B1(n9600), .B2(keyinput63), 
        .ZN(n8378) );
  AOI221_X1 U9896 ( .B1(n8379), .B2(keyinput3), .C1(keyinput63), .C2(n9600), 
        .A(n8378), .ZN(n8384) );
  OAI22_X1 U9897 ( .A1(n8382), .A2(keyinput40), .B1(n8381), .B2(keyinput23), 
        .ZN(n8380) );
  AOI221_X1 U9898 ( .B1(n8382), .B2(keyinput40), .C1(keyinput23), .C2(n8381), 
        .A(n8380), .ZN(n8383) );
  NAND3_X1 U9899 ( .A1(n8385), .A2(n8384), .A3(n8383), .ZN(n8386) );
  NOR3_X1 U9900 ( .A1(n8388), .A2(n8387), .A3(n8386), .ZN(n8389) );
  XOR2_X1 U9901 ( .A(n8390), .B(n8389), .Z(P2_U3558) );
  MUX2_X1 U9902 ( .A(n8391), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8395), .Z(
        P2_U3557) );
  MUX2_X1 U9903 ( .A(n8392), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8395), .Z(
        P2_U3556) );
  MUX2_X1 U9904 ( .A(n8393), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8395), .Z(
        P2_U3555) );
  MUX2_X1 U9905 ( .A(n8394), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8395), .Z(
        P2_U3554) );
  MUX2_X1 U9906 ( .A(n6697), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8395), .Z(
        P2_U3553) );
  MUX2_X1 U9907 ( .A(n6502), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8395), .Z(
        P2_U3552) );
  OAI211_X1 U9908 ( .C1(n8398), .C2(n8397), .A(n9803), .B(n8396), .ZN(n8409)
         );
  NOR2_X1 U9909 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8399), .ZN(n8400) );
  AOI21_X1 U9910 ( .B1(n9809), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8400), .ZN(
        n8408) );
  NAND2_X1 U9911 ( .A1(n9620), .A2(n8401), .ZN(n8407) );
  AOI21_X1 U9912 ( .B1(n8404), .B2(n8403), .A(n8402), .ZN(n8405) );
  NAND2_X1 U9913 ( .A1(n9804), .A2(n8405), .ZN(n8406) );
  NAND4_X1 U9914 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(
        P2_U3248) );
  OAI211_X1 U9915 ( .C1(n8412), .C2(n8411), .A(n9803), .B(n8410), .ZN(n8422)
         );
  AND2_X1 U9916 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8413) );
  AOI21_X1 U9917 ( .B1(n9809), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8413), .ZN(
        n8421) );
  NAND2_X1 U9918 ( .A1(n9620), .A2(n8414), .ZN(n8420) );
  AOI21_X1 U9919 ( .B1(n8417), .B2(n8416), .A(n8415), .ZN(n8418) );
  NAND2_X1 U9920 ( .A1(n9804), .A2(n8418), .ZN(n8419) );
  NAND4_X1 U9921 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(
        P2_U3249) );
  OAI211_X1 U9922 ( .C1(n8425), .C2(n8424), .A(n9803), .B(n8423), .ZN(n8436)
         );
  NOR2_X1 U9923 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8426), .ZN(n8427) );
  AOI21_X1 U9924 ( .B1(n9809), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8427), .ZN(
        n8435) );
  NAND2_X1 U9925 ( .A1(n9620), .A2(n8428), .ZN(n8434) );
  AOI21_X1 U9926 ( .B1(n8431), .B2(n8430), .A(n8429), .ZN(n8432) );
  NAND2_X1 U9927 ( .A1(n9804), .A2(n8432), .ZN(n8433) );
  NAND4_X1 U9928 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(
        P2_U3250) );
  OAI211_X1 U9929 ( .C1(n8439), .C2(n8438), .A(n9803), .B(n8437), .ZN(n8449)
         );
  INV_X1 U9930 ( .A(n8440), .ZN(n8441) );
  AOI21_X1 U9931 ( .B1(n9809), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8441), .ZN(
        n8448) );
  NAND2_X1 U9932 ( .A1(n9620), .A2(n8442), .ZN(n8447) );
  OAI211_X1 U9933 ( .C1(n8445), .C2(n8444), .A(n9804), .B(n8443), .ZN(n8446)
         );
  NAND4_X1 U9934 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(
        P2_U3251) );
  OAI211_X1 U9935 ( .C1(n8452), .C2(n8451), .A(n9803), .B(n8450), .ZN(n8462)
         );
  AOI21_X1 U9936 ( .B1(n9809), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8453), .ZN(
        n8461) );
  NAND2_X1 U9937 ( .A1(n9620), .A2(n8454), .ZN(n8460) );
  NAND2_X1 U9938 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  NAND3_X1 U9939 ( .A1(n9804), .A2(n8458), .A3(n8457), .ZN(n8459) );
  NAND4_X1 U9940 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(
        P2_U3252) );
  OAI211_X1 U9941 ( .C1(n8465), .C2(n8464), .A(n9803), .B(n8463), .ZN(n8474)
         );
  NOR2_X1 U9942 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8466), .ZN(n8467) );
  AOI21_X1 U9943 ( .B1(n9809), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8467), .ZN(
        n8473) );
  NAND2_X1 U9944 ( .A1(n9620), .A2(n4539), .ZN(n8472) );
  OAI211_X1 U9945 ( .C1(n8470), .C2(n8469), .A(n9804), .B(n8468), .ZN(n8471)
         );
  NAND4_X1 U9946 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(
        P2_U3253) );
  OAI211_X1 U9947 ( .C1(n8477), .C2(n8476), .A(n9803), .B(n8475), .ZN(n8487)
         );
  AOI21_X1 U9948 ( .B1(n9809), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8478), .ZN(
        n8486) );
  NAND2_X1 U9949 ( .A1(n9620), .A2(n8479), .ZN(n8485) );
  INV_X1 U9950 ( .A(n8480), .ZN(n8481) );
  OAI211_X1 U9951 ( .C1(n8483), .C2(n8482), .A(n9804), .B(n8481), .ZN(n8484)
         );
  NAND4_X1 U9952 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(
        P2_U3254) );
  MUX2_X1 U9953 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8488), .S(n8494), .Z(n8490)
         );
  OAI211_X1 U9954 ( .C1(n8491), .C2(n8490), .A(n9803), .B(n8489), .ZN(n8503)
         );
  INV_X1 U9955 ( .A(n8492), .ZN(n8493) );
  AOI21_X1 U9956 ( .B1(n9809), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8493), .ZN(
        n8502) );
  NAND2_X1 U9957 ( .A1(n9620), .A2(n8494), .ZN(n8501) );
  NAND2_X1 U9958 ( .A1(n8496), .A2(n8495), .ZN(n8497) );
  NAND2_X1 U9959 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U9960 ( .A1(n9804), .A2(n8499), .ZN(n8500) );
  NAND4_X1 U9961 ( .A1(n8503), .A2(n8502), .A3(n8501), .A4(n8500), .ZN(
        P2_U3257) );
  NOR2_X1 U9962 ( .A1(n8505), .A2(n8504), .ZN(n8507) );
  NOR2_X1 U9963 ( .A1(n8507), .A2(n8506), .ZN(n8510) );
  XNOR2_X1 U9964 ( .A(n8532), .B(n8508), .ZN(n8509) );
  OAI21_X1 U9965 ( .B1(n8510), .B2(n8509), .A(n8531), .ZN(n8511) );
  NAND2_X1 U9966 ( .A1(n8511), .A2(n9804), .ZN(n8524) );
  AOI21_X1 U9967 ( .B1(n9809), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8512), .ZN(
        n8523) );
  NOR2_X1 U9968 ( .A1(n8514), .A2(n8513), .ZN(n8516) );
  NOR2_X1 U9969 ( .A1(n8516), .A2(n8515), .ZN(n8520) );
  NAND2_X1 U9970 ( .A1(n8532), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8526) );
  INV_X1 U9971 ( .A(n8526), .ZN(n8517) );
  AOI21_X1 U9972 ( .B1(n5622), .B2(n8518), .A(n8517), .ZN(n8519) );
  NAND2_X1 U9973 ( .A1(n8519), .A2(n8520), .ZN(n8525) );
  OAI211_X1 U9974 ( .C1(n8520), .C2(n8519), .A(n9803), .B(n8525), .ZN(n8522)
         );
  NAND2_X1 U9975 ( .A1(n9620), .A2(n8532), .ZN(n8521) );
  NAND4_X1 U9976 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(
        P2_U3261) );
  NAND2_X1 U9977 ( .A1(n8526), .A2(n8525), .ZN(n8529) );
  NAND2_X1 U9978 ( .A1(n8546), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8541) );
  INV_X1 U9979 ( .A(n8541), .ZN(n8527) );
  AOI21_X1 U9980 ( .B1(n8809), .B2(n8539), .A(n8527), .ZN(n8528) );
  NAND2_X1 U9981 ( .A1(n8528), .A2(n8529), .ZN(n8540) );
  OAI211_X1 U9982 ( .C1(n8529), .C2(n8528), .A(n9803), .B(n8540), .ZN(n8538)
         );
  NOR2_X1 U9983 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8530), .ZN(n8536) );
  XNOR2_X1 U9984 ( .A(n8546), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8533) );
  NOR2_X1 U9985 ( .A1(n8533), .A2(n8534), .ZN(n8545) );
  AOI211_X1 U9986 ( .C1(n8534), .C2(n8533), .A(n8545), .B(n9614), .ZN(n8535)
         );
  AOI211_X1 U9987 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9809), .A(n8536), .B(
        n8535), .ZN(n8537) );
  OAI211_X1 U9988 ( .C1(n9806), .C2(n8539), .A(n8538), .B(n8537), .ZN(P2_U3262) );
  NAND2_X1 U9989 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NOR2_X1 U9990 ( .A1(n8542), .A2(n8551), .ZN(n8555) );
  AOI21_X1 U9991 ( .B1(n8542), .B2(n8551), .A(n8555), .ZN(n8543) );
  INV_X1 U9992 ( .A(n8543), .ZN(n8544) );
  NOR2_X1 U9993 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8544), .ZN(n8554) );
  AOI21_X1 U9994 ( .B1(n8544), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8554), .ZN(
        n8553) );
  XOR2_X1 U9995 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8551), .Z(n8560) );
  AOI21_X1 U9996 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8546), .A(n8545), .ZN(
        n8559) );
  XNOR2_X1 U9997 ( .A(n8560), .B(n8559), .ZN(n8547) );
  NAND2_X1 U9998 ( .A1(n9804), .A2(n8547), .ZN(n8549) );
  OAI211_X1 U9999 ( .C1(n9602), .C2(n9978), .A(n8549), .B(n8548), .ZN(n8550)
         );
  AOI21_X1 U10000 ( .B1(n8551), .B2(n9620), .A(n8550), .ZN(n8552) );
  OAI21_X1 U10001 ( .B1(n8553), .B2(n9807), .A(n8552), .ZN(P2_U3263) );
  NOR2_X1 U10002 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  XOR2_X1 U10003 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8556), .Z(n8563) );
  AOI22_X1 U10004 ( .A1(n8560), .A2(n8559), .B1(n8558), .B2(n8557), .ZN(n8561)
         );
  XNOR2_X1 U10005 ( .A(n8561), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8565) );
  INV_X1 U10006 ( .A(n8565), .ZN(n8562) );
  NOR2_X1 U10007 ( .A1(n8563), .A2(n9807), .ZN(n8564) );
  AOI211_X1 U10008 ( .C1(n9804), .C2(n8565), .A(n9620), .B(n8564), .ZN(n8566)
         );
  INV_X1 U10009 ( .A(n8567), .ZN(n8568) );
  OAI211_X1 U10010 ( .C1(n9602), .C2(n8570), .A(n8569), .B(n8568), .ZN(
        P2_U3264) );
  NAND2_X1 U10011 ( .A1(n8842), .A2(n8830), .ZN(n8825) );
  INV_X1 U10012 ( .A(n8914), .ZN(n8752) );
  INV_X1 U10013 ( .A(n8899), .ZN(n8703) );
  INV_X1 U10014 ( .A(n8891), .ZN(n8672) );
  NAND2_X1 U10015 ( .A1(n8681), .A2(n8672), .ZN(n8655) );
  XNOR2_X1 U10016 ( .A(n8571), .B(n8575), .ZN(n8860) );
  NAND2_X1 U10017 ( .A1(n8860), .A2(n8858), .ZN(n8574) );
  AOI21_X1 U10018 ( .B1(n4476), .B2(P2_B_REG_SCAN_IN), .A(n8806), .ZN(n8603)
         );
  NAND2_X1 U10019 ( .A1(n8572), .A2(n8603), .ZN(n8865) );
  NOR2_X1 U10020 ( .A1(n8846), .A2(n8865), .ZN(n8577) );
  AOI21_X1 U10021 ( .B1(n9837), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8577), .ZN(
        n8573) );
  OAI211_X1 U10022 ( .C1(n8862), .C2(n8848), .A(n8574), .B(n8573), .ZN(
        P2_U3265) );
  INV_X1 U10023 ( .A(n8575), .ZN(n8864) );
  NAND2_X1 U10024 ( .A1(n4332), .A2(n8576), .ZN(n8863) );
  NAND3_X1 U10025 ( .A1(n8864), .A2(n8858), .A3(n8863), .ZN(n8579) );
  AOI21_X1 U10026 ( .B1(n8846), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8577), .ZN(
        n8578) );
  OAI211_X1 U10027 ( .C1(n8867), .C2(n8848), .A(n8579), .B(n8578), .ZN(
        P2_U3266) );
  OAI22_X1 U10028 ( .A1(n8583), .A2(n8582), .B1(n8581), .B2(n8580), .ZN(n8840)
         );
  NAND2_X1 U10029 ( .A1(n8923), .A2(n8765), .ZN(n8587) );
  INV_X1 U10030 ( .A(n8923), .ZN(n8787) );
  INV_X1 U10031 ( .A(n8909), .ZN(n8736) );
  OAI21_X1 U10032 ( .B1(n8756), .B2(n8909), .A(n8590), .ZN(n8713) );
  INV_X1 U10033 ( .A(n8904), .ZN(n8719) );
  AOI22_X1 U10034 ( .A1(n8648), .A2(n8650), .B1(n8659), .B2(n8594), .ZN(n8629)
         );
  OAI22_X1 U10035 ( .A1(n8629), .A2(n8638), .B1(n8880), .B2(n8619), .ZN(n8615)
         );
  NAND2_X1 U10036 ( .A1(n8615), .A2(n8616), .ZN(n8597) );
  NAND2_X1 U10037 ( .A1(n8597), .A2(n8596), .ZN(n8599) );
  INV_X1 U10038 ( .A(n8600), .ZN(n8598) );
  XNOR2_X1 U10039 ( .A(n8599), .B(n8598), .ZN(n8868) );
  INV_X1 U10040 ( .A(n8868), .ZN(n8613) );
  XNOR2_X1 U10041 ( .A(n8601), .B(n8598), .ZN(n8605) );
  AOI22_X1 U10042 ( .A1(n8641), .A2(n8819), .B1(n8603), .B2(n8602), .ZN(n8604)
         );
  OAI21_X1 U10043 ( .B1(n8605), .B2(n9815), .A(n8604), .ZN(n8872) );
  OAI21_X1 U10044 ( .B1(n8620), .B2(n8869), .A(n4332), .ZN(n8870) );
  OAI22_X1 U10045 ( .A1(n8607), .A2(n9827), .B1(n8606), .B2(n4316), .ZN(n8608)
         );
  AOI21_X1 U10046 ( .B1(n8609), .B2(n9831), .A(n8608), .ZN(n8610) );
  OAI21_X1 U10047 ( .B1(n8870), .B2(n9833), .A(n8610), .ZN(n8611) );
  AOI21_X1 U10048 ( .B1(n8872), .B2(n4316), .A(n8611), .ZN(n8612) );
  OAI21_X1 U10049 ( .B1(n8613), .B2(n9825), .A(n8612), .ZN(P2_U3267) );
  XNOR2_X1 U10050 ( .A(n8615), .B(n8614), .ZN(n8879) );
  OR2_X1 U10051 ( .A1(n8878), .A2(n8846), .ZN(n8627) );
  AOI21_X1 U10052 ( .B1(n8875), .B2(n8630), .A(n8620), .ZN(n8876) );
  NOR2_X1 U10053 ( .A1(n8621), .A2(n8848), .ZN(n8625) );
  OAI22_X1 U10054 ( .A1(n8623), .A2(n9827), .B1(n8622), .B2(n4316), .ZN(n8624)
         );
  AOI211_X1 U10055 ( .C1(n8876), .C2(n8858), .A(n8625), .B(n8624), .ZN(n8626)
         );
  OAI211_X1 U10056 ( .C1(n8879), .C2(n9825), .A(n8627), .B(n8626), .ZN(
        P2_U3268) );
  XNOR2_X1 U10057 ( .A(n8629), .B(n8628), .ZN(n8884) );
  INV_X1 U10058 ( .A(n8654), .ZN(n8632) );
  INV_X1 U10059 ( .A(n8630), .ZN(n8631) );
  AOI21_X1 U10060 ( .B1(n8880), .B2(n8632), .A(n8631), .ZN(n8881) );
  INV_X1 U10061 ( .A(n8633), .ZN(n8634) );
  AOI22_X1 U10062 ( .A1(n8634), .A2(n8844), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9837), .ZN(n8635) );
  OAI21_X1 U10063 ( .B1(n8636), .B2(n8848), .A(n8635), .ZN(n8645) );
  OAI211_X1 U10064 ( .C1(n8639), .C2(n8638), .A(n8637), .B(n8824), .ZN(n8643)
         );
  AOI22_X1 U10065 ( .A1(n8641), .A2(n8821), .B1(n8819), .B2(n8640), .ZN(n8642)
         );
  AND2_X1 U10066 ( .A1(n8643), .A2(n8642), .ZN(n8883) );
  NOR2_X1 U10067 ( .A1(n8883), .A2(n9837), .ZN(n8644) );
  AOI211_X1 U10068 ( .C1(n8858), .C2(n8881), .A(n8645), .B(n8644), .ZN(n8646)
         );
  OAI21_X1 U10069 ( .B1(n8884), .B2(n9825), .A(n8646), .ZN(P2_U3269) );
  XNOR2_X1 U10070 ( .A(n8648), .B(n8647), .ZN(n8889) );
  NAND2_X1 U10071 ( .A1(n8671), .A2(n8649), .ZN(n8651) );
  XNOR2_X1 U10072 ( .A(n8651), .B(n8650), .ZN(n8653) );
  AOI21_X1 U10073 ( .B1(n8653), .B2(n8824), .A(n8652), .ZN(n8888) );
  AOI211_X1 U10074 ( .C1(n8886), .C2(n8655), .A(n9917), .B(n8654), .ZN(n8885)
         );
  AOI22_X1 U10075 ( .A1(n8885), .A2(n8807), .B1(n8844), .B2(n8656), .ZN(n8657)
         );
  AOI21_X1 U10076 ( .B1(n8888), .B2(n8657), .A(n8846), .ZN(n8661) );
  OAI22_X1 U10077 ( .A1(n8659), .A2(n8848), .B1(n4316), .B2(n8658), .ZN(n8660)
         );
  NOR2_X1 U10078 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  OAI21_X1 U10079 ( .B1(n8889), .B2(n9825), .A(n8662), .ZN(P2_U3270) );
  XNOR2_X1 U10080 ( .A(n8663), .B(n4679), .ZN(n8893) );
  OAI22_X1 U10081 ( .A1(n4316), .A2(n8665), .B1(n8664), .B2(n9827), .ZN(n8677)
         );
  NOR2_X1 U10082 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  AOI21_X1 U10083 ( .B1(n8686), .B2(n8668), .A(n9815), .ZN(n8670) );
  AOI21_X1 U10084 ( .B1(n8671), .B2(n8670), .A(n8669), .ZN(n8675) );
  XNOR2_X1 U10085 ( .A(n8681), .B(n8672), .ZN(n8673) );
  OAI21_X1 U10086 ( .B1(n9917), .B2(n8673), .A(n8675), .ZN(n8890) );
  INV_X1 U10087 ( .A(n8890), .ZN(n8674) );
  AOI211_X1 U10088 ( .C1(n5654), .C2(n8675), .A(n8846), .B(n8674), .ZN(n8676)
         );
  AOI211_X1 U10089 ( .C1(n9831), .C2(n8891), .A(n8677), .B(n8676), .ZN(n8678)
         );
  OAI21_X1 U10090 ( .B1(n8893), .B2(n9825), .A(n8678), .ZN(P2_U3271) );
  AOI21_X1 U10091 ( .B1(n8687), .B2(n8680), .A(n8679), .ZN(n8898) );
  AOI21_X1 U10092 ( .B1(n8894), .B2(n8698), .A(n8681), .ZN(n8895) );
  INV_X1 U10093 ( .A(n8682), .ZN(n8683) );
  AOI22_X1 U10094 ( .A1(n8683), .A2(n8844), .B1(n8846), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8684) );
  OAI21_X1 U10095 ( .B1(n8685), .B2(n8848), .A(n8684), .ZN(n8694) );
  OAI211_X1 U10096 ( .C1(n8688), .C2(n8687), .A(n8686), .B(n8824), .ZN(n8692)
         );
  AOI22_X1 U10097 ( .A1(n8690), .A2(n8821), .B1(n8819), .B2(n8689), .ZN(n8691)
         );
  AND2_X1 U10098 ( .A1(n8692), .A2(n8691), .ZN(n8897) );
  NOR2_X1 U10099 ( .A1(n8897), .A2(n9837), .ZN(n8693) );
  AOI211_X1 U10100 ( .C1(n8895), .C2(n8858), .A(n8694), .B(n8693), .ZN(n8695)
         );
  OAI21_X1 U10101 ( .B1(n8898), .B2(n9825), .A(n8695), .ZN(P2_U3272) );
  OAI21_X1 U10102 ( .B1(n8697), .B2(n8706), .A(n8696), .ZN(n8903) );
  INV_X1 U10103 ( .A(n8698), .ZN(n8699) );
  AOI21_X1 U10104 ( .B1(n8899), .B2(n4564), .A(n8699), .ZN(n8900) );
  INV_X1 U10105 ( .A(n8700), .ZN(n8701) );
  AOI22_X1 U10106 ( .A1(n8846), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8701), .B2(
        n8844), .ZN(n8702) );
  OAI21_X1 U10107 ( .B1(n8703), .B2(n8848), .A(n8702), .ZN(n8711) );
  AOI21_X1 U10108 ( .B1(n8706), .B2(n8705), .A(n8704), .ZN(n8707) );
  INV_X1 U10109 ( .A(n8707), .ZN(n8709) );
  AOI222_X1 U10110 ( .A1(n8824), .A2(n8709), .B1(n8740), .B2(n8819), .C1(n8708), .C2(n8821), .ZN(n8902) );
  NOR2_X1 U10111 ( .A1(n8902), .A2(n8846), .ZN(n8710) );
  AOI211_X1 U10112 ( .C1(n8900), .C2(n8858), .A(n8711), .B(n8710), .ZN(n8712)
         );
  OAI21_X1 U10113 ( .B1(n9825), .B2(n8903), .A(n8712), .ZN(P2_U3273) );
  XNOR2_X1 U10114 ( .A(n8713), .B(n8721), .ZN(n8908) );
  AOI21_X1 U10115 ( .B1(n8904), .B2(n8715), .A(n8714), .ZN(n8905) );
  INV_X1 U10116 ( .A(n8716), .ZN(n8717) );
  AOI22_X1 U10117 ( .A1(n8846), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8717), .B2(
        n8844), .ZN(n8718) );
  OAI21_X1 U10118 ( .B1(n8719), .B2(n8848), .A(n8718), .ZN(n8730) );
  INV_X1 U10119 ( .A(n8720), .ZN(n8724) );
  AOI21_X1 U10120 ( .B1(n8737), .B2(n8722), .A(n8721), .ZN(n8723) );
  NOR3_X1 U10121 ( .A1(n8724), .A2(n8723), .A3(n9815), .ZN(n8728) );
  OAI22_X1 U10122 ( .A1(n8726), .A2(n8806), .B1(n8725), .B2(n8804), .ZN(n8727)
         );
  NOR2_X1 U10123 ( .A1(n8728), .A2(n8727), .ZN(n8907) );
  NOR2_X1 U10124 ( .A1(n8907), .A2(n8846), .ZN(n8729) );
  AOI211_X1 U10125 ( .C1(n8905), .C2(n8858), .A(n8730), .B(n8729), .ZN(n8731)
         );
  OAI21_X1 U10126 ( .B1(n8908), .B2(n9825), .A(n8731), .ZN(P2_U3274) );
  XNOR2_X1 U10127 ( .A(n8732), .B(n8738), .ZN(n8913) );
  XNOR2_X1 U10128 ( .A(n8747), .B(n8736), .ZN(n8910) );
  INV_X1 U10129 ( .A(n8733), .ZN(n8734) );
  AOI22_X1 U10130 ( .A1(n8846), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8734), .B2(
        n8844), .ZN(n8735) );
  OAI21_X1 U10131 ( .B1(n8736), .B2(n8848), .A(n8735), .ZN(n8743) );
  OAI21_X1 U10132 ( .B1(n8739), .B2(n8738), .A(n8737), .ZN(n8741) );
  AOI222_X1 U10133 ( .A1(n8824), .A2(n8741), .B1(n8740), .B2(n8821), .C1(n8766), .C2(n8819), .ZN(n8912) );
  NOR2_X1 U10134 ( .A1(n8912), .A2(n9837), .ZN(n8742) );
  AOI211_X1 U10135 ( .C1(n8910), .C2(n8858), .A(n8743), .B(n8742), .ZN(n8744)
         );
  OAI21_X1 U10136 ( .B1(n9825), .B2(n8913), .A(n8744), .ZN(P2_U3275) );
  XNOR2_X1 U10137 ( .A(n8745), .B(n8755), .ZN(n8918) );
  INV_X1 U10138 ( .A(n8746), .ZN(n8768) );
  INV_X1 U10139 ( .A(n8747), .ZN(n8748) );
  AOI21_X1 U10140 ( .B1(n8914), .B2(n8768), .A(n8748), .ZN(n8915) );
  INV_X1 U10141 ( .A(n8749), .ZN(n8750) );
  AOI22_X1 U10142 ( .A1(n8846), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8750), .B2(
        n8844), .ZN(n8751) );
  OAI21_X1 U10143 ( .B1(n8752), .B2(n8848), .A(n8751), .ZN(n8759) );
  NAND2_X1 U10144 ( .A1(n8762), .A2(n8753), .ZN(n8754) );
  XOR2_X1 U10145 ( .A(n8755), .B(n8754), .Z(n8757) );
  AOI222_X1 U10146 ( .A1(n8824), .A2(n8757), .B1(n8756), .B2(n8821), .C1(n8793), .C2(n8819), .ZN(n8917) );
  NOR2_X1 U10147 ( .A1(n8917), .A2(n8846), .ZN(n8758) );
  AOI211_X1 U10148 ( .C1(n8915), .C2(n8858), .A(n8759), .B(n8758), .ZN(n8760)
         );
  OAI21_X1 U10149 ( .B1(n9825), .B2(n8918), .A(n8760), .ZN(P2_U3276) );
  XNOR2_X1 U10150 ( .A(n8761), .B(n8764), .ZN(n8771) );
  INV_X1 U10151 ( .A(n8771), .ZN(n8922) );
  OAI21_X1 U10152 ( .B1(n8764), .B2(n8763), .A(n8762), .ZN(n8767) );
  AOI222_X1 U10153 ( .A1(n8824), .A2(n8767), .B1(n8766), .B2(n8821), .C1(n8765), .C2(n8819), .ZN(n8774) );
  OAI211_X1 U10154 ( .C1(n8769), .C2(n8783), .A(n8768), .B(n9868), .ZN(n8770)
         );
  NAND2_X1 U10155 ( .A1(n8774), .A2(n8770), .ZN(n8919) );
  AOI21_X1 U10156 ( .B1(n8772), .B2(n8771), .A(n8919), .ZN(n8773) );
  AOI211_X1 U10157 ( .C1(n5654), .C2(n8774), .A(n8846), .B(n8773), .ZN(n8775)
         );
  INV_X1 U10158 ( .A(n8775), .ZN(n8780) );
  OAI22_X1 U10159 ( .A1(n4316), .A2(n8777), .B1(n8776), .B2(n9827), .ZN(n8778)
         );
  AOI21_X1 U10160 ( .B1(n8920), .B2(n9831), .A(n8778), .ZN(n8779) );
  OAI211_X1 U10161 ( .C1(n8922), .C2(n8781), .A(n8780), .B(n8779), .ZN(
        P2_U3277) );
  XNOR2_X1 U10162 ( .A(n8782), .B(n8791), .ZN(n8927) );
  AOI21_X1 U10163 ( .B1(n8923), .B2(n8798), .A(n8783), .ZN(n8924) );
  INV_X1 U10164 ( .A(n8784), .ZN(n8785) );
  AOI22_X1 U10165 ( .A1(n8846), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8785), .B2(
        n8844), .ZN(n8786) );
  OAI21_X1 U10166 ( .B1(n8787), .B2(n8848), .A(n8786), .ZN(n8796) );
  AND2_X1 U10167 ( .A1(n8789), .A2(n8788), .ZN(n8792) );
  OAI21_X1 U10168 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8794) );
  AOI222_X1 U10169 ( .A1(n8824), .A2(n8794), .B1(n8793), .B2(n8821), .C1(n8822), .C2(n8819), .ZN(n8926) );
  NOR2_X1 U10170 ( .A1(n8926), .A2(n8846), .ZN(n8795) );
  AOI211_X1 U10171 ( .C1(n8924), .C2(n8858), .A(n8796), .B(n8795), .ZN(n8797)
         );
  OAI21_X1 U10172 ( .B1(n8927), .B2(n9825), .A(n8797), .ZN(P2_U3278) );
  INV_X1 U10173 ( .A(n8798), .ZN(n8799) );
  AOI211_X1 U10174 ( .C1(n8930), .C2(n8825), .A(n9917), .B(n8799), .ZN(n8929)
         );
  XNOR2_X1 U10175 ( .A(n8801), .B(n8800), .ZN(n8802) );
  OAI222_X1 U10176 ( .A1(n8806), .A2(n8805), .B1(n8804), .B2(n8803), .C1(n9815), .C2(n8802), .ZN(n8928) );
  AOI21_X1 U10177 ( .B1(n8929), .B2(n8807), .A(n8928), .ZN(n8817) );
  OAI22_X1 U10178 ( .A1(n4316), .A2(n8809), .B1(n8808), .B2(n9827), .ZN(n8815)
         );
  OAI21_X1 U10179 ( .B1(n8812), .B2(n8811), .A(n8810), .ZN(n8813) );
  INV_X1 U10180 ( .A(n8813), .ZN(n8932) );
  NOR2_X1 U10181 ( .A1(n8932), .A2(n9825), .ZN(n8814) );
  AOI211_X1 U10182 ( .C1(n9831), .C2(n8930), .A(n8815), .B(n8814), .ZN(n8816)
         );
  OAI21_X1 U10183 ( .B1(n8817), .B2(n9837), .A(n8816), .ZN(P2_U3279) );
  XNOR2_X1 U10184 ( .A(n8818), .B(n8833), .ZN(n8823) );
  AOI222_X1 U10185 ( .A1(n8824), .A2(n8823), .B1(n8822), .B2(n8821), .C1(n8820), .C2(n8819), .ZN(n8936) );
  INV_X1 U10186 ( .A(n8842), .ZN(n8827) );
  INV_X1 U10187 ( .A(n8825), .ZN(n8826) );
  AOI21_X1 U10188 ( .B1(n8933), .B2(n8827), .A(n8826), .ZN(n8934) );
  AOI22_X1 U10189 ( .A1(n8846), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8828), .B2(
        n8844), .ZN(n8829) );
  OAI21_X1 U10190 ( .B1(n8830), .B2(n8848), .A(n8829), .ZN(n8836) );
  AOI21_X1 U10191 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n8834) );
  INV_X1 U10192 ( .A(n8834), .ZN(n8937) );
  NOR2_X1 U10193 ( .A1(n8937), .A2(n9825), .ZN(n8835) );
  AOI211_X1 U10194 ( .C1(n8934), .C2(n8858), .A(n8836), .B(n8835), .ZN(n8837)
         );
  OAI21_X1 U10195 ( .B1(n8936), .B2(n9837), .A(n8837), .ZN(P2_U3280) );
  OAI21_X1 U10196 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8841) );
  INV_X1 U10197 ( .A(n8841), .ZN(n8942) );
  AOI21_X1 U10198 ( .B1(n8938), .B2(n4331), .A(n8842), .ZN(n8939) );
  INV_X1 U10199 ( .A(n8843), .ZN(n8845) );
  AOI22_X1 U10200 ( .A1(n8846), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8845), .B2(
        n8844), .ZN(n8847) );
  OAI21_X1 U10201 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8857) );
  NOR2_X1 U10202 ( .A1(n4840), .A2(n4837), .ZN(n8853) );
  AOI211_X1 U10203 ( .C1(n8853), .C2(n8852), .A(n9815), .B(n8851), .ZN(n8855)
         );
  NOR2_X1 U10204 ( .A1(n8855), .A2(n8854), .ZN(n8941) );
  NOR2_X1 U10205 ( .A1(n8941), .A2(n9837), .ZN(n8856) );
  AOI211_X1 U10206 ( .C1(n8939), .C2(n8858), .A(n8857), .B(n8856), .ZN(n8859)
         );
  OAI21_X1 U10207 ( .B1(n8942), .B2(n9825), .A(n8859), .ZN(P2_U3281) );
  NAND2_X1 U10208 ( .A1(n8860), .A2(n9868), .ZN(n8861) );
  OAI211_X1 U10209 ( .C1(n8862), .C2(n9915), .A(n8861), .B(n8865), .ZN(n8955)
         );
  MUX2_X1 U10210 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8955), .S(n9939), .Z(
        P2_U3551) );
  NAND3_X1 U10211 ( .A1(n8864), .A2(n9868), .A3(n8863), .ZN(n8866) );
  OAI211_X1 U10212 ( .C1(n8867), .C2(n9915), .A(n8866), .B(n8865), .ZN(n8956)
         );
  MUX2_X1 U10213 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8956), .S(n9939), .Z(
        P2_U3550) );
  NAND2_X1 U10214 ( .A1(n8868), .A2(n9921), .ZN(n8874) );
  OAI22_X1 U10215 ( .A1(n8870), .A2(n9917), .B1(n8869), .B2(n9915), .ZN(n8871)
         );
  NOR2_X1 U10216 ( .A1(n8872), .A2(n8871), .ZN(n8873) );
  NAND2_X1 U10217 ( .A1(n8874), .A2(n8873), .ZN(n8957) );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8957), .S(n9939), .Z(
        P2_U3549) );
  AOI22_X1 U10219 ( .A1(n8876), .A2(n9868), .B1(n9886), .B2(n8875), .ZN(n8877)
         );
  OAI211_X1 U10220 ( .C1(n8879), .C2(n9889), .A(n8878), .B(n8877), .ZN(n8958)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8958), .S(n9939), .Z(
        P2_U3548) );
  AOI22_X1 U10222 ( .A1(n8881), .A2(n9868), .B1(n9886), .B2(n8880), .ZN(n8882)
         );
  OAI211_X1 U10223 ( .C1(n8884), .C2(n9889), .A(n8883), .B(n8882), .ZN(n8959)
         );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8959), .S(n9939), .Z(
        P2_U3547) );
  AOI21_X1 U10225 ( .B1(n9886), .B2(n8886), .A(n8885), .ZN(n8887) );
  OAI211_X1 U10226 ( .C1(n8889), .C2(n9889), .A(n8888), .B(n8887), .ZN(n8960)
         );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8960), .S(n9939), .Z(
        P2_U3546) );
  AOI21_X1 U10228 ( .B1(n9886), .B2(n8891), .A(n8890), .ZN(n8892) );
  OAI21_X1 U10229 ( .B1(n9889), .B2(n8893), .A(n8892), .ZN(n8961) );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8961), .S(n9939), .Z(
        P2_U3545) );
  AOI22_X1 U10231 ( .A1(n8895), .A2(n9868), .B1(n9886), .B2(n8894), .ZN(n8896)
         );
  OAI211_X1 U10232 ( .C1(n8898), .C2(n9889), .A(n8897), .B(n8896), .ZN(n8962)
         );
  MUX2_X1 U10233 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8962), .S(n9939), .Z(
        P2_U3544) );
  AOI22_X1 U10234 ( .A1(n8900), .A2(n9868), .B1(n9886), .B2(n8899), .ZN(n8901)
         );
  OAI211_X1 U10235 ( .C1(n9889), .C2(n8903), .A(n8902), .B(n8901), .ZN(n8963)
         );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8963), .S(n9939), .Z(
        P2_U3543) );
  AOI22_X1 U10237 ( .A1(n8905), .A2(n9868), .B1(n9886), .B2(n8904), .ZN(n8906)
         );
  OAI211_X1 U10238 ( .C1(n9889), .C2(n8908), .A(n8907), .B(n8906), .ZN(n8964)
         );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8964), .S(n9939), .Z(
        P2_U3542) );
  AOI22_X1 U10240 ( .A1(n8910), .A2(n9868), .B1(n9886), .B2(n8909), .ZN(n8911)
         );
  OAI211_X1 U10241 ( .C1(n9889), .C2(n8913), .A(n8912), .B(n8911), .ZN(n8965)
         );
  MUX2_X1 U10242 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8965), .S(n9939), .Z(
        P2_U3541) );
  AOI22_X1 U10243 ( .A1(n8915), .A2(n9868), .B1(n9886), .B2(n8914), .ZN(n8916)
         );
  OAI211_X1 U10244 ( .C1(n9889), .C2(n8918), .A(n8917), .B(n8916), .ZN(n8966)
         );
  MUX2_X1 U10245 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8966), .S(n9939), .Z(
        P2_U3540) );
  AOI21_X1 U10246 ( .B1(n9886), .B2(n8920), .A(n8919), .ZN(n8921) );
  OAI21_X1 U10247 ( .B1(n9889), .B2(n8922), .A(n8921), .ZN(n8967) );
  MUX2_X1 U10248 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8967), .S(n9939), .Z(
        P2_U3539) );
  AOI22_X1 U10249 ( .A1(n8924), .A2(n9868), .B1(n9886), .B2(n8923), .ZN(n8925)
         );
  OAI211_X1 U10250 ( .C1(n9889), .C2(n8927), .A(n8926), .B(n8925), .ZN(n8968)
         );
  MUX2_X1 U10251 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8968), .S(n9939), .Z(
        P2_U3538) );
  AOI211_X1 U10252 ( .C1(n9886), .C2(n8930), .A(n8929), .B(n8928), .ZN(n8931)
         );
  OAI21_X1 U10253 ( .B1(n9889), .B2(n8932), .A(n8931), .ZN(n8969) );
  MUX2_X1 U10254 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8969), .S(n9939), .Z(
        P2_U3537) );
  AOI22_X1 U10255 ( .A1(n8934), .A2(n9868), .B1(n9886), .B2(n8933), .ZN(n8935)
         );
  OAI211_X1 U10256 ( .C1(n9889), .C2(n8937), .A(n8936), .B(n8935), .ZN(n8970)
         );
  MUX2_X1 U10257 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8970), .S(n9939), .Z(
        P2_U3536) );
  AOI22_X1 U10258 ( .A1(n8939), .A2(n9868), .B1(n9886), .B2(n8938), .ZN(n8940)
         );
  OAI211_X1 U10259 ( .C1(n9889), .C2(n8942), .A(n8941), .B(n8940), .ZN(n8971)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8971), .S(n9939), .Z(
        P2_U3535) );
  AOI22_X1 U10261 ( .A1(n8944), .A2(n9868), .B1(n9886), .B2(n8943), .ZN(n8945)
         );
  OAI211_X1 U10262 ( .C1(n9867), .C2(n8947), .A(n8946), .B(n8945), .ZN(n8972)
         );
  MUX2_X1 U10263 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8972), .S(n9939), .Z(
        P2_U3533) );
  INV_X1 U10264 ( .A(n8948), .ZN(n8949) );
  OAI22_X1 U10265 ( .A1(n8950), .A2(n9917), .B1(n8949), .B2(n9915), .ZN(n8951)
         );
  INV_X1 U10266 ( .A(n8951), .ZN(n8952) );
  OAI211_X1 U10267 ( .C1(n9889), .C2(n8954), .A(n8953), .B(n8952), .ZN(n8973)
         );
  MUX2_X1 U10268 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8973), .S(n9939), .Z(
        P2_U3531) );
  MUX2_X1 U10269 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8955), .S(n9924), .Z(
        P2_U3519) );
  MUX2_X1 U10270 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8956), .S(n9924), .Z(
        P2_U3518) );
  MUX2_X1 U10271 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8957), .S(n9924), .Z(
        P2_U3517) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8958), .S(n9924), .Z(
        P2_U3516) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8959), .S(n9924), .Z(
        P2_U3515) );
  MUX2_X1 U10274 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8960), .S(n9924), .Z(
        P2_U3514) );
  MUX2_X1 U10275 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8961), .S(n9924), .Z(
        P2_U3513) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8962), .S(n9924), .Z(
        P2_U3512) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8963), .S(n9924), .Z(
        P2_U3511) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8964), .S(n9924), .Z(
        P2_U3510) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8965), .S(n9924), .Z(
        P2_U3509) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8966), .S(n9924), .Z(
        P2_U3508) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8967), .S(n9924), .Z(
        P2_U3507) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8968), .S(n9924), .Z(
        P2_U3505) );
  MUX2_X1 U10283 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8969), .S(n9924), .Z(
        P2_U3502) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8970), .S(n9924), .Z(
        P2_U3499) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8971), .S(n9924), .Z(
        P2_U3496) );
  MUX2_X1 U10286 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8972), .S(n9924), .Z(
        P2_U3490) );
  MUX2_X1 U10287 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8973), .S(n9924), .Z(
        P2_U3484) );
  NAND3_X1 U10288 ( .A1(n8974), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8976) );
  OAI22_X1 U10289 ( .A1(n8977), .A2(n8976), .B1(n8975), .B2(n8987), .ZN(n8978)
         );
  AOI21_X1 U10290 ( .B1(n9586), .B2(n8979), .A(n8978), .ZN(n8980) );
  INV_X1 U10291 ( .A(n8980), .ZN(P2_U3327) );
  OAI222_X1 U10292 ( .A1(n6866), .A2(n8983), .B1(P2_U3152), .B2(n8982), .C1(
        n8981), .C2(n8987), .ZN(P2_U3329) );
  INV_X1 U10293 ( .A(n8984), .ZN(n9598) );
  OAI222_X1 U10294 ( .A1(n8987), .A2(n8986), .B1(n6866), .B2(n9598), .C1(n8985), .C2(P2_U3152), .ZN(P2_U3331) );
  MUX2_X1 U10295 ( .A(n8988), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AOI21_X1 U10296 ( .B1(n8991), .B2(n8990), .A(n8989), .ZN(n8993) );
  OAI21_X1 U10297 ( .B1(n8993), .B2(n8992), .A(n9678), .ZN(n8997) );
  AOI22_X1 U10298 ( .A1(n9111), .A2(n9272), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8994) );
  OAI21_X1 U10299 ( .B1(n9096), .B2(n9235), .A(n8994), .ZN(n8995) );
  AOI21_X1 U10300 ( .B1(n9267), .B2(n9100), .A(n8995), .ZN(n8996) );
  OAI211_X1 U10301 ( .C1(n9269), .C2(n9056), .A(n8997), .B(n8996), .ZN(
        P1_U3212) );
  NAND2_X1 U10302 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  XOR2_X1 U10303 ( .A(n9001), .B(n9000), .Z(n9008) );
  OAI22_X1 U10304 ( .A1(n9003), .A2(n9667), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9002), .ZN(n9005) );
  NOR2_X1 U10305 ( .A1(n9642), .A2(n9056), .ZN(n9004) );
  AOI211_X1 U10306 ( .C1(n9006), .C2(n9100), .A(n9005), .B(n9004), .ZN(n9007)
         );
  OAI21_X1 U10307 ( .B1(n9008), .B2(n9117), .A(n9007), .ZN(P1_U3213) );
  INV_X1 U10308 ( .A(n9009), .ZN(n9011) );
  XNOR2_X1 U10309 ( .A(n9011), .B(n9010), .ZN(n9012) );
  XNOR2_X1 U10310 ( .A(n9013), .B(n9012), .ZN(n9019) );
  OAI22_X1 U10311 ( .A1(n6830), .A2(n9356), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9014), .ZN(n9017) );
  INV_X1 U10312 ( .A(n9324), .ZN(n9015) );
  OAI22_X1 U10313 ( .A1(n9096), .A2(n9330), .B1(n9683), .B2(n9015), .ZN(n9016)
         );
  AOI211_X1 U10314 ( .C1(n9513), .C2(n9115), .A(n9017), .B(n9016), .ZN(n9018)
         );
  OAI21_X1 U10315 ( .B1(n9019), .B2(n9117), .A(n9018), .ZN(P1_U3214) );
  NAND2_X1 U10316 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  XNOR2_X1 U10317 ( .A(n9023), .B(n9022), .ZN(n9028) );
  NAND2_X1 U10318 ( .A1(n9100), .A2(n9359), .ZN(n9025) );
  AOI22_X1 U10319 ( .A1(n9394), .A2(n9111), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9024) );
  OAI211_X1 U10320 ( .C1(n9356), .C2(n9096), .A(n9025), .B(n9024), .ZN(n9026)
         );
  AOI21_X1 U10321 ( .B1(n9525), .B2(n9115), .A(n9026), .ZN(n9027) );
  OAI21_X1 U10322 ( .B1(n9028), .B2(n9117), .A(n9027), .ZN(P1_U3221) );
  OAI21_X1 U10323 ( .B1(n9030), .B2(n9029), .A(n5538), .ZN(n9031) );
  NAND2_X1 U10324 ( .A1(n9031), .A2(n9678), .ZN(n9035) );
  AOI22_X1 U10325 ( .A1(n9207), .A2(n9111), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9032) );
  OAI21_X1 U10326 ( .B1(n9096), .B2(n9295), .A(n9032), .ZN(n9033) );
  AOI21_X1 U10327 ( .B1(n9297), .B2(n9100), .A(n9033), .ZN(n9034) );
  OAI211_X1 U10328 ( .C1(n9208), .C2(n9056), .A(n9035), .B(n9034), .ZN(
        P1_U3223) );
  XOR2_X1 U10329 ( .A(n9037), .B(n9036), .Z(n9043) );
  OAI22_X1 U10330 ( .A1(n6830), .A2(n9437), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9038), .ZN(n9041) );
  INV_X1 U10331 ( .A(n9445), .ZN(n9039) );
  OAI22_X1 U10332 ( .A1(n9096), .A2(n9439), .B1(n9683), .B2(n9039), .ZN(n9040)
         );
  AOI211_X1 U10333 ( .C1(n9552), .C2(n9115), .A(n9041), .B(n9040), .ZN(n9042)
         );
  OAI21_X1 U10334 ( .B1(n9043), .B2(n9117), .A(n9042), .ZN(P1_U3224) );
  XOR2_X1 U10335 ( .A(n9045), .B(n9044), .Z(n9051) );
  NAND2_X1 U10336 ( .A1(n9100), .A2(n9419), .ZN(n9047) );
  AOI22_X1 U10337 ( .A1(n9424), .A2(n9111), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n9046) );
  OAI211_X1 U10338 ( .C1(n9048), .C2(n9096), .A(n9047), .B(n9046), .ZN(n9049)
         );
  AOI21_X1 U10339 ( .B1(n9545), .B2(n9115), .A(n9049), .ZN(n9050) );
  OAI21_X1 U10340 ( .B1(n9051), .B2(n9117), .A(n9050), .ZN(P1_U3226) );
  AOI21_X1 U10341 ( .B1(n9053), .B2(n9052), .A(n4362), .ZN(n9060) );
  AOI22_X1 U10342 ( .A1(n9345), .A2(n9111), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9055) );
  OAI21_X1 U10343 ( .B1(n9096), .B2(n9310), .A(n9055), .ZN(n9058) );
  NOR2_X1 U10344 ( .A1(n9206), .A2(n9056), .ZN(n9057) );
  AOI211_X1 U10345 ( .C1(n9313), .C2(n9100), .A(n9058), .B(n9057), .ZN(n9059)
         );
  OAI21_X1 U10346 ( .B1(n9060), .B2(n9117), .A(n9059), .ZN(P1_U3227) );
  INV_X1 U10347 ( .A(n9061), .ZN(n9062) );
  NOR2_X1 U10348 ( .A1(n9063), .A2(n9062), .ZN(n9064) );
  XNOR2_X1 U10349 ( .A(n9065), .B(n9064), .ZN(n9070) );
  NOR2_X1 U10350 ( .A1(n9683), .A2(n9371), .ZN(n9068) );
  AOI22_X1 U10351 ( .A1(n9111), .A2(n9402), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9066) );
  OAI21_X1 U10352 ( .B1(n9201), .B2(n9096), .A(n9066), .ZN(n9067) );
  AOI211_X1 U10353 ( .C1(n9528), .C2(n9115), .A(n9068), .B(n9067), .ZN(n9069)
         );
  OAI21_X1 U10354 ( .B1(n9070), .B2(n9117), .A(n9069), .ZN(P1_U3231) );
  XOR2_X1 U10355 ( .A(n9072), .B(n9071), .Z(n9073) );
  XNOR2_X1 U10356 ( .A(n9074), .B(n9073), .ZN(n9079) );
  INV_X1 U10357 ( .A(n9201), .ZN(n9369) );
  AOI22_X1 U10358 ( .A1(n9369), .A2(n9111), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9076) );
  NAND2_X1 U10359 ( .A1(n9100), .A2(n9339), .ZN(n9075) );
  OAI211_X1 U10360 ( .C1(n9309), .C2(n9096), .A(n9076), .B(n9075), .ZN(n9077)
         );
  AOI21_X1 U10361 ( .B1(n9519), .B2(n9115), .A(n9077), .ZN(n9078) );
  OAI21_X1 U10362 ( .B1(n9079), .B2(n9117), .A(n9078), .ZN(P1_U3233) );
  NAND2_X1 U10363 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  XOR2_X1 U10364 ( .A(n9083), .B(n9082), .Z(n9089) );
  NAND2_X1 U10365 ( .A1(n9100), .A2(n9406), .ZN(n9086) );
  NOR2_X1 U10366 ( .A1(n9084), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9697) );
  AOI21_X1 U10367 ( .B1(n9403), .B2(n9111), .A(n9697), .ZN(n9085) );
  OAI211_X1 U10368 ( .C1(n9199), .C2(n9096), .A(n9086), .B(n9085), .ZN(n9087)
         );
  AOI21_X1 U10369 ( .B1(n9539), .B2(n9115), .A(n9087), .ZN(n9088) );
  OAI21_X1 U10370 ( .B1(n9089), .B2(n9117), .A(n9088), .ZN(P1_U3236) );
  INV_X1 U10371 ( .A(n9090), .ZN(n9094) );
  NOR3_X1 U10372 ( .A1(n9092), .A2(n4776), .A3(n9091), .ZN(n9093) );
  OAI21_X1 U10373 ( .B1(n9094), .B2(n9093), .A(n9678), .ZN(n9103) );
  NOR2_X1 U10374 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  AOI211_X1 U10375 ( .C1(n9111), .C2(n9129), .A(n9098), .B(n9097), .ZN(n9102)
         );
  AOI22_X1 U10376 ( .A1(n9100), .A2(n9099), .B1(n9115), .B2(n4315), .ZN(n9101)
         );
  NAND3_X1 U10377 ( .A1(n9103), .A2(n9102), .A3(n9101), .ZN(P1_U3237) );
  NAND2_X1 U10378 ( .A1(n9104), .A2(n9105), .ZN(n9106) );
  XOR2_X1 U10379 ( .A(n9107), .B(n9106), .Z(n9118) );
  NOR2_X1 U10380 ( .A1(n9096), .A2(n9108), .ZN(n9109) );
  AOI211_X1 U10381 ( .C1(n9111), .C2(n9121), .A(n9110), .B(n9109), .ZN(n9112)
         );
  OAI21_X1 U10382 ( .B1(n9683), .B2(n9113), .A(n9112), .ZN(n9114) );
  AOI21_X1 U10383 ( .B1(n9197), .B2(n9115), .A(n9114), .ZN(n9116) );
  OAI21_X1 U10384 ( .B1(n9118), .B2(n9117), .A(n9116), .ZN(P1_U3239) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9119), .S(n9132), .Z(
        P1_U3586) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9120), .S(n9132), .Z(
        P1_U3585) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9258), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9273), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9286), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9272), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9209), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9207), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9345), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9202), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9369), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9394), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9402), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9425), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9403), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9424), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9196), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9121), .S(n9132), .Z(
        P1_U3569) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9122), .S(n9132), .Z(
        P1_U3568) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9123), .S(n9132), .Z(
        P1_U3567) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9124), .S(n9132), .Z(
        P1_U3566) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9125), .S(n9132), .Z(
        P1_U3565) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9126), .S(n9132), .Z(
        P1_U3564) );
  MUX2_X1 U10408 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9127), .S(n9132), .Z(
        P1_U3563) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9128), .S(n9132), .Z(
        P1_U3562) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9457), .S(n9132), .Z(
        P1_U3561) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9129), .S(n9132), .Z(
        P1_U3560) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9455), .S(n9132), .Z(
        P1_U3559) );
  MUX2_X1 U10413 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9130), .S(n9132), .Z(
        P1_U3558) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9131), .S(n9132), .Z(
        P1_U3557) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9133), .S(n9132), .Z(
        P1_U3556) );
  OAI211_X1 U10416 ( .C1(n9136), .C2(n9135), .A(n9157), .B(n9134), .ZN(n9146)
         );
  AOI21_X1 U10417 ( .B1(n9698), .B2(n9138), .A(n9137), .ZN(n9145) );
  OAI21_X1 U10418 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(n9142) );
  NAND2_X1 U10419 ( .A1(n9142), .A2(n9704), .ZN(n9144) );
  NAND2_X1 U10420 ( .A1(n9703), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n9143) );
  NAND4_X1 U10421 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(
        P1_U3250) );
  INV_X1 U10422 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9162) );
  AND2_X1 U10423 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9152) );
  AOI21_X1 U10424 ( .B1(n9148), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9147), .ZN(
        n9150) );
  XNOR2_X1 U10425 ( .A(n9171), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9149) );
  NOR2_X1 U10426 ( .A1(n9150), .A2(n9149), .ZN(n9170) );
  AOI211_X1 U10427 ( .C1(n9150), .C2(n9149), .A(n9170), .B(n9173), .ZN(n9151)
         );
  AOI211_X1 U10428 ( .C1(n9698), .C2(n9171), .A(n9152), .B(n9151), .ZN(n9161)
         );
  INV_X1 U10429 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9153) );
  XNOR2_X1 U10430 ( .A(n9171), .B(n9153), .ZN(n9159) );
  INV_X1 U10431 ( .A(n9154), .ZN(n9155) );
  NAND2_X1 U10432 ( .A1(n9156), .A2(n9155), .ZN(n9158) );
  NAND2_X1 U10433 ( .A1(n9158), .A2(n9159), .ZN(n9164) );
  OAI211_X1 U10434 ( .C1(n9159), .C2(n9158), .A(n9157), .B(n9164), .ZN(n9160)
         );
  OAI211_X1 U10435 ( .C1(n9184), .C2(n9162), .A(n9161), .B(n9160), .ZN(
        P1_U3258) );
  NAND2_X1 U10436 ( .A1(n9171), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U10437 ( .A1(n9164), .A2(n9163), .ZN(n9692) );
  OR2_X1 U10438 ( .A1(n9699), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U10439 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9699), .ZN(n9165) );
  AND2_X1 U10440 ( .A1(n9166), .A2(n9165), .ZN(n9691) );
  XNOR2_X1 U10441 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9167), .ZN(n9178) );
  INV_X1 U10442 ( .A(n9178), .ZN(n9174) );
  INV_X1 U10443 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9168) );
  AOI22_X1 U10444 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9699), .B1(n9169), .B2(
        n9168), .ZN(n9701) );
  AOI21_X1 U10445 ( .B1(n9171), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9170), .ZN(
        n9702) );
  NAND2_X1 U10446 ( .A1(n9701), .A2(n9702), .ZN(n9700) );
  OAI21_X1 U10447 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9699), .A(n9700), .ZN(
        n9172) );
  XOR2_X1 U10448 ( .A(n9172), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9175) );
  OAI22_X1 U10449 ( .A1(n9174), .A2(n9695), .B1(n9175), .B2(n9173), .ZN(n9180)
         );
  AOI21_X1 U10450 ( .B1(n9175), .B2(n9704), .A(n9698), .ZN(n9176) );
  OAI21_X1 U10451 ( .B1(n9178), .B2(n9177), .A(n9176), .ZN(n9179) );
  MUX2_X1 U10452 ( .A(n9180), .B(n9179), .S(n9315), .Z(n9181) );
  INV_X1 U10453 ( .A(n9181), .ZN(n9183) );
  OAI211_X1 U10454 ( .C1(n4581), .C2(n9184), .A(n9183), .B(n9182), .ZN(
        P1_U3260) );
  NAND2_X1 U10455 ( .A1(n9405), .A2(n9388), .ZN(n9382) );
  NAND2_X1 U10456 ( .A1(n9278), .A2(n9269), .ZN(n9264) );
  NOR2_X2 U10457 ( .A1(n9237), .A2(n9248), .ZN(n9236) );
  NAND2_X1 U10458 ( .A1(n9192), .A2(n9236), .ZN(n9185) );
  XNOR2_X1 U10459 ( .A(n9185), .B(n9476), .ZN(n9478) );
  NAND2_X1 U10460 ( .A1(n9186), .A2(P1_B_REG_SCAN_IN), .ZN(n9187) );
  NAND2_X1 U10461 ( .A1(n9456), .A2(n9187), .ZN(n9234) );
  NOR2_X1 U10462 ( .A1(n9188), .A2(n9234), .ZN(n9479) );
  INV_X1 U10463 ( .A(n9479), .ZN(n9189) );
  NOR2_X1 U10464 ( .A1(n9189), .A2(n9305), .ZN(n9194) );
  AOI21_X1 U10465 ( .B1(n9305), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9194), .ZN(
        n9191) );
  NAND2_X1 U10466 ( .A1(n9476), .A2(n9374), .ZN(n9190) );
  OAI211_X1 U10467 ( .C1(n9478), .C2(n9376), .A(n9191), .B(n9190), .ZN(
        P1_U3261) );
  XNOR2_X1 U10468 ( .A(n9192), .B(n9236), .ZN(n9482) );
  NOR2_X1 U10469 ( .A1(n9192), .A2(n9467), .ZN(n9193) );
  AOI211_X1 U10470 ( .C1(n9305), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9194), .B(
        n9193), .ZN(n9195) );
  OAI21_X1 U10471 ( .B1(n9376), .B2(n9482), .A(n9195), .ZN(P1_U3262) );
  INV_X1 U10472 ( .A(n9525), .ZN(n9362) );
  NOR2_X1 U10473 ( .A1(n9411), .A2(n9410), .ZN(n9544) );
  NOR2_X1 U10474 ( .A1(n9533), .A2(n9402), .ZN(n9200) );
  OAI22_X1 U10475 ( .A1(n9381), .A2(n9200), .B1(n9199), .B2(n9388), .ZN(n9365)
         );
  NAND2_X1 U10476 ( .A1(n9326), .A2(n9309), .ZN(n9205) );
  OAI21_X1 U10477 ( .B1(n9252), .B2(n9235), .A(n9245), .ZN(n9211) );
  XNOR2_X1 U10478 ( .A(n9211), .B(n9231), .ZN(n9483) );
  INV_X1 U10479 ( .A(n9483), .ZN(n9243) );
  INV_X1 U10480 ( .A(n9351), .ZN(n9353) );
  INV_X1 U10481 ( .A(n9224), .ZN(n9225) );
  NAND3_X1 U10482 ( .A1(n9254), .A2(n9256), .A3(n9253), .ZN(n9255) );
  INV_X1 U10483 ( .A(n9231), .ZN(n9232) );
  AOI21_X1 U10484 ( .B1(n9237), .B2(n9248), .A(n9236), .ZN(n9486) );
  NAND2_X1 U10485 ( .A1(n9486), .A2(n9429), .ZN(n9240) );
  AOI22_X1 U10486 ( .A1(n9305), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9238), .B2(
        n9444), .ZN(n9239) );
  OAI211_X1 U10487 ( .C1(n9484), .C2(n9467), .A(n9240), .B(n9239), .ZN(n9241)
         );
  AOI21_X1 U10488 ( .B1(n9485), .B2(n9460), .A(n9241), .ZN(n9242) );
  OAI21_X1 U10489 ( .B1(n9243), .B2(n9450), .A(n9242), .ZN(P1_U3355) );
  INV_X1 U10490 ( .A(n9244), .ZN(n9247) );
  OAI21_X1 U10491 ( .B1(n9247), .B2(n9246), .A(n9245), .ZN(n9492) );
  INV_X1 U10492 ( .A(n9248), .ZN(n9249) );
  AOI21_X1 U10493 ( .B1(n9488), .B2(n9264), .A(n9249), .ZN(n9489) );
  AOI22_X1 U10494 ( .A1(n9305), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9250), .B2(
        n9444), .ZN(n9251) );
  OAI21_X1 U10495 ( .B1(n9252), .B2(n9467), .A(n9251), .ZN(n9261) );
  AND2_X1 U10496 ( .A1(n9254), .A2(n9253), .ZN(n9257) );
  OAI21_X1 U10497 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9259) );
  AOI211_X1 U10498 ( .C1(n9489), .C2(n9429), .A(n9261), .B(n9260), .ZN(n9262)
         );
  OAI21_X1 U10499 ( .B1(n9492), .B2(n9450), .A(n9262), .ZN(P1_U3263) );
  XOR2_X1 U10500 ( .A(n9263), .B(n9271), .Z(n9497) );
  INV_X1 U10501 ( .A(n9278), .ZN(n9266) );
  INV_X1 U10502 ( .A(n9264), .ZN(n9265) );
  AOI21_X1 U10503 ( .B1(n9493), .B2(n9266), .A(n9265), .ZN(n9494) );
  AOI22_X1 U10504 ( .A1(n9305), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9267), .B2(
        n9444), .ZN(n9268) );
  OAI21_X1 U10505 ( .B1(n9269), .B2(n9467), .A(n9268), .ZN(n9276) );
  XOR2_X1 U10506 ( .A(n9271), .B(n9270), .Z(n9274) );
  AOI211_X1 U10507 ( .C1(n9429), .C2(n9494), .A(n9276), .B(n9275), .ZN(n9277)
         );
  OAI21_X1 U10508 ( .B1(n9497), .B2(n9450), .A(n9277), .ZN(P1_U3264) );
  XNOR2_X1 U10509 ( .A(n4381), .B(n9284), .ZN(n9502) );
  AOI21_X1 U10510 ( .B1(n9498), .B2(n4575), .A(n9278), .ZN(n9499) );
  AOI22_X1 U10511 ( .A1(n9305), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9279), .B2(
        n9444), .ZN(n9280) );
  OAI21_X1 U10512 ( .B1(n9281), .B2(n9467), .A(n9280), .ZN(n9289) );
  NAND2_X1 U10513 ( .A1(n9283), .A2(n9282), .ZN(n9285) );
  XNOR2_X1 U10514 ( .A(n9285), .B(n9284), .ZN(n9287) );
  AOI222_X1 U10515 ( .A1(n9459), .A2(n9287), .B1(n9286), .B2(n9456), .C1(n9209), .C2(n9454), .ZN(n9501) );
  NOR2_X1 U10516 ( .A1(n9501), .A2(n9305), .ZN(n9288) );
  AOI211_X1 U10517 ( .C1(n9499), .C2(n9429), .A(n9289), .B(n9288), .ZN(n9290)
         );
  OAI21_X1 U10518 ( .B1(n9502), .B2(n9450), .A(n9290), .ZN(P1_U3265) );
  XOR2_X1 U10519 ( .A(n9293), .B(n9291), .Z(n9507) );
  AOI22_X1 U10520 ( .A1(n9505), .A2(n9374), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9305), .ZN(n9302) );
  XOR2_X1 U10521 ( .A(n9293), .B(n9292), .Z(n9294) );
  OAI222_X1 U10522 ( .A1(n9440), .A2(n9295), .B1(n9438), .B2(n9330), .C1(n9436), .C2(n9294), .ZN(n9503) );
  AOI211_X1 U10523 ( .C1(n9505), .C2(n9311), .A(n9775), .B(n9296), .ZN(n9504)
         );
  INV_X1 U10524 ( .A(n9504), .ZN(n9299) );
  INV_X1 U10525 ( .A(n9297), .ZN(n9298) );
  OAI22_X1 U10526 ( .A1(n9299), .A2(n9315), .B1(n9298), .B2(n9465), .ZN(n9300)
         );
  OAI21_X1 U10527 ( .B1(n9503), .B2(n9300), .A(n9460), .ZN(n9301) );
  OAI211_X1 U10528 ( .C1(n9507), .C2(n9450), .A(n9302), .B(n9301), .ZN(
        P1_U3266) );
  XNOR2_X1 U10529 ( .A(n9304), .B(n9303), .ZN(n9512) );
  AOI22_X1 U10530 ( .A1(n9510), .A2(n9374), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9305), .ZN(n9319) );
  XNOR2_X1 U10531 ( .A(n9307), .B(n9306), .ZN(n9308) );
  OAI222_X1 U10532 ( .A1(n9440), .A2(n9310), .B1(n9438), .B2(n9309), .C1(n9308), .C2(n9436), .ZN(n9508) );
  INV_X1 U10533 ( .A(n9311), .ZN(n9312) );
  AOI211_X1 U10534 ( .C1(n9510), .C2(n9321), .A(n9775), .B(n9312), .ZN(n9509)
         );
  INV_X1 U10535 ( .A(n9509), .ZN(n9316) );
  INV_X1 U10536 ( .A(n9313), .ZN(n9314) );
  OAI22_X1 U10537 ( .A1(n9316), .A2(n9315), .B1(n9314), .B2(n9465), .ZN(n9317)
         );
  OAI21_X1 U10538 ( .B1(n9508), .B2(n9317), .A(n9460), .ZN(n9318) );
  OAI211_X1 U10539 ( .C1(n9512), .C2(n9450), .A(n9319), .B(n9318), .ZN(
        P1_U3267) );
  XNOR2_X1 U10540 ( .A(n9320), .B(n9329), .ZN(n9517) );
  INV_X1 U10541 ( .A(n9337), .ZN(n9323) );
  INV_X1 U10542 ( .A(n9321), .ZN(n9322) );
  AOI21_X1 U10543 ( .B1(n9513), .B2(n9323), .A(n9322), .ZN(n9514) );
  AOI22_X1 U10544 ( .A1(n9305), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9324), .B2(
        n9444), .ZN(n9325) );
  OAI21_X1 U10545 ( .B1(n9326), .B2(n9467), .A(n9325), .ZN(n9334) );
  AOI211_X1 U10546 ( .C1(n9329), .C2(n9328), .A(n9436), .B(n9327), .ZN(n9332)
         );
  OAI22_X1 U10547 ( .A1(n9356), .A2(n9438), .B1(n9330), .B2(n9440), .ZN(n9331)
         );
  NOR2_X1 U10548 ( .A1(n9332), .A2(n9331), .ZN(n9516) );
  NOR2_X1 U10549 ( .A1(n9516), .A2(n9305), .ZN(n9333) );
  AOI211_X1 U10550 ( .C1(n9514), .C2(n9429), .A(n9334), .B(n9333), .ZN(n9335)
         );
  OAI21_X1 U10551 ( .B1(n9517), .B2(n9450), .A(n9335), .ZN(P1_U3268) );
  XOR2_X1 U10552 ( .A(n9336), .B(n9344), .Z(n9522) );
  INV_X1 U10553 ( .A(n9358), .ZN(n9338) );
  AOI211_X1 U10554 ( .C1(n9519), .C2(n9338), .A(n9775), .B(n9337), .ZN(n9518)
         );
  AOI22_X1 U10555 ( .A1(n9305), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9339), .B2(
        n9444), .ZN(n9340) );
  OAI21_X1 U10556 ( .B1(n9341), .B2(n9467), .A(n9340), .ZN(n9348) );
  OAI21_X1 U10557 ( .B1(n9344), .B2(n9343), .A(n9342), .ZN(n9346) );
  AOI222_X1 U10558 ( .A1(n9459), .A2(n9346), .B1(n9369), .B2(n9454), .C1(n9345), .C2(n9456), .ZN(n9521) );
  NOR2_X1 U10559 ( .A1(n9521), .A2(n9305), .ZN(n9347) );
  AOI211_X1 U10560 ( .C1(n9518), .C2(n9469), .A(n9348), .B(n9347), .ZN(n9349)
         );
  OAI21_X1 U10561 ( .B1(n9522), .B2(n9450), .A(n9349), .ZN(P1_U3269) );
  OAI21_X1 U10562 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9527) );
  XNOR2_X1 U10563 ( .A(n9354), .B(n9353), .ZN(n9355) );
  OAI222_X1 U10564 ( .A1(n9438), .A2(n9357), .B1(n9440), .B2(n9356), .C1(n9436), .C2(n9355), .ZN(n9523) );
  AOI211_X1 U10565 ( .C1(n9525), .C2(n9373), .A(n9775), .B(n9358), .ZN(n9524)
         );
  NAND2_X1 U10566 ( .A1(n9524), .A2(n9469), .ZN(n9361) );
  AOI22_X1 U10567 ( .A1(n9305), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9359), .B2(
        n9444), .ZN(n9360) );
  OAI211_X1 U10568 ( .C1(n9362), .C2(n9467), .A(n9361), .B(n9360), .ZN(n9363)
         );
  AOI21_X1 U10569 ( .B1(n9523), .B2(n9460), .A(n9363), .ZN(n9364) );
  OAI21_X1 U10570 ( .B1(n9527), .B2(n9450), .A(n9364), .ZN(P1_U3270) );
  XOR2_X1 U10571 ( .A(n9368), .B(n9365), .Z(n9532) );
  NOR2_X1 U10572 ( .A1(n9390), .A2(n9366), .ZN(n9367) );
  XOR2_X1 U10573 ( .A(n9368), .B(n9367), .Z(n9370) );
  AOI222_X1 U10574 ( .A1(n9459), .A2(n9370), .B1(n9369), .B2(n9456), .C1(n9402), .C2(n9454), .ZN(n9531) );
  OAI21_X1 U10575 ( .B1(n9371), .B2(n9465), .A(n9531), .ZN(n9379) );
  NAND2_X1 U10576 ( .A1(n9382), .A2(n9528), .ZN(n9372) );
  AND2_X1 U10577 ( .A1(n9373), .A2(n9372), .ZN(n9529) );
  INV_X1 U10578 ( .A(n9529), .ZN(n9377) );
  AOI22_X1 U10579 ( .A1(n9528), .A2(n9374), .B1(n9305), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9375) );
  OAI21_X1 U10580 ( .B1(n9377), .B2(n9376), .A(n9375), .ZN(n9378) );
  AOI21_X1 U10581 ( .B1(n9379), .B2(n9460), .A(n9378), .ZN(n9380) );
  OAI21_X1 U10582 ( .B1(n9532), .B2(n9450), .A(n9380), .ZN(P1_U3271) );
  XNOR2_X1 U10583 ( .A(n9381), .B(n9393), .ZN(n9537) );
  INV_X1 U10584 ( .A(n9405), .ZN(n9384) );
  INV_X1 U10585 ( .A(n9382), .ZN(n9383) );
  AOI21_X1 U10586 ( .B1(n9533), .B2(n9384), .A(n9383), .ZN(n9534) );
  INV_X1 U10587 ( .A(n9385), .ZN(n9386) );
  AOI22_X1 U10588 ( .A1(n9305), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9386), .B2(
        n9444), .ZN(n9387) );
  OAI21_X1 U10589 ( .B1(n9388), .B2(n9467), .A(n9387), .ZN(n9397) );
  INV_X1 U10590 ( .A(n9389), .ZN(n9392) );
  INV_X1 U10591 ( .A(n9390), .ZN(n9391) );
  OAI21_X1 U10592 ( .B1(n9393), .B2(n9392), .A(n9391), .ZN(n9395) );
  AOI222_X1 U10593 ( .A1(n9459), .A2(n9395), .B1(n9394), .B2(n9456), .C1(n9425), .C2(n9454), .ZN(n9536) );
  NOR2_X1 U10594 ( .A1(n9536), .A2(n9305), .ZN(n9396) );
  AOI211_X1 U10595 ( .C1(n9534), .C2(n9429), .A(n9397), .B(n9396), .ZN(n9398)
         );
  OAI21_X1 U10596 ( .B1(n9450), .B2(n9537), .A(n9398), .ZN(P1_U3272) );
  NAND2_X1 U10597 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  XOR2_X1 U10598 ( .A(n9410), .B(n9401), .Z(n9404) );
  AOI222_X1 U10599 ( .A1(n9459), .A2(n9404), .B1(n9403), .B2(n9454), .C1(n9402), .C2(n9456), .ZN(n9542) );
  AOI21_X1 U10600 ( .B1(n9539), .B2(n9417), .A(n9405), .ZN(n9540) );
  AOI22_X1 U10601 ( .A1(n9305), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9406), .B2(
        n9444), .ZN(n9407) );
  OAI21_X1 U10602 ( .B1(n9408), .B2(n9467), .A(n9407), .ZN(n9409) );
  AOI21_X1 U10603 ( .B1(n9540), .B2(n9429), .A(n9409), .ZN(n9414) );
  INV_X1 U10604 ( .A(n9544), .ZN(n9412) );
  NAND2_X1 U10605 ( .A1(n9411), .A2(n9410), .ZN(n9538) );
  NAND3_X1 U10606 ( .A1(n9412), .A2(n9472), .A3(n9538), .ZN(n9413) );
  OAI211_X1 U10607 ( .C1(n9542), .C2(n9305), .A(n9414), .B(n9413), .ZN(
        P1_U3273) );
  XNOR2_X1 U10608 ( .A(n9416), .B(n9415), .ZN(n9549) );
  INV_X1 U10609 ( .A(n9417), .ZN(n9418) );
  AOI21_X1 U10610 ( .B1(n9545), .B2(n9441), .A(n9418), .ZN(n9546) );
  AOI22_X1 U10611 ( .A1(n9305), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9419), .B2(
        n9444), .ZN(n9420) );
  OAI21_X1 U10612 ( .B1(n9421), .B2(n9467), .A(n9420), .ZN(n9428) );
  XNOR2_X1 U10613 ( .A(n9423), .B(n9422), .ZN(n9426) );
  AOI222_X1 U10614 ( .A1(n9459), .A2(n9426), .B1(n9425), .B2(n9456), .C1(n9424), .C2(n9454), .ZN(n9548) );
  NOR2_X1 U10615 ( .A1(n9548), .A2(n9305), .ZN(n9427) );
  AOI211_X1 U10616 ( .C1(n9546), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9430)
         );
  OAI21_X1 U10617 ( .B1(n9450), .B2(n9549), .A(n9430), .ZN(P1_U3274) );
  XNOR2_X1 U10618 ( .A(n9431), .B(n9433), .ZN(n9554) );
  AOI21_X1 U10619 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9435) );
  OAI222_X1 U10620 ( .A1(n9440), .A2(n9439), .B1(n9438), .B2(n9437), .C1(n9436), .C2(n9435), .ZN(n9550) );
  INV_X1 U10621 ( .A(n9441), .ZN(n9442) );
  AOI211_X1 U10622 ( .C1(n9552), .C2(n9443), .A(n9775), .B(n9442), .ZN(n9551)
         );
  NAND2_X1 U10623 ( .A1(n9551), .A2(n9469), .ZN(n9447) );
  AOI22_X1 U10624 ( .A1(n9305), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9445), .B2(
        n9444), .ZN(n9446) );
  OAI211_X1 U10625 ( .C1(n4569), .C2(n9467), .A(n9447), .B(n9446), .ZN(n9448)
         );
  AOI21_X1 U10626 ( .B1(n9550), .B2(n9460), .A(n9448), .ZN(n9449) );
  OAI21_X1 U10627 ( .B1(n9450), .B2(n9554), .A(n9449), .ZN(P1_U3275) );
  NAND2_X1 U10628 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  XOR2_X1 U10629 ( .A(n9470), .B(n9453), .Z(n9458) );
  AOI222_X1 U10630 ( .A1(n9459), .A2(n9458), .B1(n9457), .B2(n9456), .C1(n9455), .C2(n9454), .ZN(n9745) );
  MUX2_X1 U10631 ( .A(n6256), .B(n9745), .S(n9460), .Z(n9475) );
  INV_X1 U10632 ( .A(n9461), .ZN(n9462) );
  AOI211_X1 U10633 ( .C1(n9740), .C2(n9463), .A(n9775), .B(n9462), .ZN(n9739)
         );
  OAI22_X1 U10634 ( .A1(n9467), .A2(n9466), .B1(n9465), .B2(n9464), .ZN(n9468)
         );
  AOI21_X1 U10635 ( .B1(n9739), .B2(n9469), .A(n9468), .ZN(n9474) );
  NAND2_X1 U10636 ( .A1(n9471), .A2(n9470), .ZN(n9741) );
  NAND3_X1 U10637 ( .A1(n9742), .A2(n9741), .A3(n9472), .ZN(n9473) );
  NAND3_X1 U10638 ( .A1(n9475), .A2(n9474), .A3(n9473), .ZN(P1_U3286) );
  AOI21_X1 U10639 ( .B1(n9476), .B2(n9748), .A(n9479), .ZN(n9477) );
  OAI21_X1 U10640 ( .B1(n9478), .B2(n9775), .A(n9477), .ZN(n9563) );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9563), .S(n9802), .Z(
        P1_U3554) );
  AOI21_X1 U10642 ( .B1(n9480), .B2(n9748), .A(n9479), .ZN(n9481) );
  OAI21_X1 U10643 ( .B1(n9482), .B2(n9775), .A(n9481), .ZN(n9564) );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9564), .S(n9802), .Z(
        P1_U3553) );
  NAND2_X1 U10645 ( .A1(n9483), .A2(n9770), .ZN(n9487) );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9565), .S(n9802), .Z(
        P1_U3552) );
  AOI22_X1 U10647 ( .A1(n9489), .A2(n9749), .B1(n9748), .B2(n9488), .ZN(n9490)
         );
  OAI211_X1 U10648 ( .C1(n9492), .C2(n9655), .A(n9491), .B(n9490), .ZN(n9566)
         );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9566), .S(n9802), .Z(
        P1_U3551) );
  AOI22_X1 U10650 ( .A1(n9494), .A2(n9749), .B1(n9748), .B2(n9493), .ZN(n9495)
         );
  OAI211_X1 U10651 ( .C1(n9497), .C2(n9655), .A(n9496), .B(n9495), .ZN(n9567)
         );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9567), .S(n9802), .Z(
        P1_U3550) );
  AOI22_X1 U10653 ( .A1(n9499), .A2(n9749), .B1(n9748), .B2(n9498), .ZN(n9500)
         );
  OAI211_X1 U10654 ( .C1(n9502), .C2(n9655), .A(n9501), .B(n9500), .ZN(n9568)
         );
  MUX2_X1 U10655 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9568), .S(n9802), .Z(
        P1_U3549) );
  AOI211_X1 U10656 ( .C1(n9748), .C2(n9505), .A(n9504), .B(n9503), .ZN(n9506)
         );
  OAI21_X1 U10657 ( .B1(n9507), .B2(n9655), .A(n9506), .ZN(n9569) );
  MUX2_X1 U10658 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9569), .S(n9802), .Z(
        P1_U3548) );
  AOI211_X1 U10659 ( .C1(n9748), .C2(n9510), .A(n9509), .B(n9508), .ZN(n9511)
         );
  OAI21_X1 U10660 ( .B1(n9512), .B2(n9655), .A(n9511), .ZN(n9570) );
  MUX2_X1 U10661 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9570), .S(n9802), .Z(
        P1_U3547) );
  AOI22_X1 U10662 ( .A1(n9514), .A2(n9749), .B1(n9748), .B2(n9513), .ZN(n9515)
         );
  OAI211_X1 U10663 ( .C1(n9517), .C2(n9655), .A(n9516), .B(n9515), .ZN(n9571)
         );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9571), .S(n9802), .Z(
        P1_U3546) );
  AOI21_X1 U10665 ( .B1(n9748), .B2(n9519), .A(n9518), .ZN(n9520) );
  OAI211_X1 U10666 ( .C1(n9522), .C2(n9655), .A(n9521), .B(n9520), .ZN(n9572)
         );
  MUX2_X1 U10667 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9572), .S(n9802), .Z(
        P1_U3545) );
  AOI211_X1 U10668 ( .C1(n9748), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9526)
         );
  OAI21_X1 U10669 ( .B1(n9527), .B2(n9655), .A(n9526), .ZN(n9573) );
  MUX2_X1 U10670 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9573), .S(n9802), .Z(
        P1_U3544) );
  AOI22_X1 U10671 ( .A1(n9529), .A2(n9749), .B1(n9748), .B2(n9528), .ZN(n9530)
         );
  OAI211_X1 U10672 ( .C1(n9532), .C2(n9655), .A(n9531), .B(n9530), .ZN(n9574)
         );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9574), .S(n9802), .Z(
        P1_U3543) );
  AOI22_X1 U10674 ( .A1(n9534), .A2(n9749), .B1(n9748), .B2(n9533), .ZN(n9535)
         );
  OAI211_X1 U10675 ( .C1(n9537), .C2(n9655), .A(n9536), .B(n9535), .ZN(n9575)
         );
  MUX2_X1 U10676 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9575), .S(n9802), .Z(
        P1_U3542) );
  NAND2_X1 U10677 ( .A1(n9538), .A2(n9770), .ZN(n9543) );
  AOI22_X1 U10678 ( .A1(n9540), .A2(n9749), .B1(n9748), .B2(n9539), .ZN(n9541)
         );
  OAI211_X1 U10679 ( .C1(n9544), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9576)
         );
  MUX2_X1 U10680 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9576), .S(n9802), .Z(
        P1_U3541) );
  AOI22_X1 U10681 ( .A1(n9546), .A2(n9749), .B1(n9748), .B2(n9545), .ZN(n9547)
         );
  OAI211_X1 U10682 ( .C1(n9549), .C2(n9655), .A(n9548), .B(n9547), .ZN(n9577)
         );
  MUX2_X1 U10683 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9577), .S(n9802), .Z(
        P1_U3540) );
  AOI211_X1 U10684 ( .C1(n9748), .C2(n9552), .A(n9551), .B(n9550), .ZN(n9553)
         );
  OAI21_X1 U10685 ( .B1(n9655), .B2(n9554), .A(n9553), .ZN(n9578) );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9578), .S(n9802), .Z(
        P1_U3539) );
  AOI21_X1 U10687 ( .B1(n9748), .B2(n9556), .A(n9555), .ZN(n9557) );
  OAI211_X1 U10688 ( .C1(n9559), .C2(n9753), .A(n9558), .B(n9557), .ZN(n9579)
         );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9579), .S(n9802), .Z(
        P1_U3533) );
  OAI21_X1 U10690 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9580) );
  MUX2_X1 U10691 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9580), .S(n9802), .Z(
        P1_U3523) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9563), .S(n9784), .Z(
        P1_U3522) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9564), .S(n9784), .Z(
        P1_U3521) );
  MUX2_X1 U10694 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9565), .S(n9784), .Z(
        P1_U3520) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9566), .S(n9784), .Z(
        P1_U3519) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9567), .S(n9784), .Z(
        P1_U3518) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9568), .S(n9784), .Z(
        P1_U3517) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9569), .S(n9784), .Z(
        P1_U3516) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9570), .S(n9784), .Z(
        P1_U3515) );
  MUX2_X1 U10700 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9571), .S(n9784), .Z(
        P1_U3514) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9572), .S(n9784), .Z(
        P1_U3513) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9573), .S(n9784), .Z(
        P1_U3512) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9574), .S(n9784), .Z(
        P1_U3511) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9575), .S(n9784), .Z(
        P1_U3510) );
  MUX2_X1 U10705 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9576), .S(n9784), .Z(
        P1_U3508) );
  MUX2_X1 U10706 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9577), .S(n9784), .Z(
        P1_U3505) );
  MUX2_X1 U10707 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9578), .S(n9784), .Z(
        P1_U3502) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9579), .S(n9784), .Z(
        P1_U3484) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_0__SCAN_IN), .B(n9580), .S(n9784), .Z(
        P1_U3454) );
  MUX2_X1 U10710 ( .A(n9581), .B(P1_D_REG_0__SCAN_IN), .S(n9711), .Z(P1_U3440)
         );
  INV_X1 U10711 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9582) );
  NAND3_X1 U10712 ( .A1(n9582), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9583) );
  OAI22_X1 U10713 ( .A1(n9584), .A2(n9583), .B1(n6304), .B2(n9593), .ZN(n9585)
         );
  AOI21_X1 U10714 ( .B1(n9586), .B2(n9588), .A(n9585), .ZN(n9587) );
  INV_X1 U10715 ( .A(n9587), .ZN(P1_U3322) );
  NAND2_X1 U10716 ( .A1(n9589), .A2(n9588), .ZN(n9591) );
  OAI211_X1 U10717 ( .C1(n9593), .C2(n9592), .A(n9591), .B(n9590), .ZN(
        P1_U3325) );
  AOI21_X1 U10718 ( .B1(n9595), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9594), .ZN(
        n9596) );
  OAI21_X1 U10719 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(P1_U3326) );
  INV_X1 U10720 ( .A(n9599), .ZN(n9608) );
  OAI22_X1 U10721 ( .A1(n9602), .A2(n9601), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9600), .ZN(n9607) );
  NAND2_X1 U10722 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9605) );
  AOI211_X1 U10723 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9614), .ZN(n9606)
         );
  AOI211_X1 U10724 ( .C1(n9620), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9613)
         );
  NOR2_X1 U10725 ( .A1(n9812), .A2(n5672), .ZN(n9611) );
  OAI211_X1 U10726 ( .C1(n9611), .C2(n9610), .A(n9803), .B(n9609), .ZN(n9612)
         );
  NAND2_X1 U10727 ( .A1(n9613), .A2(n9612), .ZN(P2_U3246) );
  AOI22_X1 U10728 ( .A1(n9809), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9626) );
  AOI211_X1 U10729 ( .C1(n9617), .C2(n9616), .A(n9615), .B(n9614), .ZN(n9618)
         );
  AOI21_X1 U10730 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9625) );
  OAI211_X1 U10731 ( .C1(n9623), .C2(n9622), .A(n9803), .B(n9621), .ZN(n9624)
         );
  NAND3_X1 U10732 ( .A1(n9626), .A2(n9625), .A3(n9624), .ZN(P2_U3247) );
  OAI22_X1 U10733 ( .A1(n9628), .A2(n9917), .B1(n9627), .B2(n9915), .ZN(n9630)
         );
  AOI211_X1 U10734 ( .C1(n9631), .C2(n9921), .A(n9630), .B(n9629), .ZN(n9633)
         );
  AOI22_X1 U10735 ( .A1(n9939), .A2(n9633), .B1(n5896), .B2(n9937), .ZN(
        P2_U3534) );
  INV_X1 U10736 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9632) );
  AOI22_X1 U10737 ( .A1(n9924), .A2(n9633), .B1(n9632), .B2(n9923), .ZN(
        P2_U3493) );
  OAI22_X1 U10738 ( .A1(n9635), .A2(n9775), .B1(n9634), .B2(n9773), .ZN(n9636)
         );
  AOI21_X1 U10739 ( .B1(n9637), .B2(n9781), .A(n9636), .ZN(n9638) );
  AND2_X1 U10740 ( .A1(n9639), .A2(n9638), .ZN(n9660) );
  AOI22_X1 U10741 ( .A1(n9802), .A2(n9660), .B1(n9640), .B2(n9799), .ZN(
        P1_U3538) );
  OAI21_X1 U10742 ( .B1(n9642), .B2(n9773), .A(n9641), .ZN(n9643) );
  AOI211_X1 U10743 ( .C1(n9645), .C2(n9770), .A(n9644), .B(n9643), .ZN(n9662)
         );
  AOI22_X1 U10744 ( .A1(n9802), .A2(n9662), .B1(n6852), .B2(n9799), .ZN(
        P1_U3537) );
  OAI22_X1 U10745 ( .A1(n9647), .A2(n9775), .B1(n9646), .B2(n9773), .ZN(n9649)
         );
  AOI211_X1 U10746 ( .C1(n9781), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9664)
         );
  AOI22_X1 U10747 ( .A1(n9802), .A2(n9664), .B1(n6572), .B2(n9799), .ZN(
        P1_U3536) );
  AOI22_X1 U10748 ( .A1(n9652), .A2(n9749), .B1(n9748), .B2(n9651), .ZN(n9653)
         );
  OAI211_X1 U10749 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9657)
         );
  INV_X1 U10750 ( .A(n9657), .ZN(n9666) );
  AOI22_X1 U10751 ( .A1(n9802), .A2(n9666), .B1(n9658), .B2(n9799), .ZN(
        P1_U3534) );
  INV_X1 U10752 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9659) );
  INV_X1 U10753 ( .A(n9784), .ZN(n9782) );
  AOI22_X1 U10754 ( .A1(n9784), .A2(n9660), .B1(n9659), .B2(n9782), .ZN(
        P1_U3499) );
  INV_X1 U10755 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9661) );
  AOI22_X1 U10756 ( .A1(n9784), .A2(n9662), .B1(n9661), .B2(n9782), .ZN(
        P1_U3496) );
  INV_X1 U10757 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U10758 ( .A1(n9784), .A2(n9664), .B1(n9663), .B2(n9782), .ZN(
        P1_U3493) );
  INV_X1 U10759 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U10760 ( .A1(n9784), .A2(n9666), .B1(n9665), .B2(n9782), .ZN(
        P1_U3487) );
  XNOR2_X1 U10761 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10762 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10763 ( .A(n9667), .ZN(n9670) );
  INV_X1 U10764 ( .A(n9668), .ZN(n9669) );
  AOI21_X1 U10765 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9681) );
  NAND2_X1 U10766 ( .A1(n9673), .A2(n9672), .ZN(n9675) );
  XNOR2_X1 U10767 ( .A(n9675), .B(n9674), .ZN(n9679) );
  NOR2_X1 U10768 ( .A1(n9676), .A2(n9773), .ZN(n9764) );
  AOI22_X1 U10769 ( .A1(n9679), .A2(n9678), .B1(n9764), .B2(n9677), .ZN(n9680)
         );
  OAI211_X1 U10770 ( .C1(n9683), .C2(n9682), .A(n9681), .B(n9680), .ZN(
        P1_U3219) );
  AOI22_X1 U10771 ( .A1(n9703), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9690) );
  OAI22_X1 U10772 ( .A1(n6268), .A2(n6258), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9687), .ZN(n9685) );
  OAI211_X1 U10773 ( .C1(n9686), .C2(n9685), .A(P1_U3083), .B(n9684), .ZN(
        n9689) );
  NAND3_X1 U10774 ( .A1(n9704), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9687), .ZN(
        n9688) );
  NAND3_X1 U10775 ( .A1(n9690), .A2(n9689), .A3(n9688), .ZN(P1_U3241) );
  NOR2_X1 U10776 ( .A1(n9692), .A2(n9691), .ZN(n9693) );
  NOR3_X1 U10777 ( .A1(n9695), .A2(n9694), .A3(n9693), .ZN(n9696) );
  AOI211_X1 U10778 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(n9707)
         );
  OAI21_X1 U10779 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9705) );
  AOI22_X1 U10780 ( .A1(n9705), .A2(n9704), .B1(n9703), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U10781 ( .A1(n9707), .A2(n9706), .ZN(P1_U3259) );
  AND2_X1 U10782 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9711), .ZN(P1_U3292) );
  AND2_X1 U10783 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9711), .ZN(P1_U3293) );
  AND2_X1 U10784 ( .A1(n9711), .A2(P1_D_REG_29__SCAN_IN), .ZN(P1_U3294) );
  AND2_X1 U10785 ( .A1(n9711), .A2(P1_D_REG_28__SCAN_IN), .ZN(P1_U3295) );
  AND2_X1 U10786 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9711), .ZN(P1_U3296) );
  AND2_X1 U10787 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9711), .ZN(P1_U3297) );
  AND2_X1 U10788 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9711), .ZN(P1_U3298) );
  AND2_X1 U10789 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9711), .ZN(P1_U3299) );
  INV_X1 U10790 ( .A(n9711), .ZN(n9710) );
  NOR2_X1 U10791 ( .A1(n9710), .A2(n9708), .ZN(P1_U3300) );
  AND2_X1 U10792 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9711), .ZN(P1_U3301) );
  AND2_X1 U10793 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9711), .ZN(P1_U3302) );
  AND2_X1 U10794 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9711), .ZN(P1_U3303) );
  AND2_X1 U10795 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9711), .ZN(P1_U3304) );
  AND2_X1 U10796 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9711), .ZN(P1_U3305) );
  AND2_X1 U10797 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9711), .ZN(P1_U3306) );
  AND2_X1 U10798 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9711), .ZN(P1_U3307) );
  AND2_X1 U10799 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9711), .ZN(P1_U3308) );
  AND2_X1 U10800 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9711), .ZN(P1_U3309) );
  NOR2_X1 U10801 ( .A1(n9710), .A2(n9709), .ZN(P1_U3310) );
  AND2_X1 U10802 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9711), .ZN(P1_U3311) );
  AND2_X1 U10803 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9711), .ZN(P1_U3312) );
  AND2_X1 U10804 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9711), .ZN(P1_U3313) );
  AND2_X1 U10805 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9711), .ZN(P1_U3314) );
  AND2_X1 U10806 ( .A1(n9711), .A2(P1_D_REG_8__SCAN_IN), .ZN(P1_U3315) );
  AND2_X1 U10807 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9711), .ZN(P1_U3316) );
  AND2_X1 U10808 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9711), .ZN(P1_U3317) );
  AND2_X1 U10809 ( .A1(n9711), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3318) );
  AND2_X1 U10810 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9711), .ZN(P1_U3319) );
  AND2_X1 U10811 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9711), .ZN(P1_U3320) );
  AND2_X1 U10812 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9711), .ZN(P1_U3321) );
  INV_X1 U10813 ( .A(n9712), .ZN(n9716) );
  INV_X1 U10814 ( .A(n9713), .ZN(n9715) );
  AOI211_X1 U10815 ( .C1(n9781), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9786)
         );
  INV_X1 U10816 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9717) );
  AOI22_X1 U10817 ( .A1(n9784), .A2(n9786), .B1(n9717), .B2(n9782), .ZN(
        P1_U3457) );
  OAI22_X1 U10818 ( .A1(n9719), .A2(n9775), .B1(n9718), .B2(n9773), .ZN(n9722)
         );
  INV_X1 U10819 ( .A(n9720), .ZN(n9721) );
  AOI211_X1 U10820 ( .C1(n9781), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9788)
         );
  INV_X1 U10821 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9724) );
  AOI22_X1 U10822 ( .A1(n9784), .A2(n9788), .B1(n9724), .B2(n9782), .ZN(
        P1_U3460) );
  AOI22_X1 U10823 ( .A1(n9726), .A2(n9749), .B1(n9748), .B2(n9725), .ZN(n9729)
         );
  NAND2_X1 U10824 ( .A1(n9727), .A2(n9770), .ZN(n9728) );
  AND3_X1 U10825 ( .A1(n9730), .A2(n9729), .A3(n9728), .ZN(n9789) );
  AOI22_X1 U10826 ( .A1(n9784), .A2(n9789), .B1(n9731), .B2(n9782), .ZN(
        P1_U3463) );
  OAI22_X1 U10827 ( .A1(n9733), .A2(n9775), .B1(n9732), .B2(n9773), .ZN(n9734)
         );
  AOI21_X1 U10828 ( .B1(n9735), .B2(n9781), .A(n9734), .ZN(n9736) );
  AOI22_X1 U10829 ( .A1(n9784), .A2(n9790), .B1(n9738), .B2(n9782), .ZN(
        P1_U3466) );
  AOI21_X1 U10830 ( .B1(n9748), .B2(n9740), .A(n9739), .ZN(n9744) );
  NAND3_X1 U10831 ( .A1(n9742), .A2(n9741), .A3(n9770), .ZN(n9743) );
  AND3_X1 U10832 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(n9792) );
  INV_X1 U10833 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U10834 ( .A1(n9784), .A2(n9792), .B1(n9746), .B2(n9782), .ZN(
        P1_U3469) );
  AOI22_X1 U10835 ( .A1(n9750), .A2(n9749), .B1(n9748), .B2(n4315), .ZN(n9751)
         );
  OAI211_X1 U10836 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n9751), .ZN(n9755)
         );
  INV_X1 U10837 ( .A(n9755), .ZN(n9794) );
  INV_X1 U10838 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9756) );
  AOI22_X1 U10839 ( .A1(n9784), .A2(n9794), .B1(n9756), .B2(n9782), .ZN(
        P1_U3472) );
  OAI211_X1 U10840 ( .C1(n9759), .C2(n9773), .A(n9758), .B(n9757), .ZN(n9760)
         );
  AOI21_X1 U10841 ( .B1(n9770), .B2(n9761), .A(n9760), .ZN(n9796) );
  INV_X1 U10842 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9762) );
  AOI22_X1 U10843 ( .A1(n9784), .A2(n9796), .B1(n9762), .B2(n9782), .ZN(
        P1_U3475) );
  INV_X1 U10844 ( .A(n9763), .ZN(n9771) );
  INV_X1 U10845 ( .A(n9764), .ZN(n9765) );
  OAI21_X1 U10846 ( .B1(n9766), .B2(n9775), .A(n9765), .ZN(n9769) );
  INV_X1 U10847 ( .A(n9767), .ZN(n9768) );
  AOI211_X1 U10848 ( .C1(n9771), .C2(n9770), .A(n9769), .B(n9768), .ZN(n9798)
         );
  INV_X1 U10849 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10850 ( .A1(n9784), .A2(n9798), .B1(n9772), .B2(n9782), .ZN(
        P1_U3478) );
  OAI22_X1 U10851 ( .A1(n9776), .A2(n9775), .B1(n9774), .B2(n9773), .ZN(n9779)
         );
  INV_X1 U10852 ( .A(n9777), .ZN(n9778) );
  AOI211_X1 U10853 ( .C1(n9781), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9801)
         );
  INV_X1 U10854 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10855 ( .A1(n9784), .A2(n9801), .B1(n9783), .B2(n9782), .ZN(
        P1_U3481) );
  AOI22_X1 U10856 ( .A1(n9802), .A2(n9786), .B1(n9785), .B2(n9799), .ZN(
        P1_U3524) );
  AOI22_X1 U10857 ( .A1(n9802), .A2(n9788), .B1(n9787), .B2(n9799), .ZN(
        P1_U3525) );
  AOI22_X1 U10858 ( .A1(n9802), .A2(n9789), .B1(n5116), .B2(n9799), .ZN(
        P1_U3526) );
  AOI22_X1 U10859 ( .A1(n9802), .A2(n9790), .B1(n5133), .B2(n9799), .ZN(
        P1_U3527) );
  INV_X1 U10860 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9791) );
  AOI22_X1 U10861 ( .A1(n9802), .A2(n9792), .B1(n9791), .B2(n9799), .ZN(
        P1_U3528) );
  INV_X1 U10862 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10863 ( .A1(n9802), .A2(n9794), .B1(n9793), .B2(n9799), .ZN(
        P1_U3529) );
  INV_X1 U10864 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U10865 ( .A1(n9802), .A2(n9796), .B1(n9795), .B2(n9799), .ZN(
        P1_U3530) );
  INV_X1 U10866 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U10867 ( .A1(n9802), .A2(n9798), .B1(n9797), .B2(n9799), .ZN(
        P1_U3531) );
  INV_X1 U10868 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U10869 ( .A1(n9802), .A2(n9801), .B1(n9800), .B2(n9799), .ZN(
        P1_U3532) );
  AOI22_X1 U10870 ( .A1(n9803), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9804), .ZN(n9813) );
  NAND2_X1 U10871 ( .A1(n9804), .A2(n9925), .ZN(n9805) );
  OAI211_X1 U10872 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9807), .A(n9806), .B(
        n9805), .ZN(n9808) );
  INV_X1 U10873 ( .A(n9808), .ZN(n9811) );
  AOI22_X1 U10874 ( .A1(n9809), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9810) );
  OAI221_X1 U10875 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9813), .C1(n9812), .C2(
        n9811), .A(n9810), .ZN(P2_U3245) );
  AOI21_X1 U10876 ( .B1(n9816), .B2(n9823), .A(n9815), .ZN(n9819) );
  AOI21_X1 U10877 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(n9878) );
  NAND2_X1 U10878 ( .A1(n7008), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U10879 ( .A1(n9822), .A2(n9821), .ZN(n9824) );
  XNOR2_X1 U10880 ( .A(n9824), .B(n9823), .ZN(n9881) );
  INV_X1 U10881 ( .A(n9825), .ZN(n9835) );
  XNOR2_X1 U10882 ( .A(n9826), .B(n9830), .ZN(n9877) );
  OAI22_X1 U10883 ( .A1(n4316), .A2(n6532), .B1(n9828), .B2(n9827), .ZN(n9829)
         );
  AOI21_X1 U10884 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9832) );
  OAI21_X1 U10885 ( .B1(n9833), .B2(n9877), .A(n9832), .ZN(n9834) );
  AOI21_X1 U10886 ( .B1(n9881), .B2(n9835), .A(n9834), .ZN(n9836) );
  OAI21_X1 U10887 ( .B1(n9837), .B2(n9878), .A(n9836), .ZN(P2_U3292) );
  AND2_X1 U10888 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9844), .ZN(P2_U3297) );
  AND2_X1 U10889 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9844), .ZN(P2_U3298) );
  AND2_X1 U10890 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9844), .ZN(P2_U3299) );
  AND2_X1 U10891 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9844), .ZN(P2_U3300) );
  AND2_X1 U10892 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9844), .ZN(P2_U3301) );
  AND2_X1 U10893 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9844), .ZN(P2_U3302) );
  AND2_X1 U10894 ( .A1(n9844), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3303) );
  AND2_X1 U10895 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9844), .ZN(P2_U3304) );
  AND2_X1 U10896 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9844), .ZN(P2_U3305) );
  AND2_X1 U10897 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9844), .ZN(P2_U3306) );
  AND2_X1 U10898 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9844), .ZN(P2_U3307) );
  AND2_X1 U10899 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9844), .ZN(P2_U3308) );
  AND2_X1 U10900 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9844), .ZN(P2_U3309) );
  AND2_X1 U10901 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9844), .ZN(P2_U3310) );
  AND2_X1 U10902 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9844), .ZN(P2_U3311) );
  AND2_X1 U10903 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9844), .ZN(P2_U3312) );
  AND2_X1 U10904 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9844), .ZN(P2_U3313) );
  AND2_X1 U10905 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9844), .ZN(P2_U3314) );
  AND2_X1 U10906 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9844), .ZN(P2_U3315) );
  AND2_X1 U10907 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9844), .ZN(P2_U3316) );
  AND2_X1 U10908 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9844), .ZN(P2_U3317) );
  AND2_X1 U10909 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9844), .ZN(P2_U3318) );
  AND2_X1 U10910 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9844), .ZN(P2_U3319) );
  AND2_X1 U10911 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9844), .ZN(P2_U3320) );
  AND2_X1 U10912 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9844), .ZN(P2_U3321) );
  NOR2_X1 U10913 ( .A1(n9841), .A2(n9840), .ZN(P2_U3322) );
  AND2_X1 U10914 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9844), .ZN(P2_U3323) );
  AND2_X1 U10915 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9844), .ZN(P2_U3324) );
  AND2_X1 U10916 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9844), .ZN(P2_U3325) );
  AND2_X1 U10917 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9844), .ZN(P2_U3326) );
  AOI22_X1 U10918 ( .A1(n9847), .A2(n9843), .B1(n9842), .B2(n9844), .ZN(
        P2_U3437) );
  AOI22_X1 U10919 ( .A1(n9847), .A2(n9846), .B1(n9845), .B2(n9844), .ZN(
        P2_U3438) );
  OAI21_X1 U10920 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  AOI21_X1 U10921 ( .B1(n9921), .B2(n9852), .A(n9851), .ZN(n9926) );
  AOI22_X1 U10922 ( .A1(n9924), .A2(n9926), .B1(n5671), .B2(n9923), .ZN(
        P2_U3451) );
  INV_X1 U10923 ( .A(n9853), .ZN(n9860) );
  NAND3_X1 U10924 ( .A1(n9855), .A2(n9868), .A3(n9854), .ZN(n9856) );
  OAI211_X1 U10925 ( .C1(n9858), .C2(n9915), .A(n9857), .B(n9856), .ZN(n9859)
         );
  AOI21_X1 U10926 ( .B1(n9921), .B2(n9860), .A(n9859), .ZN(n9927) );
  INV_X1 U10927 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U10928 ( .A1(n9924), .A2(n9927), .B1(n9861), .B2(n9923), .ZN(
        P2_U3454) );
  OAI22_X1 U10929 ( .A1(n9863), .A2(n9917), .B1(n9862), .B2(n9915), .ZN(n9865)
         );
  AOI211_X1 U10930 ( .C1(n9921), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9928)
         );
  AOI22_X1 U10931 ( .A1(n9924), .A2(n9928), .B1(n5691), .B2(n9923), .ZN(
        P2_U3457) );
  INV_X1 U10932 ( .A(n9867), .ZN(n9913) );
  NAND2_X1 U10933 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  OAI21_X1 U10934 ( .B1(n9871), .B2(n9915), .A(n9870), .ZN(n9873) );
  AOI211_X1 U10935 ( .C1(n9913), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9929)
         );
  INV_X1 U10936 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U10937 ( .A1(n9924), .A2(n9929), .B1(n9875), .B2(n9923), .ZN(
        P2_U3460) );
  OAI22_X1 U10938 ( .A1(n9877), .A2(n9917), .B1(n9876), .B2(n9915), .ZN(n9880)
         );
  INV_X1 U10939 ( .A(n9878), .ZN(n9879) );
  AOI211_X1 U10940 ( .C1(n9921), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9930)
         );
  INV_X1 U10941 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U10942 ( .A1(n9924), .A2(n9930), .B1(n9882), .B2(n9923), .ZN(
        P2_U3463) );
  AOI211_X1 U10943 ( .C1(n9886), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9887)
         );
  OAI21_X1 U10944 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n9890) );
  INV_X1 U10945 ( .A(n9890), .ZN(n9932) );
  INV_X1 U10946 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9891) );
  AOI22_X1 U10947 ( .A1(n9924), .A2(n9932), .B1(n9891), .B2(n9923), .ZN(
        P2_U3466) );
  INV_X1 U10948 ( .A(n9892), .ZN(n9898) );
  INV_X1 U10949 ( .A(n9893), .ZN(n9895) );
  OAI22_X1 U10950 ( .A1(n9895), .A2(n9917), .B1(n9894), .B2(n9915), .ZN(n9897)
         );
  AOI211_X1 U10951 ( .C1(n9898), .C2(n9921), .A(n9897), .B(n9896), .ZN(n9933)
         );
  INV_X1 U10952 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U10953 ( .A1(n9924), .A2(n9933), .B1(n9899), .B2(n9923), .ZN(
        P2_U3469) );
  OAI22_X1 U10954 ( .A1(n9901), .A2(n9917), .B1(n9900), .B2(n9915), .ZN(n9903)
         );
  AOI211_X1 U10955 ( .C1(n9913), .C2(n9904), .A(n9903), .B(n9902), .ZN(n9934)
         );
  INV_X1 U10956 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U10957 ( .A1(n9924), .A2(n9934), .B1(n9905), .B2(n9923), .ZN(
        P2_U3475) );
  INV_X1 U10958 ( .A(n9906), .ZN(n9912) );
  INV_X1 U10959 ( .A(n9907), .ZN(n9908) );
  OAI22_X1 U10960 ( .A1(n9909), .A2(n9917), .B1(n9908), .B2(n9915), .ZN(n9911)
         );
  AOI211_X1 U10961 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n9910), .ZN(n9936)
         );
  INV_X1 U10962 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U10963 ( .A1(n9924), .A2(n9936), .B1(n9914), .B2(n9923), .ZN(
        P2_U3481) );
  OAI22_X1 U10964 ( .A1(n9918), .A2(n9917), .B1(n9916), .B2(n9915), .ZN(n9920)
         );
  AOI211_X1 U10965 ( .C1(n9922), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9938)
         );
  AOI22_X1 U10966 ( .A1(n9924), .A2(n9938), .B1(n5862), .B2(n9923), .ZN(
        P2_U3487) );
  AOI22_X1 U10967 ( .A1(n9939), .A2(n9926), .B1(n9925), .B2(n9937), .ZN(
        P2_U3520) );
  AOI22_X1 U10968 ( .A1(n9939), .A2(n9927), .B1(n6511), .B2(n9937), .ZN(
        P2_U3521) );
  AOI22_X1 U10969 ( .A1(n9939), .A2(n9928), .B1(n6512), .B2(n9937), .ZN(
        P2_U3522) );
  AOI22_X1 U10970 ( .A1(n9939), .A2(n9929), .B1(n5705), .B2(n9937), .ZN(
        P2_U3523) );
  AOI22_X1 U10971 ( .A1(n9939), .A2(n9930), .B1(n5720), .B2(n9937), .ZN(
        P2_U3524) );
  INV_X1 U10972 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U10973 ( .A1(n9939), .A2(n9932), .B1(n9931), .B2(n9937), .ZN(
        P2_U3525) );
  AOI22_X1 U10974 ( .A1(n9939), .A2(n9933), .B1(n5756), .B2(n9937), .ZN(
        P2_U3526) );
  AOI22_X1 U10975 ( .A1(n9939), .A2(n9934), .B1(n5795), .B2(n9937), .ZN(
        P2_U3528) );
  INV_X1 U10976 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U10977 ( .A1(n9939), .A2(n9936), .B1(n9935), .B2(n9937), .ZN(
        P2_U3530) );
  AOI22_X1 U10978 ( .A1(n9939), .A2(n9938), .B1(n5861), .B2(n9937), .ZN(
        P2_U3532) );
  INV_X1 U10979 ( .A(n9940), .ZN(n9941) );
  NAND2_X1 U10980 ( .A1(n9942), .A2(n9941), .ZN(n9943) );
  XNOR2_X1 U10981 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9943), .ZN(ADD_1071_U5) );
  XOR2_X1 U10982 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10983 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(ADD_1071_U56) );
  OAI21_X1 U10984 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(ADD_1071_U57) );
  OAI21_X1 U10985 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(ADD_1071_U58) );
  OAI21_X1 U10986 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(ADD_1071_U59) );
  OAI21_X1 U10987 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(ADD_1071_U60) );
  OAI21_X1 U10988 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(ADD_1071_U61) );
  AOI21_X1 U10989 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(ADD_1071_U62) );
  AOI21_X1 U10990 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(ADD_1071_U63) );
  XOR2_X1 U10991 ( .A(n9968), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  AOI21_X1 U10992 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(ADD_1071_U47) );
  XOR2_X1 U10993 ( .A(n9972), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U10994 ( .A1(n9974), .A2(n9973), .ZN(n9975) );
  XOR2_X1 U10995 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9975), .Z(ADD_1071_U51) );
  OAI21_X1 U10996 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9979) );
  XNOR2_X1 U10997 ( .A(n9979), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U10998 ( .A(n9981), .B(n9980), .Z(ADD_1071_U54) );
  XOR2_X1 U10999 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9982), .Z(ADD_1071_U48) );
  XOR2_X1 U11000 ( .A(n9984), .B(n9983), .Z(ADD_1071_U53) );
  XNOR2_X1 U11001 ( .A(n9986), .B(n9985), .ZN(ADD_1071_U52) );
  OR2_X2 U5807 ( .A1(n9917), .A2(n5654), .ZN(n5678) );
endmodule

