

module b14_C_gen_AntiSAT_k_256_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109;

  NAND4_X1 U2466 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n2982)
         );
  INV_X1 U2467 ( .A(n2954), .ZN(n3518) );
  INV_X2 U2468 ( .A(n3538), .ZN(n2923) );
  AND2_X1 U2469 ( .A1(n2957), .A2(n3040), .ZN(n3536) );
  INV_X2 U2470 ( .A(n3518), .ZN(n2224) );
  NOR2_X1 U2472 ( .A1(n4409), .A2(n3765), .ZN(n2864) );
  AND4_X1 U2473 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n2955)
         );
  MUX2_X1 U2474 ( .A(REG1_REG_29__SCAN_IN), .B(n2868), .S(n4729), .Z(n2863) );
  INV_X1 U2476 ( .A(n3072), .ZN(n3859) );
  OAI21_X2 U2479 ( .B1(n2311), .B2(n3816), .A(n2312), .ZN(n4087) );
  XNOR2_X2 U2480 ( .A(n3938), .B(n3937), .ZN(n4560) );
  NAND2_X2 U2481 ( .A1(n2844), .A2(n2843), .ZN(n2917) );
  NAND2_X2 U2482 ( .A1(n2788), .A2(n3765), .ZN(n3040) );
  BUF_X2 U2483 ( .A(n2518), .Z(n3707) );
  NAND2_X1 U2484 ( .A1(n2499), .A2(n2385), .ZN(n2524) );
  INV_X2 U2485 ( .A(IR_REG_31__SCAN_IN), .ZN(n2823) );
  MUX2_X1 U2486 ( .A(REG1_REG_28__SCAN_IN), .B(n4348), .S(n4729), .Z(n4233) );
  MUX2_X1 U2487 ( .A(REG0_REG_28__SCAN_IN), .B(n4348), .S(n4708), .Z(n4349) );
  NAND2_X1 U2488 ( .A1(n2343), .A2(n2342), .ZN(n3661) );
  OAI21_X1 U2489 ( .B1(n3578), .B2(n2339), .A(n2259), .ZN(n2338) );
  NAND2_X1 U2490 ( .A1(n4010), .A2(n3824), .ZN(n3992) );
  NOR2_X1 U2491 ( .A1(n3326), .A2(n3324), .ZN(n3321) );
  NAND2_X1 U2492 ( .A1(n4522), .A2(n3931), .ZN(n4534) );
  AND2_X1 U2493 ( .A1(n2318), .A2(n2263), .ZN(n2316) );
  NAND2_X1 U2494 ( .A1(n2307), .A2(n2306), .ZN(n4608) );
  AOI21_X1 U2495 ( .B1(REG1_REG_5__SCAN_IN), .B2(n3920), .A(n4442), .ZN(n3921)
         );
  AND4_X1 U2496 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n3072)
         );
  NAND4_X1 U2497 ( .A1(n2548), .A2(n2547), .A3(n2546), .A4(n2545), .ZN(n3858)
         );
  BUF_X2 U2498 ( .A(n2978), .Z(n3508) );
  INV_X2 U2499 ( .A(n3536), .ZN(n3526) );
  NAND3_X1 U2500 ( .A1(n2514), .A2(n2236), .A3(n2513), .ZN(n4611) );
  NAND2_X1 U2501 ( .A1(n2494), .A2(REG2_REG_1__SCAN_IN), .ZN(n2496) );
  CLKBUF_X3 U2502 ( .A(n2512), .Z(n3703) );
  NOR2_X1 U2503 ( .A1(n2912), .A2(n4718), .ZN(n3918) );
  OAI22_X1 U2504 ( .A1(n3891), .A2(n3890), .B1(n3889), .B2(n2295), .ZN(n4448)
         );
  NOR2_X1 U2505 ( .A1(n2938), .A2(n4414), .ZN(n4610) );
  OAI211_X1 U2506 ( .C1(n2298), .C2(n2295), .A(n2246), .B(n2293), .ZN(n2912)
         );
  CLKBUF_X3 U2507 ( .A(n2509), .Z(n2544) );
  NAND2_X2 U2508 ( .A1(n2481), .A2(n2278), .ZN(n3702) );
  INV_X1 U2509 ( .A(n2490), .ZN(n2880) );
  XNOR2_X1 U2510 ( .A(n2778), .B(n2781), .ZN(n3949) );
  XNOR2_X1 U2511 ( .A(n2786), .B(IR_REG_22__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U2512 ( .A1(n2703), .A2(IR_REG_31__SCAN_IN), .ZN(n2778) );
  XNOR2_X1 U2513 ( .A(n2315), .B(n2314), .ZN(n2490) );
  OR2_X1 U2514 ( .A1(n3443), .A2(n2823), .ZN(n2485) );
  NOR2_X1 U2515 ( .A1(n2702), .A2(IR_REG_18__SCAN_IN), .ZN(n2783) );
  NOR2_X1 U2516 ( .A1(n2635), .A2(n2376), .ZN(n2690) );
  NAND2_X1 U2517 ( .A1(n2301), .A2(n2299), .ZN(n2899) );
  AND2_X1 U2518 ( .A1(n2476), .A2(n2453), .ZN(n2451) );
  NOR2_X1 U2519 ( .A1(n2454), .A2(n2235), .ZN(n2453) );
  AND2_X1 U2520 ( .A1(n2467), .A2(n2469), .ZN(n2409) );
  AND3_X1 U2521 ( .A1(n2468), .A2(n2615), .A3(n2623), .ZN(n2469) );
  INV_X1 U2522 ( .A(IR_REG_20__SCAN_IN), .ZN(n2782) );
  INV_X1 U2523 ( .A(IR_REG_10__SCAN_IN), .ZN(n2615) );
  INV_X1 U2524 ( .A(IR_REG_3__SCAN_IN), .ZN(n2532) );
  INV_X1 U2525 ( .A(IR_REG_11__SCAN_IN), .ZN(n2623) );
  INV_X1 U2526 ( .A(IR_REG_13__SCAN_IN), .ZN(n2470) );
  INV_X2 U2527 ( .A(n2978), .ZN(n2922) );
  NAND2_X1 U2528 ( .A1(n4485), .A2(n3926), .ZN(n3927) );
  INV_X1 U2529 ( .A(n2428), .ZN(n2426) );
  INV_X1 U2530 ( .A(n2461), .ZN(n2427) );
  INV_X1 U2531 ( .A(n2812), .ZN(n4049) );
  AOI21_X1 U2532 ( .B1(n3432), .B2(n2463), .A(n2657), .ZN(n4188) );
  INV_X1 U2533 ( .A(n2656), .ZN(n2657) );
  INV_X1 U2534 ( .A(n2635), .ZN(n2471) );
  OR2_X1 U2535 ( .A1(n2482), .A2(IR_REG_28__SCAN_IN), .ZN(n2278) );
  NOR2_X1 U2536 ( .A1(n2358), .A2(n2357), .ZN(n2356) );
  INV_X1 U2537 ( .A(n3511), .ZN(n2358) );
  OAI22_X1 U2538 ( .A1(n4331), .A2(n3538), .B1(n2224), .B2(n4323), .ZN(n3412)
         );
  AND2_X1 U2539 ( .A1(n2487), .A2(n2880), .ZN(n2512) );
  NAND2_X1 U2540 ( .A1(n4407), .A2(n2490), .ZN(n2518) );
  XNOR2_X1 U2541 ( .A(n3903), .B(n4654), .ZN(n4518) );
  NOR2_X1 U2542 ( .A1(n2446), .A2(n2234), .ZN(n2445) );
  INV_X1 U2543 ( .A(n2448), .ZN(n2446) );
  AND2_X1 U2544 ( .A1(n4015), .A2(n4034), .ZN(n2734) );
  NAND2_X1 U2545 ( .A1(n4056), .A2(n4038), .ZN(n2733) );
  AND2_X1 U2546 ( .A1(n2726), .A2(REG3_REG_24__SCAN_IN), .ZN(n2745) );
  NAND2_X1 U2547 ( .A1(n2309), .A2(n2308), .ZN(n3396) );
  INV_X1 U2548 ( .A(n3800), .ZN(n2308) );
  INV_X1 U2549 ( .A(n3782), .ZN(n2321) );
  OAI21_X1 U2550 ( .B1(n2421), .B2(n2418), .A(n2417), .ZN(n3294) );
  NOR2_X1 U2551 ( .A1(n2415), .A2(n2413), .ZN(n2417) );
  OAI22_X1 U2552 ( .A1(n2418), .A2(n3280), .B1(n3195), .B2(n3854), .ZN(n2415)
         );
  AND2_X1 U2553 ( .A1(n2414), .A2(n2564), .ZN(n2413) );
  AOI21_X1 U2554 ( .B1(n2830), .B2(n4621), .A(n2829), .ZN(n3453) );
  AND2_X1 U2555 ( .A1(n3954), .A2(n3845), .ZN(n2829) );
  AOI21_X1 U2556 ( .B1(n3961), .B2(n2817), .A(n3748), .ZN(n2818) );
  INV_X1 U2557 ( .A(IR_REG_18__SCAN_IN), .ZN(n2472) );
  INV_X1 U2558 ( .A(IR_REG_24__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U2559 ( .A1(n2470), .A2(n2455), .ZN(n2454) );
  INV_X1 U2560 ( .A(IR_REG_5__SCAN_IN), .ZN(n2466) );
  INV_X1 U2561 ( .A(IR_REG_8__SCAN_IN), .ZN(n2465) );
  AND2_X1 U2562 ( .A1(n2359), .A2(n2357), .ZN(n2355) );
  AND2_X1 U2563 ( .A1(n4425), .A2(n4423), .ZN(n2373) );
  NOR2_X1 U2564 ( .A1(n2425), .A2(n2725), .ZN(n2424) );
  NOR2_X1 U2565 ( .A1(n2232), .A2(n2426), .ZN(n2425) );
  NAND2_X1 U2566 ( .A1(n3394), .A2(n2638), .ZN(n3432) );
  NOR2_X1 U2567 ( .A1(n2402), .A2(n2401), .ZN(n2400) );
  NAND2_X1 U2568 ( .A1(n2604), .A2(n2627), .ZN(n2401) );
  NOR2_X1 U2569 ( .A1(n2403), .A2(n2399), .ZN(n2398) );
  INV_X1 U2570 ( .A(n2627), .ZN(n2399) );
  NAND2_X1 U2571 ( .A1(n2955), .A2(n4625), .ZN(n3766) );
  AND2_X1 U2572 ( .A1(n4239), .A2(n3962), .ZN(n3748) );
  NOR2_X1 U2573 ( .A1(n2270), .A2(n4071), .ZN(n2269) );
  INV_X1 U2574 ( .A(n2271), .ZN(n2270) );
  AND2_X1 U2575 ( .A1(n2229), .A2(n4290), .ZN(n2286) );
  INV_X1 U2576 ( .A(n4625), .ZN(n2959) );
  AND2_X1 U2577 ( .A1(n3559), .A2(n3557), .ZN(n2359) );
  XNOR2_X1 U2578 ( .A(n2981), .B(n3536), .ZN(n3077) );
  NAND2_X1 U2579 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  OAI21_X1 U2580 ( .B1(n3661), .B2(n3659), .A(n3657), .ZN(n3542) );
  OAI21_X1 U2581 ( .B1(n3170), .B2(n2363), .A(n2361), .ZN(n3225) );
  INV_X1 U2582 ( .A(n2362), .ZN(n2361) );
  OAI21_X1 U2583 ( .B1(n2365), .B2(n2363), .A(n3179), .ZN(n2362) );
  INV_X1 U2584 ( .A(n2364), .ZN(n2363) );
  OR2_X1 U2585 ( .A1(n2355), .A2(n2352), .ZN(n2350) );
  AND2_X1 U2586 ( .A1(n2359), .A2(n3614), .ZN(n2352) );
  INV_X1 U2587 ( .A(n2338), .ZN(n3636) );
  AND2_X1 U2588 ( .A1(n3576), .A2(n3495), .ZN(n2339) );
  NOR2_X1 U2589 ( .A1(n2354), .A2(n2243), .ZN(n2349) );
  INV_X1 U2590 ( .A(n3614), .ZN(n2351) );
  AOI21_X1 U2591 ( .B1(n2346), .B2(n2349), .A(n3587), .ZN(n2345) );
  INV_X1 U2592 ( .A(n2350), .ZN(n2346) );
  OR2_X1 U2593 ( .A1(n2911), .A2(n2294), .ZN(n2293) );
  NAND2_X1 U2594 ( .A1(n2233), .A2(n2295), .ZN(n2294) );
  NAND2_X1 U2595 ( .A1(n4447), .A2(n3892), .ZN(n3894) );
  NAND2_X1 U2596 ( .A1(n4470), .A2(n3896), .ZN(n3897) );
  NAND2_X1 U2597 ( .A1(n4497), .A2(n3928), .ZN(n4507) );
  NAND2_X1 U2598 ( .A1(n4507), .A2(n4508), .ZN(n4506) );
  NAND2_X1 U2599 ( .A1(n4509), .A2(n3902), .ZN(n3903) );
  NAND2_X1 U2600 ( .A1(n4518), .A2(REG2_REG_12__SCAN_IN), .ZN(n4517) );
  XNOR2_X1 U2601 ( .A(n2384), .B(n3933), .ZN(n4540) );
  INV_X1 U2602 ( .A(n3905), .ZN(n2384) );
  OR2_X1 U2603 ( .A1(n4540), .A2(n2641), .ZN(n2382) );
  NAND2_X1 U2604 ( .A1(n4565), .A2(n2392), .ZN(n2391) );
  NAND2_X1 U2605 ( .A1(n4648), .A2(n4173), .ZN(n2392) );
  NOR2_X1 U2606 ( .A1(n2391), .A2(n4576), .ZN(n4575) );
  NOR2_X1 U2607 ( .A1(n2442), .A2(n2436), .ZN(n2435) );
  INV_X1 U2608 ( .A(n2743), .ZN(n2436) );
  INV_X1 U2609 ( .A(n2445), .ZN(n2439) );
  NOR2_X1 U2610 ( .A1(n2449), .A2(n2234), .ZN(n2443) );
  AND2_X1 U2611 ( .A1(n2450), .A2(n2761), .ZN(n2449) );
  NOR2_X1 U2612 ( .A1(n2231), .A2(n2742), .ZN(n2448) );
  NAND2_X1 U2613 ( .A1(n4270), .A2(n4071), .ZN(n2428) );
  NAND2_X1 U2614 ( .A1(n2719), .A2(n2232), .ZN(n2429) );
  NOR2_X1 U2615 ( .A1(n4049), .A2(n2720), .ZN(n4068) );
  NOR2_X1 U2616 ( .A1(n4150), .A2(n4138), .ZN(n4115) );
  AND4_X1 U2617 ( .A1(n2688), .A2(n2687), .A3(n2686), .A4(n2685), .ZN(n4291)
         );
  AND4_X1 U2618 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(n3375)
         );
  NAND2_X1 U2619 ( .A1(n2404), .A2(n2254), .ZN(n2403) );
  INV_X1 U2620 ( .A(n2405), .ZN(n2404) );
  AOI21_X1 U2621 ( .B1(n2604), .B2(n2605), .A(n2406), .ZN(n2405) );
  INV_X1 U2622 ( .A(n4588), .ZN(n2406) );
  INV_X1 U2623 ( .A(n2254), .ZN(n2402) );
  INV_X1 U2624 ( .A(n2604), .ZN(n2397) );
  OAI21_X1 U2625 ( .B1(n3294), .B2(n2595), .A(n2594), .ZN(n3303) );
  NAND2_X1 U2626 ( .A1(n2798), .A2(n3792), .ZN(n4589) );
  AOI21_X1 U2627 ( .B1(n3782), .B2(n2320), .A(n2319), .ZN(n2318) );
  INV_X1 U2628 ( .A(n3788), .ZN(n2320) );
  INV_X1 U2629 ( .A(n3787), .ZN(n2319) );
  NAND2_X1 U2630 ( .A1(n2329), .A2(n2325), .ZN(n2324) );
  NOR2_X1 U2631 ( .A1(n2563), .A2(n2462), .ZN(n2564) );
  NAND2_X1 U2632 ( .A1(n2789), .A2(n4614), .ZN(n4616) );
  NAND2_X1 U2633 ( .A1(n2820), .A2(n2819), .ZN(n4621) );
  INV_X1 U2634 ( .A(n4621), .ZN(n4598) );
  NAND2_X1 U2635 ( .A1(n3967), .A2(n3732), .ZN(n4225) );
  AND2_X1 U2636 ( .A1(n4040), .A2(n2280), .ZN(n3967) );
  NOR2_X1 U2637 ( .A1(n2281), .A2(n3962), .ZN(n2280) );
  INV_X1 U2638 ( .A(n2282), .ZN(n2281) );
  NAND2_X1 U2639 ( .A1(n4040), .A2(n2284), .ZN(n3997) );
  INV_X1 U2640 ( .A(n3847), .ZN(n4248) );
  AND2_X1 U2641 ( .A1(n4059), .A2(n4038), .ZN(n4040) );
  INV_X1 U2642 ( .A(n3858), .ZN(n3132) );
  NAND2_X1 U2643 ( .A1(n2864), .A2(n2788), .ZN(n4693) );
  NAND2_X1 U2644 ( .A1(n2842), .A2(n4408), .ZN(n2885) );
  AND2_X1 U2645 ( .A1(n2451), .A2(n2250), .ZN(n2333) );
  AND2_X1 U2646 ( .A1(n3414), .A2(n2341), .ZN(n2340) );
  INV_X1 U2647 ( .A(n4415), .ZN(n3675) );
  INV_X1 U2648 ( .A(n3665), .ZN(n4421) );
  INV_X1 U2649 ( .A(n4002), .ZN(n4245) );
  OAI21_X1 U2650 ( .B1(n4041), .B2(n2732), .A(n2731), .ZN(n4015) );
  INV_X1 U2651 ( .A(n4331), .ZN(n3851) );
  INV_X1 U2652 ( .A(n4322), .ZN(n4595) );
  NAND2_X1 U2653 ( .A1(n4448), .A2(n4449), .ZN(n4447) );
  XNOR2_X1 U2654 ( .A(n3894), .B(n4661), .ZN(n4459) );
  NAND2_X1 U2655 ( .A1(n4471), .A2(n4472), .ZN(n4470) );
  XNOR2_X1 U2656 ( .A(n3897), .B(n2378), .ZN(n4479) );
  NAND2_X1 U2657 ( .A1(n4489), .A2(n4490), .ZN(n4488) );
  OAI21_X1 U2658 ( .B1(n4560), .B2(n2303), .A(n2302), .ZN(n4570) );
  NAND2_X1 U2659 ( .A1(n2305), .A2(n2304), .ZN(n2303) );
  NAND2_X1 U2660 ( .A1(n3939), .A2(n2305), .ZN(n2302) );
  INV_X1 U2661 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2304) );
  AOI21_X1 U2662 ( .B1(n4578), .B2(ADDR_REG_18__SCAN_IN), .A(n4577), .ZN(n2388) );
  AOI21_X1 U2663 ( .B1(n2391), .B2(n4576), .A(n4574), .ZN(n2389) );
  INV_X1 U2664 ( .A(n4575), .ZN(n2390) );
  INV_X1 U2665 ( .A(n4235), .ZN(n3985) );
  NAND2_X1 U2666 ( .A1(n4187), .A2(n2670), .ZN(n4169) );
  AND4_X1 U2667 ( .A1(n2664), .A2(n2663), .A3(n2662), .A4(n2661), .ZN(n4292)
         );
  NAND2_X1 U2668 ( .A1(n3453), .A2(n2322), .ZN(n2868) );
  INV_X1 U2669 ( .A(n2323), .ZN(n2322) );
  OAI21_X1 U2670 ( .B1(n3456), .B2(n4337), .A(n2831), .ZN(n2323) );
  OAI21_X1 U2671 ( .B1(n3967), .B2(n3732), .A(n4225), .ZN(n3448) );
  INV_X1 U2672 ( .A(n2844), .ZN(n2887) );
  AND2_X1 U2673 ( .A1(n3395), .A2(n3393), .ZN(n3799) );
  NAND2_X1 U2674 ( .A1(n2974), .A2(n2959), .ZN(n3763) );
  INV_X1 U2675 ( .A(IR_REG_4__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U2676 ( .A1(n4030), .A2(n3818), .ZN(n4010) );
  INV_X1 U2677 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U2678 ( .A1(n2247), .A2(n2574), .ZN(n2418) );
  NOR2_X1 U2679 ( .A1(n2566), .A2(n5006), .ZN(n2575) );
  INV_X1 U2680 ( .A(n3283), .ZN(n3172) );
  OAI22_X1 U2681 ( .A1(n3018), .A2(n2526), .B1(n3772), .B2(n2525), .ZN(n3060)
         );
  XNOR2_X1 U2682 ( .A(n2982), .B(n3771), .ZN(n3021) );
  NOR2_X1 U2683 ( .A1(n2283), .A2(n4235), .ZN(n2282) );
  INV_X1 U2684 ( .A(n2284), .ZN(n2283) );
  NOR2_X1 U2685 ( .A1(n4244), .A2(n4014), .ZN(n2284) );
  NOR2_X1 U2686 ( .A1(n4269), .A2(n4116), .ZN(n2271) );
  OAI21_X1 U2687 ( .B1(n4136), .B2(n3688), .A(n3687), .ZN(n4110) );
  INV_X1 U2688 ( .A(n3195), .ZN(n3160) );
  AND2_X1 U2689 ( .A1(n2408), .A2(n4623), .ZN(n2274) );
  OR2_X1 U2690 ( .A1(n2885), .A2(n2858), .ZN(n2934) );
  AND2_X1 U2691 ( .A1(n2838), .A2(n2335), .ZN(n2334) );
  INV_X1 U2692 ( .A(IR_REG_25__SCAN_IN), .ZN(n2335) );
  NOR2_X1 U2693 ( .A1(n2475), .A2(n2474), .ZN(n2476) );
  INV_X1 U2694 ( .A(n2453), .ZN(n2376) );
  INV_X1 U2695 ( .A(n2454), .ZN(n2452) );
  INV_X2 U2696 ( .A(n2524), .ZN(n2268) );
  INV_X1 U2697 ( .A(IR_REG_6__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U2698 ( .A1(n3168), .A2(n3169), .ZN(n2364) );
  NAND2_X1 U2699 ( .A1(n2367), .A2(n2366), .ZN(n2365) );
  INV_X1 U2700 ( .A(n3168), .ZN(n2367) );
  INV_X1 U2701 ( .A(n3169), .ZN(n2366) );
  OR2_X1 U2702 ( .A1(n2763), .A2(n2762), .ZN(n2771) );
  XOR2_X1 U2703 ( .A(n3545), .B(n3546), .Z(n3543) );
  AND2_X1 U2704 ( .A1(n2919), .A2(n2918), .ZN(n2960) );
  AOI21_X1 U2705 ( .B1(n2373), .B2(n2371), .A(n3474), .ZN(n2370) );
  INV_X1 U2706 ( .A(n3083), .ZN(n3081) );
  NAND2_X1 U2707 ( .A1(n2337), .A2(n2926), .ZN(n2962) );
  NAND2_X1 U2708 ( .A1(n3625), .A2(n3626), .ZN(n3624) );
  NAND2_X1 U2709 ( .A1(n3566), .A2(n3488), .ZN(n3625) );
  NAND2_X1 U2710 ( .A1(n3487), .A2(n3486), .ZN(n3488) );
  INV_X1 U2711 ( .A(n3485), .ZN(n3486) );
  INV_X1 U2712 ( .A(n3484), .ZN(n3487) );
  OR2_X1 U2713 ( .A1(n2711), .A2(n3580), .ZN(n2713) );
  INV_X1 U2714 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2607) );
  OAI22_X1 U2715 ( .A1(n2955), .A2(n2954), .B1(n3508), .B2(n2959), .ZN(n2958)
         );
  NOR2_X1 U2716 ( .A1(n2370), .A2(n2264), .ZN(n2369) );
  INV_X1 U2717 ( .A(n3460), .ZN(n3461) );
  NOR2_X1 U2718 ( .A1(n2373), .A2(n2255), .ZN(n2372) );
  NAND2_X1 U2719 ( .A1(n3473), .A2(n3472), .ZN(n4422) );
  NOR2_X1 U2720 ( .A1(n2639), .A2(n4993), .ZN(n2649) );
  AND2_X1 U2721 ( .A1(n4409), .A2(n3949), .ZN(n2956) );
  OR2_X1 U2722 ( .A1(n2753), .A2(n2746), .ZN(n3662) );
  NAND2_X1 U2723 ( .A1(n4476), .A2(n3925), .ZN(n4486) );
  NAND2_X1 U2724 ( .A1(n4486), .A2(n4487), .ZN(n4485) );
  XNOR2_X1 U2725 ( .A(n3927), .B(n2377), .ZN(n4498) );
  NAND2_X1 U2726 ( .A1(n4488), .A2(n3899), .ZN(n3900) );
  NAND2_X1 U2727 ( .A1(n4506), .A2(n2266), .ZN(n3930) );
  NAND2_X1 U2728 ( .A1(n4533), .A2(n3932), .ZN(n3934) );
  INV_X1 U2729 ( .A(n4569), .ZN(n2305) );
  AOI21_X1 U2730 ( .B1(n3992), .B2(n3750), .A(n3829), .ZN(n3975) );
  NAND2_X1 U2731 ( .A1(n2423), .A2(n2422), .ZN(n4028) );
  AOI21_X1 U2732 ( .B1(n2424), .B2(n2426), .A(n2260), .ZN(n2422) );
  AND2_X1 U2733 ( .A1(n3702), .A2(DATAI_22_), .ZN(n4071) );
  AOI21_X1 U2734 ( .B1(n2811), .B2(n3811), .A(n2313), .ZN(n2312) );
  INV_X1 U2735 ( .A(n3815), .ZN(n2313) );
  NAND2_X1 U2736 ( .A1(n2311), .A2(n2805), .ZN(n4104) );
  NOR2_X1 U2737 ( .A1(n2682), .A2(n2681), .ZN(n2696) );
  AND4_X1 U2738 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(n4158)
         );
  INV_X1 U2739 ( .A(n2432), .ZN(n2431) );
  OAI21_X1 U2740 ( .B1(n2670), .B2(n2433), .A(n2680), .ZN(n2432) );
  NAND2_X1 U2741 ( .A1(n4188), .A2(n2669), .ZN(n4187) );
  AND2_X1 U2742 ( .A1(n2649), .A2(REG3_REG_15__SCAN_IN), .ZN(n2658) );
  NOR2_X1 U2743 ( .A1(n2398), .A2(n2256), .ZN(n2393) );
  OR2_X1 U2744 ( .A1(n3311), .A2(n3351), .ZN(n4604) );
  NAND2_X1 U2745 ( .A1(n2796), .A2(n3788), .ZN(n3154) );
  NAND2_X1 U2746 ( .A1(n2421), .A2(n2420), .ZN(n2416) );
  NOR2_X1 U2747 ( .A1(n2564), .A2(n3719), .ZN(n2420) );
  AND2_X1 U2748 ( .A1(n3277), .A2(n3172), .ZN(n3278) );
  AND4_X1 U2749 ( .A1(n2572), .A2(n2571), .A3(n2570), .A4(n2569), .ZN(n3249)
         );
  NAND2_X1 U2750 ( .A1(n3774), .A2(n3776), .ZN(n3693) );
  OR2_X1 U2751 ( .A1(n2506), .A2(n2408), .ZN(n3767) );
  NAND2_X1 U2752 ( .A1(n4608), .A2(n3766), .ZN(n2790) );
  NOR2_X1 U2753 ( .A1(n2507), .A2(n3718), .ZN(n2515) );
  AND2_X1 U2754 ( .A1(n2934), .A2(n2933), .ZN(n3038) );
  OR2_X1 U2755 ( .A1(n2885), .A2(D_REG_1__SCAN_IN), .ZN(n3035) );
  NOR2_X1 U2756 ( .A1(n4225), .A2(n4228), .ZN(n4224) );
  AND2_X1 U2757 ( .A1(n3702), .A2(DATAI_27_), .ZN(n4235) );
  NAND2_X1 U2758 ( .A1(n4040), .A2(n4020), .ZN(n4019) );
  AND2_X1 U2759 ( .A1(n4115), .A2(n2230), .ZN(n4059) );
  NAND2_X1 U2760 ( .A1(n4115), .A2(n2271), .ZN(n4090) );
  INV_X1 U2761 ( .A(n4131), .ZN(n4138) );
  NAND2_X1 U2762 ( .A1(n4207), .A2(n2267), .ZN(n4150) );
  NAND2_X1 U2763 ( .A1(n4207), .A2(n2286), .ZN(n4171) );
  INV_X1 U2764 ( .A(n4305), .ZN(n3437) );
  NOR2_X1 U2765 ( .A1(n4206), .A2(n4313), .ZN(n4207) );
  OR2_X1 U2766 ( .A1(n3400), .A2(n3406), .ZN(n4206) );
  AND4_X1 U2767 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), .ZN(n4322)
         );
  NOR2_X1 U2768 ( .A1(n4604), .A2(n4605), .ZN(n4603) );
  OR2_X1 U2769 ( .A1(n3161), .A2(n3357), .ZN(n3311) );
  NOR2_X1 U2770 ( .A1(n3142), .A2(n3246), .ZN(n3277) );
  AND2_X1 U2771 ( .A1(n4617), .A2(n4669), .ZN(n4337) );
  INV_X1 U2772 ( .A(n4609), .ZN(n4590) );
  NAND3_X1 U2773 ( .A1(n2273), .A2(n3143), .A3(n2525), .ZN(n3142) );
  AND3_X1 U2774 ( .A1(n2408), .A2(n4623), .A3(n3071), .ZN(n2273) );
  AND2_X1 U2775 ( .A1(n2274), .A2(n2525), .ZN(n3059) );
  INV_X1 U2776 ( .A(n4613), .ZN(n4596) );
  INV_X1 U2777 ( .A(n4610), .ZN(n4592) );
  AND2_X1 U2778 ( .A1(n2959), .A2(n3092), .ZN(n4623) );
  NAND2_X1 U2779 ( .A1(n2408), .A2(n4623), .ZN(n3047) );
  INV_X1 U2780 ( .A(n4693), .ZN(n4701) );
  OR2_X1 U2781 ( .A1(n4409), .A2(n3093), .ZN(n4669) );
  NAND2_X1 U2782 ( .A1(n2275), .A2(n2334), .ZN(n2840) );
  INV_X1 U2783 ( .A(n2832), .ZN(n2275) );
  NAND2_X1 U2784 ( .A1(n2486), .A2(IR_REG_31__SCAN_IN), .ZN(n2315) );
  AND2_X1 U2785 ( .A1(n2479), .A2(n2478), .ZN(n2822) );
  NAND2_X1 U2786 ( .A1(n2840), .A2(n2480), .ZN(n2821) );
  AND2_X1 U2787 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2480)
         );
  XNOR2_X1 U2788 ( .A(n2845), .B(n2846), .ZN(n2998) );
  NAND2_X1 U2789 ( .A1(n2779), .A2(IR_REG_31__SCAN_IN), .ZN(n2780) );
  NOR2_X1 U2790 ( .A1(n2499), .A2(n2300), .ZN(n2299) );
  NAND2_X1 U2791 ( .A1(n2248), .A2(IR_REG_1__SCAN_IN), .ZN(n2301) );
  NOR2_X1 U2792 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2300)
         );
  NAND2_X1 U2793 ( .A1(n2360), .A2(n2364), .ZN(n3180) );
  NAND2_X1 U2794 ( .A1(n3170), .A2(n2365), .ZN(n2360) );
  AND3_X1 U2795 ( .A1(n2493), .A2(n2492), .A3(n2491), .ZN(n4095) );
  OAI21_X1 U2796 ( .B1(n3649), .B2(n3645), .A(n3646), .ZN(n3567) );
  NAND2_X1 U2797 ( .A1(n3624), .A2(n3627), .ZN(n3578) );
  OR2_X1 U2798 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  NAND2_X1 U2799 ( .A1(n3635), .A2(n2350), .ZN(n2344) );
  NAND2_X1 U2800 ( .A1(n3558), .A2(n2356), .ZN(n3613) );
  OAI21_X1 U2801 ( .B1(n3384), .B2(n3383), .A(n3382), .ZN(n3413) );
  OR2_X1 U2802 ( .A1(n2964), .A2(n2950), .ZN(n4415) );
  AND2_X1 U2803 ( .A1(n2760), .A2(n2759), .ZN(n4002) );
  OR2_X1 U2804 ( .A1(n2964), .A2(n2951), .ZN(n3665) );
  AOI21_X1 U2805 ( .B1(n2345), .B2(n2347), .A(n2257), .ZN(n2342) );
  INV_X1 U2806 ( .A(n2349), .ZN(n2347) );
  AND2_X1 U2807 ( .A1(n3468), .A2(n3467), .ZN(n4423) );
  NAND2_X1 U2808 ( .A1(n2741), .A2(n2740), .ZN(n3847) );
  INV_X1 U2809 ( .A(n4291), .ZN(n4133) );
  INV_X1 U2810 ( .A(n4158), .ZN(n4420) );
  INV_X1 U2811 ( .A(n4292), .ZN(n4306) );
  INV_X1 U2812 ( .A(n3375), .ZN(n4334) );
  INV_X1 U2813 ( .A(n3249), .ZN(n3855) );
  NAND4_X1 U2814 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n3857)
         );
  CLKBUF_X1 U2815 ( .A(U4043), .Z(n3856) );
  NAND3_X1 U2816 ( .A1(n2505), .A2(n2504), .A3(n2503), .ZN(n2506) );
  OR2_X1 U2817 ( .A1(n2518), .A2(n2502), .ZN(n2504) );
  NAND2_X1 U2818 ( .A1(n2512), .A2(REG1_REG_2__SCAN_IN), .ZN(n2503) );
  AND2_X1 U2819 ( .A1(n2501), .A2(n2500), .ZN(n2505) );
  XNOR2_X1 U2820 ( .A(n2899), .B(REG1_REG_1__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U2821 ( .A1(n3863), .A2(n3862), .ZN(n3861) );
  NOR2_X1 U2822 ( .A1(n3918), .A2(n2296), .ZN(n4444) );
  NAND2_X1 U2823 ( .A1(n4458), .A2(n3895), .ZN(n4471) );
  NAND2_X1 U2824 ( .A1(n4478), .A2(n3898), .ZN(n4489) );
  XNOR2_X1 U2825 ( .A(n3900), .B(n2377), .ZN(n4500) );
  AND2_X1 U2826 ( .A1(n4438), .A2(n3839), .ZN(n4527) );
  XNOR2_X1 U2827 ( .A(n3930), .B(n4654), .ZN(n4523) );
  NAND2_X1 U2828 ( .A1(n4517), .A2(n3904), .ZN(n4529) );
  NAND2_X1 U2829 ( .A1(n4534), .A2(n4535), .ZN(n4533) );
  XNOR2_X1 U2830 ( .A(n3934), .B(n4652), .ZN(n4544) );
  INV_X1 U2831 ( .A(n2382), .ZN(n4539) );
  OAI21_X1 U2832 ( .B1(n4540), .B2(n2380), .A(n2379), .ZN(n4547) );
  NAND2_X1 U2833 ( .A1(n2383), .A2(REG2_REG_14__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U2834 ( .A1(n3906), .A2(n2383), .ZN(n2379) );
  INV_X1 U2835 ( .A(n4548), .ZN(n2383) );
  INV_X1 U2836 ( .A(n3906), .ZN(n2381) );
  NOR2_X1 U2837 ( .A1(n4560), .A2(REG1_REG_16__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U2838 ( .A1(n2434), .A2(n2438), .ZN(n2777) );
  AOI21_X1 U2839 ( .B1(n2441), .B2(n2439), .A(n2244), .ZN(n2438) );
  NAND2_X1 U2840 ( .A1(n4008), .A2(n2435), .ZN(n2434) );
  NOR2_X1 U2841 ( .A1(n3454), .A2(n2290), .ZN(n2289) );
  AND2_X1 U2842 ( .A1(n4175), .A2(n3455), .ZN(n2290) );
  NAND2_X1 U2843 ( .A1(n2444), .A2(n2440), .ZN(n3959) );
  INV_X1 U2844 ( .A(n2443), .ZN(n2440) );
  NAND2_X1 U2845 ( .A1(n2437), .A2(n2445), .ZN(n2444) );
  AOI21_X1 U2846 ( .B1(n2437), .B2(n2448), .A(n2752), .ZN(n3980) );
  INV_X1 U2847 ( .A(n2742), .ZN(n2447) );
  OR2_X1 U2848 ( .A1(n2745), .A2(n2727), .ZN(n4041) );
  AND2_X1 U2849 ( .A1(n2429), .A2(n2428), .ZN(n4047) );
  NAND2_X1 U2850 ( .A1(n2719), .A2(n2461), .ZN(n4067) );
  NAND2_X1 U2851 ( .A1(n4115), .A2(n3717), .ZN(n4278) );
  NAND2_X1 U2852 ( .A1(n4207), .A2(n2229), .ZN(n4300) );
  AND4_X1 U2853 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n4324)
         );
  AND4_X1 U2854 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(n4331)
         );
  INV_X1 U2855 ( .A(n4324), .ZN(n3850) );
  AND2_X1 U2856 ( .A1(n3399), .A2(n4621), .ZN(n4327) );
  INV_X1 U2857 ( .A(n2309), .ZN(n3371) );
  AND2_X1 U2858 ( .A1(n4205), .A2(n4609), .ZN(n4175) );
  NAND2_X1 U2859 ( .A1(n2395), .A2(n2403), .ZN(n3370) );
  NAND2_X1 U2860 ( .A1(n3303), .A2(n2396), .ZN(n2395) );
  NOR2_X1 U2861 ( .A1(n2397), .A2(n2402), .ZN(n2396) );
  NAND2_X1 U2862 ( .A1(n2317), .A2(n2318), .ZN(n3292) );
  AND2_X1 U2863 ( .A1(n2421), .A2(n2419), .ZN(n3287) );
  INV_X1 U2864 ( .A(n2564), .ZN(n2419) );
  NAND2_X1 U2865 ( .A1(n3061), .A2(n2331), .ZN(n2328) );
  NAND2_X1 U2866 ( .A1(n2332), .A2(n3776), .ZN(n3144) );
  OR2_X1 U2867 ( .A1(n3061), .A2(n2792), .ZN(n2332) );
  NAND2_X1 U2868 ( .A1(n4205), .A2(n3245), .ZN(n4165) );
  INV_X1 U2869 ( .A(n3949), .ZN(n4161) );
  INV_X1 U2870 ( .A(n2506), .ZN(n2516) );
  INV_X1 U2871 ( .A(n4629), .ZN(n4180) );
  NAND2_X1 U2872 ( .A1(n2947), .A2(n2946), .ZN(n4190) );
  INV_X1 U2873 ( .A(n2945), .ZN(n2946) );
  AND2_X1 U2874 ( .A1(n4205), .A2(n3041), .ZN(n4631) );
  INV_X1 U2875 ( .A(n4190), .ZN(n4622) );
  OR2_X1 U2876 ( .A1(n2867), .A2(n3036), .ZN(n4726) );
  INV_X2 U2877 ( .A(n4726), .ZN(n4729) );
  OAI21_X1 U2878 ( .B1(n3982), .B2(n3985), .A(n2285), .ZN(n4355) );
  AND2_X1 U2879 ( .A1(n4298), .A2(n4297), .ZN(n4386) );
  INV_X1 U2880 ( .A(n4644), .ZN(n2890) );
  NAND2_X1 U2881 ( .A1(n2836), .A2(IR_REG_31__SCAN_IN), .ZN(n2336) );
  AND2_X1 U2882 ( .A1(n2998), .A2(STATE_REG_SCAN_IN), .ZN(n4644) );
  NOR2_X1 U2883 ( .A1(n2499), .A2(n2823), .ZN(n2386) );
  AOI21_X1 U2884 ( .B1(n2390), .B2(n2389), .A(n2387), .ZN(n4584) );
  INV_X1 U2885 ( .A(n2388), .ZN(n2387) );
  NAND2_X1 U2886 ( .A1(n2291), .A2(n2287), .ZN(U3354) );
  INV_X1 U2887 ( .A(n2288), .ZN(n2287) );
  NAND2_X1 U2888 ( .A1(n2292), .A2(n4205), .ZN(n2291) );
  OAI21_X1 U2889 ( .B1(n3456), .B2(n4165), .A(n2289), .ZN(n2288) );
  OAI21_X1 U2890 ( .B1(n2868), .B2(n4706), .A(n2265), .ZN(n2870) );
  NAND2_X1 U2891 ( .A1(n2917), .A2(n3040), .ZN(n2978) );
  INV_X1 U2892 ( .A(n4410), .ZN(n2295) );
  AND2_X1 U2893 ( .A1(n2459), .A2(n2374), .ZN(n2225) );
  INV_X1 U2894 ( .A(n2354), .ZN(n2353) );
  NOR2_X1 U2895 ( .A1(n3511), .A2(n3510), .ZN(n2354) );
  AND2_X1 U2896 ( .A1(n2471), .A2(n2333), .ZN(n2484) );
  NAND2_X1 U2897 ( .A1(n2917), .A2(n2916), .ZN(n2954) );
  AND2_X1 U2898 ( .A1(n2225), .A2(n2835), .ZN(n2226) );
  INV_X1 U2899 ( .A(n3472), .ZN(n2371) );
  INV_X1 U2900 ( .A(n3762), .ZN(n2306) );
  NAND2_X1 U2901 ( .A1(n2237), .A2(n2457), .ZN(n2412) );
  NAND2_X1 U2902 ( .A1(n2471), .A2(n2470), .ZN(n2646) );
  NOR2_X1 U2903 ( .A1(n2372), .A2(n2264), .ZN(n2227) );
  AND2_X1 U2904 ( .A1(n2471), .A2(n2452), .ZN(n2228) );
  INV_X2 U2905 ( .A(n4706), .ZN(n4708) );
  AND2_X1 U2906 ( .A1(n3437), .A2(n4417), .ZN(n2229) );
  AND2_X1 U2907 ( .A1(n2269), .A2(n4057), .ZN(n2230) );
  XNOR2_X1 U2908 ( .A(n2780), .B(n2782), .ZN(n2788) );
  AND2_X1 U2909 ( .A1(n4236), .A2(n4244), .ZN(n2231) );
  NOR2_X1 U2910 ( .A1(n4068), .A2(n2427), .ZN(n2232) );
  NAND2_X1 U2911 ( .A1(n2910), .A2(n4411), .ZN(n2233) );
  NOR2_X1 U2912 ( .A1(n4002), .A2(n3985), .ZN(n2234) );
  OR2_X1 U2913 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2235)
         );
  AND2_X1 U2914 ( .A1(n2511), .A2(n2510), .ZN(n2236) );
  AND4_X1 U2915 ( .A1(n2466), .A2(n2558), .A3(n2581), .A4(n2465), .ZN(n2237)
         );
  AND2_X1 U2916 ( .A1(n2344), .A2(n2349), .ZN(n2238) );
  XNOR2_X1 U2917 ( .A(n2784), .B(IR_REG_21__SCAN_IN), .ZN(n3765) );
  INV_X1 U2918 ( .A(IR_REG_28__SCAN_IN), .ZN(n2824) );
  OR2_X1 U2919 ( .A1(n2832), .A2(IR_REG_25__SCAN_IN), .ZN(n2239) );
  NOR2_X1 U2920 ( .A1(n4561), .A2(n3939), .ZN(n2240) );
  NOR2_X2 U2921 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2499)
         );
  INV_X1 U2922 ( .A(n3050), .ZN(n2408) );
  INV_X1 U2923 ( .A(n2325), .ZN(n2331) );
  INV_X1 U2924 ( .A(IR_REG_2__SCAN_IN), .ZN(n2385) );
  INV_X1 U2925 ( .A(n2442), .ZN(n2441) );
  OR2_X1 U2926 ( .A1(n3960), .A2(n2443), .ZN(n2442) );
  AND2_X1 U2927 ( .A1(n3081), .A2(n3078), .ZN(n2241) );
  NAND2_X1 U2928 ( .A1(n2783), .A2(n2225), .ZN(n2242) );
  NOR2_X1 U2929 ( .A1(n2356), .A2(n2351), .ZN(n2243) );
  NOR2_X1 U2930 ( .A1(n4239), .A2(n3969), .ZN(n2244) );
  AND2_X1 U2931 ( .A1(n2348), .A2(n2353), .ZN(n2245) );
  XNOR2_X1 U2932 ( .A(n2958), .B(n3536), .ZN(n2985) );
  INV_X1 U2933 ( .A(IR_REG_21__SCAN_IN), .ZN(n2374) );
  OR2_X1 U2934 ( .A1(n2233), .A2(n2295), .ZN(n2246) );
  NAND2_X1 U2935 ( .A1(n3854), .A2(n3195), .ZN(n2247) );
  AND2_X1 U2936 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2248)
         );
  AND2_X1 U2937 ( .A1(n2437), .A2(n2447), .ZN(n2249) );
  AND2_X1 U2938 ( .A1(n2334), .A2(n2477), .ZN(n2250) );
  AND2_X1 U2939 ( .A1(n2382), .A2(n2381), .ZN(n2251) );
  NAND2_X1 U2940 ( .A1(n4207), .A2(n3437), .ZN(n2252) );
  NAND2_X1 U2941 ( .A1(n3858), .A2(n3143), .ZN(n2253) );
  OR2_X1 U2942 ( .A1(n4334), .A2(n4605), .ZN(n2254) );
  INV_X1 U2943 ( .A(n3510), .ZN(n2357) );
  NAND2_X1 U2944 ( .A1(n4040), .A2(n2282), .ZN(n2285) );
  NOR2_X1 U2945 ( .A1(n2411), .A2(n2412), .ZN(n2602) );
  NAND2_X1 U2946 ( .A1(n2394), .A2(n2393), .ZN(n3394) );
  OAI22_X1 U2947 ( .A1(n3413), .A2(n2340), .B1(n2341), .B2(n3414), .ZN(n3459)
         );
  OAI21_X1 U2948 ( .B1(n3473), .B2(n2372), .A(n2370), .ZN(n3604) );
  INV_X1 U2949 ( .A(n4035), .ZN(n4074) );
  OAI211_X1 U2950 ( .C1(n4060), .C2(n2732), .A(n2724), .B(n2723), .ZN(n4035)
         );
  AND2_X1 U2951 ( .A1(n4425), .A2(n2371), .ZN(n2255) );
  INV_X1 U2952 ( .A(n3785), .ZN(n2330) );
  INV_X1 U2953 ( .A(n3811), .ZN(n2805) );
  AND2_X1 U2954 ( .A1(n4595), .A2(n3378), .ZN(n2256) );
  NAND2_X1 U2955 ( .A1(n4115), .A2(n2269), .ZN(n2272) );
  NOR2_X1 U2956 ( .A1(n3517), .A2(n3516), .ZN(n2257) );
  INV_X1 U2957 ( .A(n2679), .ZN(n2433) );
  OR2_X1 U2958 ( .A1(n2369), .A2(n3605), .ZN(n2258) );
  INV_X1 U2959 ( .A(IR_REG_22__SCAN_IN), .ZN(n2835) );
  NAND2_X1 U2960 ( .A1(n3496), .A2(n3575), .ZN(n2259) );
  INV_X1 U2961 ( .A(n2752), .ZN(n2450) );
  NOR2_X1 U2962 ( .A1(n4236), .A2(n4244), .ZN(n2752) );
  AND2_X1 U2963 ( .A1(n4035), .A2(n4053), .ZN(n2260) );
  AND2_X1 U2964 ( .A1(n2669), .A2(n2679), .ZN(n2261) );
  AND2_X1 U2965 ( .A1(n2410), .A2(n2268), .ZN(n2262) );
  NAND2_X1 U2966 ( .A1(n2375), .A2(IR_REG_31__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U2967 ( .A1(n3763), .A2(n3766), .ZN(n2789) );
  INV_X1 U2968 ( .A(n2789), .ZN(n2307) );
  NAND2_X1 U2969 ( .A1(n3853), .A2(n3295), .ZN(n2263) );
  XNOR2_X1 U2970 ( .A(n2336), .B(IR_REG_24__SCAN_IN), .ZN(n2844) );
  OAI21_X1 U2971 ( .B1(n3303), .B2(n2605), .A(n2604), .ZN(n4587) );
  NAND2_X1 U2972 ( .A1(n2416), .A2(n2574), .ZN(n3153) );
  INV_X1 U2973 ( .A(n3798), .ZN(n2310) );
  AND2_X1 U2974 ( .A1(n3477), .A2(n3476), .ZN(n2264) );
  INV_X1 U2975 ( .A(n2326), .ZN(n2329) );
  NAND2_X1 U2976 ( .A1(n3079), .A2(n3078), .ZN(n3080) );
  NAND3_X1 U2977 ( .A1(n2410), .A2(n2409), .A3(n2268), .ZN(n2635) );
  NAND2_X1 U2978 ( .A1(n2690), .A2(n2689), .ZN(n2702) );
  OR2_X1 U2979 ( .A1(REG0_REG_29__SCAN_IN), .A2(n4708), .ZN(n2265) );
  OR2_X1 U2980 ( .A1(n4655), .A2(n4727), .ZN(n2266) );
  AND2_X1 U2981 ( .A1(n2286), .A2(n4151), .ZN(n2267) );
  NAND2_X1 U2982 ( .A1(n3702), .A2(DATAI_25_), .ZN(n4020) );
  NAND2_X1 U2983 ( .A1(n3702), .A2(DATAI_23_), .ZN(n4057) );
  INV_X1 U2984 ( .A(n2407), .ZN(n3718) );
  NAND2_X1 U2985 ( .A1(n3767), .A2(n3769), .ZN(n2407) );
  INV_X1 U2986 ( .A(IR_REG_0__SCAN_IN), .ZN(n2277) );
  INV_X1 U2987 ( .A(IR_REG_17__SCAN_IN), .ZN(n2689) );
  INV_X1 U2988 ( .A(n4496), .ZN(n2377) );
  INV_X1 U2989 ( .A(n4475), .ZN(n2378) );
  INV_X1 U2990 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2585) );
  INV_X1 U2991 ( .A(IR_REG_14__SCAN_IN), .ZN(n2455) );
  INV_X1 U2992 ( .A(IR_REG_29__SCAN_IN), .ZN(n2314) );
  INV_X1 U2993 ( .A(IR_REG_23__SCAN_IN), .ZN(n2846) );
  NOR2_X1 U2994 ( .A1(n2486), .A2(IR_REG_29__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U2995 ( .A1(n2268), .A2(n2457), .ZN(n2549) );
  NAND2_X1 U2996 ( .A1(n2268), .A2(n2467), .ZN(n2411) );
  INV_X1 U2997 ( .A(n2272), .ZN(n4075) );
  NAND3_X1 U2998 ( .A1(n2274), .A2(n2525), .A3(n3071), .ZN(n3140) );
  OAI21_X1 U2999 ( .B1(n3702), .B2(n2277), .A(n2276), .ZN(n4624) );
  NAND2_X1 U3000 ( .A1(n3702), .A2(DATAI_0_), .ZN(n2276) );
  OAI21_X1 U3001 ( .B1(n3702), .B2(n2899), .A(n2279), .ZN(n4625) );
  NAND2_X1 U3002 ( .A1(n3702), .A2(DATAI_1_), .ZN(n2279) );
  INV_X1 U3003 ( .A(n2285), .ZN(n3981) );
  NAND3_X1 U3004 ( .A1(n3452), .A2(n3451), .A3(n3453), .ZN(n2292) );
  NAND2_X1 U3005 ( .A1(n2298), .A2(n2233), .ZN(n2297) );
  AND2_X1 U3006 ( .A1(n2297), .A2(n4410), .ZN(n2296) );
  INV_X1 U3007 ( .A(n2911), .ZN(n2298) );
  AND2_X2 U3008 ( .A1(n3975), .A2(n3979), .ZN(n3977) );
  AOI21_X2 U3009 ( .B1(n4589), .B2(n3797), .A(n2310), .ZN(n2309) );
  INV_X1 U3010 ( .A(n4123), .ZN(n2311) );
  NAND2_X1 U3011 ( .A1(n2317), .A2(n2316), .ZN(n2797) );
  OR2_X2 U3012 ( .A1(n2796), .A2(n2321), .ZN(n2317) );
  OAI211_X1 U3013 ( .C1(n3061), .C2(n2326), .A(n2324), .B(n3786), .ZN(n2794)
         );
  NAND2_X1 U3014 ( .A1(n2253), .A2(n3776), .ZN(n2325) );
  NAND2_X1 U3015 ( .A1(n3785), .A2(n2327), .ZN(n2326) );
  NAND3_X1 U3016 ( .A1(n2253), .A2(n3776), .A3(n2792), .ZN(n2327) );
  NAND2_X1 U3017 ( .A1(n2328), .A2(n2329), .ZN(n3129) );
  NAND2_X1 U3018 ( .A1(n2471), .A2(n2451), .ZN(n2832) );
  NAND2_X1 U3019 ( .A1(n2790), .A2(n3718), .ZN(n3020) );
  NAND2_X2 U3020 ( .A1(n3737), .A2(n4199), .ZN(n4200) );
  NAND2_X2 U3021 ( .A1(n2803), .A2(n3809), .ZN(n4123) );
  NAND2_X1 U3022 ( .A1(n3023), .A2(n3773), .ZN(n3061) );
  NAND2_X1 U3023 ( .A1(n2799), .A2(n3802), .ZN(n3737) );
  INV_X1 U3024 ( .A(n2822), .ZN(n2482) );
  OAI21_X1 U3025 ( .B1(n2926), .B2(n2337), .A(n2962), .ZN(n2973) );
  NAND2_X1 U3026 ( .A1(n2924), .A2(n2925), .ZN(n2337) );
  INV_X1 U3027 ( .A(n3459), .ZN(n3462) );
  INV_X1 U3028 ( .A(n3412), .ZN(n2341) );
  NAND2_X1 U3029 ( .A1(n3635), .A2(n2345), .ZN(n2343) );
  NAND2_X1 U3030 ( .A1(n3635), .A2(n2355), .ZN(n2348) );
  NAND2_X1 U3031 ( .A1(n3635), .A2(n2359), .ZN(n3558) );
  NAND2_X1 U3032 ( .A1(n3102), .A2(n3101), .ZN(n3595) );
  NAND2_X1 U3033 ( .A1(n2241), .A2(n3079), .ZN(n3102) );
  INV_X1 U3034 ( .A(n3473), .ZN(n2368) );
  AOI21_X2 U3035 ( .B1(n2368), .B2(n2227), .A(n2258), .ZN(n3649) );
  NOR2_X1 U3036 ( .A1(n3473), .A2(n3472), .ZN(n3671) );
  NAND2_X1 U3037 ( .A1(n2783), .A2(n2459), .ZN(n2785) );
  NAND2_X1 U3038 ( .A1(n2783), .A2(n2226), .ZN(n2375) );
  XNOR2_X2 U3039 ( .A(n2386), .B(n2385), .ZN(n4412) );
  NAND2_X1 U3040 ( .A1(n3303), .A2(n2400), .ZN(n2394) );
  INV_X1 U3041 ( .A(n2412), .ZN(n2410) );
  INV_X1 U3042 ( .A(n2418), .ZN(n2414) );
  NAND2_X1 U3043 ( .A1(n2565), .A2(n2458), .ZN(n2421) );
  NAND2_X1 U3044 ( .A1(n2719), .A2(n2424), .ZN(n2423) );
  INV_X1 U3045 ( .A(n2429), .ZN(n4066) );
  NAND2_X1 U3046 ( .A1(n4188), .A2(n2261), .ZN(n2430) );
  NAND2_X1 U3047 ( .A1(n2430), .A2(n2431), .ZN(n4148) );
  NAND2_X1 U3048 ( .A1(n4008), .A2(n2743), .ZN(n2437) );
  NAND2_X1 U3049 ( .A1(n2821), .A2(IR_REG_28__SCAN_IN), .ZN(n2481) );
  OAI21_X1 U3050 ( .B1(n3321), .B2(n3322), .A(n3320), .ZN(n3328) );
  NAND2_X1 U3051 ( .A1(n3449), .A2(n4629), .ZN(n3452) );
  OAI22_X1 U3052 ( .A1(n2516), .A2(n2954), .B1(n3508), .B2(n2408), .ZN(n2990)
         );
  AND2_X1 U3053 ( .A1(n3702), .A2(DATAI_28_), .ZN(n3962) );
  AOI21_X2 U3054 ( .B1(n3462), .B2(n2460), .A(n3461), .ZN(n3473) );
  AND3_X1 U3055 ( .A1(n3550), .A2(n3549), .A3(n4426), .ZN(n2456) );
  NAND2_X2 U3056 ( .A1(n3039), .A2(n4190), .ZN(n4205) );
  AND2_X1 U3057 ( .A1(n2532), .A2(n2464), .ZN(n2457) );
  NOR2_X1 U3058 ( .A1(n3125), .A2(n2462), .ZN(n2458) );
  AND2_X1 U3059 ( .A1(n2782), .A2(n2781), .ZN(n2459) );
  INV_X1 U3060 ( .A(IR_REG_9__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3061 ( .A1(n3416), .A2(n3417), .ZN(n2460) );
  OR2_X1 U3062 ( .A1(n4107), .A2(n4269), .ZN(n2461) );
  INV_X1 U3063 ( .A(n4153), .ZN(n2692) );
  INV_X1 U3064 ( .A(n4269), .ZN(n4091) );
  AND2_X1 U3065 ( .A1(n3702), .A2(DATAI_21_), .ZN(n4269) );
  OAI21_X1 U3066 ( .B1(n3662), .B2(n2732), .A(n2751), .ZN(n4236) );
  AND2_X1 U3067 ( .A1(n3812), .A2(n3809), .ZN(n3695) );
  INV_X1 U3068 ( .A(n3695), .ZN(n2669) );
  AND2_X1 U3069 ( .A1(n3857), .A2(n3246), .ZN(n2462) );
  AND3_X1 U3070 ( .A1(n4202), .A2(n3431), .A3(n2655), .ZN(n2463) );
  INV_X1 U3071 ( .A(n3640), .ZN(n4107) );
  NAND2_X1 U3072 ( .A1(n3702), .A2(DATAI_26_), .ZN(n4001) );
  INV_X1 U3073 ( .A(n4001), .ZN(n4244) );
  INV_X1 U3074 ( .A(IR_REG_12__SCAN_IN), .ZN(n2468) );
  OR2_X1 U3075 ( .A1(n4102), .A2(n2810), .ZN(n3816) );
  INV_X1 U3076 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2628) );
  AND2_X1 U3077 ( .A1(n3682), .A2(n4029), .ZN(n3818) );
  OR2_X1 U3078 ( .A1(n2629), .A2(n2628), .ZN(n2639) );
  NAND2_X1 U3079 ( .A1(n4107), .A2(n4269), .ZN(n2718) );
  OR2_X1 U3080 ( .A1(n4669), .A2(n3765), .ZN(n2945) );
  AND2_X1 U3081 ( .A1(n2696), .A2(REG3_REG_19__SCAN_IN), .ZN(n2704) );
  AND3_X1 U3082 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2551) );
  NOR2_X1 U3083 ( .A1(n2886), .A2(n2872), .ZN(n2843) );
  OR2_X1 U3084 ( .A1(n2596), .A2(n4820), .ZN(n2608) );
  AND2_X2 U3085 ( .A1(n4407), .A2(n2880), .ZN(n2508) );
  NAND2_X1 U3086 ( .A1(n3450), .A2(n4622), .ZN(n3451) );
  AND2_X1 U3087 ( .A1(n2754), .A2(n2763), .ZN(n3983) );
  OR2_X1 U3088 ( .A1(n2672), .A2(n2671), .ZN(n2682) );
  NOR2_X1 U3089 ( .A1(n2608), .A2(n2607), .ZN(n2617) );
  OR2_X1 U3090 ( .A1(n2586), .A2(n2585), .ZN(n2596) );
  NAND2_X1 U3091 ( .A1(n3702), .A2(DATAI_20_), .ZN(n3717) );
  INV_X1 U3092 ( .A(n3086), .ZN(n3071) );
  INV_X1 U3093 ( .A(n4189), .ZN(n4417) );
  NAND2_X1 U3094 ( .A1(n2704), .A2(REG3_REG_20__SCAN_IN), .ZN(n2711) );
  OR2_X1 U3095 ( .A1(n2713), .A2(n3639), .ZN(n2721) );
  AND2_X1 U3096 ( .A1(n2745), .A2(n2744), .ZN(n2753) );
  NAND2_X1 U3097 ( .A1(n3703), .A2(REG1_REG_3__SCAN_IN), .ZN(n2521) );
  INV_X1 U3098 ( .A(n4661), .ZN(n3893) );
  INV_X1 U3099 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4820) );
  AND2_X1 U3100 ( .A1(n3846), .A2(n3969), .ZN(n3728) );
  AOI22_X1 U3101 ( .A1(n4110), .A2(n2710), .B1(n4116), .B2(n3849), .ZN(n4085)
         );
  OR2_X1 U3102 ( .A1(n2885), .A2(D_REG_0__SCAN_IN), .ZN(n2862) );
  NAND2_X1 U3103 ( .A1(n3702), .A2(DATAI_24_), .ZN(n4038) );
  INV_X1 U3104 ( .A(n4323), .ZN(n3406) );
  NAND2_X1 U3105 ( .A1(n2917), .A2(n4644), .ZN(n3034) );
  NOR2_X1 U3106 ( .A1(n2721), .A2(n4816), .ZN(n2726) );
  AND2_X1 U3107 ( .A1(n2771), .A2(n2764), .ZN(n3970) );
  NAND2_X1 U3108 ( .A1(n2658), .A2(REG3_REG_16__SCAN_IN), .ZN(n2672) );
  AND2_X1 U3109 ( .A1(n2770), .A2(n2769), .ZN(n4239) );
  AND4_X1 U3110 ( .A1(n2717), .A2(n2716), .A3(n2715), .A4(n2714), .ZN(n3640)
         );
  NAND2_X1 U3111 ( .A1(n2512), .A2(REG1_REG_0__SCAN_IN), .ZN(n2513) );
  AND2_X1 U3112 ( .A1(n2896), .A2(n2895), .ZN(n4438) );
  AND2_X1 U3113 ( .A1(n4438), .A2(n2927), .ZN(n4580) );
  NOR2_X1 U3114 ( .A1(n3748), .A2(n3728), .ZN(n3960) );
  AND2_X1 U3115 ( .A1(n4127), .A2(n4128), .ZN(n4153) );
  INV_X1 U3116 ( .A(n4202), .ZN(n4199) );
  INV_X1 U3117 ( .A(n4165), .ZN(n4194) );
  AND2_X1 U3118 ( .A1(n4205), .A2(n3046), .ZN(n4629) );
  NAND2_X1 U3119 ( .A1(n2862), .A2(n2861), .ZN(n3036) );
  INV_X1 U3120 ( .A(n3962), .ZN(n3969) );
  INV_X1 U3121 ( .A(n4337), .ZN(n4686) );
  INV_X1 U3122 ( .A(n3036), .ZN(n2935) );
  INV_X1 U3123 ( .A(n3034), .ZN(n2947) );
  AND2_X1 U3124 ( .A1(n2896), .A2(n2884), .ZN(n4578) );
  AND2_X1 U3125 ( .A1(n3002), .A2(n3001), .ZN(n4431) );
  INV_X1 U3126 ( .A(n4239), .ZN(n3846) );
  INV_X1 U3127 ( .A(n4095), .ZN(n4270) );
  NAND2_X1 U3128 ( .A1(n4438), .A2(n4414), .ZN(n4586) );
  INV_X1 U3129 ( .A(n4527), .ZN(n4574) );
  OR2_X1 U3130 ( .A1(n3448), .A2(n4714), .ZN(n2865) );
  NAND2_X1 U3131 ( .A1(n4729), .A2(n4701), .ZN(n4714) );
  OR2_X1 U3132 ( .A1(n3448), .A2(n4677), .ZN(n2869) );
  NAND2_X1 U3133 ( .A1(n4708), .A2(n4701), .ZN(n4677) );
  OR2_X1 U3134 ( .A1(n2867), .A2(n2935), .ZN(n4706) );
  AND2_X2 U3135 ( .A1(n2885), .A2(n2947), .ZN(n4643) );
  XNOR2_X1 U3136 ( .A(n2825), .B(n2824), .ZN(n4414) );
  INV_X1 U3137 ( .A(n3915), .ZN(n4653) );
  OR2_X1 U3138 ( .A1(n2561), .A2(n2560), .ZN(n4661) );
  INV_X2 U3139 ( .A(IR_REG_7__SCAN_IN), .ZN(n2581) );
  INV_X2 U3140 ( .A(IR_REG_19__SCAN_IN), .ZN(n2781) );
  NAND4_X1 U3141 ( .A1(n2473), .A2(n2472), .A3(n2781), .A4(n2689), .ZN(n2475)
         );
  NAND4_X1 U3142 ( .A1(n2846), .A2(n2374), .A3(n2782), .A4(n2835), .ZN(n2474)
         );
  INV_X1 U3143 ( .A(n2484), .ZN(n2479) );
  INV_X1 U3144 ( .A(IR_REG_27__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3145 ( .A1(n2823), .A2(n2477), .ZN(n2478) );
  NAND2_X1 U3146 ( .A1(n2551), .A2(REG3_REG_6__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U3147 ( .A1(n2575), .A2(REG3_REG_8__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U31480 ( .A1(n2617), .A2(REG3_REG_12__SCAN_IN), .ZN(n2629) );
  INV_X1 U31490 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2671) );
  INV_X1 U3150 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2681) );
  INV_X1 U3151 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3580) );
  INV_X1 U3152 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U3153 ( .A1(n2713), .A2(n3639), .ZN(n2483) );
  AND2_X1 U3154 ( .A1(n2721), .A2(n2483), .ZN(n4078) );
  NAND2_X1 U3155 ( .A1(n2484), .A2(n2824), .ZN(n2486) );
  XNOR2_X2 U3156 ( .A(n2485), .B(IR_REG_30__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U3157 ( .A1(n4078), .A2(n2606), .ZN(n2493) );
  NOR2_X2 U3158 ( .A1(n4407), .A2(n2880), .ZN(n2509) );
  NAND2_X1 U3159 ( .A1(n2544), .A2(REG0_REG_22__SCAN_IN), .ZN(n2489) );
  INV_X1 U3160 ( .A(n4407), .ZN(n2487) );
  NAND2_X1 U3161 ( .A1(n3703), .A2(REG1_REG_22__SCAN_IN), .ZN(n2488) );
  AND2_X1 U3162 ( .A1(n2489), .A2(n2488), .ZN(n2492) );
  INV_X1 U3163 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4080) );
  OR2_X1 U3164 ( .A1(n3707), .A2(n4080), .ZN(n2491) );
  NAND2_X1 U3165 ( .A1(n2512), .A2(REG1_REG_1__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3166 ( .A1(n2508), .A2(REG3_REG_1__SCAN_IN), .ZN(n2497) );
  INV_X1 U3167 ( .A(n2518), .ZN(n2494) );
  NAND2_X1 U3168 ( .A1(n2509), .A2(REG0_REG_1__SCAN_IN), .ZN(n2495) );
  INV_X1 U3169 ( .A(n2899), .ZN(n4413) );
  OR2_X1 U3170 ( .A1(n2955), .A2(n2959), .ZN(n3042) );
  INV_X1 U3171 ( .A(n3042), .ZN(n2507) );
  NAND2_X1 U3172 ( .A1(n2508), .A2(REG3_REG_2__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3173 ( .A1(n2509), .A2(REG0_REG_2__SCAN_IN), .ZN(n2500) );
  INV_X1 U3174 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2502) );
  MUX2_X1 U3175 ( .A(n4412), .B(DATAI_2_), .S(n3702), .Z(n3050) );
  NAND2_X1 U3176 ( .A1(n2506), .A2(n2408), .ZN(n3769) );
  INV_X1 U3177 ( .A(n2955), .ZN(n2974) );
  INV_X1 U3178 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2928) );
  OR2_X1 U3179 ( .A1(n2518), .A2(n2928), .ZN(n2514) );
  NAND2_X1 U3180 ( .A1(n2508), .A2(REG3_REG_0__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U3181 ( .A1(n2509), .A2(REG0_REG_0__SCAN_IN), .ZN(n2510) );
  AND2_X1 U3182 ( .A1(n4611), .A2(n4624), .ZN(n4614) );
  NAND2_X1 U3183 ( .A1(n2515), .A2(n4616), .ZN(n3045) );
  NAND2_X1 U3184 ( .A1(n2516), .A2(n2408), .ZN(n2517) );
  NAND2_X1 U3185 ( .A1(n3045), .A2(n2517), .ZN(n3018) );
  INV_X1 U3186 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3204) );
  OR2_X1 U3187 ( .A1(n3707), .A2(n3204), .ZN(n2523) );
  INV_X1 U3188 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3189 ( .A1(n2508), .A2(n2519), .ZN(n2522) );
  NAND2_X1 U3190 ( .A1(n2544), .A2(REG0_REG_3__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U3191 ( .A1(n2524), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  XNOR2_X1 U3192 ( .A(n2533), .B(IR_REG_3__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U3193 ( .A(n4411), .B(DATAI_3_), .S(n3702), .Z(n3771) );
  NOR2_X1 U3194 ( .A1(n2982), .A2(n3771), .ZN(n2526) );
  INV_X1 U3195 ( .A(n2982), .ZN(n3772) );
  INV_X1 U3196 ( .A(n3771), .ZN(n2525) );
  NAND2_X1 U3197 ( .A1(n2544), .A2(REG0_REG_4__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U3198 ( .A1(n3703), .A2(REG1_REG_4__SCAN_IN), .ZN(n2530) );
  INV_X1 U3199 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2527) );
  XNOR2_X1 U3200 ( .A(n2527), .B(REG3_REG_3__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3201 ( .A1(n2508), .A2(n3084), .ZN(n2529) );
  INV_X1 U3202 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3890) );
  OR2_X1 U3203 ( .A1(n3707), .A2(n3890), .ZN(n2528) );
  NAND2_X1 U3204 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  NAND2_X1 U3205 ( .A1(n2534), .A2(IR_REG_31__SCAN_IN), .ZN(n2535) );
  XNOR2_X1 U3206 ( .A(n2535), .B(IR_REG_4__SCAN_IN), .ZN(n4410) );
  MUX2_X1 U3207 ( .A(n4410), .B(DATAI_4_), .S(n3702), .Z(n3086) );
  NAND2_X1 U3208 ( .A1(n3072), .A2(n3086), .ZN(n3774) );
  NAND2_X1 U3209 ( .A1(n3859), .A2(n3071), .ZN(n3776) );
  NAND2_X1 U32100 ( .A1(n3060), .A2(n3693), .ZN(n2537) );
  NAND2_X1 U32110 ( .A1(n3859), .A2(n3086), .ZN(n2536) );
  NAND2_X1 U32120 ( .A1(n2537), .A2(n2536), .ZN(n3124) );
  INV_X1 U32130 ( .A(n3124), .ZN(n2565) );
  INV_X1 U32140 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2538) );
  OR2_X1 U32150 ( .A1(n3707), .A2(n2538), .ZN(n2548) );
  INV_X1 U32160 ( .A(n2551), .ZN(n2542) );
  INV_X1 U32170 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32180 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2539) );
  NAND2_X1 U32190 ( .A1(n2540), .A2(n2539), .ZN(n2541) );
  NAND2_X1 U32200 ( .A1(n2542), .A2(n2541), .ZN(n3599) );
  INV_X1 U32210 ( .A(n3599), .ZN(n2543) );
  NAND2_X1 U32220 ( .A1(n2508), .A2(n2543), .ZN(n2547) );
  NAND2_X1 U32230 ( .A1(n3703), .A2(REG1_REG_5__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32240 ( .A1(n2544), .A2(REG0_REG_5__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32250 ( .A1(n2549), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  XNOR2_X1 U32260 ( .A(n2550), .B(IR_REG_5__SCAN_IN), .ZN(n3920) );
  MUX2_X1 U32270 ( .A(n3920), .B(DATAI_5_), .S(n3702), .Z(n3598) );
  AND2_X1 U32280 ( .A1(n3858), .A2(n3598), .ZN(n3125) );
  INV_X1 U32290 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3248) );
  OR2_X1 U32300 ( .A1(n3707), .A2(n3248), .ZN(n2556) );
  NAND2_X1 U32310 ( .A1(n2544), .A2(REG0_REG_6__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32320 ( .A1(n3703), .A2(REG1_REG_6__SCAN_IN), .ZN(n2554) );
  OAI21_X1 U32330 ( .B1(n2551), .B2(REG3_REG_6__SCAN_IN), .A(n2566), .ZN(n3247) );
  INV_X1 U32340 ( .A(n3247), .ZN(n2552) );
  NAND2_X1 U32350 ( .A1(n2606), .A2(n2552), .ZN(n2553) );
  NOR2_X1 U32360 ( .A1(n2549), .A2(IR_REG_5__SCAN_IN), .ZN(n2559) );
  NOR2_X1 U32370 ( .A1(n2559), .A2(n2823), .ZN(n2557) );
  MUX2_X1 U32380 ( .A(n2823), .B(n2557), .S(IR_REG_6__SCAN_IN), .Z(n2561) );
  NAND2_X1 U32390 ( .A1(n2559), .A2(n2558), .ZN(n2573) );
  INV_X1 U32400 ( .A(n2573), .ZN(n2560) );
  MUX2_X1 U32410 ( .A(n3893), .B(DATAI_6_), .S(n3702), .Z(n3246) );
  INV_X1 U32420 ( .A(n3598), .ZN(n3143) );
  NAND2_X1 U32430 ( .A1(n3132), .A2(n3143), .ZN(n3126) );
  OR2_X1 U32440 ( .A1(n3857), .A2(n3246), .ZN(n2562) );
  AND2_X1 U32450 ( .A1(n3126), .A2(n2562), .ZN(n2563) );
  NAND2_X1 U32460 ( .A1(n2544), .A2(REG0_REG_7__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U32470 ( .A1(n3703), .A2(REG1_REG_7__SCAN_IN), .ZN(n2571) );
  AND2_X1 U32480 ( .A1(n2566), .A2(n5006), .ZN(n2567) );
  NOR2_X1 U32490 ( .A1(n2575), .A2(n2567), .ZN(n3173) );
  NAND2_X1 U32500 ( .A1(n2606), .A2(n3173), .ZN(n2570) );
  INV_X1 U32510 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2568) );
  OR2_X1 U32520 ( .A1(n3707), .A2(n2568), .ZN(n2569) );
  NAND2_X1 U32530 ( .A1(n2573), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  XNOR2_X1 U32540 ( .A(n2582), .B(IR_REG_7__SCAN_IN), .ZN(n3923) );
  MUX2_X1 U32550 ( .A(n3923), .B(DATAI_7_), .S(n3702), .Z(n3283) );
  NAND2_X1 U32560 ( .A1(n3249), .A2(n3283), .ZN(n3779) );
  NAND2_X1 U32570 ( .A1(n3855), .A2(n3172), .ZN(n3788) );
  NAND2_X1 U32580 ( .A1(n3779), .A2(n3788), .ZN(n3280) );
  NAND2_X1 U32590 ( .A1(n3855), .A2(n3283), .ZN(n2574) );
  INV_X1 U32600 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3163) );
  OR2_X1 U32610 ( .A1(n3707), .A2(n3163), .ZN(n2580) );
  NAND2_X1 U32620 ( .A1(n2544), .A2(REG0_REG_8__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32630 ( .A1(n3703), .A2(REG1_REG_8__SCAN_IN), .ZN(n2578) );
  OR2_X1 U32640 ( .A1(n2575), .A2(REG3_REG_8__SCAN_IN), .ZN(n2576) );
  AND2_X1 U32650 ( .A1(n2586), .A2(n2576), .ZN(n3162) );
  NAND2_X1 U32660 ( .A1(n2606), .A2(n3162), .ZN(n2577) );
  NAND4_X1 U32670 ( .A1(n2580), .A2(n2579), .A3(n2578), .A4(n2577), .ZN(n3854)
         );
  NAND2_X1 U32680 ( .A1(n2582), .A2(n2581), .ZN(n2583) );
  NAND2_X1 U32690 ( .A1(n2583), .A2(IR_REG_31__SCAN_IN), .ZN(n2584) );
  XNOR2_X1 U32700 ( .A(n2584), .B(IR_REG_8__SCAN_IN), .ZN(n4475) );
  MUX2_X1 U32710 ( .A(n4475), .B(DATAI_8_), .S(n3702), .Z(n3195) );
  OR2_X1 U32720 ( .A1(n3707), .A2(n3887), .ZN(n2592) );
  NAND2_X1 U32730 ( .A1(n3703), .A2(REG1_REG_9__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U32740 ( .A1(n2544), .A2(REG0_REG_9__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U32750 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  NAND2_X1 U32760 ( .A1(n2596), .A2(n2587), .ZN(n3296) );
  INV_X1 U32770 ( .A(n3296), .ZN(n2588) );
  NAND2_X1 U32780 ( .A1(n2508), .A2(n2588), .ZN(n2589) );
  NAND4_X1 U32790 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n3853)
         );
  OR2_X1 U32800 ( .A1(n2262), .A2(n2823), .ZN(n2593) );
  XNOR2_X1 U32810 ( .A(n2593), .B(IR_REG_9__SCAN_IN), .ZN(n3917) );
  MUX2_X1 U32820 ( .A(n3917), .B(DATAI_9_), .S(n3702), .Z(n3357) );
  NOR2_X1 U32830 ( .A1(n3853), .A2(n3357), .ZN(n2595) );
  NAND2_X1 U32840 ( .A1(n3853), .A2(n3357), .ZN(n2594) );
  INV_X1 U32850 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3315) );
  OR2_X1 U32860 ( .A1(n3707), .A2(n3315), .ZN(n2601) );
  NAND2_X1 U32870 ( .A1(n2544), .A2(REG0_REG_10__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U32880 ( .A1(n3703), .A2(REG1_REG_10__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U32890 ( .A1(n2596), .A2(n4820), .ZN(n2597) );
  AND2_X1 U32900 ( .A1(n2608), .A2(n2597), .ZN(n3314) );
  NAND2_X1 U32910 ( .A1(n2606), .A2(n3314), .ZN(n2598) );
  NAND4_X1 U32920 ( .A1(n2601), .A2(n2600), .A3(n2599), .A4(n2598), .ZN(n3852)
         );
  OR2_X1 U32930 ( .A1(n2602), .A2(n2823), .ZN(n2603) );
  XNOR2_X1 U32940 ( .A(n2603), .B(IR_REG_10__SCAN_IN), .ZN(n4496) );
  MUX2_X1 U32950 ( .A(n4496), .B(DATAI_10_), .S(n3702), .Z(n3351) );
  AND2_X1 U32960 ( .A1(n3852), .A2(n3351), .ZN(n2605) );
  INV_X1 U32970 ( .A(n3852), .ZN(n4593) );
  INV_X1 U32980 ( .A(n3351), .ZN(n3312) );
  NAND2_X1 U32990 ( .A1(n4593), .A2(n3312), .ZN(n2604) );
  AND2_X1 U33000 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  OR2_X1 U33010 ( .A1(n2609), .A2(n2617), .ZN(n3240) );
  INV_X1 U33020 ( .A(n3240), .ZN(n4602) );
  NAND2_X1 U33030 ( .A1(n2606), .A2(n4602), .ZN(n2614) );
  NAND2_X1 U33040 ( .A1(n3703), .A2(REG1_REG_11__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33050 ( .A1(n2544), .A2(REG0_REG_11__SCAN_IN), .ZN(n2612) );
  INV_X1 U33060 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2610) );
  OR2_X1 U33070 ( .A1(n3707), .A2(n2610), .ZN(n2611) );
  NAND2_X1 U33080 ( .A1(n2602), .A2(n2615), .ZN(n2616) );
  NAND2_X1 U33090 ( .A1(n2616), .A2(IR_REG_31__SCAN_IN), .ZN(n2624) );
  XNOR2_X1 U33100 ( .A(n2624), .B(IR_REG_11__SCAN_IN), .ZN(n3916) );
  MUX2_X1 U33110 ( .A(n3916), .B(DATAI_11_), .S(n3702), .Z(n4605) );
  NAND2_X1 U33120 ( .A1(n3375), .A2(n4605), .ZN(n3798) );
  INV_X1 U33130 ( .A(n4605), .ZN(n4591) );
  NAND2_X1 U33140 ( .A1(n4334), .A2(n4591), .ZN(n3797) );
  NAND2_X1 U33150 ( .A1(n3798), .A2(n3797), .ZN(n4588) );
  NAND2_X1 U33160 ( .A1(n2544), .A2(REG0_REG_12__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U33170 ( .A1(n3703), .A2(REG1_REG_12__SCAN_IN), .ZN(n2621) );
  OR2_X1 U33180 ( .A1(n2617), .A2(REG3_REG_12__SCAN_IN), .ZN(n2618) );
  AND2_X1 U33190 ( .A1(n2618), .A2(n2629), .ZN(n3336) );
  NAND2_X1 U33200 ( .A1(n2606), .A2(n3336), .ZN(n2620) );
  INV_X1 U33210 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3374) );
  OR2_X1 U33220 ( .A1(n3707), .A2(n3374), .ZN(n2619) );
  NAND2_X1 U33230 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
  NAND2_X1 U33240 ( .A1(n2625), .A2(IR_REG_31__SCAN_IN), .ZN(n2626) );
  XNOR2_X1 U33250 ( .A(n2626), .B(IR_REG_12__SCAN_IN), .ZN(n3929) );
  INV_X1 U33260 ( .A(n3929), .ZN(n4654) );
  INV_X1 U33270 ( .A(DATAI_12_), .ZN(n5082) );
  MUX2_X1 U33280 ( .A(n4654), .B(n5082), .S(n3702), .Z(n4330) );
  NAND2_X1 U33290 ( .A1(n4322), .A2(n4330), .ZN(n2627) );
  INV_X1 U33300 ( .A(n4330), .ZN(n3378) );
  NAND2_X1 U33310 ( .A1(n2544), .A2(REG0_REG_13__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U33320 ( .A1(n3703), .A2(REG1_REG_13__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U33330 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
  AND2_X1 U33340 ( .A1(n2639), .A2(n2630), .ZN(n3387) );
  NAND2_X1 U33350 ( .A1(n2606), .A2(n3387), .ZN(n2632) );
  INV_X1 U33360 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3403) );
  OR2_X1 U33370 ( .A1(n3707), .A2(n3403), .ZN(n2631) );
  NAND2_X1 U33380 ( .A1(n2635), .A2(IR_REG_31__SCAN_IN), .ZN(n2636) );
  XNOR2_X1 U33390 ( .A(n2636), .B(IR_REG_13__SCAN_IN), .ZN(n3915) );
  INV_X1 U33400 ( .A(DATAI_13_), .ZN(n2637) );
  MUX2_X1 U33410 ( .A(n4653), .B(n2637), .S(n3702), .Z(n4323) );
  NAND2_X1 U33420 ( .A1(n4331), .A2(n4323), .ZN(n2638) );
  NAND2_X1 U33430 ( .A1(n2544), .A2(REG0_REG_14__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U33440 ( .A1(n3703), .A2(REG1_REG_14__SCAN_IN), .ZN(n2644) );
  AND2_X1 U33450 ( .A1(n2639), .A2(n4993), .ZN(n2640) );
  NOR2_X1 U33460 ( .A1(n2649), .A2(n2640), .ZN(n4210) );
  NAND2_X1 U33470 ( .A1(n2606), .A2(n4210), .ZN(n2643) );
  INV_X1 U33480 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2641) );
  OR2_X1 U33490 ( .A1(n3707), .A2(n2641), .ZN(n2642) );
  NAND2_X1 U33500 ( .A1(n2646), .A2(IR_REG_31__SCAN_IN), .ZN(n2647) );
  XNOR2_X1 U33510 ( .A(n2647), .B(IR_REG_14__SCAN_IN), .ZN(n3933) );
  MUX2_X1 U33520 ( .A(n3933), .B(DATAI_14_), .S(n3702), .Z(n4313) );
  NAND2_X1 U3353 ( .A1(n4324), .A2(n4313), .ZN(n3803) );
  INV_X1 U33540 ( .A(n4313), .ZN(n4212) );
  NAND2_X1 U3355 ( .A1(n3850), .A2(n4212), .ZN(n3735) );
  NAND2_X1 U3356 ( .A1(n3803), .A2(n3735), .ZN(n4202) );
  NAND2_X1 U3357 ( .A1(n3851), .A2(n3406), .ZN(n3431) );
  INV_X1 U3358 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2648) );
  OR2_X1 U3359 ( .A1(n3707), .A2(n2648), .ZN(n2654) );
  NAND2_X1 U3360 ( .A1(n2544), .A2(REG0_REG_15__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3361 ( .A1(n3703), .A2(REG1_REG_15__SCAN_IN), .ZN(n2652) );
  NOR2_X1 U3362 ( .A1(n2649), .A2(REG3_REG_15__SCAN_IN), .ZN(n2650) );
  OR2_X1 U3363 ( .A1(n2658), .A2(n2650), .ZN(n3678) );
  INV_X1 U3364 ( .A(n3678), .ZN(n3435) );
  NAND2_X1 U3365 ( .A1(n2606), .A2(n3435), .ZN(n2651) );
  NAND4_X1 U3366 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .ZN(n4314)
         );
  OR2_X1 U3367 ( .A1(n2228), .A2(n2823), .ZN(n2666) );
  XNOR2_X1 U3368 ( .A(n2666), .B(IR_REG_15__SCAN_IN), .ZN(n3913) );
  MUX2_X1 U3369 ( .A(n3913), .B(DATAI_15_), .S(n3702), .Z(n4305) );
  NAND2_X1 U3370 ( .A1(n4314), .A2(n4305), .ZN(n2655) );
  NOR2_X1 U3371 ( .A1(n3850), .A2(n4313), .ZN(n3433) );
  INV_X1 U3372 ( .A(n4314), .ZN(n4416) );
  AOI22_X1 U3373 ( .A1(n3433), .A2(n2655), .B1(n4416), .B2(n3437), .ZN(n2656)
         );
  OR2_X1 U3374 ( .A1(n2658), .A2(REG3_REG_16__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3375 ( .A1(n2672), .A2(n2659), .ZN(n4430) );
  INV_X1 U3376 ( .A(n4430), .ZN(n2660) );
  NAND2_X1 U3377 ( .A1(n2606), .A2(n2660), .ZN(n2664) );
  NAND2_X1 U3378 ( .A1(n3703), .A2(REG1_REG_16__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3379 ( .A1(n2544), .A2(REG0_REG_16__SCAN_IN), .ZN(n2662) );
  INV_X1 U3380 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4191) );
  OR2_X1 U3381 ( .A1(n3707), .A2(n4191), .ZN(n2661) );
  INV_X1 U3382 ( .A(IR_REG_15__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3383 ( .A1(n2666), .A2(n2665), .ZN(n2667) );
  NAND2_X1 U3384 ( .A1(n2667), .A2(IR_REG_31__SCAN_IN), .ZN(n2668) );
  XNOR2_X1 U3385 ( .A(n2668), .B(IR_REG_16__SCAN_IN), .ZN(n3937) );
  MUX2_X1 U3386 ( .A(n3937), .B(DATAI_16_), .S(n3702), .Z(n4189) );
  NAND2_X1 U3387 ( .A1(n4292), .A2(n4189), .ZN(n3812) );
  NAND2_X1 U3388 ( .A1(n4306), .A2(n4417), .ZN(n3809) );
  NAND2_X1 U3389 ( .A1(n4306), .A2(n4189), .ZN(n2670) );
  NAND2_X1 U3390 ( .A1(n2672), .A2(n2671), .ZN(n2673) );
  AND2_X1 U3391 ( .A1(n2682), .A2(n2673), .ZN(n3607) );
  NAND2_X1 U3392 ( .A1(n2606), .A2(n3607), .ZN(n2677) );
  NAND2_X1 U3393 ( .A1(n3703), .A2(REG1_REG_17__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3394 ( .A1(n2544), .A2(REG0_REG_17__SCAN_IN), .ZN(n2675) );
  INV_X1 U3395 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4173) );
  OR2_X1 U3396 ( .A1(n3707), .A2(n4173), .ZN(n2674) );
  OR2_X1 U3397 ( .A1(n2690), .A2(n2823), .ZN(n2678) );
  XNOR2_X1 U3398 ( .A(n2678), .B(IR_REG_17__SCAN_IN), .ZN(n3941) );
  MUX2_X1 U3399 ( .A(n3941), .B(DATAI_17_), .S(n3702), .Z(n4176) );
  INV_X1 U3400 ( .A(n4176), .ZN(n4290) );
  NAND2_X1 U3401 ( .A1(n4158), .A2(n4290), .ZN(n2679) );
  NAND2_X1 U3402 ( .A1(n4420), .A2(n4176), .ZN(n2680) );
  INV_X1 U3403 ( .A(n4148), .ZN(n2693) );
  NAND2_X1 U3404 ( .A1(n2544), .A2(REG0_REG_18__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U3405 ( .A1(n3703), .A2(REG1_REG_18__SCAN_IN), .ZN(n2687) );
  AND2_X1 U3406 ( .A1(n2682), .A2(n2681), .ZN(n2683) );
  NOR2_X1 U3407 ( .A1(n2696), .A2(n2683), .ZN(n4149) );
  NAND2_X1 U3408 ( .A1(n2606), .A2(n4149), .ZN(n2686) );
  INV_X1 U3409 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2684) );
  OR2_X1 U3410 ( .A1(n3707), .A2(n2684), .ZN(n2685) );
  NAND2_X1 U3411 ( .A1(n2702), .A2(IR_REG_31__SCAN_IN), .ZN(n2691) );
  XNOR2_X1 U3412 ( .A(n2691), .B(IR_REG_18__SCAN_IN), .ZN(n4645) );
  MUX2_X1 U3413 ( .A(n4645), .B(DATAI_18_), .S(n3702), .Z(n4155) );
  NAND2_X1 U3414 ( .A1(n4291), .A2(n4155), .ZN(n4127) );
  INV_X1 U3415 ( .A(n4155), .ZN(n4151) );
  NAND2_X1 U3416 ( .A1(n4133), .A2(n4151), .ZN(n4128) );
  NAND2_X1 U3417 ( .A1(n2693), .A2(n2692), .ZN(n4146) );
  NAND2_X1 U3418 ( .A1(n4291), .A2(n4151), .ZN(n2694) );
  NAND2_X1 U3419 ( .A1(n4146), .A2(n2694), .ZN(n4136) );
  INV_X1 U3420 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2695) );
  OR2_X1 U3421 ( .A1(n3707), .A2(n2695), .ZN(n2701) );
  NAND2_X1 U3422 ( .A1(n3703), .A2(REG1_REG_19__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3423 ( .A1(n2544), .A2(REG0_REG_19__SCAN_IN), .ZN(n2699) );
  NOR2_X1 U3424 ( .A1(n2696), .A2(REG3_REG_19__SCAN_IN), .ZN(n2697) );
  OR2_X1 U3425 ( .A1(n2704), .A2(n2697), .ZN(n3571) );
  INV_X1 U3426 ( .A(n3571), .ZN(n4141) );
  NAND2_X1 U3427 ( .A1(n2606), .A2(n4141), .ZN(n2698) );
  NAND4_X1 U3428 ( .A1(n2701), .A2(n2700), .A3(n2699), .A4(n2698), .ZN(n4156)
         );
  INV_X1 U3429 ( .A(n2783), .ZN(n2703) );
  INV_X1 U3430 ( .A(DATAI_19_), .ZN(n2873) );
  MUX2_X1 U3431 ( .A(n3949), .B(n2873), .S(n3702), .Z(n4131) );
  NOR2_X1 U3432 ( .A1(n4156), .A2(n4138), .ZN(n3688) );
  NAND2_X1 U3433 ( .A1(n4156), .A2(n4138), .ZN(n3687) );
  INV_X1 U3434 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4118) );
  OR2_X1 U3435 ( .A1(n3707), .A2(n4118), .ZN(n2709) );
  NAND2_X1 U3436 ( .A1(n2544), .A2(REG0_REG_20__SCAN_IN), .ZN(n2708) );
  NAND2_X1 U3437 ( .A1(n3703), .A2(REG1_REG_20__SCAN_IN), .ZN(n2707) );
  OR2_X1 U3438 ( .A1(n2704), .A2(REG3_REG_20__SCAN_IN), .ZN(n2705) );
  AND2_X1 U3439 ( .A1(n2711), .A2(n2705), .ZN(n3622) );
  NAND2_X1 U3440 ( .A1(n2606), .A2(n3622), .ZN(n2706) );
  NAND4_X1 U3441 ( .A1(n2709), .A2(n2708), .A3(n2707), .A4(n2706), .ZN(n3849)
         );
  INV_X1 U3442 ( .A(n3849), .ZN(n4272) );
  NAND2_X1 U3443 ( .A1(n4272), .A2(n3717), .ZN(n2710) );
  INV_X1 U3444 ( .A(n3717), .ZN(n4116) );
  NAND2_X1 U3445 ( .A1(n2711), .A2(n3580), .ZN(n2712) );
  AND2_X1 U3446 ( .A1(n2713), .A2(n2712), .ZN(n3579) );
  NAND2_X1 U3447 ( .A1(n3579), .A2(n2606), .ZN(n2717) );
  NAND2_X1 U3448 ( .A1(n2544), .A2(REG0_REG_21__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3449 ( .A1(n3703), .A2(REG1_REG_21__SCAN_IN), .ZN(n2715) );
  INV_X1 U3450 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4094) );
  OR2_X1 U3451 ( .A1(n3707), .A2(n4094), .ZN(n2714) );
  NAND2_X1 U3452 ( .A1(n4085), .A2(n2718), .ZN(n2719) );
  NAND2_X1 U3453 ( .A1(n4095), .A2(n4071), .ZN(n2812) );
  INV_X1 U3454 ( .A(n4071), .ZN(n4076) );
  NAND2_X1 U3455 ( .A1(n4270), .A2(n4076), .ZN(n2813) );
  INV_X1 U3456 ( .A(n2813), .ZN(n2720) );
  INV_X1 U3457 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4816) );
  AND2_X1 U34580 ( .A1(n2721), .A2(n4816), .ZN(n2722) );
  OR2_X1 U34590 ( .A1(n2722), .A2(n2726), .ZN(n4060) );
  AOI22_X1 U3460 ( .A1(n3703), .A2(REG1_REG_23__SCAN_IN), .B1(n2544), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2724) );
  INV_X1 U3461 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4061) );
  OR2_X1 U3462 ( .A1(n3707), .A2(n4061), .ZN(n2723) );
  INV_X1 U3463 ( .A(n4057), .ZN(n4053) );
  NOR2_X1 U3464 ( .A1(n4035), .A2(n4053), .ZN(n2725) );
  NOR2_X1 U3465 ( .A1(n2726), .A2(REG3_REG_24__SCAN_IN), .ZN(n2727) );
  INV_X1 U3466 ( .A(n2606), .ZN(n2732) );
  INV_X1 U34670 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4042) );
  NAND2_X1 U3468 ( .A1(n2544), .A2(REG0_REG_24__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U34690 ( .A1(n3703), .A2(REG1_REG_24__SCAN_IN), .ZN(n2728) );
  OAI211_X1 U3470 ( .C1(n4042), .C2(n3707), .A(n2729), .B(n2728), .ZN(n2730)
         );
  INV_X1 U34710 ( .A(n2730), .ZN(n2731) );
  INV_X1 U3472 ( .A(n4038), .ZN(n4034) );
  INV_X1 U34730 ( .A(n4015), .ZN(n4056) );
  OAI21_X1 U3474 ( .B1(n4028), .B2(n2734), .A(n2733), .ZN(n2735) );
  INV_X1 U34750 ( .A(n2735), .ZN(n4008) );
  INV_X1 U3476 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2736) );
  XNOR2_X1 U34770 ( .A(n2745), .B(n2736), .ZN(n4021) );
  NAND2_X1 U3478 ( .A1(n4021), .A2(n2606), .ZN(n2741) );
  INV_X1 U34790 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U3480 ( .A1(n3703), .A2(REG1_REG_25__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U34810 ( .A1(n2544), .A2(REG0_REG_25__SCAN_IN), .ZN(n2737) );
  OAI211_X1 U3482 ( .C1(n4023), .C2(n3707), .A(n2738), .B(n2737), .ZN(n2739)
         );
  INV_X1 U34830 ( .A(n2739), .ZN(n2740) );
  NAND2_X1 U3484 ( .A1(n4248), .A2(n4020), .ZN(n2743) );
  NOR2_X1 U34850 ( .A1(n4248), .A2(n4020), .ZN(n2742) );
  AND2_X1 U3486 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2744) );
  AOI21_X1 U34870 ( .B1(n2745), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2746) );
  INV_X1 U3488 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U34890 ( .A1(n2544), .A2(REG0_REG_26__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U3490 ( .A1(n3703), .A2(REG1_REG_26__SCAN_IN), .ZN(n2747) );
  OAI211_X1 U34910 ( .C1(n2749), .C2(n3707), .A(n2748), .B(n2747), .ZN(n2750)
         );
  INV_X1 U3492 ( .A(n2750), .ZN(n2751) );
  INV_X1 U34930 ( .A(n4236), .ZN(n4018) );
  OR2_X1 U3494 ( .A1(n2753), .A2(REG3_REG_27__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U34950 ( .A1(n2753), .A2(REG3_REG_27__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U3496 ( .A1(n3983), .A2(n2606), .ZN(n2760) );
  INV_X1 U34970 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U3498 ( .A1(n3703), .A2(REG1_REG_27__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U34990 ( .A1(n2544), .A2(REG0_REG_27__SCAN_IN), .ZN(n2755) );
  OAI211_X1 U3500 ( .C1(n2757), .C2(n3707), .A(n2756), .B(n2755), .ZN(n2758)
         );
  INV_X1 U35010 ( .A(n2758), .ZN(n2759) );
  NAND2_X1 U3502 ( .A1(n4002), .A2(n3985), .ZN(n2761) );
  INV_X1 U35030 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U3504 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  NAND2_X1 U35050 ( .A1(n3970), .A2(n2606), .ZN(n2770) );
  INV_X1 U35060 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2767) );
  NAND2_X1 U35070 ( .A1(n2544), .A2(REG0_REG_28__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U35080 ( .A1(n3703), .A2(REG1_REG_28__SCAN_IN), .ZN(n2765) );
  OAI211_X1 U35090 ( .C1(n2767), .C2(n3707), .A(n2766), .B(n2765), .ZN(n2768)
         );
  INV_X1 U35100 ( .A(n2768), .ZN(n2769) );
  INV_X1 U35110 ( .A(n2771), .ZN(n3450) );
  NAND2_X1 U35120 ( .A1(n3450), .A2(n2606), .ZN(n2776) );
  INV_X1 U35130 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U35140 ( .A1(n2544), .A2(REG0_REG_29__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U35150 ( .A1(n3703), .A2(REG1_REG_29__SCAN_IN), .ZN(n2772) );
  OAI211_X1 U35160 ( .C1(n3447), .C2(n3707), .A(n2773), .B(n2772), .ZN(n2774)
         );
  INV_X1 U35170 ( .A(n2774), .ZN(n2775) );
  NAND2_X1 U35180 ( .A1(n2776), .A2(n2775), .ZN(n3963) );
  NAND2_X1 U35190 ( .A1(n3702), .A2(DATAI_29_), .ZN(n3732) );
  XNOR2_X1 U35200 ( .A(n3963), .B(n3732), .ZN(n3724) );
  XNOR2_X1 U35210 ( .A(n2777), .B(n3724), .ZN(n3456) );
  NAND2_X1 U35220 ( .A1(n2778), .A2(n2781), .ZN(n2779) );
  NAND2_X1 U35230 ( .A1(n2785), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U35240 ( .A1(n2242), .A2(IR_REG_31__SCAN_IN), .ZN(n2786) );
  XNOR2_X1 U35250 ( .A(n3040), .B(n4409), .ZN(n2787) );
  NAND2_X1 U35260 ( .A1(n2787), .A2(n3949), .ZN(n4617) );
  NAND2_X1 U35270 ( .A1(n2788), .A2(n4161), .ZN(n3093) );
  INV_X1 U35280 ( .A(n4611), .ZN(n2952) );
  NAND2_X1 U35290 ( .A1(n2952), .A2(n4624), .ZN(n3762) );
  NAND2_X1 U35300 ( .A1(n3020), .A2(n3767), .ZN(n2791) );
  NAND2_X1 U35310 ( .A1(n2791), .A2(n3021), .ZN(n3023) );
  NAND2_X1 U35320 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  INV_X1 U35330 ( .A(n3774), .ZN(n2792) );
  NAND2_X1 U35340 ( .A1(n3132), .A2(n3598), .ZN(n3785) );
  INV_X1 U35350 ( .A(n3246), .ZN(n2793) );
  NAND2_X1 U35360 ( .A1(n3857), .A2(n2793), .ZN(n3786) );
  INV_X1 U35370 ( .A(n3857), .ZN(n3286) );
  NAND2_X1 U35380 ( .A1(n3286), .A2(n3246), .ZN(n3778) );
  NAND2_X1 U35390 ( .A1(n2794), .A2(n3778), .ZN(n3281) );
  INV_X1 U35400 ( .A(n3779), .ZN(n2795) );
  OR2_X2 U35410 ( .A1(n3281), .A2(n2795), .ZN(n2796) );
  INV_X1 U35420 ( .A(n3854), .ZN(n3360) );
  NAND2_X1 U35430 ( .A1(n3360), .A2(n3195), .ZN(n3782) );
  NAND2_X1 U35440 ( .A1(n3854), .A2(n3160), .ZN(n3787) );
  INV_X1 U35450 ( .A(n3357), .ZN(n3295) );
  INV_X1 U35460 ( .A(n3853), .ZN(n3306) );
  NAND2_X1 U35470 ( .A1(n3306), .A2(n3357), .ZN(n3783) );
  NAND2_X1 U35480 ( .A1(n2797), .A2(n3783), .ZN(n3304) );
  NAND2_X1 U35490 ( .A1(n3852), .A2(n3312), .ZN(n3796) );
  NAND2_X1 U35500 ( .A1(n3304), .A2(n3796), .ZN(n2798) );
  NAND2_X1 U35510 ( .A1(n4593), .A2(n3351), .ZN(n3792) );
  NOR2_X1 U35520 ( .A1(n4595), .A2(n4330), .ZN(n3800) );
  NAND2_X1 U35530 ( .A1(n4595), .A2(n4330), .ZN(n3395) );
  NAND2_X1 U35540 ( .A1(n3851), .A2(n4323), .ZN(n3393) );
  NAND2_X1 U35550 ( .A1(n3396), .A2(n3799), .ZN(n2799) );
  NAND2_X1 U35560 ( .A1(n4331), .A2(n3406), .ZN(n3802) );
  NAND2_X1 U35570 ( .A1(n4416), .A2(n4305), .ZN(n3801) );
  NAND2_X1 U35580 ( .A1(n4314), .A2(n3437), .ZN(n3736) );
  NAND2_X1 U35590 ( .A1(n3801), .A2(n3736), .ZN(n3428) );
  INV_X1 U35600 ( .A(n3803), .ZN(n2800) );
  NOR2_X1 U35610 ( .A1(n3428), .A2(n2800), .ZN(n2801) );
  NAND2_X1 U35620 ( .A1(n4200), .A2(n2801), .ZN(n2802) );
  NAND2_X1 U35630 ( .A1(n2802), .A2(n3736), .ZN(n4183) );
  NAND2_X1 U35640 ( .A1(n4183), .A2(n3695), .ZN(n2803) );
  NAND2_X1 U35650 ( .A1(n4420), .A2(n4290), .ZN(n4124) );
  NAND2_X1 U35660 ( .A1(n4156), .A2(n4131), .ZN(n2804) );
  AND2_X1 U35670 ( .A1(n4128), .A2(n2804), .ZN(n2806) );
  NAND2_X1 U35680 ( .A1(n4124), .A2(n2806), .ZN(n3811) );
  NAND2_X1 U35690 ( .A1(n4158), .A2(n4176), .ZN(n4125) );
  NAND2_X1 U35700 ( .A1(n4127), .A2(n4125), .ZN(n2807) );
  NAND2_X1 U35710 ( .A1(n2807), .A2(n2806), .ZN(n2809) );
  INV_X1 U35720 ( .A(n4156), .ZN(n4109) );
  NAND2_X1 U35730 ( .A1(n4109), .A2(n4138), .ZN(n2808) );
  NAND2_X1 U35740 ( .A1(n2809), .A2(n2808), .ZN(n4102) );
  NOR2_X1 U35750 ( .A1(n3849), .A2(n3717), .ZN(n2810) );
  INV_X1 U35760 ( .A(n3816), .ZN(n2811) );
  NAND2_X1 U35770 ( .A1(n3849), .A2(n3717), .ZN(n3815) );
  NAND2_X1 U35780 ( .A1(n3640), .A2(n4269), .ZN(n4048) );
  AND2_X1 U35790 ( .A1(n2812), .A2(n4048), .ZN(n3820) );
  NAND2_X1 U35800 ( .A1(n4087), .A2(n3820), .ZN(n2816) );
  NAND2_X1 U35810 ( .A1(n4035), .A2(n4057), .ZN(n2814) );
  NAND2_X1 U3582 ( .A1(n2814), .A2(n2813), .ZN(n3821) );
  NAND2_X1 U3583 ( .A1(n4107), .A2(n4091), .ZN(n3814) );
  NOR2_X1 U3584 ( .A1(n4049), .A2(n3814), .ZN(n2815) );
  NOR2_X1 U3585 ( .A1(n3821), .A2(n2815), .ZN(n3745) );
  NAND2_X1 U3586 ( .A1(n2816), .A2(n3745), .ZN(n4030) );
  OR2_X1 U3587 ( .A1(n4015), .A2(n4038), .ZN(n3682) );
  OR2_X1 U3588 ( .A1(n4035), .A2(n4057), .ZN(n4029) );
  NAND2_X1 U3589 ( .A1(n3847), .A2(n4020), .ZN(n3723) );
  NAND2_X1 U3590 ( .A1(n4015), .A2(n4038), .ZN(n4009) );
  AND2_X1 U3591 ( .A1(n3723), .A2(n4009), .ZN(n3824) );
  OR2_X1 U3592 ( .A1(n4236), .A2(n4001), .ZN(n3716) );
  OR2_X1 U3593 ( .A1(n3847), .A2(n4020), .ZN(n3991) );
  NAND2_X1 U3594 ( .A1(n3716), .A2(n3991), .ZN(n3822) );
  INV_X1 U3595 ( .A(n3822), .ZN(n3750) );
  AND2_X1 U3596 ( .A1(n4236), .A2(n4001), .ZN(n3829) );
  XNOR2_X1 U3597 ( .A(n4245), .B(n4235), .ZN(n3979) );
  AND2_X1 U3598 ( .A1(n4002), .A2(n4235), .ZN(n3747) );
  OR2_X2 U3599 ( .A1(n3977), .A2(n3747), .ZN(n3961) );
  INV_X1 U3600 ( .A(n3728), .ZN(n2817) );
  XNOR2_X1 U3601 ( .A(n2818), .B(n3724), .ZN(n2830) );
  NAND2_X1 U3602 ( .A1(n4409), .A2(n4161), .ZN(n2820) );
  INV_X1 U3603 ( .A(n2788), .ZN(n2876) );
  NAND2_X1 U3604 ( .A1(n2876), .A2(n3765), .ZN(n2819) );
  AND2_X1 U3605 ( .A1(n2822), .A2(n2821), .ZN(n4436) );
  NAND2_X1 U3606 ( .A1(n4409), .A2(n3765), .ZN(n2938) );
  INV_X1 U3607 ( .A(n2938), .ZN(n2882) );
  OR2_X1 U3608 ( .A1(n2484), .A2(n2823), .ZN(n2825) );
  NAND2_X1 U3609 ( .A1(n2882), .A2(n4414), .ZN(n4613) );
  AOI21_X1 U3610 ( .B1(B_REG_SCAN_IN), .B2(n4436), .A(n4613), .ZN(n3954) );
  INV_X1 U3611 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U3612 ( .A1(n3703), .A2(REG1_REG_30__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3613 ( .A1(n2544), .A2(REG0_REG_30__SCAN_IN), .ZN(n2826) );
  OAI211_X1 U3614 ( .C1(n3707), .C2(n2828), .A(n2827), .B(n2826), .ZN(n3845)
         );
  AND2_X2 U3615 ( .A1(n2864), .A2(n2876), .ZN(n4609) );
  INV_X1 U3616 ( .A(n3732), .ZN(n3455) );
  AOI22_X1 U3617 ( .A1(n3846), .A2(n4610), .B1(n4609), .B2(n3455), .ZN(n2831)
         );
  NAND2_X1 U3618 ( .A1(n2832), .A2(IR_REG_31__SCAN_IN), .ZN(n2833) );
  MUX2_X1 U3619 ( .A(IR_REG_31__SCAN_IN), .B(n2833), .S(IR_REG_25__SCAN_IN), 
        .Z(n2834) );
  NAND2_X1 U3620 ( .A1(n2834), .A2(n2239), .ZN(n2872) );
  NAND2_X1 U3621 ( .A1(n2872), .A2(B_REG_SCAN_IN), .ZN(n2837) );
  NAND2_X1 U3622 ( .A1(n2845), .A2(n2846), .ZN(n2836) );
  MUX2_X1 U3623 ( .A(n2837), .B(B_REG_SCAN_IN), .S(n2844), .Z(n2842) );
  NAND2_X1 U3624 ( .A1(n2239), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  INV_X1 U3625 ( .A(IR_REG_26__SCAN_IN), .ZN(n2838) );
  MUX2_X1 U3626 ( .A(n2839), .B(IR_REG_31__SCAN_IN), .S(n2838), .Z(n2841) );
  NAND2_X1 U3627 ( .A1(n2841), .A2(n2840), .ZN(n2886) );
  INV_X1 U3628 ( .A(n2886), .ZN(n4408) );
  NAND2_X1 U3629 ( .A1(n2886), .A2(n2872), .ZN(n2933) );
  NAND2_X1 U3630 ( .A1(n3035), .A2(n2933), .ZN(n2860) );
  AND2_X1 U3631 ( .A1(n2788), .A2(n3949), .ZN(n2936) );
  OR2_X1 U3632 ( .A1(n2938), .A2(n2936), .ZN(n3032) );
  NAND2_X1 U3633 ( .A1(n3032), .A2(n2945), .ZN(n2847) );
  NOR2_X1 U3634 ( .A1(n3034), .A2(n2847), .ZN(n2859) );
  NOR2_X1 U3635 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .ZN(n2851)
         );
  NOR4_X1 U3636 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2850) );
  NOR4_X1 U3637 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2849) );
  NOR4_X1 U3638 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2848) );
  NAND4_X1 U3639 ( .A1(n2851), .A2(n2850), .A3(n2849), .A4(n2848), .ZN(n2857)
         );
  NOR4_X1 U3640 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2855) );
  NOR4_X1 U3641 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2854) );
  NOR4_X1 U3642 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2853) );
  NOR4_X1 U3643 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2852) );
  NAND4_X1 U3644 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .ZN(n2856)
         );
  NOR2_X1 U3645 ( .A1(n2857), .A2(n2856), .ZN(n2858) );
  NAND3_X1 U3646 ( .A1(n2860), .A2(n2859), .A3(n2934), .ZN(n2867) );
  NAND2_X1 U3647 ( .A1(n2887), .A2(n2886), .ZN(n2861) );
  INV_X1 U3648 ( .A(n2863), .ZN(n2866) );
  INV_X1 U3649 ( .A(n4624), .ZN(n3092) );
  NAND2_X1 U3650 ( .A1(n3278), .A2(n3160), .ZN(n3161) );
  NAND2_X1 U3651 ( .A1(n4603), .A2(n4330), .ZN(n3400) );
  NAND2_X1 U3652 ( .A1(n2866), .A2(n2865), .ZN(U3547) );
  NAND2_X1 U3653 ( .A1(n2870), .A2(n2869), .ZN(U3515) );
  NOR2_X2 U3654 ( .A1(n2890), .A2(n2917), .ZN(U4043) );
  INV_X2 U3655 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3656 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2871) );
  OAI21_X1 U3657 ( .B1(n2872), .B2(U3149), .A(n2871), .ZN(U3327) );
  MUX2_X1 U3658 ( .A(n2873), .B(n3949), .S(STATE_REG_SCAN_IN), .Z(n2874) );
  INV_X1 U3659 ( .A(n2874), .ZN(U3333) );
  INV_X1 U3660 ( .A(DATAI_21_), .ZN(n5055) );
  NAND2_X1 U3661 ( .A1(n3765), .A2(STATE_REG_SCAN_IN), .ZN(n2875) );
  OAI21_X1 U3662 ( .B1(STATE_REG_SCAN_IN), .B2(n5055), .A(n2875), .ZN(U3331)
         );
  INV_X1 U3663 ( .A(DATAI_20_), .ZN(n2878) );
  NAND2_X1 U3664 ( .A1(n2876), .A2(STATE_REG_SCAN_IN), .ZN(n2877) );
  OAI21_X1 U3665 ( .B1(STATE_REG_SCAN_IN), .B2(n2878), .A(n2877), .ZN(U3332)
         );
  INV_X1 U3666 ( .A(DATAI_27_), .ZN(n5052) );
  NAND2_X1 U3667 ( .A1(n4436), .A2(STATE_REG_SCAN_IN), .ZN(n2879) );
  OAI21_X1 U3668 ( .B1(STATE_REG_SCAN_IN), .B2(n5052), .A(n2879), .ZN(U3325)
         );
  INV_X1 U3669 ( .A(DATAI_29_), .ZN(n4985) );
  NAND2_X1 U3670 ( .A1(n2880), .A2(STATE_REG_SCAN_IN), .ZN(n2881) );
  OAI21_X1 U3671 ( .B1(STATE_REG_SCAN_IN), .B2(n4985), .A(n2881), .ZN(U3323)
         );
  OR2_X1 U3672 ( .A1(n2998), .A2(U3149), .ZN(n3843) );
  NAND2_X1 U3673 ( .A1(n3034), .A2(n3843), .ZN(n2896) );
  NAND2_X1 U3674 ( .A1(n2882), .A2(n2998), .ZN(n2883) );
  AND2_X1 U3675 ( .A1(n2883), .A2(n3702), .ZN(n2895) );
  INV_X1 U3676 ( .A(n2895), .ZN(n2884) );
  NOR2_X1 U3677 ( .A1(n4578), .A2(U4043), .ZN(U3148) );
  NAND3_X1 U3678 ( .A1(n2887), .A2(n4644), .A3(n2886), .ZN(n2888) );
  OAI21_X1 U3679 ( .B1(n4643), .B2(D_REG_0__SCAN_IN), .A(n2888), .ZN(n2889) );
  INV_X1 U3680 ( .A(n2889), .ZN(U3458) );
  OAI22_X1 U3681 ( .A1(n4643), .A2(D_REG_1__SCAN_IN), .B1(n2933), .B2(n2890), 
        .ZN(n2891) );
  INV_X1 U3682 ( .A(n2891), .ZN(U3459) );
  INV_X1 U3683 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2898) );
  AND2_X1 U3684 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3862)
         );
  NAND2_X1 U3685 ( .A1(n4413), .A2(REG1_REG_1__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U3686 ( .A1(n3861), .A2(n2892), .ZN(n3880) );
  INV_X1 U3687 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2893) );
  MUX2_X1 U3688 ( .A(REG1_REG_2__SCAN_IN), .B(n2893), .S(n4412), .Z(n3881) );
  NAND2_X1 U3689 ( .A1(n3880), .A2(n3881), .ZN(n3879) );
  NAND2_X1 U3690 ( .A1(n4412), .A2(REG1_REG_2__SCAN_IN), .ZN(n2894) );
  NAND2_X1 U3691 ( .A1(n3879), .A2(n2894), .ZN(n2910) );
  XNOR2_X1 U3692 ( .A(n2910), .B(n4411), .ZN(n2897) );
  NOR2_X1 U3693 ( .A1(n2898), .A2(n2897), .ZN(n2911) );
  INV_X1 U3694 ( .A(n4436), .ZN(n2927) );
  INV_X1 U3695 ( .A(n4580), .ZN(n4452) );
  AOI211_X1 U3696 ( .C1(n2898), .C2(n2897), .A(n2911), .B(n4452), .ZN(n2905)
         );
  INV_X1 U3697 ( .A(n4411), .ZN(n2907) );
  INV_X1 U3698 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2900) );
  MUX2_X1 U3699 ( .A(n2900), .B(REG2_REG_1__SCAN_IN), .S(n2899), .Z(n3864) );
  NAND3_X1 U3700 ( .A1(n3864), .A2(REG2_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n3876) );
  NAND2_X1 U3701 ( .A1(n4413), .A2(REG2_REG_1__SCAN_IN), .ZN(n3875) );
  MUX2_X1 U3702 ( .A(n2502), .B(REG2_REG_2__SCAN_IN), .S(n4412), .Z(n3874) );
  AOI21_X1 U3703 ( .B1(n3876), .B2(n3875), .A(n3874), .ZN(n3873) );
  AOI21_X1 U3704 ( .B1(n4412), .B2(REG2_REG_2__SCAN_IN), .A(n3873), .ZN(n2908)
         );
  XNOR2_X1 U3705 ( .A(n2908), .B(n4411), .ZN(n2901) );
  NOR2_X1 U3706 ( .A1(n2927), .A2(n4414), .ZN(n3839) );
  NAND2_X1 U3707 ( .A1(REG2_REG_3__SCAN_IN), .A2(n2901), .ZN(n2906) );
  OAI211_X1 U3708 ( .C1(REG2_REG_3__SCAN_IN), .C2(n2901), .A(n4527), .B(n2906), 
        .ZN(n2903) );
  NOR2_X1 U3709 ( .A1(STATE_REG_SCAN_IN), .A2(n2519), .ZN(n3003) );
  AOI21_X1 U3710 ( .B1(n4578), .B2(ADDR_REG_3__SCAN_IN), .A(n3003), .ZN(n2902)
         );
  OAI211_X1 U3711 ( .C1(n4586), .C2(n2907), .A(n2903), .B(n2902), .ZN(n2904)
         );
  OR2_X1 U3712 ( .A1(n2905), .A2(n2904), .ZN(U3243) );
  OAI21_X1 U3713 ( .B1(n2908), .B2(n2907), .A(n2906), .ZN(n3888) );
  XNOR2_X1 U3714 ( .A(n3888), .B(n4410), .ZN(n3891) );
  XNOR2_X1 U3715 ( .A(n3891), .B(REG2_REG_4__SCAN_IN), .ZN(n2915) );
  NOR2_X1 U3716 ( .A1(STATE_REG_SCAN_IN), .A2(n2527), .ZN(n3085) );
  AOI21_X1 U3717 ( .B1(n4578), .B2(ADDR_REG_4__SCAN_IN), .A(n3085), .ZN(n2909)
         );
  OAI21_X1 U3718 ( .B1(n4586), .B2(n2295), .A(n2909), .ZN(n2914) );
  INV_X1 U3719 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4718) );
  AOI211_X1 U3720 ( .C1(n4718), .C2(n2912), .A(n3918), .B(n4452), .ZN(n2913)
         );
  AOI211_X1 U3721 ( .C1(n4527), .C2(n2915), .A(n2914), .B(n2913), .ZN(n2932)
         );
  INV_X1 U3722 ( .A(n3040), .ZN(n2916) );
  INV_X1 U3723 ( .A(n2954), .ZN(n3463) );
  NAND2_X1 U3724 ( .A1(n4611), .A2(n3463), .ZN(n2919) );
  NAND2_X1 U3725 ( .A1(n2922), .A2(n4624), .ZN(n2918) );
  INV_X1 U3726 ( .A(n2917), .ZN(n2921) );
  NAND2_X1 U3727 ( .A1(n2921), .A2(REG1_REG_0__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3728 ( .A1(n2960), .A2(n2920), .ZN(n2926) );
  AOI22_X1 U3729 ( .A1(n3463), .A2(n4624), .B1(n2921), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2925) );
  NAND2_X4 U3730 ( .A1(n2922), .A2(n4693), .ZN(n3538) );
  NAND2_X1 U3731 ( .A1(n2923), .A2(n4611), .ZN(n2924) );
  INV_X1 U3732 ( .A(n4414), .ZN(n2949) );
  NAND3_X1 U3733 ( .A1(n2973), .A2(n2949), .A3(n2927), .ZN(n2931) );
  AND2_X1 U3734 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3865)
         );
  NAND2_X1 U3735 ( .A1(n4436), .A2(n2928), .ZN(n2929) );
  NAND2_X1 U3736 ( .A1(n2949), .A2(n2929), .ZN(n4437) );
  AOI22_X1 U3737 ( .A1(n3839), .A2(n3865), .B1(n4437), .B2(n2277), .ZN(n2930)
         );
  NAND3_X1 U3738 ( .A1(n2931), .A2(U4043), .A3(n2930), .ZN(n3885) );
  NAND2_X1 U3739 ( .A1(n2932), .A2(n3885), .ZN(U3244) );
  NAND3_X1 U3740 ( .A1(n2935), .A2(n3038), .A3(n3035), .ZN(n2964) );
  INV_X1 U3741 ( .A(n2936), .ZN(n2937) );
  NAND2_X1 U3742 ( .A1(n2864), .A2(n2937), .ZN(n2939) );
  NAND2_X1 U3743 ( .A1(n2939), .A2(n2938), .ZN(n2965) );
  NAND2_X1 U3744 ( .A1(n4590), .A2(n2965), .ZN(n2940) );
  NAND2_X1 U3745 ( .A1(n2964), .A2(n2940), .ZN(n2941) );
  NAND2_X1 U3746 ( .A1(n2941), .A2(n3032), .ZN(n3000) );
  INV_X1 U3747 ( .A(n3000), .ZN(n2943) );
  NAND2_X1 U3748 ( .A1(n4644), .A2(n2956), .ZN(n2942) );
  NOR2_X1 U3749 ( .A1(n2224), .A2(n2942), .ZN(n3840) );
  NAND2_X1 U3750 ( .A1(n2964), .A2(n3840), .ZN(n3001) );
  NAND3_X1 U3751 ( .A1(n2943), .A2(n2947), .A3(n3001), .ZN(n3015) );
  INV_X1 U3752 ( .A(n3015), .ZN(n2972) );
  INV_X1 U3753 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3754 ( .A1(n2947), .A2(n4609), .ZN(n2944) );
  OR2_X1 U3755 ( .A1(n2964), .A2(n2944), .ZN(n2948) );
  NAND2_X2 U3756 ( .A1(n2948), .A2(n4190), .ZN(n3674) );
  NAND2_X1 U3757 ( .A1(n3840), .A2(n2949), .ZN(n2950) );
  NAND2_X1 U3758 ( .A1(n3840), .A2(n4414), .ZN(n2951) );
  OAI22_X1 U3759 ( .A1(n2952), .A2(n4415), .B1(n3665), .B2(n2516), .ZN(n2953)
         );
  AOI21_X1 U3760 ( .B1(n4625), .B2(n3674), .A(n2953), .ZN(n2970) );
  INV_X1 U3761 ( .A(n2956), .ZN(n2957) );
  OAI22_X1 U3762 ( .A1(n2955), .A2(n3538), .B1(n2954), .B2(n2959), .ZN(n2986)
         );
  XNOR2_X1 U3763 ( .A(n2985), .B(n2986), .ZN(n2963) );
  NAND2_X1 U3764 ( .A1(n2960), .A2(n3536), .ZN(n2961) );
  NAND2_X1 U3765 ( .A1(n2962), .A2(n2961), .ZN(n2968) );
  NAND2_X1 U3766 ( .A1(n2968), .A2(n2963), .ZN(n2989) );
  INV_X1 U3767 ( .A(n2964), .ZN(n2967) );
  NOR2_X1 U3768 ( .A1(n3034), .A2(n2965), .ZN(n2966) );
  AND2_X2 U3769 ( .A1(n2967), .A2(n2966), .ZN(n4426) );
  OAI211_X1 U3770 ( .C1(n2963), .C2(n2968), .A(n2989), .B(n4426), .ZN(n2969)
         );
  OAI211_X1 U3771 ( .C1(n2972), .C2(n2971), .A(n2970), .B(n2969), .ZN(U3219)
         );
  INV_X1 U3772 ( .A(n3674), .ZN(n4418) );
  NAND2_X1 U3773 ( .A1(n3015), .A2(REG3_REG_0__SCAN_IN), .ZN(n2977) );
  INV_X1 U3774 ( .A(n2973), .ZN(n2975) );
  AOI22_X1 U3775 ( .A1(n4426), .A2(n2975), .B1(n4421), .B2(n2974), .ZN(n2976)
         );
  OAI211_X1 U3776 ( .C1(n4418), .C2(n3092), .A(n2977), .B(n2976), .ZN(U3229)
         );
  NAND2_X1 U3777 ( .A1(n2982), .A2(n3518), .ZN(n2980) );
  NAND2_X1 U3778 ( .A1(n2922), .A2(n3771), .ZN(n2979) );
  NAND2_X1 U3779 ( .A1(n2923), .A2(n2982), .ZN(n2984) );
  NAND2_X1 U3780 ( .A1(n3518), .A2(n3771), .ZN(n2983) );
  NAND2_X1 U3781 ( .A1(n2984), .A2(n2983), .ZN(n3075) );
  XNOR2_X1 U3782 ( .A(n3077), .B(n3075), .ZN(n3073) );
  INV_X1 U3783 ( .A(n2985), .ZN(n2987) );
  NAND2_X1 U3784 ( .A1(n2987), .A2(n2986), .ZN(n2988) );
  NAND2_X1 U3785 ( .A1(n2989), .A2(n2988), .ZN(n3010) );
  INV_X1 U3786 ( .A(n3010), .ZN(n2992) );
  XNOR2_X1 U3787 ( .A(n2990), .B(n3526), .ZN(n2993) );
  OAI22_X1 U3788 ( .A1(n2516), .A2(n3538), .B1(n3525), .B2(n2408), .ZN(n2994)
         );
  XNOR2_X1 U3789 ( .A(n2993), .B(n2994), .ZN(n3009) );
  INV_X1 U3790 ( .A(n3009), .ZN(n2991) );
  NAND2_X1 U3791 ( .A1(n2992), .A2(n2991), .ZN(n3011) );
  INV_X1 U3792 ( .A(n2993), .ZN(n2996) );
  INV_X1 U3793 ( .A(n2994), .ZN(n2995) );
  NAND2_X1 U3794 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  NAND2_X1 U3795 ( .A1(n3011), .A2(n2997), .ZN(n3074) );
  XNOR2_X1 U3796 ( .A(n3073), .B(n3074), .ZN(n3007) );
  NAND2_X1 U3797 ( .A1(n2917), .A2(n2998), .ZN(n2999) );
  OAI21_X1 U3798 ( .B1(n3000), .B2(n2999), .A(STATE_REG_SCAN_IN), .ZN(n3002)
         );
  AOI21_X1 U3799 ( .B1(n4421), .B2(n3859), .A(n3003), .ZN(n3005) );
  AOI22_X1 U3800 ( .A1(n3675), .A2(n2506), .B1(n3674), .B2(n3771), .ZN(n3004)
         );
  OAI211_X1 U3801 ( .C1(n4431), .C2(REG3_REG_3__SCAN_IN), .A(n3005), .B(n3004), 
        .ZN(n3006) );
  AOI21_X1 U3802 ( .B1(n3007), .B2(n4426), .A(n3006), .ZN(n3008) );
  INV_X1 U3803 ( .A(n3008), .ZN(U3215) );
  INV_X1 U3804 ( .A(n3011), .ZN(n3012) );
  AOI21_X1 U3805 ( .B1(n3009), .B2(n3010), .A(n3012), .ZN(n3017) );
  INV_X1 U3806 ( .A(n4426), .ZN(n3669) );
  AOI22_X1 U3807 ( .A1(n4421), .A2(n2982), .B1(n3675), .B2(n2974), .ZN(n3013)
         );
  OAI21_X1 U3808 ( .B1(n4418), .B2(n2408), .A(n3013), .ZN(n3014) );
  AOI21_X1 U3809 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3015), .A(n3014), .ZN(n3016)
         );
  OAI21_X1 U3810 ( .B1(n3017), .B2(n3669), .A(n3016), .ZN(U3234) );
  INV_X1 U3811 ( .A(n4669), .ZN(n4702) );
  XNOR2_X1 U3812 ( .A(n3018), .B(n3021), .ZN(n3025) );
  INV_X1 U3813 ( .A(n3025), .ZN(n3209) );
  AOI22_X1 U3814 ( .A1(n3859), .A2(n4596), .B1(n4609), .B2(n3771), .ZN(n3019)
         );
  OAI21_X1 U3815 ( .B1(n2516), .B2(n4592), .A(n3019), .ZN(n3026) );
  INV_X1 U3816 ( .A(n3021), .ZN(n3714) );
  NAND3_X1 U3817 ( .A1(n3020), .A2(n3767), .A3(n3714), .ZN(n3022) );
  AND2_X1 U3818 ( .A1(n3023), .A2(n3022), .ZN(n3024) );
  OAI22_X1 U3819 ( .A1(n3025), .A2(n4617), .B1(n3024), .B2(n4598), .ZN(n3202)
         );
  AOI211_X1 U3820 ( .C1(n4702), .C2(n3209), .A(n3026), .B(n3202), .ZN(n3031)
         );
  INV_X1 U3821 ( .A(n4677), .ZN(n3135) );
  AND2_X1 U3822 ( .A1(n3047), .A2(n3771), .ZN(n3027) );
  NOR2_X1 U3823 ( .A1(n3059), .A2(n3027), .ZN(n3203) );
  AOI22_X1 U3824 ( .A1(n3135), .A2(n3203), .B1(REG0_REG_3__SCAN_IN), .B2(n4706), .ZN(n3028) );
  OAI21_X1 U3825 ( .B1(n3031), .B2(n4706), .A(n3028), .ZN(U3473) );
  NAND2_X1 U3826 ( .A1(n4726), .A2(REG1_REG_3__SCAN_IN), .ZN(n3030) );
  INV_X1 U3827 ( .A(n4714), .ZN(n3137) );
  NAND2_X1 U3828 ( .A1(n3137), .A2(n3203), .ZN(n3029) );
  OAI211_X1 U3829 ( .C1(n3031), .C2(n4726), .A(n3030), .B(n3029), .ZN(U3521)
         );
  INV_X1 U3830 ( .A(n3032), .ZN(n3033) );
  NOR2_X1 U3831 ( .A1(n3034), .A2(n3033), .ZN(n3037) );
  NAND4_X1 U3832 ( .A1(n3038), .A2(n3037), .A3(n3036), .A4(n3035), .ZN(n3039)
         );
  OR2_X1 U3833 ( .A1(n3040), .A2(n3949), .ZN(n3244) );
  INV_X1 U3834 ( .A(n3244), .ZN(n3041) );
  NAND2_X1 U3835 ( .A1(n4616), .A2(n3042), .ZN(n3043) );
  NAND2_X1 U3836 ( .A1(n3043), .A2(n3718), .ZN(n3044) );
  NAND2_X1 U3837 ( .A1(n3045), .A2(n3044), .ZN(n4675) );
  AND2_X1 U3838 ( .A1(n4701), .A2(n3949), .ZN(n3046) );
  OAI21_X1 U3839 ( .B1(n4623), .B2(n2408), .A(n3047), .ZN(n4713) );
  INV_X1 U3840 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3048) );
  OAI22_X1 U3841 ( .A1(n4180), .A2(n4713), .B1(n3048), .B2(n4190), .ZN(n3057)
         );
  NAND3_X1 U3842 ( .A1(n2407), .A2(n3766), .A3(n4608), .ZN(n3049) );
  NAND2_X1 U3843 ( .A1(n3020), .A2(n3049), .ZN(n3053) );
  AOI22_X1 U3844 ( .A1(n2982), .A2(n4596), .B1(n3050), .B2(n4609), .ZN(n3051)
         );
  OAI21_X1 U3845 ( .B1(n2955), .B2(n4592), .A(n3051), .ZN(n3052) );
  AOI21_X1 U3846 ( .B1(n3053), .B2(n4621), .A(n3052), .ZN(n3055) );
  INV_X1 U3847 ( .A(n4617), .ZN(n4601) );
  NAND2_X1 U3848 ( .A1(n4675), .A2(n4601), .ZN(n3054) );
  NAND2_X1 U3849 ( .A1(n3055), .A2(n3054), .ZN(n4674) );
  MUX2_X1 U3850 ( .A(REG2_REG_2__SCAN_IN), .B(n4674), .S(n4205), .Z(n3056) );
  AOI211_X1 U3851 ( .C1(n4631), .C2(n4675), .A(n3057), .B(n3056), .ZN(n3058)
         );
  INV_X1 U3852 ( .A(n3058), .ZN(U3288) );
  OAI211_X1 U3853 ( .C1(n3059), .C2(n3071), .A(n3140), .B(n4701), .ZN(n4680)
         );
  NOR2_X1 U3854 ( .A1(n4680), .A2(n4161), .ZN(n3066) );
  XNOR2_X1 U3855 ( .A(n3060), .B(n3693), .ZN(n3067) );
  XOR2_X1 U3856 ( .A(n3693), .B(n3061), .Z(n3064) );
  AOI22_X1 U3857 ( .A1(n3858), .A2(n4596), .B1(n3086), .B2(n4609), .ZN(n3062)
         );
  OAI21_X1 U3858 ( .B1(n3772), .B2(n4592), .A(n3062), .ZN(n3063) );
  AOI21_X1 U3859 ( .B1(n3064), .B2(n4621), .A(n3063), .ZN(n3065) );
  OAI21_X1 U3860 ( .B1(n3067), .B2(n4617), .A(n3065), .ZN(n4681) );
  AOI211_X1 U3861 ( .C1(n4622), .C2(n3084), .A(n3066), .B(n4681), .ZN(n3069)
         );
  INV_X2 U3862 ( .A(n4205), .ZN(n4634) );
  INV_X1 U3863 ( .A(n3067), .ZN(n4683) );
  AOI22_X1 U3864 ( .A1(n4683), .A2(n4631), .B1(REG2_REG_4__SCAN_IN), .B2(n4634), .ZN(n3068) );
  OAI21_X1 U3865 ( .B1(n3069), .B2(n4634), .A(n3068), .ZN(U3286) );
  INV_X1 U3866 ( .A(n3463), .ZN(n3525) );
  OAI22_X1 U3867 ( .A1(n3072), .A2(n3525), .B1(n3508), .B2(n3071), .ZN(n3070)
         );
  XNOR2_X1 U3868 ( .A(n3070), .B(n3526), .ZN(n3100) );
  OAI22_X1 U3869 ( .A1(n3072), .A2(n3538), .B1(n3525), .B2(n3071), .ZN(n3099)
         );
  XNOR2_X1 U3870 ( .A(n3100), .B(n3099), .ZN(n3083) );
  NAND2_X1 U3871 ( .A1(n3074), .A2(n3073), .ZN(n3079) );
  INV_X1 U3872 ( .A(n3075), .ZN(n3076) );
  NAND2_X1 U3873 ( .A1(n3077), .A2(n3076), .ZN(n3078) );
  INV_X1 U3874 ( .A(n3102), .ZN(n3082) );
  AOI211_X1 U3875 ( .C1(n3083), .C2(n3080), .A(n3669), .B(n3082), .ZN(n3091)
         );
  INV_X1 U3876 ( .A(n3084), .ZN(n3089) );
  AOI21_X1 U3877 ( .B1(n4421), .B2(n3858), .A(n3085), .ZN(n3088) );
  AOI22_X1 U3878 ( .A1(n3675), .A2(n2982), .B1(n3674), .B2(n3086), .ZN(n3087)
         );
  OAI211_X1 U3879 ( .C1(n4431), .C2(n3089), .A(n3088), .B(n3087), .ZN(n3090)
         );
  OR2_X1 U3880 ( .A1(n3091), .A2(n3090), .ZN(U3227) );
  NAND2_X1 U3881 ( .A1(n4611), .A2(n3092), .ZN(n3764) );
  AND2_X1 U3882 ( .A1(n3762), .A2(n3764), .ZN(n4665) );
  INV_X1 U3883 ( .A(n4631), .ZN(n4221) );
  INV_X1 U3884 ( .A(n3093), .ZN(n3095) );
  NAND2_X1 U3885 ( .A1(n4624), .A2(n2864), .ZN(n4663) );
  AOI21_X1 U3886 ( .B1(n4598), .B2(n4617), .A(n4665), .ZN(n3094) );
  AOI21_X1 U3887 ( .B1(n4596), .B2(n2974), .A(n3094), .ZN(n4664) );
  OAI21_X1 U3888 ( .B1(n3095), .B2(n4663), .A(n4664), .ZN(n3096) );
  AOI22_X1 U3889 ( .A1(n3096), .A2(n4205), .B1(REG3_REG_0__SCAN_IN), .B2(n4622), .ZN(n3098) );
  NAND2_X1 U3890 ( .A1(n4634), .A2(REG2_REG_0__SCAN_IN), .ZN(n3097) );
  OAI211_X1 U3891 ( .C1(n4665), .C2(n4221), .A(n3098), .B(n3097), .ZN(U3290)
         );
  NAND2_X1 U3892 ( .A1(n3100), .A2(n3099), .ZN(n3101) );
  NAND2_X1 U3893 ( .A1(n3858), .A2(n3463), .ZN(n3104) );
  NAND2_X1 U3894 ( .A1(n2922), .A2(n3598), .ZN(n3103) );
  NAND2_X1 U3895 ( .A1(n3104), .A2(n3103), .ZN(n3105) );
  XNOR2_X1 U3896 ( .A(n3105), .B(n3536), .ZN(n3108) );
  NAND2_X1 U3897 ( .A1(n2923), .A2(n3858), .ZN(n3107) );
  NAND2_X1 U3898 ( .A1(n3518), .A2(n3598), .ZN(n3106) );
  NAND2_X1 U3899 ( .A1(n3107), .A2(n3106), .ZN(n3109) );
  XNOR2_X1 U3900 ( .A(n3108), .B(n3109), .ZN(n3597) );
  NAND2_X1 U3901 ( .A1(n3595), .A2(n3597), .ZN(n3596) );
  INV_X1 U3902 ( .A(n3108), .ZN(n3110) );
  NAND2_X1 U3903 ( .A1(n3110), .A2(n3109), .ZN(n3111) );
  NAND2_X1 U3904 ( .A1(n3596), .A2(n3111), .ZN(n3170) );
  NAND2_X1 U3905 ( .A1(n3857), .A2(n3518), .ZN(n3113) );
  NAND2_X1 U3906 ( .A1(n2922), .A2(n3246), .ZN(n3112) );
  NAND2_X1 U3907 ( .A1(n3113), .A2(n3112), .ZN(n3114) );
  XNOR2_X1 U3908 ( .A(n3114), .B(n3526), .ZN(n3168) );
  NAND2_X1 U3909 ( .A1(n2923), .A2(n3857), .ZN(n3116) );
  NAND2_X1 U3910 ( .A1(n3518), .A2(n3246), .ZN(n3115) );
  NAND2_X1 U3911 ( .A1(n3116), .A2(n3115), .ZN(n3169) );
  XNOR2_X1 U3912 ( .A(n3168), .B(n3169), .ZN(n3117) );
  XNOR2_X1 U3913 ( .A(n3170), .B(n3117), .ZN(n3122) );
  INV_X1 U3914 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3118) );
  NOR2_X1 U3915 ( .A1(STATE_REG_SCAN_IN), .A2(n3118), .ZN(n4456) );
  AOI21_X1 U3916 ( .B1(n3675), .B2(n3858), .A(n4456), .ZN(n3120) );
  AOI22_X1 U3917 ( .A1(n4421), .A2(n3855), .B1(n3674), .B2(n3246), .ZN(n3119)
         );
  OAI211_X1 U3918 ( .C1(n4431), .C2(n3247), .A(n3120), .B(n3119), .ZN(n3121)
         );
  AOI21_X1 U3919 ( .B1(n3122), .B2(n4426), .A(n3121), .ZN(n3123) );
  INV_X1 U3920 ( .A(n3123), .ZN(U3236) );
  OR2_X1 U3921 ( .A1(n3124), .A2(n3125), .ZN(n3127) );
  NAND2_X1 U3922 ( .A1(n3127), .A2(n3126), .ZN(n3128) );
  NAND2_X1 U3923 ( .A1(n3778), .A2(n3786), .ZN(n3696) );
  XNOR2_X1 U3924 ( .A(n3128), .B(n3696), .ZN(n3257) );
  XOR2_X1 U3925 ( .A(n3696), .B(n3129), .Z(n3130) );
  NAND2_X1 U3926 ( .A1(n3130), .A2(n4621), .ZN(n3255) );
  AOI22_X1 U3927 ( .A1(n3855), .A2(n4596), .B1(n3246), .B2(n4609), .ZN(n3131)
         );
  OAI211_X1 U3928 ( .C1(n3132), .C2(n4592), .A(n3255), .B(n3131), .ZN(n3133)
         );
  AOI21_X1 U3929 ( .B1(n4686), .B2(n3257), .A(n3133), .ZN(n3139) );
  AND2_X1 U3930 ( .A1(n3142), .A2(n3246), .ZN(n3134) );
  NOR2_X1 U3931 ( .A1(n3277), .A2(n3134), .ZN(n3252) );
  AOI22_X1 U3932 ( .A1(n3252), .A2(n3135), .B1(n4706), .B2(REG0_REG_6__SCAN_IN), .ZN(n3136) );
  OAI21_X1 U3933 ( .B1(n3139), .B2(n4706), .A(n3136), .ZN(U3479) );
  AOI22_X1 U3934 ( .A1(n3252), .A2(n3137), .B1(n4726), .B2(REG1_REG_6__SCAN_IN), .ZN(n3138) );
  OAI21_X1 U3935 ( .B1(n3139), .B2(n4726), .A(n3138), .ZN(U3524) );
  NAND2_X1 U3936 ( .A1(n3140), .A2(n3598), .ZN(n3141) );
  NAND2_X1 U3937 ( .A1(n3142), .A2(n3141), .ZN(n3261) );
  NAND2_X1 U3938 ( .A1(n2253), .A2(n3785), .ZN(n3694) );
  XNOR2_X1 U3939 ( .A(n3124), .B(n3694), .ZN(n3266) );
  OAI22_X1 U3940 ( .A1(n3286), .A2(n4613), .B1(n4590), .B2(n3143), .ZN(n3146)
         );
  XOR2_X1 U3941 ( .A(n3694), .B(n3144), .Z(n3145) );
  NOR2_X1 U3942 ( .A1(n3145), .A2(n4598), .ZN(n3264) );
  AOI211_X1 U3943 ( .C1(n4610), .C2(n3859), .A(n3146), .B(n3264), .ZN(n3147)
         );
  OAI21_X1 U3944 ( .B1(n4337), .B2(n3266), .A(n3147), .ZN(n3150) );
  NAND2_X1 U3945 ( .A1(n3150), .A2(n4729), .ZN(n3149) );
  NAND2_X1 U3946 ( .A1(n4726), .A2(REG1_REG_5__SCAN_IN), .ZN(n3148) );
  OAI211_X1 U3947 ( .C1(n4714), .C2(n3261), .A(n3149), .B(n3148), .ZN(U3523)
         );
  NAND2_X1 U3948 ( .A1(n3150), .A2(n4708), .ZN(n3152) );
  NAND2_X1 U3949 ( .A1(n4706), .A2(REG0_REG_5__SCAN_IN), .ZN(n3151) );
  OAI211_X1 U3950 ( .C1(n3261), .C2(n4677), .A(n3152), .B(n3151), .ZN(U3477)
         );
  NAND2_X1 U3951 ( .A1(n3782), .A2(n3787), .ZN(n3697) );
  XNOR2_X1 U3952 ( .A(n3153), .B(n3697), .ZN(n3159) );
  XNOR2_X1 U3953 ( .A(n3154), .B(n3697), .ZN(n3157) );
  AOI22_X1 U3954 ( .A1(n3853), .A2(n4596), .B1(n3195), .B2(n4609), .ZN(n3155)
         );
  OAI21_X1 U3955 ( .B1(n3249), .B2(n4592), .A(n3155), .ZN(n3156) );
  AOI21_X1 U3956 ( .B1(n3157), .B2(n4621), .A(n3156), .ZN(n3158) );
  OAI21_X1 U3957 ( .B1(n3159), .B2(n4617), .A(n3158), .ZN(n4690) );
  INV_X1 U3958 ( .A(n4690), .ZN(n3167) );
  INV_X1 U3959 ( .A(n3159), .ZN(n4692) );
  NOR2_X1 U3960 ( .A1(n3278), .A2(n3160), .ZN(n4689) );
  INV_X1 U3961 ( .A(n3161), .ZN(n4688) );
  NOR3_X1 U3962 ( .A1(n4689), .A2(n4688), .A3(n4180), .ZN(n3165) );
  INV_X1 U3963 ( .A(n3162), .ZN(n3198) );
  OAI22_X1 U3964 ( .A1(n4205), .A2(n3163), .B1(n3198), .B2(n4190), .ZN(n3164)
         );
  AOI211_X1 U3965 ( .C1(n4692), .C2(n4631), .A(n3165), .B(n3164), .ZN(n3166)
         );
  OAI21_X1 U3966 ( .B1(n3167), .B2(n4634), .A(n3166), .ZN(U3282) );
  OAI22_X1 U3967 ( .A1(n3249), .A2(n2224), .B1(n3508), .B2(n3172), .ZN(n3171)
         );
  XNOR2_X1 U3968 ( .A(n3171), .B(n3536), .ZN(n3181) );
  OAI22_X1 U3969 ( .A1(n3249), .A2(n3538), .B1(n2224), .B2(n3172), .ZN(n3182)
         );
  XNOR2_X1 U3970 ( .A(n3181), .B(n3182), .ZN(n3179) );
  XOR2_X1 U3971 ( .A(n3180), .B(n3179), .Z(n3177) );
  INV_X1 U3972 ( .A(n3173), .ZN(n3288) );
  INV_X1 U3973 ( .A(REG3_REG_7__SCAN_IN), .ZN(n5006) );
  NOR2_X1 U3974 ( .A1(STATE_REG_SCAN_IN), .A2(n5006), .ZN(n4468) );
  AOI21_X1 U3975 ( .B1(n4421), .B2(n3854), .A(n4468), .ZN(n3175) );
  AOI22_X1 U3976 ( .A1(n3675), .A2(n3857), .B1(n3674), .B2(n3283), .ZN(n3174)
         );
  OAI211_X1 U3977 ( .C1(n4431), .C2(n3288), .A(n3175), .B(n3174), .ZN(n3176)
         );
  AOI21_X1 U3978 ( .B1(n3177), .B2(n4426), .A(n3176), .ZN(n3178) );
  INV_X1 U3979 ( .A(n3178), .ZN(U3210) );
  INV_X1 U3980 ( .A(n3181), .ZN(n3183) );
  NAND2_X1 U3981 ( .A1(n3183), .A2(n3182), .ZN(n3222) );
  NAND2_X1 U3982 ( .A1(n3225), .A2(n3222), .ZN(n3344) );
  NAND2_X1 U3983 ( .A1(n3854), .A2(n3518), .ZN(n3185) );
  NAND2_X1 U3984 ( .A1(n2922), .A2(n3195), .ZN(n3184) );
  NAND2_X1 U3985 ( .A1(n3185), .A2(n3184), .ZN(n3186) );
  XNOR2_X1 U3986 ( .A(n3186), .B(n3526), .ZN(n3189) );
  NAND2_X1 U3987 ( .A1(n2923), .A2(n3854), .ZN(n3188) );
  NAND2_X1 U3988 ( .A1(n3518), .A2(n3195), .ZN(n3187) );
  NAND2_X1 U3989 ( .A1(n3188), .A2(n3187), .ZN(n3190) );
  AND2_X1 U3990 ( .A1(n3189), .A2(n3190), .ZN(n3267) );
  INV_X1 U3991 ( .A(n3267), .ZN(n3193) );
  INV_X1 U3992 ( .A(n3189), .ZN(n3192) );
  INV_X1 U3993 ( .A(n3190), .ZN(n3191) );
  NAND2_X1 U3994 ( .A1(n3192), .A2(n3191), .ZN(n3268) );
  NAND2_X1 U3995 ( .A1(n3193), .A2(n3268), .ZN(n3194) );
  XNOR2_X1 U3996 ( .A(n3344), .B(n3194), .ZN(n3200) );
  INV_X1 U3997 ( .A(REG3_REG_8__SCAN_IN), .ZN(n5084) );
  NOR2_X1 U3998 ( .A1(STATE_REG_SCAN_IN), .A2(n5084), .ZN(n4483) );
  AOI21_X1 U3999 ( .B1(n4421), .B2(n3853), .A(n4483), .ZN(n3197) );
  AOI22_X1 U4000 ( .A1(n3675), .A2(n3855), .B1(n3674), .B2(n3195), .ZN(n3196)
         );
  OAI211_X1 U4001 ( .C1(n4431), .C2(n3198), .A(n3197), .B(n3196), .ZN(n3199)
         );
  AOI21_X1 U4002 ( .B1(n3200), .B2(n4426), .A(n3199), .ZN(n3201) );
  INV_X1 U4003 ( .A(n3201), .ZN(U3218) );
  INV_X1 U4004 ( .A(n3202), .ZN(n3211) );
  NAND2_X1 U4005 ( .A1(n4205), .A2(n4610), .ZN(n4215) );
  NAND2_X1 U4006 ( .A1(n4205), .A2(n4596), .ZN(n4214) );
  INV_X1 U4007 ( .A(n4214), .ZN(n3407) );
  AOI22_X1 U4008 ( .A1(n3407), .A2(n3859), .B1(n4629), .B2(n3203), .ZN(n3207)
         );
  OAI22_X1 U4009 ( .A1(n4205), .A2(n3204), .B1(n4190), .B2(REG3_REG_3__SCAN_IN), .ZN(n3205) );
  AOI21_X1 U4010 ( .B1(n3771), .B2(n4175), .A(n3205), .ZN(n3206) );
  OAI211_X1 U4011 ( .C1(n2516), .C2(n4215), .A(n3207), .B(n3206), .ZN(n3208)
         );
  AOI21_X1 U4012 ( .B1(n3209), .B2(n4631), .A(n3208), .ZN(n3210) );
  OAI21_X1 U4013 ( .B1(n3211), .B2(n4634), .A(n3210), .ZN(U3287) );
  NAND2_X1 U4014 ( .A1(n3853), .A2(n3518), .ZN(n3213) );
  NAND2_X1 U4015 ( .A1(n2922), .A2(n3357), .ZN(n3212) );
  NAND2_X1 U4016 ( .A1(n3213), .A2(n3212), .ZN(n3214) );
  XNOR2_X1 U4017 ( .A(n3214), .B(n3536), .ZN(n3229) );
  NAND2_X1 U4018 ( .A1(n2923), .A2(n3853), .ZN(n3216) );
  NAND2_X1 U4019 ( .A1(n3518), .A2(n3357), .ZN(n3215) );
  NAND2_X1 U4020 ( .A1(n3216), .A2(n3215), .ZN(n3227) );
  XNOR2_X1 U4021 ( .A(n3229), .B(n3227), .ZN(n3270) );
  INV_X1 U4022 ( .A(n3270), .ZN(n3226) );
  OR2_X1 U4023 ( .A1(n3267), .A2(n3226), .ZN(n3343) );
  NAND2_X1 U4024 ( .A1(n3852), .A2(n3518), .ZN(n3218) );
  NAND2_X1 U4025 ( .A1(n2922), .A2(n3351), .ZN(n3217) );
  NAND2_X1 U4026 ( .A1(n3218), .A2(n3217), .ZN(n3219) );
  XNOR2_X1 U4027 ( .A(n3219), .B(n3526), .ZN(n3233) );
  NAND2_X1 U4028 ( .A1(n2923), .A2(n3852), .ZN(n3221) );
  NAND2_X1 U4029 ( .A1(n3518), .A2(n3351), .ZN(n3220) );
  NAND2_X1 U4030 ( .A1(n3221), .A2(n3220), .ZN(n3232) );
  AND2_X1 U4031 ( .A1(n3233), .A2(n3232), .ZN(n3235) );
  NOR2_X1 U4032 ( .A1(n3343), .A2(n3235), .ZN(n3223) );
  AND2_X1 U4033 ( .A1(n3223), .A2(n3222), .ZN(n3224) );
  OR2_X1 U4034 ( .A1(n3226), .A2(n3268), .ZN(n3231) );
  INV_X1 U4035 ( .A(n3227), .ZN(n3228) );
  NAND2_X1 U4036 ( .A1(n3229), .A2(n3228), .ZN(n3230) );
  AND2_X1 U4037 ( .A1(n3231), .A2(n3230), .ZN(n3345) );
  XNOR2_X1 U4038 ( .A(n3233), .B(n3232), .ZN(n3350) );
  INV_X1 U4039 ( .A(n3350), .ZN(n3234) );
  AND2_X1 U4040 ( .A1(n3345), .A2(n3234), .ZN(n3346) );
  NOR2_X1 U4041 ( .A1(n3235), .A2(n3346), .ZN(n3324) );
  OAI22_X1 U4042 ( .A1(n3375), .A2(n2224), .B1(n3508), .B2(n4591), .ZN(n3236)
         );
  XNOR2_X1 U40430 ( .A(n3236), .B(n3526), .ZN(n3320) );
  OAI22_X1 U4044 ( .A1(n3375), .A2(n3538), .B1(n2224), .B2(n4591), .ZN(n3322)
         );
  XNOR2_X1 U4045 ( .A(n3320), .B(n3322), .ZN(n3237) );
  XNOR2_X1 U4046 ( .A(n3321), .B(n3237), .ZN(n3242) );
  AND2_X1 U4047 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4515) );
  AOI21_X1 U4048 ( .B1(n4421), .B2(n4595), .A(n4515), .ZN(n3239) );
  AOI22_X1 U4049 ( .A1(n3675), .A2(n3852), .B1(n3674), .B2(n4605), .ZN(n3238)
         );
  OAI211_X1 U4050 ( .C1(n4431), .C2(n3240), .A(n3239), .B(n3238), .ZN(n3241)
         );
  AOI21_X1 U4051 ( .B1(n3242), .B2(n4426), .A(n3241), .ZN(n3243) );
  INV_X1 U4052 ( .A(n3243), .ZN(U3233) );
  NAND2_X1 U4053 ( .A1(n4617), .A2(n3244), .ZN(n3245) );
  INV_X1 U4054 ( .A(n4215), .ZN(n3405) );
  AOI22_X1 U4055 ( .A1(n3405), .A2(n3858), .B1(n4175), .B2(n3246), .ZN(n3254)
         );
  OAI22_X1 U4056 ( .A1(n4205), .A2(n3248), .B1(n3247), .B2(n4190), .ZN(n3251)
         );
  NOR2_X1 U4057 ( .A1(n4214), .A2(n3249), .ZN(n3250) );
  AOI211_X1 U4058 ( .C1(n3252), .C2(n4629), .A(n3251), .B(n3250), .ZN(n3253)
         );
  OAI211_X1 U4059 ( .C1(n3255), .C2(n4634), .A(n3254), .B(n3253), .ZN(n3256)
         );
  AOI21_X1 U4060 ( .B1(n4194), .B2(n3257), .A(n3256), .ZN(n3258) );
  INV_X1 U4061 ( .A(n3258), .ZN(U3284) );
  OAI22_X1 U4062 ( .A1(n3599), .A2(n4190), .B1(n2538), .B2(n4205), .ZN(n3263)
         );
  AOI22_X1 U4063 ( .A1(n3405), .A2(n3859), .B1(n3407), .B2(n3857), .ZN(n3260)
         );
  NAND2_X1 U4064 ( .A1(n4175), .A2(n3598), .ZN(n3259) );
  OAI211_X1 U4065 ( .C1(n3261), .C2(n4180), .A(n3260), .B(n3259), .ZN(n3262)
         );
  AOI211_X1 U4066 ( .C1(n3264), .C2(n4205), .A(n3263), .B(n3262), .ZN(n3265)
         );
  OAI21_X1 U4067 ( .B1(n4165), .B2(n3266), .A(n3265), .ZN(U3285) );
  OR2_X1 U4068 ( .A1(n3344), .A2(n3267), .ZN(n3269) );
  NAND2_X1 U4069 ( .A1(n3269), .A2(n3268), .ZN(n3271) );
  XNOR2_X1 U4070 ( .A(n3271), .B(n3270), .ZN(n3275) );
  NOR2_X1 U4071 ( .A1(STATE_REG_SCAN_IN), .A2(n2585), .ZN(n4494) );
  AOI21_X1 U4072 ( .B1(n4421), .B2(n3852), .A(n4494), .ZN(n3273) );
  AOI22_X1 U4073 ( .A1(n3675), .A2(n3854), .B1(n3674), .B2(n3357), .ZN(n3272)
         );
  OAI211_X1 U4074 ( .C1(n4431), .C2(n3296), .A(n3273), .B(n3272), .ZN(n3274)
         );
  AOI21_X1 U4075 ( .B1(n3275), .B2(n4426), .A(n3274), .ZN(n3276) );
  INV_X1 U4076 ( .A(n3276), .ZN(U3228) );
  INV_X1 U4077 ( .A(n3277), .ZN(n3279) );
  AOI211_X1 U4078 ( .C1(n3283), .C2(n3279), .A(n4693), .B(n3278), .ZN(n4685)
         );
  INV_X1 U4079 ( .A(n3280), .ZN(n3719) );
  XNOR2_X1 U4080 ( .A(n3281), .B(n3719), .ZN(n3282) );
  NAND2_X1 U4081 ( .A1(n3282), .A2(n4621), .ZN(n3285) );
  AOI22_X1 U4082 ( .A1(n3854), .A2(n4596), .B1(n4609), .B2(n3283), .ZN(n3284)
         );
  OAI211_X1 U4083 ( .C1(n3286), .C2(n4592), .A(n3285), .B(n3284), .ZN(n4684)
         );
  AOI21_X1 U4084 ( .B1(n4685), .B2(n3949), .A(n4684), .ZN(n3291) );
  XNOR2_X1 U4085 ( .A(n3287), .B(n3719), .ZN(n4687) );
  OAI22_X1 U4086 ( .A1(n4205), .A2(n2568), .B1(n3288), .B2(n4190), .ZN(n3289)
         );
  AOI21_X1 U4087 ( .B1(n4687), .B2(n4194), .A(n3289), .ZN(n3290) );
  OAI21_X1 U4088 ( .B1(n3291), .B2(n4634), .A(n3290), .ZN(U3283) );
  AND2_X1 U4089 ( .A1(n2263), .A2(n3783), .ZN(n3684) );
  XOR2_X1 U4090 ( .A(n3292), .B(n3684), .Z(n3293) );
  NAND2_X1 U4091 ( .A1(n3293), .A2(n4621), .ZN(n3359) );
  XOR2_X1 U4092 ( .A(n3294), .B(n3684), .Z(n3362) );
  NAND2_X1 U4093 ( .A1(n3362), .A2(n4194), .ZN(n3302) );
  OAI21_X1 U4094 ( .B1(n4688), .B2(n3295), .A(n3311), .ZN(n3368) );
  INV_X1 U4095 ( .A(n3368), .ZN(n3300) );
  INV_X1 U4096 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3887) );
  OAI22_X1 U4097 ( .A1(n3296), .A2(n4190), .B1(n3887), .B2(n4205), .ZN(n3299)
         );
  AOI22_X1 U4098 ( .A1(n3407), .A2(n3852), .B1(n4175), .B2(n3357), .ZN(n3297)
         );
  OAI21_X1 U4099 ( .B1(n3360), .B2(n4215), .A(n3297), .ZN(n3298) );
  AOI211_X1 U4100 ( .C1(n3300), .C2(n4629), .A(n3299), .B(n3298), .ZN(n3301)
         );
  OAI211_X1 U4101 ( .C1(n4634), .C2(n3359), .A(n3302), .B(n3301), .ZN(U3281)
         );
  NAND2_X1 U4102 ( .A1(n3792), .A2(n3796), .ZN(n3690) );
  XNOR2_X1 U4103 ( .A(n3303), .B(n3690), .ZN(n3310) );
  XOR2_X1 U4104 ( .A(n3690), .B(n3304), .Z(n3308) );
  AOI22_X1 U4105 ( .A1(n4334), .A2(n4596), .B1(n4609), .B2(n3351), .ZN(n3305)
         );
  OAI21_X1 U4106 ( .B1(n3306), .B2(n4592), .A(n3305), .ZN(n3307) );
  AOI21_X1 U4107 ( .B1(n3308), .B2(n4621), .A(n3307), .ZN(n3309) );
  OAI21_X1 U4108 ( .B1(n3310), .B2(n4617), .A(n3309), .ZN(n4696) );
  INV_X1 U4109 ( .A(n4696), .ZN(n3319) );
  INV_X1 U4110 ( .A(n3310), .ZN(n4698) );
  INV_X1 U4111 ( .A(n3311), .ZN(n3313) );
  NOR2_X1 U4112 ( .A1(n3313), .A2(n3312), .ZN(n4695) );
  INV_X1 U4113 ( .A(n4604), .ZN(n4694) );
  NOR3_X1 U4114 ( .A1(n4695), .A2(n4694), .A3(n4180), .ZN(n3317) );
  INV_X1 U4115 ( .A(n3314), .ZN(n3354) );
  OAI22_X1 U4116 ( .A1(n4205), .A2(n3315), .B1(n3354), .B2(n4190), .ZN(n3316)
         );
  AOI211_X1 U4117 ( .C1(n4698), .C2(n4631), .A(n3317), .B(n3316), .ZN(n3318)
         );
  OAI21_X1 U4118 ( .B1(n3319), .B2(n4634), .A(n3318), .ZN(U3280) );
  INV_X1 U4119 ( .A(n3322), .ZN(n3323) );
  OR2_X1 U4120 ( .A1(n3324), .A2(n3323), .ZN(n3325) );
  NAND2_X1 U4121 ( .A1(n3328), .A2(n3327), .ZN(n3384) );
  OAI22_X1 U4122 ( .A1(n4322), .A2(n2224), .B1(n3508), .B2(n4330), .ZN(n3329)
         );
  XNOR2_X1 U4123 ( .A(n3329), .B(n3526), .ZN(n3330) );
  OAI22_X1 U4124 ( .A1(n4322), .A2(n3538), .B1(n2224), .B2(n4330), .ZN(n3331)
         );
  AND2_X1 U4125 ( .A1(n3330), .A2(n3331), .ZN(n3383) );
  INV_X1 U4126 ( .A(n3383), .ZN(n3334) );
  INV_X1 U4127 ( .A(n3330), .ZN(n3333) );
  INV_X1 U4128 ( .A(n3331), .ZN(n3332) );
  NAND2_X1 U4129 ( .A1(n3333), .A2(n3332), .ZN(n3382) );
  NAND2_X1 U4130 ( .A1(n3334), .A2(n3382), .ZN(n3335) );
  XNOR2_X1 U4131 ( .A(n3384), .B(n3335), .ZN(n3341) );
  INV_X1 U4132 ( .A(n3336), .ZN(n3373) );
  NAND2_X1 U4133 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4519) );
  OAI21_X1 U4134 ( .B1(n4415), .B2(n3375), .A(n4519), .ZN(n3337) );
  INV_X1 U4135 ( .A(n3337), .ZN(n3339) );
  AOI22_X1 U4136 ( .A1(n4421), .A2(n3851), .B1(n3674), .B2(n3378), .ZN(n3338)
         );
  OAI211_X1 U4137 ( .C1(n4431), .C2(n3373), .A(n3339), .B(n3338), .ZN(n3340)
         );
  AOI21_X1 U4138 ( .B1(n3341), .B2(n4426), .A(n3340), .ZN(n3342) );
  INV_X1 U4139 ( .A(n3342), .ZN(U3221) );
  OR2_X1 U4140 ( .A1(n3344), .A2(n3343), .ZN(n3347) );
  NAND2_X1 U4141 ( .A1(n3347), .A2(n3345), .ZN(n3349) );
  AND2_X1 U4142 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  AOI211_X1 U4143 ( .C1(n3350), .C2(n3349), .A(n3669), .B(n3348), .ZN(n3356)
         );
  NOR2_X1 U4144 ( .A1(STATE_REG_SCAN_IN), .A2(n4820), .ZN(n4504) );
  AOI21_X1 U4145 ( .B1(n3675), .B2(n3853), .A(n4504), .ZN(n3353) );
  AOI22_X1 U4146 ( .A1(n4421), .A2(n4334), .B1(n3674), .B2(n3351), .ZN(n3352)
         );
  OAI211_X1 U4147 ( .C1(n4431), .C2(n3354), .A(n3353), .B(n3352), .ZN(n3355)
         );
  OR2_X1 U4148 ( .A1(n3356), .A2(n3355), .ZN(U3214) );
  INV_X1 U4149 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4150 ( .A1(n3852), .A2(n4596), .B1(n4609), .B2(n3357), .ZN(n3358)
         );
  OAI211_X1 U4151 ( .C1(n3360), .C2(n4592), .A(n3359), .B(n3358), .ZN(n3361)
         );
  AOI21_X1 U4152 ( .B1(n4686), .B2(n3362), .A(n3361), .ZN(n3365) );
  MUX2_X1 U4153 ( .A(n3363), .B(n3365), .S(n4708), .Z(n3364) );
  OAI21_X1 U4154 ( .B1(n3368), .B2(n4677), .A(n3364), .ZN(U3485) );
  INV_X1 U4155 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3366) );
  MUX2_X1 U4156 ( .A(n3366), .B(n3365), .S(n4729), .Z(n3367) );
  OAI21_X1 U4157 ( .B1(n4714), .B2(n3368), .A(n3367), .ZN(U3527) );
  INV_X1 U4158 ( .A(n3395), .ZN(n3369) );
  OR2_X1 U4159 ( .A1(n3369), .A2(n3800), .ZN(n3683) );
  XNOR2_X1 U4160 ( .A(n3370), .B(n3683), .ZN(n4336) );
  XNOR2_X1 U4161 ( .A(n3371), .B(n3683), .ZN(n3372) );
  NOR2_X1 U4162 ( .A1(n3372), .A2(n4598), .ZN(n4332) );
  OAI21_X1 U4163 ( .B1(n4603), .B2(n4330), .A(n3400), .ZN(n4406) );
  OAI22_X1 U4164 ( .A1(n4205), .A2(n3374), .B1(n3373), .B2(n4190), .ZN(n3377)
         );
  OAI22_X1 U4165 ( .A1(n3375), .A2(n4215), .B1(n4214), .B2(n4331), .ZN(n3376)
         );
  AOI211_X1 U4166 ( .C1(n3378), .C2(n4175), .A(n3377), .B(n3376), .ZN(n3379)
         );
  OAI21_X1 U4167 ( .B1(n4406), .B2(n4180), .A(n3379), .ZN(n3380) );
  AOI21_X1 U4168 ( .B1(n4332), .B2(n4205), .A(n3380), .ZN(n3381) );
  OAI21_X1 U4169 ( .B1(n4336), .B2(n4165), .A(n3381), .ZN(U3278) );
  OAI22_X1 U4170 ( .A1(n4331), .A2(n2224), .B1(n3508), .B2(n4323), .ZN(n3385)
         );
  XNOR2_X1 U4171 ( .A(n3385), .B(n3536), .ZN(n3414) );
  XNOR2_X1 U4172 ( .A(n3414), .B(n3412), .ZN(n3386) );
  XNOR2_X1 U4173 ( .A(n3413), .B(n3386), .ZN(n3391) );
  INV_X1 U4174 ( .A(n3387), .ZN(n3402) );
  NOR2_X1 U4175 ( .A1(STATE_REG_SCAN_IN), .A2(n2628), .ZN(n4532) );
  AOI21_X1 U4176 ( .B1(n3675), .B2(n4595), .A(n4532), .ZN(n3389) );
  AOI22_X1 U4177 ( .A1(n4421), .A2(n3850), .B1(n3674), .B2(n3406), .ZN(n3388)
         );
  OAI211_X1 U4178 ( .C1(n4431), .C2(n3402), .A(n3389), .B(n3388), .ZN(n3390)
         );
  AOI21_X1 U4179 ( .B1(n3391), .B2(n4426), .A(n3390), .ZN(n3392) );
  INV_X1 U4180 ( .A(n3392), .ZN(U3231) );
  AND2_X1 U4181 ( .A1(n3802), .A2(n3393), .ZN(n3685) );
  XOR2_X1 U4182 ( .A(n3685), .B(n3394), .Z(n4321) );
  NAND2_X1 U4183 ( .A1(n3396), .A2(n3395), .ZN(n3398) );
  INV_X1 U4184 ( .A(n3685), .ZN(n3397) );
  XNOR2_X1 U4185 ( .A(n3398), .B(n3397), .ZN(n3399) );
  NAND2_X1 U4186 ( .A1(n3400), .A2(n3406), .ZN(n3401) );
  OAI22_X1 U4187 ( .A1(n4205), .A2(n3403), .B1(n3402), .B2(n4190), .ZN(n3404)
         );
  AOI21_X1 U4188 ( .B1(n3405), .B2(n4595), .A(n3404), .ZN(n3409) );
  AOI22_X1 U4189 ( .A1(n3407), .A2(n3850), .B1(n4175), .B2(n3406), .ZN(n3408)
         );
  OAI211_X1 U4190 ( .C1(n4402), .C2(n4180), .A(n3409), .B(n3408), .ZN(n3410)
         );
  AOI21_X1 U4191 ( .B1(n4327), .B2(n4205), .A(n3410), .ZN(n3411) );
  OAI21_X1 U4192 ( .B1(n4321), .B2(n4165), .A(n3411), .ZN(U3277) );
  OAI22_X1 U4193 ( .A1(n4324), .A2(n2224), .B1(n3508), .B2(n4212), .ZN(n3415)
         );
  XNOR2_X1 U4194 ( .A(n3415), .B(n3526), .ZN(n3416) );
  OAI22_X1 U4195 ( .A1(n4324), .A2(n3538), .B1(n2224), .B2(n4212), .ZN(n3417)
         );
  INV_X1 U4196 ( .A(n3416), .ZN(n3419) );
  INV_X1 U4197 ( .A(n3417), .ZN(n3418) );
  NAND2_X1 U4198 ( .A1(n3419), .A2(n3418), .ZN(n3460) );
  NAND2_X1 U4199 ( .A1(n2460), .A2(n3460), .ZN(n3420) );
  XNOR2_X1 U4200 ( .A(n3459), .B(n3420), .ZN(n3426) );
  INV_X1 U4201 ( .A(n4210), .ZN(n3424) );
  NAND2_X1 U4202 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4538) );
  OAI21_X1 U4203 ( .B1(n3665), .B2(n4416), .A(n4538), .ZN(n3421) );
  INV_X1 U4204 ( .A(n3421), .ZN(n3423) );
  AOI22_X1 U4205 ( .A1(n3675), .A2(n3851), .B1(n3674), .B2(n4313), .ZN(n3422)
         );
  OAI211_X1 U4206 ( .C1(n4431), .C2(n3424), .A(n3423), .B(n3422), .ZN(n3425)
         );
  AOI21_X1 U4207 ( .B1(n3426), .B2(n4426), .A(n3425), .ZN(n3427) );
  INV_X1 U4208 ( .A(n3427), .ZN(U3212) );
  NAND2_X1 U4209 ( .A1(n4200), .A2(n3803), .ZN(n3429) );
  INV_X1 U4210 ( .A(n3428), .ZN(n3711) );
  XNOR2_X1 U4211 ( .A(n3429), .B(n3711), .ZN(n3430) );
  NAND2_X1 U4212 ( .A1(n3430), .A2(n4621), .ZN(n4308) );
  NAND2_X1 U4213 ( .A1(n3432), .A2(n3431), .ZN(n4198) );
  NOR2_X1 U4214 ( .A1(n4198), .A2(n4199), .ZN(n4197) );
  NOR2_X1 U4215 ( .A1(n4197), .A2(n3433), .ZN(n3434) );
  XNOR2_X1 U4216 ( .A(n3434), .B(n3711), .ZN(n4310) );
  NAND2_X1 U4217 ( .A1(n4310), .A2(n4194), .ZN(n3442) );
  OAI21_X1 U4218 ( .B1(n4207), .B2(n3437), .A(n2252), .ZN(n4394) );
  INV_X1 U4219 ( .A(n4394), .ZN(n3440) );
  INV_X1 U4220 ( .A(n4175), .ZN(n4213) );
  AOI22_X1 U4221 ( .A1(n4634), .A2(REG2_REG_15__SCAN_IN), .B1(n3435), .B2(
        n4622), .ZN(n3436) );
  OAI21_X1 U4222 ( .B1(n4213), .B2(n3437), .A(n3436), .ZN(n3439) );
  OAI22_X1 U4223 ( .A1(n4324), .A2(n4215), .B1(n4214), .B2(n4292), .ZN(n3438)
         );
  AOI211_X1 U4224 ( .C1(n3440), .C2(n4629), .A(n3439), .B(n3438), .ZN(n3441)
         );
  OAI211_X1 U4225 ( .C1(n4634), .C2(n4308), .A(n3442), .B(n3441), .ZN(U3275)
         );
  INV_X1 U4226 ( .A(n3443), .ZN(n3446) );
  INV_X1 U4227 ( .A(IR_REG_30__SCAN_IN), .ZN(n3444) );
  NAND3_X1 U4228 ( .A1(n3444), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3445) );
  INV_X1 U4229 ( .A(DATAI_31_), .ZN(n4986) );
  OAI22_X1 U4230 ( .A1(n3446), .A2(n3445), .B1(STATE_REG_SCAN_IN), .B2(n4986), 
        .ZN(U3321) );
  OAI22_X1 U4231 ( .A1(n4239), .A2(n4215), .B1(n4205), .B2(n3447), .ZN(n3454)
         );
  INV_X1 U4232 ( .A(n3448), .ZN(n3449) );
  OAI22_X1 U4233 ( .A1(n3640), .A2(n2224), .B1(n3508), .B2(n4091), .ZN(n3457)
         );
  XNOR2_X1 U4234 ( .A(n3457), .B(n3536), .ZN(n3576) );
  NOR2_X1 U4235 ( .A1(n2224), .A2(n4091), .ZN(n3458) );
  AOI21_X1 U4236 ( .B1(n4107), .B2(n2923), .A(n3458), .ZN(n3495) );
  NAND2_X1 U4237 ( .A1(n4314), .A2(n3463), .ZN(n3465) );
  NAND2_X1 U4238 ( .A1(n2922), .A2(n4305), .ZN(n3464) );
  NAND2_X1 U4239 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  XNOR2_X1 U4240 ( .A(n3466), .B(n3526), .ZN(n3472) );
  NAND2_X1 U4241 ( .A1(n2923), .A2(n4314), .ZN(n3468) );
  NAND2_X1 U4242 ( .A1(n3518), .A2(n4305), .ZN(n3467) );
  OAI22_X1 U4243 ( .A1(n4292), .A2(n2224), .B1(n3508), .B2(n4417), .ZN(n3469)
         );
  XNOR2_X1 U4244 ( .A(n3469), .B(n3526), .ZN(n3471) );
  OAI22_X1 U4245 ( .A1(n4292), .A2(n3538), .B1(n2224), .B2(n4417), .ZN(n3470)
         );
  NOR2_X1 U4246 ( .A1(n3471), .A2(n3470), .ZN(n3474) );
  AOI21_X1 U4247 ( .B1(n3471), .B2(n3470), .A(n3474), .ZN(n4425) );
  OAI22_X1 U4248 ( .A1(n4158), .A2(n3525), .B1(n3508), .B2(n4290), .ZN(n3475)
         );
  XNOR2_X1 U4249 ( .A(n3475), .B(n3526), .ZN(n3477) );
  OAI22_X1 U4250 ( .A1(n4158), .A2(n3538), .B1(n3525), .B2(n4290), .ZN(n3476)
         );
  NOR2_X1 U4251 ( .A1(n3477), .A2(n3476), .ZN(n3605) );
  OAI22_X1 U4252 ( .A1(n4291), .A2(n2224), .B1(n3508), .B2(n4151), .ZN(n3478)
         );
  XNOR2_X1 U4253 ( .A(n3478), .B(n3526), .ZN(n3480) );
  OAI22_X1 U4254 ( .A1(n4291), .A2(n3538), .B1(n2224), .B2(n4151), .ZN(n3479)
         );
  AND2_X1 U4255 ( .A1(n3480), .A2(n3479), .ZN(n3645) );
  OR2_X1 U4256 ( .A1(n3480), .A2(n3479), .ZN(n3646) );
  NAND2_X1 U4257 ( .A1(n4156), .A2(n3518), .ZN(n3482) );
  NAND2_X1 U4258 ( .A1(n2922), .A2(n4138), .ZN(n3481) );
  NAND2_X1 U4259 ( .A1(n3482), .A2(n3481), .ZN(n3483) );
  XNOR2_X1 U4260 ( .A(n3483), .B(n3526), .ZN(n3484) );
  OAI22_X1 U4261 ( .A1(n4109), .A2(n3538), .B1(n2224), .B2(n4131), .ZN(n3485)
         );
  XOR2_X1 U4262 ( .A(n3484), .B(n3485), .Z(n3568) );
  NAND2_X1 U4263 ( .A1(n3567), .A2(n3568), .ZN(n3566) );
  NAND2_X1 U4264 ( .A1(n3849), .A2(n3518), .ZN(n3490) );
  NAND2_X1 U4265 ( .A1(n2922), .A2(n4116), .ZN(n3489) );
  NAND2_X1 U4266 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  XNOR2_X1 U4267 ( .A(n3491), .B(n3536), .ZN(n3494) );
  NOR2_X1 U4268 ( .A1(n2224), .A2(n3717), .ZN(n3492) );
  AOI21_X1 U4269 ( .B1(n2923), .B2(n3849), .A(n3492), .ZN(n3493) );
  OR2_X1 U4270 ( .A1(n3494), .A2(n3493), .ZN(n3626) );
  NAND2_X1 U4271 ( .A1(n3494), .A2(n3493), .ZN(n3627) );
  INV_X1 U4272 ( .A(n3576), .ZN(n3496) );
  INV_X1 U4273 ( .A(n3495), .ZN(n3575) );
  OAI22_X1 U4274 ( .A1(n4095), .A2(n3538), .B1(n2224), .B2(n4076), .ZN(n3501)
         );
  OAI22_X1 U4275 ( .A1(n4095), .A2(n2224), .B1(n3508), .B2(n4076), .ZN(n3497)
         );
  XNOR2_X1 U4276 ( .A(n3497), .B(n3526), .ZN(n3500) );
  XOR2_X1 U4277 ( .A(n3501), .B(n3500), .Z(n3637) );
  NAND2_X1 U4278 ( .A1(n3636), .A2(n3637), .ZN(n3635) );
  OAI22_X1 U4279 ( .A1(n4074), .A2(n2224), .B1(n3508), .B2(n4057), .ZN(n3498)
         );
  XNOR2_X1 U4280 ( .A(n3498), .B(n3526), .ZN(n3505) );
  NOR2_X1 U4281 ( .A1(n2224), .A2(n4057), .ZN(n3499) );
  AOI21_X1 U4282 ( .B1(n4035), .B2(n2923), .A(n3499), .ZN(n3506) );
  XNOR2_X1 U4283 ( .A(n3505), .B(n3506), .ZN(n3559) );
  INV_X1 U4284 ( .A(n3500), .ZN(n3503) );
  INV_X1 U4285 ( .A(n3501), .ZN(n3502) );
  NAND2_X1 U4286 ( .A1(n3503), .A2(n3502), .ZN(n3557) );
  NOR2_X1 U4287 ( .A1(n2224), .A2(n4038), .ZN(n3504) );
  AOI21_X1 U4288 ( .B1(n4015), .B2(n2923), .A(n3504), .ZN(n3510) );
  INV_X1 U4289 ( .A(n3505), .ZN(n3507) );
  OR2_X1 U4290 ( .A1(n3507), .A2(n3506), .ZN(n3511) );
  OAI22_X1 U4291 ( .A1(n4056), .A2(n2224), .B1(n3508), .B2(n4038), .ZN(n3509)
         );
  XNOR2_X1 U4292 ( .A(n3509), .B(n3526), .ZN(n3614) );
  NAND2_X1 U4293 ( .A1(n3847), .A2(n3518), .ZN(n3513) );
  INV_X1 U4294 ( .A(n4020), .ZN(n4014) );
  NAND2_X1 U4295 ( .A1(n2922), .A2(n4014), .ZN(n3512) );
  NAND2_X1 U4296 ( .A1(n3513), .A2(n3512), .ZN(n3514) );
  XNOR2_X1 U4297 ( .A(n3514), .B(n3536), .ZN(n3517) );
  NOR2_X1 U4298 ( .A1(n2224), .A2(n4020), .ZN(n3515) );
  AOI21_X1 U4299 ( .B1(n3847), .B2(n2923), .A(n3515), .ZN(n3516) );
  AND2_X1 U4300 ( .A1(n3517), .A2(n3516), .ZN(n3587) );
  NAND2_X1 U4301 ( .A1(n4236), .A2(n3518), .ZN(n3520) );
  NAND2_X1 U4302 ( .A1(n2922), .A2(n4244), .ZN(n3519) );
  NAND2_X1 U4303 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  XNOR2_X1 U4304 ( .A(n3521), .B(n3536), .ZN(n3524) );
  NOR2_X1 U4305 ( .A1(n2224), .A2(n4001), .ZN(n3522) );
  AOI21_X1 U4306 ( .B1(n4236), .B2(n2923), .A(n3522), .ZN(n3523) );
  NOR2_X1 U4307 ( .A1(n3524), .A2(n3523), .ZN(n3659) );
  NAND2_X1 U4308 ( .A1(n3524), .A2(n3523), .ZN(n3657) );
  OAI22_X1 U4309 ( .A1(n4002), .A2(n3538), .B1(n3985), .B2(n2224), .ZN(n3545)
         );
  OAI22_X1 U4310 ( .A1(n4002), .A2(n3525), .B1(n3985), .B2(n3508), .ZN(n3527)
         );
  XNOR2_X1 U4311 ( .A(n3527), .B(n3526), .ZN(n3546) );
  XNOR2_X1 U4312 ( .A(n3542), .B(n3543), .ZN(n3528) );
  NAND2_X1 U4313 ( .A1(n3528), .A2(n4426), .ZN(n3535) );
  INV_X1 U4314 ( .A(n3983), .ZN(n3529) );
  NOR2_X1 U4315 ( .A1(n4431), .A2(n3529), .ZN(n3533) );
  AOI22_X1 U4316 ( .A1(n3675), .A2(n4236), .B1(n3674), .B2(n4235), .ZN(n3531)
         );
  NAND2_X1 U4317 ( .A1(U3149), .A2(REG3_REG_27__SCAN_IN), .ZN(n3530) );
  OAI211_X1 U4318 ( .C1(n4239), .C2(n3665), .A(n3531), .B(n3530), .ZN(n3532)
         );
  NOR2_X1 U4319 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  NAND2_X1 U4320 ( .A1(n3535), .A2(n3534), .ZN(U3211) );
  OAI22_X1 U4321 ( .A1(n4239), .A2(n2224), .B1(n3508), .B2(n3969), .ZN(n3537)
         );
  XNOR2_X1 U4322 ( .A(n3537), .B(n3536), .ZN(n3540) );
  OAI22_X1 U4323 ( .A1(n4239), .A2(n3538), .B1(n2224), .B2(n3969), .ZN(n3539)
         );
  XNOR2_X1 U4324 ( .A(n3540), .B(n3539), .ZN(n3550) );
  INV_X1 U4325 ( .A(n3550), .ZN(n3541) );
  NAND2_X1 U4326 ( .A1(n3541), .A2(n4426), .ZN(n3556) );
  INV_X1 U4327 ( .A(n3542), .ZN(n3544) );
  NAND2_X1 U4328 ( .A1(n3544), .A2(n3543), .ZN(n3555) );
  NAND2_X1 U4329 ( .A1(n3546), .A2(n3545), .ZN(n3549) );
  NAND2_X1 U4330 ( .A1(n3555), .A2(n2456), .ZN(n3554) );
  INV_X1 U4331 ( .A(n4431), .ZN(n3667) );
  AOI22_X1 U4332 ( .A1(n4245), .A2(n3675), .B1(n3962), .B2(n3674), .ZN(n3548)
         );
  AOI22_X1 U4333 ( .A1(n3963), .A2(n4421), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3547) );
  NAND2_X1 U4334 ( .A1(n3548), .A2(n3547), .ZN(n3552) );
  NOR3_X1 U4335 ( .A1(n3550), .A2(n3669), .A3(n3549), .ZN(n3551) );
  AOI211_X1 U4336 ( .C1(n3970), .C2(n3667), .A(n3552), .B(n3551), .ZN(n3553)
         );
  OAI211_X1 U4337 ( .C1(n3556), .C2(n3555), .A(n3554), .B(n3553), .ZN(U3217)
         );
  AND2_X1 U4338 ( .A1(n3635), .A2(n3557), .ZN(n3560) );
  OAI211_X1 U4339 ( .C1(n3560), .C2(n3559), .A(n4426), .B(n3558), .ZN(n3565)
         );
  NAND2_X1 U4340 ( .A1(n3674), .A2(n4053), .ZN(n3561) );
  OAI21_X1 U4341 ( .B1(n4056), .B2(n3665), .A(n3561), .ZN(n3563) );
  OAI22_X1 U4342 ( .A1(n4415), .A2(n4095), .B1(STATE_REG_SCAN_IN), .B2(n4816), 
        .ZN(n3562) );
  NOR2_X1 U4343 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  OAI211_X1 U4344 ( .C1(n4431), .C2(n4060), .A(n3565), .B(n3564), .ZN(U3213)
         );
  OAI21_X1 U4345 ( .B1(n3568), .B2(n3567), .A(n3566), .ZN(n3573) );
  AND2_X1 U4346 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3947) );
  AOI21_X1 U4347 ( .B1(n3675), .B2(n4133), .A(n3947), .ZN(n3570) );
  AOI22_X1 U4348 ( .A1(n4421), .A2(n3849), .B1(n3674), .B2(n4138), .ZN(n3569)
         );
  OAI211_X1 U4349 ( .C1(n4431), .C2(n3571), .A(n3570), .B(n3569), .ZN(n3572)
         );
  AOI21_X1 U4350 ( .B1(n3573), .B2(n4426), .A(n3572), .ZN(n3574) );
  INV_X1 U4351 ( .A(n3574), .ZN(U3216) );
  XNOR2_X1 U4352 ( .A(n3576), .B(n3575), .ZN(n3577) );
  XNOR2_X1 U4353 ( .A(n3578), .B(n3577), .ZN(n3585) );
  INV_X1 U4354 ( .A(n3579), .ZN(n4093) );
  OAI22_X1 U4355 ( .A1(n4415), .A2(n4272), .B1(STATE_REG_SCAN_IN), .B2(n3580), 
        .ZN(n3581) );
  INV_X1 U4356 ( .A(n3581), .ZN(n3583) );
  AOI22_X1 U4357 ( .A1(n4421), .A2(n4270), .B1(n3674), .B2(n4269), .ZN(n3582)
         );
  OAI211_X1 U4358 ( .C1(n4431), .C2(n4093), .A(n3583), .B(n3582), .ZN(n3584)
         );
  AOI21_X1 U4359 ( .B1(n3585), .B2(n4426), .A(n3584), .ZN(n3586) );
  INV_X1 U4360 ( .A(n3586), .ZN(U3220) );
  NOR2_X1 U4361 ( .A1(n2257), .A2(n3587), .ZN(n3588) );
  XNOR2_X1 U4362 ( .A(n2238), .B(n3588), .ZN(n3593) );
  INV_X1 U4363 ( .A(n4021), .ZN(n3591) );
  AOI22_X1 U4364 ( .A1(n3675), .A2(n4015), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3590) );
  AOI22_X1 U4365 ( .A1(n4421), .A2(n4236), .B1(n3674), .B2(n4014), .ZN(n3589)
         );
  OAI211_X1 U4366 ( .C1(n4431), .C2(n3591), .A(n3590), .B(n3589), .ZN(n3592)
         );
  AOI21_X1 U4367 ( .B1(n3593), .B2(n4426), .A(n3592), .ZN(n3594) );
  INV_X1 U4368 ( .A(n3594), .ZN(U3222) );
  OAI211_X1 U4369 ( .C1(n3595), .C2(n3597), .A(n3596), .B(n4426), .ZN(n3603)
         );
  AND2_X1 U4370 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4445) );
  AOI21_X1 U4371 ( .B1(n3675), .B2(n3859), .A(n4445), .ZN(n3602) );
  AOI22_X1 U4372 ( .A1(n4421), .A2(n3857), .B1(n3674), .B2(n3598), .ZN(n3601)
         );
  OR2_X1 U4373 ( .A1(n4431), .A2(n3599), .ZN(n3600) );
  NAND4_X1 U4374 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(U3224)
         );
  NOR2_X1 U4375 ( .A1(n3605), .A2(n2264), .ZN(n3606) );
  XNOR2_X1 U4376 ( .A(n3604), .B(n3606), .ZN(n3611) );
  INV_X1 U4377 ( .A(n3607), .ZN(n4172) );
  AND2_X1 U4378 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4568) );
  AOI21_X1 U4379 ( .B1(n3675), .B2(n4306), .A(n4568), .ZN(n3609) );
  AOI22_X1 U4380 ( .A1(n4421), .A2(n4133), .B1(n3674), .B2(n4176), .ZN(n3608)
         );
  OAI211_X1 U4381 ( .C1(n4431), .C2(n4172), .A(n3609), .B(n3608), .ZN(n3610)
         );
  AOI21_X1 U4382 ( .B1(n3611), .B2(n4426), .A(n3610), .ZN(n3612) );
  INV_X1 U4383 ( .A(n3612), .ZN(U3225) );
  NAND2_X1 U4384 ( .A1(n2245), .A2(n3613), .ZN(n3615) );
  XNOR2_X1 U4385 ( .A(n3615), .B(n3614), .ZN(n3620) );
  INV_X1 U4386 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4808) );
  OAI22_X1 U4387 ( .A1(n4415), .A2(n4074), .B1(STATE_REG_SCAN_IN), .B2(n4808), 
        .ZN(n3616) );
  INV_X1 U4388 ( .A(n3616), .ZN(n3618) );
  AOI22_X1 U4389 ( .A1(n4421), .A2(n3847), .B1(n3674), .B2(n4034), .ZN(n3617)
         );
  OAI211_X1 U4390 ( .C1(n4431), .C2(n4041), .A(n3618), .B(n3617), .ZN(n3619)
         );
  AOI21_X1 U4391 ( .B1(n3620), .B2(n4426), .A(n3619), .ZN(n3621) );
  INV_X1 U4392 ( .A(n3621), .ZN(U3226) );
  INV_X1 U4393 ( .A(n3622), .ZN(n4117) );
  INV_X1 U4394 ( .A(n3627), .ZN(n3623) );
  NOR2_X1 U4395 ( .A1(n3624), .A2(n3623), .ZN(n3629) );
  AOI21_X1 U4396 ( .B1(n3627), .B2(n3626), .A(n3625), .ZN(n3628) );
  OAI21_X1 U4397 ( .B1(n3629), .B2(n3628), .A(n4426), .ZN(n3634) );
  NAND2_X1 U4398 ( .A1(n3674), .A2(n4116), .ZN(n3630) );
  OAI21_X1 U4399 ( .B1(n3640), .B2(n3665), .A(n3630), .ZN(n3632) );
  INV_X1 U4400 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4983) );
  OAI22_X1 U4401 ( .A1(n4415), .A2(n4109), .B1(STATE_REG_SCAN_IN), .B2(n4983), 
        .ZN(n3631) );
  NOR2_X1 U4402 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  OAI211_X1 U4403 ( .C1(n4431), .C2(n4117), .A(n3634), .B(n3633), .ZN(U3230)
         );
  OAI21_X1 U4404 ( .B1(n3637), .B2(n3636), .A(n3635), .ZN(n3638) );
  NAND2_X1 U4405 ( .A1(n3638), .A2(n4426), .ZN(n3644) );
  OAI22_X1 U4406 ( .A1(n3665), .A2(n4074), .B1(STATE_REG_SCAN_IN), .B2(n3639), 
        .ZN(n3642) );
  OAI22_X1 U4407 ( .A1(n4418), .A2(n4076), .B1(n3640), .B2(n4415), .ZN(n3641)
         );
  AOI211_X1 U4408 ( .C1(n3667), .C2(n4078), .A(n3642), .B(n3641), .ZN(n3643)
         );
  NAND2_X1 U4409 ( .A1(n3644), .A2(n3643), .ZN(U3232) );
  INV_X1 U4410 ( .A(n3645), .ZN(n3647) );
  NAND2_X1 U4411 ( .A1(n3647), .A2(n3646), .ZN(n3648) );
  XNOR2_X1 U4412 ( .A(n3649), .B(n3648), .ZN(n3655) );
  INV_X1 U4413 ( .A(n4149), .ZN(n3653) );
  NAND2_X1 U4414 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4573) );
  OAI21_X1 U4415 ( .B1(n3665), .B2(n4109), .A(n4573), .ZN(n3650) );
  INV_X1 U4416 ( .A(n3650), .ZN(n3652) );
  AOI22_X1 U4417 ( .A1(n3675), .A2(n4420), .B1(n3674), .B2(n4155), .ZN(n3651)
         );
  OAI211_X1 U4418 ( .C1(n4431), .C2(n3653), .A(n3652), .B(n3651), .ZN(n3654)
         );
  AOI21_X1 U4419 ( .B1(n3655), .B2(n4426), .A(n3654), .ZN(n3656) );
  INV_X1 U4420 ( .A(n3656), .ZN(U3235) );
  INV_X1 U4421 ( .A(n3657), .ZN(n3658) );
  NOR2_X1 U4422 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  XNOR2_X1 U4423 ( .A(n3661), .B(n3660), .ZN(n3670) );
  INV_X1 U4424 ( .A(n3662), .ZN(n3999) );
  AOI22_X1 U4425 ( .A1(n3675), .A2(n3847), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3664) );
  NAND2_X1 U4426 ( .A1(n3674), .A2(n4244), .ZN(n3663) );
  OAI211_X1 U4427 ( .C1(n4002), .C2(n3665), .A(n3664), .B(n3663), .ZN(n3666)
         );
  AOI21_X1 U4428 ( .B1(n3667), .B2(n3999), .A(n3666), .ZN(n3668) );
  OAI21_X1 U4429 ( .B1(n3670), .B2(n3669), .A(n3668), .ZN(U3237) );
  INV_X1 U4430 ( .A(n4422), .ZN(n3672) );
  NOR2_X1 U4431 ( .A1(n3671), .A2(n3672), .ZN(n3673) );
  XNOR2_X1 U4432 ( .A(n3673), .B(n4423), .ZN(n3680) );
  AND2_X1 U4433 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4550) );
  AOI21_X1 U4434 ( .B1(n4421), .B2(n4306), .A(n4550), .ZN(n3677) );
  AOI22_X1 U4435 ( .A1(n3675), .A2(n3850), .B1(n3674), .B2(n4305), .ZN(n3676)
         );
  OAI211_X1 U4436 ( .C1(n4431), .C2(n3678), .A(n3677), .B(n3676), .ZN(n3679)
         );
  AOI21_X1 U4437 ( .B1(n3680), .B2(n4426), .A(n3679), .ZN(n3681) );
  INV_X1 U4438 ( .A(n3681), .ZN(U3238) );
  NAND2_X1 U4439 ( .A1(n3682), .A2(n4009), .ZN(n4032) );
  AND2_X1 U4440 ( .A1(n4124), .A2(n4125), .ZN(n4168) );
  INV_X1 U4441 ( .A(n3683), .ZN(n3686) );
  NAND4_X1 U4442 ( .A1(n4168), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3692)
         );
  INV_X1 U4443 ( .A(n3687), .ZN(n3689) );
  OR2_X1 U4444 ( .A1(n3689), .A2(n3688), .ZN(n4137) );
  INV_X1 U4445 ( .A(n4137), .ZN(n3691) );
  NOR4_X1 U4446 ( .A1(n4032), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3701)
         );
  NOR4_X1 U4447 ( .A1(n2692), .A2(n3694), .A3(n4588), .A4(n3693), .ZN(n3700)
         );
  INV_X1 U4448 ( .A(n4068), .ZN(n3698) );
  NOR4_X1 U4449 ( .A1(n3698), .A2(n2669), .A3(n3697), .A4(n3696), .ZN(n3699)
         );
  NAND3_X1 U4450 ( .A1(n3701), .A2(n3700), .A3(n3699), .ZN(n3715) );
  NAND2_X1 U4451 ( .A1(n3814), .A2(n4048), .ZN(n4086) );
  INV_X1 U4452 ( .A(n4086), .ZN(n3712) );
  AND2_X1 U4453 ( .A1(n3702), .A2(DATAI_30_), .ZN(n4228) );
  INV_X1 U4454 ( .A(n4228), .ZN(n3757) );
  NAND2_X1 U4455 ( .A1(n3845), .A2(n3757), .ZN(n3734) );
  INV_X1 U4456 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4457 ( .A1(n3703), .A2(REG1_REG_31__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U4458 ( .A1(n2544), .A2(REG0_REG_31__SCAN_IN), .ZN(n3704) );
  OAI211_X1 U4459 ( .C1(n3707), .C2(n3706), .A(n3705), .B(n3704), .ZN(n3955)
         );
  NAND2_X1 U4460 ( .A1(n3702), .A2(DATAI_31_), .ZN(n3956) );
  OR2_X1 U4461 ( .A1(n3955), .A2(n3956), .ZN(n3708) );
  NAND2_X1 U4462 ( .A1(n3734), .A2(n3708), .ZN(n3834) );
  NAND2_X1 U4463 ( .A1(n3955), .A2(n3956), .ZN(n3833) );
  OR2_X1 U4464 ( .A1(n3845), .A2(n3757), .ZN(n3709) );
  NAND2_X1 U4465 ( .A1(n3833), .A2(n3709), .ZN(n3730) );
  NOR2_X1 U4466 ( .A1(n3834), .A2(n3730), .ZN(n3710) );
  NAND4_X1 U4467 ( .A1(n3712), .A2(n3711), .A3(n4665), .A4(n3710), .ZN(n3713)
         );
  NOR3_X1 U4468 ( .A1(n3715), .A2(n3714), .A3(n3713), .ZN(n3722) );
  INV_X1 U4469 ( .A(n3829), .ZN(n3729) );
  NAND2_X1 U4470 ( .A1(n3729), .A2(n3716), .ZN(n3996) );
  XNOR2_X1 U4471 ( .A(n4035), .B(n4057), .ZN(n4050) );
  XNOR2_X1 U4472 ( .A(n3849), .B(n3717), .ZN(n4111) );
  NAND4_X1 U4473 ( .A1(n2307), .A2(n4199), .A3(n3719), .A4(n3718), .ZN(n3720)
         );
  NOR4_X1 U4474 ( .A1(n3996), .A2(n4050), .A3(n4111), .A4(n3720), .ZN(n3721)
         );
  NAND3_X1 U4475 ( .A1(n3722), .A2(n3979), .A3(n3721), .ZN(n3726) );
  INV_X1 U4476 ( .A(n3960), .ZN(n3725) );
  NAND2_X1 U4477 ( .A1(n3991), .A2(n3723), .ZN(n4011) );
  NOR4_X1 U4478 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n4011), .ZN(n3761)
         );
  INV_X1 U4480 ( .A(n3956), .ZN(n3758) );
  AND2_X1 U4481 ( .A1(n3963), .A2(n3732), .ZN(n3727) );
  NOR2_X1 U4482 ( .A1(n3728), .A2(n3727), .ZN(n3825) );
  NAND3_X1 U4483 ( .A1(n3825), .A2(n3979), .A3(n3729), .ZN(n3733) );
  INV_X1 U4484 ( .A(n3730), .ZN(n3731) );
  OAI21_X1 U4485 ( .B1(n3963), .B2(n3732), .A(n3731), .ZN(n3746) );
  AOI221_X1 U4486 ( .B1(n3825), .B2(n3748), .C1(n3825), .C2(n3747), .A(n3746), 
        .ZN(n3830) );
  AND2_X1 U4487 ( .A1(n3733), .A2(n3830), .ZN(n3756) );
  AOI21_X1 U4488 ( .B1(n3734), .B2(n3955), .A(n3956), .ZN(n3755) );
  INV_X1 U4489 ( .A(n3824), .ZN(n3752) );
  NAND2_X1 U4490 ( .A1(n3736), .A2(n3735), .ZN(n3790) );
  NAND2_X1 U4491 ( .A1(n3790), .A2(n3801), .ZN(n3793) );
  INV_X1 U4492 ( .A(n3737), .ZN(n4203) );
  NAND3_X1 U4493 ( .A1(n4203), .A2(n3803), .A3(n3801), .ZN(n3738) );
  NAND2_X1 U4494 ( .A1(n3793), .A2(n3738), .ZN(n3740) );
  INV_X1 U4495 ( .A(n3809), .ZN(n3739) );
  AOI211_X1 U4496 ( .C1(n3812), .C2(n3740), .A(n3739), .B(n3811), .ZN(n3741)
         );
  OAI21_X1 U4497 ( .B1(n3741), .B2(n3816), .A(n3815), .ZN(n3742) );
  NAND2_X1 U4498 ( .A1(n3820), .A2(n3742), .ZN(n3744) );
  INV_X1 U4499 ( .A(n3818), .ZN(n3743) );
  AOI21_X1 U4500 ( .B1(n3745), .B2(n3744), .A(n3743), .ZN(n3751) );
  NOR3_X1 U4501 ( .A1(n3748), .A2(n3747), .A3(n3746), .ZN(n3749) );
  OAI211_X1 U4502 ( .C1(n3752), .C2(n3751), .A(n3750), .B(n3749), .ZN(n3753)
         );
  INV_X1 U4503 ( .A(n3753), .ZN(n3754) );
  OAI33_X1 U4504 ( .A1(1'b0), .A2(n3758), .A3(n3757), .B1(n3756), .B2(n3755), 
        .B3(n3754), .ZN(n3760) );
  MUX2_X1 U4505 ( .A(n3761), .B(n3760), .S(n3765), .Z(n3837) );
  NOR2_X1 U4506 ( .A1(n4002), .A2(n4235), .ZN(n3828) );
  OAI211_X1 U4507 ( .C1(n2306), .C2(n3765), .A(n3764), .B(n3763), .ZN(n3768)
         );
  NAND3_X1 U4508 ( .A1(n3768), .A2(n3767), .A3(n3766), .ZN(n3770) );
  OAI211_X1 U4509 ( .C1(n3772), .C2(n3771), .A(n3770), .B(n3769), .ZN(n3775)
         );
  NAND3_X1 U4510 ( .A1(n3775), .A2(n3774), .A3(n3773), .ZN(n3777) );
  NAND4_X1 U4511 ( .A1(n3777), .A2(n3776), .A3(n2253), .A4(n3786), .ZN(n3780)
         );
  NAND3_X1 U4512 ( .A1(n3780), .A2(n3779), .A3(n3778), .ZN(n3781) );
  NAND3_X1 U4513 ( .A1(n3781), .A2(n3788), .A3(n3787), .ZN(n3784) );
  AND3_X1 U4514 ( .A1(n3784), .A2(n3783), .A3(n3782), .ZN(n3791) );
  INV_X1 U4515 ( .A(n3793), .ZN(n3806) );
  NAND4_X1 U4516 ( .A1(n2330), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3789)
         );
  OAI22_X1 U4517 ( .A1(n3791), .A2(n3790), .B1(n3806), .B2(n3789), .ZN(n3795)
         );
  INV_X1 U4518 ( .A(n3792), .ZN(n3794) );
  AOI22_X1 U4519 ( .A1(n3795), .A2(n2263), .B1(n3794), .B2(n3793), .ZN(n3808)
         );
  NAND3_X1 U4520 ( .A1(n3799), .A2(n3797), .A3(n3796), .ZN(n3807) );
  OAI21_X1 U4521 ( .B1(n2310), .B2(n3800), .A(n3799), .ZN(n3804) );
  AND4_X1 U4522 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  OAI22_X1 U4523 ( .A1(n3808), .A2(n3807), .B1(n3806), .B2(n3805), .ZN(n3810)
         );
  NAND2_X1 U4524 ( .A1(n3810), .A2(n3809), .ZN(n3813) );
  AOI21_X1 U4525 ( .B1(n3813), .B2(n3812), .A(n3811), .ZN(n3817) );
  OAI211_X1 U4526 ( .C1(n3817), .C2(n3816), .A(n3815), .B(n3814), .ZN(n3819)
         );
  OAI221_X1 U4527 ( .B1(n3821), .B2(n3820), .C1(n3821), .C2(n3819), .A(n3818), 
        .ZN(n3823) );
  AOI21_X1 U4528 ( .B1(n3824), .B2(n3823), .A(n3822), .ZN(n3827) );
  INV_X1 U4529 ( .A(n3825), .ZN(n3826) );
  NOR4_X1 U4530 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3832)
         );
  INV_X1 U4531 ( .A(n3830), .ZN(n3831) );
  NOR2_X1 U4532 ( .A1(n3832), .A2(n3831), .ZN(n3835) );
  OAI21_X1 U4533 ( .B1(n3835), .B2(n3834), .A(n3833), .ZN(n3836) );
  MUX2_X1 U4534 ( .A(n3837), .B(n3836), .S(n2788), .Z(n3838) );
  XNOR2_X1 U4535 ( .A(n3838), .B(n4161), .ZN(n3844) );
  NAND2_X1 U4536 ( .A1(n3840), .A2(n3839), .ZN(n3841) );
  OAI211_X1 U4537 ( .C1(n4409), .C2(n3843), .A(n3841), .B(B_REG_SCAN_IN), .ZN(
        n3842) );
  OAI21_X1 U4538 ( .B1(n3844), .B2(n3843), .A(n3842), .ZN(U3239) );
  MUX2_X1 U4539 ( .A(DATAO_REG_31__SCAN_IN), .B(n3955), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4540 ( .A(DATAO_REG_30__SCAN_IN), .B(n3845), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4541 ( .A(DATAO_REG_29__SCAN_IN), .B(n3963), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4542 ( .A(DATAO_REG_28__SCAN_IN), .B(n3846), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4543 ( .A(DATAO_REG_27__SCAN_IN), .B(n4245), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4544 ( .A(DATAO_REG_26__SCAN_IN), .B(n4236), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4545 ( .A(DATAO_REG_25__SCAN_IN), .B(n3847), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4546 ( .A(DATAO_REG_24__SCAN_IN), .B(n4015), .S(n3856), .Z(U3574)
         );
  MUX2_X1 U4547 ( .A(DATAO_REG_23__SCAN_IN), .B(n4035), .S(n3856), .Z(U3573)
         );
  MUX2_X1 U4548 ( .A(DATAO_REG_22__SCAN_IN), .B(n4270), .S(n3856), .Z(U3572)
         );
  MUX2_X1 U4549 ( .A(DATAO_REG_21__SCAN_IN), .B(n4107), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4550 ( .A(DATAO_REG_20__SCAN_IN), .B(n3849), .S(n3856), .Z(U3570)
         );
  MUX2_X1 U4551 ( .A(DATAO_REG_19__SCAN_IN), .B(n4156), .S(n3856), .Z(U3569)
         );
  MUX2_X1 U4552 ( .A(DATAO_REG_18__SCAN_IN), .B(n4133), .S(n3856), .Z(U3568)
         );
  MUX2_X1 U4553 ( .A(DATAO_REG_17__SCAN_IN), .B(n4420), .S(n3856), .Z(U3567)
         );
  MUX2_X1 U4554 ( .A(DATAO_REG_16__SCAN_IN), .B(n4306), .S(n3856), .Z(U3566)
         );
  MUX2_X1 U4555 ( .A(DATAO_REG_15__SCAN_IN), .B(n4314), .S(n3856), .Z(U3565)
         );
  MUX2_X1 U4556 ( .A(DATAO_REG_14__SCAN_IN), .B(n3850), .S(n3856), .Z(U3564)
         );
  MUX2_X1 U4557 ( .A(DATAO_REG_13__SCAN_IN), .B(n3851), .S(n3856), .Z(U3563)
         );
  MUX2_X1 U4558 ( .A(DATAO_REG_12__SCAN_IN), .B(n4595), .S(n3856), .Z(U3562)
         );
  MUX2_X1 U4559 ( .A(DATAO_REG_11__SCAN_IN), .B(n4334), .S(n3856), .Z(U3561)
         );
  MUX2_X1 U4560 ( .A(DATAO_REG_10__SCAN_IN), .B(n3852), .S(n3856), .Z(U3560)
         );
  MUX2_X1 U4561 ( .A(DATAO_REG_9__SCAN_IN), .B(n3853), .S(n3856), .Z(U3559) );
  MUX2_X1 U4562 ( .A(DATAO_REG_8__SCAN_IN), .B(n3854), .S(n3856), .Z(U3558) );
  MUX2_X1 U4563 ( .A(DATAO_REG_7__SCAN_IN), .B(n3855), .S(n3856), .Z(U3557) );
  MUX2_X1 U4564 ( .A(DATAO_REG_6__SCAN_IN), .B(n3857), .S(n3856), .Z(U3556) );
  MUX2_X1 U4565 ( .A(DATAO_REG_5__SCAN_IN), .B(n3858), .S(U4043), .Z(U3555) );
  MUX2_X1 U4566 ( .A(DATAO_REG_4__SCAN_IN), .B(n3859), .S(U4043), .Z(U3554) );
  MUX2_X1 U4567 ( .A(DATAO_REG_3__SCAN_IN), .B(n2982), .S(U4043), .Z(U3553) );
  MUX2_X1 U4568 ( .A(DATAO_REG_2__SCAN_IN), .B(n2506), .S(U4043), .Z(U3552) );
  MUX2_X1 U4569 ( .A(DATAO_REG_1__SCAN_IN), .B(n2974), .S(U4043), .Z(U3551) );
  MUX2_X1 U4570 ( .A(DATAO_REG_0__SCAN_IN), .B(n4611), .S(U4043), .Z(U3550) );
  INV_X1 U4571 ( .A(n4586), .ZN(n3860) );
  NAND2_X1 U4572 ( .A1(n3860), .A2(n4413), .ZN(n3869) );
  OAI211_X1 U4573 ( .C1(n3863), .C2(n3862), .A(n4580), .B(n3861), .ZN(n3868)
         );
  OAI211_X1 U4574 ( .C1(n3865), .C2(n3864), .A(n4527), .B(n3876), .ZN(n3867)
         );
  AOI22_X1 U4575 ( .A1(n4578), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3866) );
  NAND4_X1 U4576 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(U3241)
         );
  INV_X1 U4577 ( .A(n4412), .ZN(n3871) );
  AOI22_X1 U4578 ( .A1(n4578), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3870) );
  OAI21_X1 U4579 ( .B1(n4586), .B2(n3871), .A(n3870), .ZN(n3872) );
  INV_X1 U4580 ( .A(n3872), .ZN(n3884) );
  INV_X1 U4581 ( .A(n3873), .ZN(n3878) );
  NAND3_X1 U4582 ( .A1(n3876), .A2(n3875), .A3(n3874), .ZN(n3877) );
  NAND3_X1 U4583 ( .A1(n4527), .A2(n3878), .A3(n3877), .ZN(n3883) );
  OAI211_X1 U4584 ( .C1(n3881), .C2(n3880), .A(n4580), .B(n3879), .ZN(n3882)
         );
  NAND4_X1 U4585 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(U3242)
         );
  MUX2_X1 U4586 ( .A(n2695), .B(REG2_REG_19__SCAN_IN), .S(n3949), .Z(n3911) );
  INV_X1 U4587 ( .A(n4645), .ZN(n4585) );
  AOI22_X1 U4588 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4585), .B1(n4645), .B2(
        n2684), .ZN(n4576) );
  NOR2_X1 U4589 ( .A1(n3941), .A2(REG2_REG_17__SCAN_IN), .ZN(n3886) );
  AOI21_X1 U4590 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3941), .A(n3886), .ZN(n4566) );
  INV_X1 U4591 ( .A(n3933), .ZN(n4652) );
  NOR2_X1 U4592 ( .A1(n3403), .A2(n4653), .ZN(n4526) );
  NAND2_X1 U4593 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3916), .ZN(n3902) );
  INV_X1 U4594 ( .A(n3916), .ZN(n4655) );
  AOI22_X1 U4595 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3916), .B1(n4655), .B2(
        n2610), .ZN(n4511) );
  NAND2_X1 U4596 ( .A1(n3917), .A2(REG2_REG_9__SCAN_IN), .ZN(n3899) );
  INV_X1 U4597 ( .A(n3917), .ZN(n4657) );
  AOI22_X1 U4598 ( .A1(n3917), .A2(REG2_REG_9__SCAN_IN), .B1(n3887), .B2(n4657), .ZN(n4490) );
  NAND2_X1 U4599 ( .A1(n3923), .A2(REG2_REG_7__SCAN_IN), .ZN(n3896) );
  INV_X1 U4600 ( .A(n3923), .ZN(n4659) );
  AOI22_X1 U4601 ( .A1(n3923), .A2(REG2_REG_7__SCAN_IN), .B1(n2568), .B2(n4659), .ZN(n4472) );
  NAND2_X1 U4602 ( .A1(n3920), .A2(REG2_REG_5__SCAN_IN), .ZN(n3892) );
  INV_X1 U4603 ( .A(n3920), .ZN(n4662) );
  AOI22_X1 U4604 ( .A1(n3920), .A2(REG2_REG_5__SCAN_IN), .B1(n2538), .B2(n4662), .ZN(n4449) );
  INV_X1 U4605 ( .A(n3888), .ZN(n3889) );
  NAND2_X1 U4606 ( .A1(n3893), .A2(n3894), .ZN(n3895) );
  NAND2_X1 U4607 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4459), .ZN(n4458) );
  NAND2_X1 U4608 ( .A1(n4475), .A2(n3897), .ZN(n3898) );
  NAND2_X1 U4609 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U4610 ( .A1(n4496), .A2(n3900), .ZN(n3901) );
  NAND2_X1 U4611 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4500), .ZN(n4499) );
  NAND2_X1 U4612 ( .A1(n3901), .A2(n4499), .ZN(n4510) );
  NAND2_X1 U4613 ( .A1(n4511), .A2(n4510), .ZN(n4509) );
  NAND2_X1 U4614 ( .A1(n3929), .A2(n3903), .ZN(n3904) );
  OAI22_X1 U4615 ( .A1(n4526), .A2(n4529), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3915), .ZN(n3905) );
  NOR2_X1 U4616 ( .A1(n4652), .A2(n3905), .ZN(n3906) );
  NAND2_X1 U4617 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3913), .ZN(n3907) );
  OAI21_X1 U4618 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3913), .A(n3907), .ZN(n4548) );
  AOI21_X1 U4619 ( .B1(n3913), .B2(REG2_REG_15__SCAN_IN), .A(n4547), .ZN(n3908) );
  INV_X1 U4620 ( .A(n3937), .ZN(n4649) );
  NAND2_X1 U4621 ( .A1(n3908), .A2(n4649), .ZN(n3909) );
  XOR2_X1 U4622 ( .A(n3908), .B(n4649), .Z(n4557) );
  NAND2_X1 U4623 ( .A1(n4557), .A2(n4191), .ZN(n4556) );
  NAND2_X1 U4624 ( .A1(n3909), .A2(n4556), .ZN(n4564) );
  NAND2_X1 U4625 ( .A1(n4566), .A2(n4564), .ZN(n4565) );
  AOI21_X1 U4626 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4645), .A(n4575), .ZN(n3910) );
  XOR2_X1 U4627 ( .A(n3911), .B(n3910), .Z(n3953) );
  INV_X1 U4628 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4629 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4645), .B1(n4585), .B2(
        n3943), .ZN(n4582) );
  NOR2_X1 U4630 ( .A1(n3941), .A2(REG1_REG_17__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4631 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3913), .ZN(n3936) );
  INV_X1 U4632 ( .A(n3913), .ZN(n4650) );
  INV_X1 U4633 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4634 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3913), .B1(n4650), .B2(
        n3912), .ZN(n4553) );
  NAND2_X1 U4635 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3915), .ZN(n3932) );
  INV_X1 U4636 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4637 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3915), .B1(n4653), .B2(
        n3914), .ZN(n4535) );
  INV_X1 U4638 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U4639 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3916), .B1(n4655), .B2(
        n4727), .ZN(n4508) );
  NAND2_X1 U4640 ( .A1(n3917), .A2(REG1_REG_9__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4641 ( .A1(n3917), .A2(REG1_REG_9__SCAN_IN), .B1(n3366), .B2(n4657), .ZN(n4487) );
  NAND2_X1 U4642 ( .A1(n3920), .A2(REG1_REG_5__SCAN_IN), .ZN(n3919) );
  OAI21_X1 U4643 ( .B1(n3920), .B2(REG1_REG_5__SCAN_IN), .A(n3919), .ZN(n4443)
         );
  NOR2_X1 U4644 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  NOR2_X1 U4645 ( .A1(n3921), .A2(n4661), .ZN(n3922) );
  INV_X1 U4646 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4455) );
  XNOR2_X1 U4647 ( .A(n3921), .B(n4661), .ZN(n4454) );
  NOR2_X1 U4648 ( .A1(n4455), .A2(n4454), .ZN(n4453) );
  NOR2_X1 U4649 ( .A1(n3922), .A2(n4453), .ZN(n4467) );
  NAND2_X1 U4650 ( .A1(n3923), .A2(REG1_REG_7__SCAN_IN), .ZN(n4463) );
  NOR2_X1 U4651 ( .A1(n3923), .A2(REG1_REG_7__SCAN_IN), .ZN(n4462) );
  AOI21_X1 U4652 ( .B1(n4467), .B2(n4463), .A(n4462), .ZN(n3924) );
  NAND2_X1 U4653 ( .A1(n4475), .A2(n3924), .ZN(n3925) );
  XOR2_X1 U4654 ( .A(n4475), .B(n3924), .Z(n4477) );
  NAND2_X1 U4655 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4477), .ZN(n4476) );
  NAND2_X1 U4656 ( .A1(n4496), .A2(n3927), .ZN(n3928) );
  NAND2_X1 U4657 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4498), .ZN(n4497) );
  NAND2_X1 U4658 ( .A1(n3929), .A2(n3930), .ZN(n3931) );
  NAND2_X1 U4659 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U4660 ( .A1(n3933), .A2(n3934), .ZN(n3935) );
  NAND2_X1 U4661 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U4662 ( .A1(n3935), .A2(n4543), .ZN(n4552) );
  NAND2_X1 U4663 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U4664 ( .A1(n3936), .A2(n4551), .ZN(n3938) );
  NOR2_X1 U4665 ( .A1(n3937), .A2(n3938), .ZN(n3939) );
  INV_X1 U4666 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3940) );
  INV_X1 U4667 ( .A(n3941), .ZN(n4648) );
  AOI22_X1 U4668 ( .A1(n3941), .A2(n3940), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4648), .ZN(n4569) );
  NOR2_X1 U4669 ( .A1(n3942), .A2(n4570), .ZN(n4581) );
  NAND2_X1 U4670 ( .A1(n4582), .A2(n4581), .ZN(n4579) );
  OAI21_X1 U4671 ( .B1(n4585), .B2(n3943), .A(n4579), .ZN(n3946) );
  INV_X1 U4672 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3944) );
  MUX2_X1 U4673 ( .A(REG1_REG_19__SCAN_IN), .B(n3944), .S(n3949), .Z(n3945) );
  XNOR2_X1 U4674 ( .A(n3946), .B(n3945), .ZN(n3951) );
  AOI21_X1 U4675 ( .B1(n4578), .B2(ADDR_REG_19__SCAN_IN), .A(n3947), .ZN(n3948) );
  OAI21_X1 U4676 ( .B1(n4586), .B2(n3949), .A(n3948), .ZN(n3950) );
  AOI21_X1 U4677 ( .B1(n3951), .B2(n4580), .A(n3950), .ZN(n3952) );
  OAI21_X1 U4678 ( .B1(n3953), .B2(n4574), .A(n3952), .ZN(U3259) );
  XNOR2_X1 U4679 ( .A(n4224), .B(n3956), .ZN(n4344) );
  NAND2_X1 U4680 ( .A1(n3955), .A2(n3954), .ZN(n4226) );
  OAI21_X1 U4681 ( .B1(n3956), .B2(n4590), .A(n4226), .ZN(n4341) );
  NAND2_X1 U4682 ( .A1(n4205), .A2(n4341), .ZN(n3958) );
  NAND2_X1 U4683 ( .A1(n4634), .A2(REG2_REG_31__SCAN_IN), .ZN(n3957) );
  OAI211_X1 U4684 ( .C1(n4344), .C2(n4180), .A(n3958), .B(n3957), .ZN(U3260)
         );
  XNOR2_X1 U4685 ( .A(n3959), .B(n3960), .ZN(n4232) );
  XNOR2_X1 U4686 ( .A(n3961), .B(n3960), .ZN(n3966) );
  AOI22_X1 U4687 ( .A1(n3963), .A2(n4596), .B1(n4609), .B2(n3962), .ZN(n3964)
         );
  OAI21_X1 U4688 ( .B1(n4002), .B2(n4592), .A(n3964), .ZN(n3965) );
  AOI21_X1 U4689 ( .B1(n3966), .B2(n4621), .A(n3965), .ZN(n4231) );
  INV_X1 U4690 ( .A(n4231), .ZN(n3973) );
  INV_X1 U4691 ( .A(n3967), .ZN(n3968) );
  OAI21_X1 U4692 ( .B1(n3981), .B2(n3969), .A(n3968), .ZN(n4351) );
  AOI22_X1 U4693 ( .A1(n3970), .A2(n4622), .B1(n4634), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3971) );
  OAI21_X1 U4694 ( .B1(n4351), .B2(n4180), .A(n3971), .ZN(n3972) );
  AOI21_X1 U4695 ( .B1(n3973), .B2(n4205), .A(n3972), .ZN(n3974) );
  OAI21_X1 U4696 ( .B1(n4232), .B2(n4165), .A(n3974), .ZN(U3262) );
  NOR2_X1 U4697 ( .A1(n3975), .A2(n3979), .ZN(n3976) );
  OR2_X1 U4698 ( .A1(n3977), .A2(n3976), .ZN(n3978) );
  NAND2_X1 U4699 ( .A1(n3978), .A2(n4621), .ZN(n4238) );
  XNOR2_X1 U4700 ( .A(n3980), .B(n3979), .ZN(n4241) );
  NAND2_X1 U4701 ( .A1(n4241), .A2(n4194), .ZN(n3990) );
  INV_X1 U4702 ( .A(n3997), .ZN(n3982) );
  INV_X1 U4703 ( .A(n4355), .ZN(n3988) );
  AOI22_X1 U4704 ( .A1(n4634), .A2(REG2_REG_27__SCAN_IN), .B1(n3983), .B2(
        n4622), .ZN(n3984) );
  OAI21_X1 U4705 ( .B1(n4213), .B2(n3985), .A(n3984), .ZN(n3987) );
  OAI22_X1 U4706 ( .A1(n4239), .A2(n4214), .B1(n4018), .B2(n4215), .ZN(n3986)
         );
  AOI211_X1 U4707 ( .C1(n3988), .C2(n4629), .A(n3987), .B(n3986), .ZN(n3989)
         );
  OAI211_X1 U4708 ( .C1(n4634), .C2(n4238), .A(n3990), .B(n3989), .ZN(U3263)
         );
  NAND2_X1 U4709 ( .A1(n3992), .A2(n3991), .ZN(n3994) );
  INV_X1 U4710 ( .A(n3996), .ZN(n3993) );
  XNOR2_X1 U4711 ( .A(n3994), .B(n3993), .ZN(n3995) );
  NAND2_X1 U4712 ( .A1(n3995), .A2(n4621), .ZN(n4247) );
  XNOR2_X1 U4713 ( .A(n2249), .B(n3996), .ZN(n4250) );
  NAND2_X1 U4714 ( .A1(n4250), .A2(n4194), .ZN(n4007) );
  INV_X1 U4715 ( .A(n4019), .ZN(n3998) );
  OAI21_X1 U4716 ( .B1(n3998), .B2(n4001), .A(n3997), .ZN(n4359) );
  INV_X1 U4717 ( .A(n4359), .ZN(n4005) );
  AOI22_X1 U4718 ( .A1(n4634), .A2(REG2_REG_26__SCAN_IN), .B1(n3999), .B2(
        n4622), .ZN(n4000) );
  OAI21_X1 U4719 ( .B1(n4213), .B2(n4001), .A(n4000), .ZN(n4004) );
  OAI22_X1 U4720 ( .A1(n4002), .A2(n4214), .B1(n4248), .B2(n4215), .ZN(n4003)
         );
  AOI211_X1 U4721 ( .C1(n4005), .C2(n4629), .A(n4004), .B(n4003), .ZN(n4006)
         );
  OAI211_X1 U4722 ( .C1(n4634), .C2(n4247), .A(n4007), .B(n4006), .ZN(U3264)
         );
  XOR2_X1 U4723 ( .A(n4011), .B(n4008), .Z(n4254) );
  INV_X1 U4724 ( .A(n4254), .ZN(n4027) );
  NAND2_X1 U4725 ( .A1(n4010), .A2(n4009), .ZN(n4012) );
  XNOR2_X1 U4726 ( .A(n4012), .B(n4011), .ZN(n4013) );
  NAND2_X1 U4727 ( .A1(n4013), .A2(n4621), .ZN(n4017) );
  AOI22_X1 U4728 ( .A1(n4015), .A2(n4610), .B1(n4014), .B2(n4609), .ZN(n4016)
         );
  OAI211_X1 U4729 ( .C1(n4018), .C2(n4613), .A(n4017), .B(n4016), .ZN(n4253)
         );
  OAI21_X1 U4730 ( .B1(n4040), .B2(n4020), .A(n4019), .ZN(n4363) );
  NOR2_X1 U4731 ( .A1(n4363), .A2(n4180), .ZN(n4025) );
  NAND2_X1 U4732 ( .A1(n4021), .A2(n4622), .ZN(n4022) );
  OAI21_X1 U4733 ( .B1(n4205), .B2(n4023), .A(n4022), .ZN(n4024) );
  AOI211_X1 U4734 ( .C1(n4253), .C2(n4205), .A(n4025), .B(n4024), .ZN(n4026)
         );
  OAI21_X1 U4735 ( .B1(n4027), .B2(n4165), .A(n4026), .ZN(U3265) );
  XOR2_X1 U4736 ( .A(n4032), .B(n4028), .Z(n4258) );
  INV_X1 U4737 ( .A(n4258), .ZN(n4046) );
  NAND2_X1 U4738 ( .A1(n4030), .A2(n4029), .ZN(n4031) );
  XOR2_X1 U4739 ( .A(n4032), .B(n4031), .Z(n4033) );
  NAND2_X1 U4740 ( .A1(n4033), .A2(n4621), .ZN(n4037) );
  AOI22_X1 U4741 ( .A1(n4035), .A2(n4610), .B1(n4609), .B2(n4034), .ZN(n4036)
         );
  OAI211_X1 U4742 ( .C1(n4248), .C2(n4613), .A(n4037), .B(n4036), .ZN(n4257)
         );
  NOR2_X1 U4743 ( .A1(n4059), .A2(n4038), .ZN(n4039) );
  OR2_X1 U4744 ( .A1(n4040), .A2(n4039), .ZN(n4367) );
  NOR2_X1 U4745 ( .A1(n4367), .A2(n4180), .ZN(n4044) );
  OAI22_X1 U4746 ( .A1(n4205), .A2(n4042), .B1(n4041), .B2(n4190), .ZN(n4043)
         );
  AOI211_X1 U4747 ( .C1(n4257), .C2(n4205), .A(n4044), .B(n4043), .ZN(n4045)
         );
  OAI21_X1 U4748 ( .B1(n4046), .B2(n4165), .A(n4045), .ZN(U3266) );
  XNOR2_X1 U4749 ( .A(n4047), .B(n4050), .ZN(n4262) );
  INV_X1 U4750 ( .A(n4262), .ZN(n4065) );
  OR2_X1 U4751 ( .A1(n4087), .A2(n4086), .ZN(n4089) );
  NAND2_X1 U4752 ( .A1(n4089), .A2(n4048), .ZN(n4069) );
  AOI21_X1 U4753 ( .B1(n4069), .B2(n4068), .A(n4049), .ZN(n4051) );
  XNOR2_X1 U4754 ( .A(n4051), .B(n4050), .ZN(n4052) );
  NAND2_X1 U4755 ( .A1(n4052), .A2(n4621), .ZN(n4055) );
  AOI22_X1 U4756 ( .A1(n4270), .A2(n4610), .B1(n4609), .B2(n4053), .ZN(n4054)
         );
  OAI211_X1 U4757 ( .C1(n4056), .C2(n4613), .A(n4055), .B(n4054), .ZN(n4261)
         );
  NOR2_X1 U4758 ( .A1(n4075), .A2(n4057), .ZN(n4058) );
  OR2_X1 U4759 ( .A1(n4059), .A2(n4058), .ZN(n4371) );
  NOR2_X1 U4760 ( .A1(n4371), .A2(n4180), .ZN(n4063) );
  OAI22_X1 U4761 ( .A1(n4205), .A2(n4061), .B1(n4060), .B2(n4190), .ZN(n4062)
         );
  AOI211_X1 U4762 ( .C1(n4261), .C2(n4205), .A(n4063), .B(n4062), .ZN(n4064)
         );
  OAI21_X1 U4763 ( .B1(n4065), .B2(n4165), .A(n4064), .ZN(U3267) );
  AOI21_X1 U4764 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n4266) );
  INV_X1 U4765 ( .A(n4266), .ZN(n4084) );
  XNOR2_X1 U4766 ( .A(n4069), .B(n4068), .ZN(n4070) );
  NAND2_X1 U4767 ( .A1(n4070), .A2(n4621), .ZN(n4073) );
  AOI22_X1 U4768 ( .A1(n4107), .A2(n4610), .B1(n4071), .B2(n4609), .ZN(n4072)
         );
  OAI211_X1 U4769 ( .C1(n4074), .C2(n4613), .A(n4073), .B(n4072), .ZN(n4265)
         );
  INV_X1 U4770 ( .A(n4090), .ZN(n4077) );
  OAI21_X1 U4771 ( .B1(n4077), .B2(n4076), .A(n2272), .ZN(n4375) );
  NOR2_X1 U4772 ( .A1(n4375), .A2(n4180), .ZN(n4082) );
  INV_X1 U4773 ( .A(n4078), .ZN(n4079) );
  OAI22_X1 U4774 ( .A1(n4205), .A2(n4080), .B1(n4079), .B2(n4190), .ZN(n4081)
         );
  AOI211_X1 U4775 ( .C1(n4265), .C2(n4205), .A(n4082), .B(n4081), .ZN(n4083)
         );
  OAI21_X1 U4776 ( .B1(n4084), .B2(n4165), .A(n4083), .ZN(U3268) );
  XNOR2_X1 U4777 ( .A(n4085), .B(n4086), .ZN(n4275) );
  INV_X1 U4778 ( .A(n4275), .ZN(n4101) );
  NAND2_X1 U4779 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  AOI21_X1 U4780 ( .B1(n4089), .B2(n4088), .A(n4598), .ZN(n4274) );
  INV_X1 U4781 ( .A(n4278), .ZN(n4092) );
  OAI21_X1 U4782 ( .B1(n4092), .B2(n4091), .A(n4090), .ZN(n4379) );
  OAI22_X1 U4783 ( .A1(n4205), .A2(n4094), .B1(n4093), .B2(n4190), .ZN(n4097)
         );
  OAI22_X1 U4784 ( .A1(n4272), .A2(n4215), .B1(n4214), .B2(n4095), .ZN(n4096)
         );
  AOI211_X1 U4785 ( .C1(n4269), .C2(n4175), .A(n4097), .B(n4096), .ZN(n4098)
         );
  OAI21_X1 U4786 ( .B1(n4379), .B2(n4180), .A(n4098), .ZN(n4099) );
  AOI21_X1 U4787 ( .B1(n4274), .B2(n4205), .A(n4099), .ZN(n4100) );
  OAI21_X1 U4788 ( .B1(n4101), .B2(n4165), .A(n4100), .ZN(U3269) );
  INV_X1 U4789 ( .A(n4102), .ZN(n4103) );
  NAND2_X1 U4790 ( .A1(n4104), .A2(n4103), .ZN(n4106) );
  INV_X1 U4791 ( .A(n4111), .ZN(n4105) );
  XNOR2_X1 U4792 ( .A(n4106), .B(n4105), .ZN(n4114) );
  AOI22_X1 U4793 ( .A1(n4107), .A2(n4596), .B1(n4609), .B2(n4116), .ZN(n4108)
         );
  OAI21_X1 U4794 ( .B1(n4109), .B2(n4592), .A(n4108), .ZN(n4113) );
  XNOR2_X1 U4795 ( .A(n4110), .B(n4111), .ZN(n4282) );
  NOR2_X1 U4796 ( .A1(n4282), .A2(n4617), .ZN(n4112) );
  AOI211_X1 U4797 ( .C1(n4114), .C2(n4621), .A(n4113), .B(n4112), .ZN(n4281)
         );
  INV_X1 U4798 ( .A(n4282), .ZN(n4121) );
  INV_X1 U4799 ( .A(n4115), .ZN(n4140) );
  NAND2_X1 U4800 ( .A1(n4140), .A2(n4116), .ZN(n4279) );
  AND3_X1 U4801 ( .A1(n4279), .A2(n4629), .A3(n4278), .ZN(n4120) );
  OAI22_X1 U4802 ( .A1(n4205), .A2(n4118), .B1(n4117), .B2(n4190), .ZN(n4119)
         );
  AOI211_X1 U4803 ( .C1(n4121), .C2(n4631), .A(n4120), .B(n4119), .ZN(n4122)
         );
  OAI21_X1 U4804 ( .B1(n4281), .B2(n4634), .A(n4122), .ZN(U3270) );
  INV_X1 U4805 ( .A(n4124), .ZN(n4126) );
  OAI21_X1 U4806 ( .B1(n4123), .B2(n4126), .A(n4125), .ZN(n4154) );
  INV_X1 U4807 ( .A(n4127), .ZN(n4129) );
  OAI21_X1 U4808 ( .B1(n4154), .B2(n4129), .A(n4128), .ZN(n4130) );
  XNOR2_X1 U4809 ( .A(n4130), .B(n4137), .ZN(n4135) );
  OAI22_X1 U4810 ( .A1(n4272), .A2(n4613), .B1(n4590), .B2(n4131), .ZN(n4132)
         );
  AOI21_X1 U4811 ( .B1(n4610), .B2(n4133), .A(n4132), .ZN(n4134) );
  OAI21_X1 U4812 ( .B1(n4135), .B2(n4598), .A(n4134), .ZN(n4283) );
  INV_X1 U4813 ( .A(n4283), .ZN(n4145) );
  XOR2_X1 U4814 ( .A(n4137), .B(n4136), .Z(n4284) );
  NAND2_X1 U4815 ( .A1(n4150), .A2(n4138), .ZN(n4139) );
  NAND2_X1 U4816 ( .A1(n4140), .A2(n4139), .ZN(n4384) );
  AOI22_X1 U4817 ( .A1(n4634), .A2(REG2_REG_19__SCAN_IN), .B1(n4141), .B2(
        n4622), .ZN(n4142) );
  OAI21_X1 U4818 ( .B1(n4384), .B2(n4180), .A(n4142), .ZN(n4143) );
  AOI21_X1 U4819 ( .B1(n4284), .B2(n4194), .A(n4143), .ZN(n4144) );
  OAI21_X1 U4820 ( .B1(n4634), .B2(n4145), .A(n4144), .ZN(U3271) );
  INV_X1 U4821 ( .A(n4146), .ZN(n4147) );
  AOI21_X1 U4822 ( .B1(n4153), .B2(n4148), .A(n4147), .ZN(n4288) );
  AOI22_X1 U4823 ( .A1(n4634), .A2(REG2_REG_18__SCAN_IN), .B1(n4149), .B2(
        n4622), .ZN(n4164) );
  INV_X1 U4824 ( .A(n4171), .ZN(n4152) );
  OAI211_X1 U4825 ( .C1(n4152), .C2(n4151), .A(n4701), .B(n4150), .ZN(n4286)
         );
  XNOR2_X1 U4826 ( .A(n4154), .B(n4153), .ZN(n4160) );
  AOI22_X1 U4827 ( .A1(n4156), .A2(n4596), .B1(n4609), .B2(n4155), .ZN(n4157)
         );
  OAI21_X1 U4828 ( .B1(n4158), .B2(n4592), .A(n4157), .ZN(n4159) );
  AOI21_X1 U4829 ( .B1(n4160), .B2(n4621), .A(n4159), .ZN(n4287) );
  OAI21_X1 U4830 ( .B1(n4161), .B2(n4286), .A(n4287), .ZN(n4162) );
  NAND2_X1 U4831 ( .A1(n4162), .A2(n4205), .ZN(n4163) );
  OAI211_X1 U4832 ( .C1(n4288), .C2(n4165), .A(n4164), .B(n4163), .ZN(U3272)
         );
  INV_X1 U4833 ( .A(n4168), .ZN(n4166) );
  XNOR2_X1 U4834 ( .A(n4123), .B(n4166), .ZN(n4167) );
  NAND2_X1 U4835 ( .A1(n4167), .A2(n4621), .ZN(n4296) );
  XNOR2_X1 U4836 ( .A(n4169), .B(n4168), .ZN(n4289) );
  NAND2_X1 U4837 ( .A1(n4300), .A2(n4176), .ZN(n4170) );
  NAND2_X1 U4838 ( .A1(n4171), .A2(n4170), .ZN(n4389) );
  OAI22_X1 U4839 ( .A1(n4205), .A2(n4173), .B1(n4172), .B2(n4190), .ZN(n4174)
         );
  AOI21_X1 U4840 ( .B1(n4176), .B2(n4175), .A(n4174), .ZN(n4179) );
  OAI22_X1 U4841 ( .A1(n4292), .A2(n4215), .B1(n4214), .B2(n4291), .ZN(n4177)
         );
  INV_X1 U4842 ( .A(n4177), .ZN(n4178) );
  OAI211_X1 U4843 ( .C1(n4389), .C2(n4180), .A(n4179), .B(n4178), .ZN(n4181)
         );
  AOI21_X1 U4844 ( .B1(n4289), .B2(n4194), .A(n4181), .ZN(n4182) );
  OAI21_X1 U4845 ( .B1(n4634), .B2(n4296), .A(n4182), .ZN(U3273) );
  XNOR2_X1 U4846 ( .A(n4183), .B(n2669), .ZN(n4186) );
  AOI22_X1 U4847 ( .A1(n4420), .A2(n4596), .B1(n4609), .B2(n4189), .ZN(n4184)
         );
  OAI21_X1 U4848 ( .B1(n4416), .B2(n4592), .A(n4184), .ZN(n4185) );
  AOI21_X1 U4849 ( .B1(n4186), .B2(n4621), .A(n4185), .ZN(n4303) );
  OAI21_X1 U4850 ( .B1(n4188), .B2(n2669), .A(n4187), .ZN(n4304) );
  INV_X1 U4851 ( .A(n4304), .ZN(n4195) );
  NAND2_X1 U4852 ( .A1(n2252), .A2(n4189), .ZN(n4301) );
  AND3_X1 U4853 ( .A1(n4301), .A2(n4629), .A3(n4300), .ZN(n4193) );
  OAI22_X1 U4854 ( .A1(n4205), .A2(n4191), .B1(n4430), .B2(n4190), .ZN(n4192)
         );
  AOI211_X1 U4855 ( .C1(n4195), .C2(n4194), .A(n4193), .B(n4192), .ZN(n4196)
         );
  OAI21_X1 U4856 ( .B1(n4634), .B2(n4303), .A(n4196), .ZN(U3274) );
  AOI21_X1 U4857 ( .B1(n4199), .B2(n4198), .A(n4197), .ZN(n4312) );
  INV_X1 U4858 ( .A(n4200), .ZN(n4201) );
  AOI21_X1 U4859 ( .B1(n4203), .B2(n4202), .A(n4201), .ZN(n4204) );
  OAI22_X1 U4860 ( .A1(n4312), .A2(n4617), .B1(n4598), .B2(n4204), .ZN(n4316)
         );
  NAND2_X1 U4861 ( .A1(n4316), .A2(n4205), .ZN(n4220) );
  INV_X1 U4862 ( .A(n4207), .ZN(n4208) );
  OAI21_X1 U4863 ( .B1(n4209), .B2(n4212), .A(n4208), .ZN(n4398) );
  INV_X1 U4864 ( .A(n4398), .ZN(n4218) );
  AOI22_X1 U4865 ( .A1(n4634), .A2(REG2_REG_14__SCAN_IN), .B1(n4210), .B2(
        n4622), .ZN(n4211) );
  OAI21_X1 U4866 ( .B1(n4213), .B2(n4212), .A(n4211), .ZN(n4217) );
  OAI22_X1 U4867 ( .A1(n4331), .A2(n4215), .B1(n4214), .B2(n4416), .ZN(n4216)
         );
  AOI211_X1 U4868 ( .C1(n4218), .C2(n4629), .A(n4217), .B(n4216), .ZN(n4219)
         );
  OAI211_X1 U4869 ( .C1(n4312), .C2(n4221), .A(n4220), .B(n4219), .ZN(U3276)
         );
  NAND2_X1 U4870 ( .A1(n4729), .A2(n4341), .ZN(n4223) );
  NAND2_X1 U4871 ( .A1(n4726), .A2(REG1_REG_31__SCAN_IN), .ZN(n4222) );
  OAI211_X1 U4872 ( .C1(n4344), .C2(n4714), .A(n4223), .B(n4222), .ZN(U3549)
         );
  AOI21_X1 U4873 ( .B1(n4228), .B2(n4225), .A(n4224), .ZN(n4432) );
  INV_X1 U4874 ( .A(n4432), .ZN(n4347) );
  INV_X1 U4875 ( .A(n4226), .ZN(n4227) );
  AOI21_X1 U4876 ( .B1(n4228), .B2(n4609), .A(n4227), .ZN(n4434) );
  INV_X1 U4877 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4229) );
  MUX2_X1 U4878 ( .A(n4434), .B(n4229), .S(n4726), .Z(n4230) );
  OAI21_X1 U4879 ( .B1(n4347), .B2(n4714), .A(n4230), .ZN(U3548) );
  OAI21_X1 U4880 ( .B1(n4232), .B2(n4337), .A(n4231), .ZN(n4348) );
  INV_X1 U4881 ( .A(n4233), .ZN(n4234) );
  OAI21_X1 U4882 ( .B1(n4714), .B2(n4351), .A(n4234), .ZN(U3546) );
  INV_X1 U4883 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U4884 ( .A1(n4236), .A2(n4610), .B1(n4235), .B2(n4609), .ZN(n4237)
         );
  OAI211_X1 U4885 ( .C1(n4239), .C2(n4613), .A(n4238), .B(n4237), .ZN(n4240)
         );
  AOI21_X1 U4886 ( .B1(n4241), .B2(n4686), .A(n4240), .ZN(n4352) );
  MUX2_X1 U4887 ( .A(n4242), .B(n4352), .S(n4729), .Z(n4243) );
  OAI21_X1 U4888 ( .B1(n4714), .B2(n4355), .A(n4243), .ZN(U3545) );
  INV_X1 U4889 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4890 ( .A1(n4245), .A2(n4596), .B1(n4609), .B2(n4244), .ZN(n4246)
         );
  OAI211_X1 U4891 ( .C1(n4248), .C2(n4592), .A(n4247), .B(n4246), .ZN(n4249)
         );
  AOI21_X1 U4892 ( .B1(n4250), .B2(n4686), .A(n4249), .ZN(n4356) );
  MUX2_X1 U4893 ( .A(n4251), .B(n4356), .S(n4729), .Z(n4252) );
  OAI21_X1 U4894 ( .B1(n4714), .B2(n4359), .A(n4252), .ZN(U3544) );
  INV_X1 U4895 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4255) );
  AOI21_X1 U4896 ( .B1(n4254), .B2(n4686), .A(n4253), .ZN(n4360) );
  MUX2_X1 U4897 ( .A(n4255), .B(n4360), .S(n4729), .Z(n4256) );
  OAI21_X1 U4898 ( .B1(n4714), .B2(n4363), .A(n4256), .ZN(U3543) );
  INV_X1 U4899 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4259) );
  AOI21_X1 U4900 ( .B1(n4258), .B2(n4686), .A(n4257), .ZN(n4364) );
  MUX2_X1 U4901 ( .A(n4259), .B(n4364), .S(n4729), .Z(n4260) );
  OAI21_X1 U4902 ( .B1(n4714), .B2(n4367), .A(n4260), .ZN(U3542) );
  INV_X1 U4903 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4263) );
  AOI21_X1 U4904 ( .B1(n4262), .B2(n4686), .A(n4261), .ZN(n4368) );
  MUX2_X1 U4905 ( .A(n4263), .B(n4368), .S(n4729), .Z(n4264) );
  OAI21_X1 U4906 ( .B1(n4714), .B2(n4371), .A(n4264), .ZN(U3541) );
  INV_X1 U4907 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4267) );
  AOI21_X1 U4908 ( .B1(n4266), .B2(n4686), .A(n4265), .ZN(n4372) );
  MUX2_X1 U4909 ( .A(n4267), .B(n4372), .S(n4729), .Z(n4268) );
  OAI21_X1 U4910 ( .B1(n4714), .B2(n4375), .A(n4268), .ZN(U3540) );
  INV_X1 U4911 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4912 ( .A1(n4270), .A2(n4596), .B1(n4609), .B2(n4269), .ZN(n4271)
         );
  OAI21_X1 U4913 ( .B1(n4272), .B2(n4592), .A(n4271), .ZN(n4273) );
  AOI211_X1 U4914 ( .C1(n4275), .C2(n4686), .A(n4274), .B(n4273), .ZN(n4376)
         );
  MUX2_X1 U4915 ( .A(n4276), .B(n4376), .S(n4729), .Z(n4277) );
  OAI21_X1 U4916 ( .B1(n4714), .B2(n4379), .A(n4277), .ZN(U3539) );
  NAND3_X1 U4917 ( .A1(n4279), .A2(n4701), .A3(n4278), .ZN(n4280) );
  OAI211_X1 U4918 ( .C1(n4282), .C2(n4669), .A(n4281), .B(n4280), .ZN(n4380)
         );
  MUX2_X1 U4919 ( .A(REG1_REG_20__SCAN_IN), .B(n4380), .S(n4729), .Z(U3538) );
  AOI21_X1 U4920 ( .B1(n4284), .B2(n4686), .A(n4283), .ZN(n4381) );
  MUX2_X1 U4921 ( .A(n3944), .B(n4381), .S(n4729), .Z(n4285) );
  OAI21_X1 U4922 ( .B1(n4714), .B2(n4384), .A(n4285), .ZN(U3537) );
  OAI211_X1 U4923 ( .C1(n4288), .C2(n4337), .A(n4287), .B(n4286), .ZN(n4385)
         );
  MUX2_X1 U4924 ( .A(REG1_REG_18__SCAN_IN), .B(n4385), .S(n4729), .Z(U3536) );
  NAND2_X1 U4925 ( .A1(n4289), .A2(n4686), .ZN(n4298) );
  OAI22_X1 U4926 ( .A1(n4291), .A2(n4613), .B1(n4590), .B2(n4290), .ZN(n4294)
         );
  NOR2_X1 U4927 ( .A1(n4292), .A2(n4592), .ZN(n4293) );
  NOR2_X1 U4928 ( .A1(n4294), .A2(n4293), .ZN(n4295) );
  AND2_X1 U4929 ( .A1(n4296), .A2(n4295), .ZN(n4297) );
  MUX2_X1 U4930 ( .A(n3940), .B(n4386), .S(n4729), .Z(n4299) );
  OAI21_X1 U4931 ( .B1(n4714), .B2(n4389), .A(n4299), .ZN(U3535) );
  NAND3_X1 U4932 ( .A1(n4301), .A2(n4701), .A3(n4300), .ZN(n4302) );
  OAI211_X1 U4933 ( .C1(n4304), .C2(n4337), .A(n4303), .B(n4302), .ZN(n4390)
         );
  MUX2_X1 U4934 ( .A(REG1_REG_16__SCAN_IN), .B(n4390), .S(n4729), .Z(U3534) );
  AOI22_X1 U4935 ( .A1(n4306), .A2(n4596), .B1(n4609), .B2(n4305), .ZN(n4307)
         );
  OAI211_X1 U4936 ( .C1(n4324), .C2(n4592), .A(n4308), .B(n4307), .ZN(n4309)
         );
  AOI21_X1 U4937 ( .B1(n4310), .B2(n4686), .A(n4309), .ZN(n4391) );
  MUX2_X1 U4938 ( .A(n3912), .B(n4391), .S(n4729), .Z(n4311) );
  OAI21_X1 U4939 ( .B1(n4714), .B2(n4394), .A(n4311), .ZN(U3533) );
  INV_X1 U4940 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4319) );
  INV_X1 U4941 ( .A(n4312), .ZN(n4318) );
  AOI22_X1 U4942 ( .A1(n4314), .A2(n4596), .B1(n4609), .B2(n4313), .ZN(n4315)
         );
  OAI21_X1 U4943 ( .B1(n4331), .B2(n4592), .A(n4315), .ZN(n4317) );
  AOI211_X1 U4944 ( .C1(n4702), .C2(n4318), .A(n4317), .B(n4316), .ZN(n4395)
         );
  MUX2_X1 U4945 ( .A(n4319), .B(n4395), .S(n4729), .Z(n4320) );
  OAI21_X1 U4946 ( .B1(n4714), .B2(n4398), .A(n4320), .ZN(U3532) );
  NOR2_X1 U4947 ( .A1(n4321), .A2(n4337), .ZN(n4328) );
  NOR2_X1 U4948 ( .A1(n4322), .A2(n4592), .ZN(n4326) );
  OAI22_X1 U4949 ( .A1(n4324), .A2(n4613), .B1(n4590), .B2(n4323), .ZN(n4325)
         );
  NOR4_X1 U4950 ( .A1(n4328), .A2(n4327), .A3(n4326), .A4(n4325), .ZN(n4399)
         );
  MUX2_X1 U4951 ( .A(n3914), .B(n4399), .S(n4729), .Z(n4329) );
  OAI21_X1 U4952 ( .B1(n4714), .B2(n4402), .A(n4329), .ZN(U3531) );
  INV_X1 U4953 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4339) );
  OAI22_X1 U4954 ( .A1(n4331), .A2(n4613), .B1(n4590), .B2(n4330), .ZN(n4333)
         );
  AOI211_X1 U4955 ( .C1(n4610), .C2(n4334), .A(n4333), .B(n4332), .ZN(n4335)
         );
  OAI21_X1 U4956 ( .B1(n4337), .B2(n4336), .A(n4335), .ZN(n4338) );
  INV_X1 U4957 ( .A(n4338), .ZN(n4403) );
  MUX2_X1 U4958 ( .A(n4339), .B(n4403), .S(n4729), .Z(n4340) );
  OAI21_X1 U4959 ( .B1(n4406), .B2(n4714), .A(n4340), .ZN(U3530) );
  NAND2_X1 U4960 ( .A1(n4708), .A2(n4341), .ZN(n4343) );
  NAND2_X1 U4961 ( .A1(n4706), .A2(REG0_REG_31__SCAN_IN), .ZN(n4342) );
  OAI211_X1 U4962 ( .C1(n4344), .C2(n4677), .A(n4343), .B(n4342), .ZN(U3517)
         );
  INV_X1 U4963 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4345) );
  MUX2_X1 U4964 ( .A(n4434), .B(n4345), .S(n4706), .Z(n4346) );
  OAI21_X1 U4965 ( .B1(n4347), .B2(n4677), .A(n4346), .ZN(U3516) );
  INV_X1 U4966 ( .A(n4349), .ZN(n4350) );
  OAI21_X1 U4967 ( .B1(n4351), .B2(n4677), .A(n4350), .ZN(U3514) );
  INV_X1 U4968 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4353) );
  MUX2_X1 U4969 ( .A(n4353), .B(n4352), .S(n4708), .Z(n4354) );
  OAI21_X1 U4970 ( .B1(n4355), .B2(n4677), .A(n4354), .ZN(U3513) );
  INV_X1 U4971 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4357) );
  MUX2_X1 U4972 ( .A(n4357), .B(n4356), .S(n4708), .Z(n4358) );
  OAI21_X1 U4973 ( .B1(n4359), .B2(n4677), .A(n4358), .ZN(U3512) );
  INV_X1 U4974 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4361) );
  MUX2_X1 U4975 ( .A(n4361), .B(n4360), .S(n4708), .Z(n4362) );
  OAI21_X1 U4976 ( .B1(n4363), .B2(n4677), .A(n4362), .ZN(U3511) );
  INV_X1 U4977 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4365) );
  MUX2_X1 U4978 ( .A(n4365), .B(n4364), .S(n4708), .Z(n4366) );
  OAI21_X1 U4979 ( .B1(n4367), .B2(n4677), .A(n4366), .ZN(U3510) );
  INV_X1 U4980 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4369) );
  MUX2_X1 U4981 ( .A(n4369), .B(n4368), .S(n4708), .Z(n4370) );
  OAI21_X1 U4982 ( .B1(n4371), .B2(n4677), .A(n4370), .ZN(U3509) );
  INV_X1 U4983 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4373) );
  MUX2_X1 U4984 ( .A(n4373), .B(n4372), .S(n4708), .Z(n4374) );
  OAI21_X1 U4985 ( .B1(n4375), .B2(n4677), .A(n4374), .ZN(U3508) );
  INV_X1 U4986 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4377) );
  MUX2_X1 U4987 ( .A(n4377), .B(n4376), .S(n4708), .Z(n4378) );
  OAI21_X1 U4988 ( .B1(n4379), .B2(n4677), .A(n4378), .ZN(U3507) );
  MUX2_X1 U4989 ( .A(REG0_REG_20__SCAN_IN), .B(n4380), .S(n4708), .Z(U3506) );
  INV_X1 U4990 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4382) );
  MUX2_X1 U4991 ( .A(n4382), .B(n4381), .S(n4708), .Z(n4383) );
  OAI21_X1 U4992 ( .B1(n4384), .B2(n4677), .A(n4383), .ZN(U3505) );
  MUX2_X1 U4993 ( .A(REG0_REG_18__SCAN_IN), .B(n4385), .S(n4708), .Z(U3503) );
  INV_X1 U4994 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4387) );
  MUX2_X1 U4995 ( .A(n4387), .B(n4386), .S(n4708), .Z(n4388) );
  OAI21_X1 U4996 ( .B1(n4389), .B2(n4677), .A(n4388), .ZN(U3501) );
  MUX2_X1 U4997 ( .A(REG0_REG_16__SCAN_IN), .B(n4390), .S(n4708), .Z(U3499) );
  INV_X1 U4998 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4392) );
  MUX2_X1 U4999 ( .A(n4392), .B(n4391), .S(n4708), .Z(n4393) );
  OAI21_X1 U5000 ( .B1(n4394), .B2(n4677), .A(n4393), .ZN(U3497) );
  INV_X1 U5001 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U5002 ( .A(n4396), .B(n4395), .S(n4708), .Z(n4397) );
  OAI21_X1 U5003 ( .B1(n4398), .B2(n4677), .A(n4397), .ZN(U3495) );
  INV_X1 U5004 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4400) );
  MUX2_X1 U5005 ( .A(n4400), .B(n4399), .S(n4708), .Z(n4401) );
  OAI21_X1 U5006 ( .B1(n4402), .B2(n4677), .A(n4401), .ZN(U3493) );
  INV_X1 U5007 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4404) );
  MUX2_X1 U5008 ( .A(n4404), .B(n4403), .S(n4708), .Z(n4405) );
  OAI21_X1 U5009 ( .B1(n4406), .B2(n4677), .A(n4405), .ZN(U3491) );
  MUX2_X1 U5010 ( .A(n4407), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5011 ( .A(n4408), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5012 ( .A(n2844), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5013 ( .A(DATAI_22_), .B(n4409), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5014 ( .A(DATAI_4_), .B(n4410), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5015 ( .A(DATAI_3_), .B(n4411), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5016 ( .A(n4412), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5017 ( .A(n4413), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5018 ( .A(DATAI_28_), .ZN(n5066) );
  AOI22_X1 U5019 ( .A1(STATE_REG_SCAN_IN), .A2(n4414), .B1(n5066), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5020 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4803) );
  NOR2_X1 U5021 ( .A1(STATE_REG_SCAN_IN), .A2(n4803), .ZN(n4559) );
  OAI22_X1 U5022 ( .A1(n4418), .A2(n4417), .B1(n4416), .B2(n4415), .ZN(n4419)
         );
  AOI211_X1 U5023 ( .C1(n4421), .C2(n4420), .A(n4559), .B(n4419), .ZN(n4429)
         );
  AOI21_X1 U5024 ( .B1(n4423), .B2(n4422), .A(n3671), .ZN(n4424) );
  XOR2_X1 U5025 ( .A(n4425), .B(n4424), .Z(n4427) );
  NAND2_X1 U5026 ( .A1(n4427), .A2(n4426), .ZN(n4428) );
  OAI211_X1 U5027 ( .C1(n4431), .C2(n4430), .A(n4429), .B(n4428), .ZN(U3223)
         );
  AOI22_X1 U5028 ( .A1(n4432), .A2(n4629), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4634), .ZN(n4433) );
  OAI21_X1 U5029 ( .B1(n4634), .B2(n4434), .A(n4433), .ZN(U3261) );
  INV_X1 U5030 ( .A(n4437), .ZN(n4435) );
  OAI211_X1 U5031 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4436), .A(n4438), .B(n4435), 
        .ZN(n4441) );
  INV_X1 U5032 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5033 ( .A1(n4438), .A2(n4437), .B1(n4580), .B2(n4709), .ZN(n4440)
         );
  AOI22_X1 U5034 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4578), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4439) );
  OAI221_X1 U5035 ( .B1(IR_REG_0__SCAN_IN), .B2(n4441), .C1(n2277), .C2(n4440), 
        .A(n4439), .ZN(U3240) );
  AOI211_X1 U5036 ( .C1(n4444), .C2(n4443), .A(n4442), .B(n4452), .ZN(n4446)
         );
  AOI211_X1 U5037 ( .C1(n4578), .C2(ADDR_REG_5__SCAN_IN), .A(n4446), .B(n4445), 
        .ZN(n4451) );
  OAI211_X1 U5038 ( .C1(n4449), .C2(n4448), .A(n4527), .B(n4447), .ZN(n4450)
         );
  OAI211_X1 U5039 ( .C1(n4586), .C2(n4662), .A(n4451), .B(n4450), .ZN(U3245)
         );
  AOI211_X1 U5040 ( .C1(n4455), .C2(n4454), .A(n4453), .B(n4452), .ZN(n4457)
         );
  AOI211_X1 U5041 ( .C1(n4578), .C2(ADDR_REG_6__SCAN_IN), .A(n4457), .B(n4456), 
        .ZN(n4461) );
  OAI211_X1 U5042 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4459), .A(n4527), .B(n4458), 
        .ZN(n4460) );
  OAI211_X1 U5043 ( .C1(n4586), .C2(n4661), .A(n4461), .B(n4460), .ZN(U3246)
         );
  INV_X1 U5044 ( .A(n4462), .ZN(n4464) );
  NAND2_X1 U5045 ( .A1(n4464), .A2(n4463), .ZN(n4466) );
  OAI21_X1 U5046 ( .B1(n4467), .B2(n4466), .A(n4580), .ZN(n4465) );
  AOI21_X1 U5047 ( .B1(n4467), .B2(n4466), .A(n4465), .ZN(n4469) );
  AOI211_X1 U5048 ( .C1(n4578), .C2(ADDR_REG_7__SCAN_IN), .A(n4469), .B(n4468), 
        .ZN(n4474) );
  OAI211_X1 U5049 ( .C1(n4472), .C2(n4471), .A(n4527), .B(n4470), .ZN(n4473)
         );
  OAI211_X1 U5050 ( .C1(n4586), .C2(n4659), .A(n4474), .B(n4473), .ZN(U3247)
         );
  OAI211_X1 U5051 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4477), .A(n4580), .B(n4476), 
        .ZN(n4481) );
  OAI211_X1 U5052 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4479), .A(n4527), .B(n4478), 
        .ZN(n4480) );
  OAI211_X1 U5053 ( .C1(n4586), .C2(n2378), .A(n4481), .B(n4480), .ZN(n4482)
         );
  AOI211_X1 U5054 ( .C1(n4578), .C2(ADDR_REG_8__SCAN_IN), .A(n4483), .B(n4482), 
        .ZN(n4484) );
  INV_X1 U5055 ( .A(n4484), .ZN(U3248) );
  OAI211_X1 U5056 ( .C1(n4487), .C2(n4486), .A(n4580), .B(n4485), .ZN(n4492)
         );
  OAI211_X1 U5057 ( .C1(n4490), .C2(n4489), .A(n4527), .B(n4488), .ZN(n4491)
         );
  OAI211_X1 U5058 ( .C1(n4586), .C2(n4657), .A(n4492), .B(n4491), .ZN(n4493)
         );
  AOI211_X1 U5059 ( .C1(n4578), .C2(ADDR_REG_9__SCAN_IN), .A(n4494), .B(n4493), 
        .ZN(n4495) );
  INV_X1 U5060 ( .A(n4495), .ZN(U3249) );
  OAI211_X1 U5061 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4498), .A(n4580), .B(n4497), .ZN(n4502) );
  OAI211_X1 U5062 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4500), .A(n4527), .B(n4499), .ZN(n4501) );
  OAI211_X1 U5063 ( .C1(n4586), .C2(n2377), .A(n4502), .B(n4501), .ZN(n4503)
         );
  AOI211_X1 U5064 ( .C1(n4578), .C2(ADDR_REG_10__SCAN_IN), .A(n4504), .B(n4503), .ZN(n4505) );
  INV_X1 U5065 ( .A(n4505), .ZN(U3250) );
  OAI211_X1 U5066 ( .C1(n4508), .C2(n4507), .A(n4580), .B(n4506), .ZN(n4513)
         );
  OAI211_X1 U5067 ( .C1(n4511), .C2(n4510), .A(n4527), .B(n4509), .ZN(n4512)
         );
  OAI211_X1 U5068 ( .C1(n4586), .C2(n4655), .A(n4513), .B(n4512), .ZN(n4514)
         );
  AOI211_X1 U5069 ( .C1(n4578), .C2(ADDR_REG_11__SCAN_IN), .A(n4515), .B(n4514), .ZN(n4516) );
  INV_X1 U5070 ( .A(n4516), .ZN(U3251) );
  OAI211_X1 U5071 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4518), .A(n4527), .B(n4517), .ZN(n4520) );
  NAND2_X1 U5072 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  AOI21_X1 U5073 ( .B1(n4578), .B2(ADDR_REG_12__SCAN_IN), .A(n4521), .ZN(n4525) );
  OAI211_X1 U5074 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4523), .A(n4580), .B(n4522), .ZN(n4524) );
  OAI211_X1 U5075 ( .C1(n4586), .C2(n4654), .A(n4525), .B(n4524), .ZN(U3252)
         );
  AOI21_X1 U5076 ( .B1(n3403), .B2(n4653), .A(n4526), .ZN(n4530) );
  OAI21_X1 U5077 ( .B1(n4530), .B2(n4529), .A(n4527), .ZN(n4528) );
  AOI21_X1 U5078 ( .B1(n4530), .B2(n4529), .A(n4528), .ZN(n4531) );
  AOI211_X1 U5079 ( .C1(n4578), .C2(ADDR_REG_13__SCAN_IN), .A(n4532), .B(n4531), .ZN(n4537) );
  OAI211_X1 U5080 ( .C1(n4535), .C2(n4534), .A(n4580), .B(n4533), .ZN(n4536)
         );
  OAI211_X1 U5081 ( .C1(n4586), .C2(n4653), .A(n4537), .B(n4536), .ZN(U3253)
         );
  INV_X1 U5082 ( .A(n4538), .ZN(n4542) );
  AOI211_X1 U5083 ( .C1(n2641), .C2(n4540), .A(n4539), .B(n4574), .ZN(n4541)
         );
  AOI211_X1 U5084 ( .C1(n4578), .C2(ADDR_REG_14__SCAN_IN), .A(n4542), .B(n4541), .ZN(n4546) );
  OAI211_X1 U5085 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4544), .A(n4580), .B(n4543), .ZN(n4545) );
  OAI211_X1 U5086 ( .C1(n4586), .C2(n4652), .A(n4546), .B(n4545), .ZN(U3254)
         );
  AOI211_X1 U5087 ( .C1(n2251), .C2(n4548), .A(n4547), .B(n4574), .ZN(n4549)
         );
  AOI211_X1 U5088 ( .C1(n4578), .C2(ADDR_REG_15__SCAN_IN), .A(n4550), .B(n4549), .ZN(n4555) );
  OAI211_X1 U5089 ( .C1(n4553), .C2(n4552), .A(n4580), .B(n4551), .ZN(n4554)
         );
  OAI211_X1 U5090 ( .C1(n4586), .C2(n4650), .A(n4555), .B(n4554), .ZN(U3255)
         );
  AOI221_X1 U5091 ( .B1(n4557), .B2(n4556), .C1(n4191), .C2(n4556), .A(n4574), 
        .ZN(n4558) );
  AOI211_X1 U5092 ( .C1(n4578), .C2(ADDR_REG_16__SCAN_IN), .A(n4559), .B(n4558), .ZN(n4563) );
  OAI221_X1 U5093 ( .B1(n4561), .B2(REG1_REG_16__SCAN_IN), .C1(n4561), .C2(
        n4560), .A(n4580), .ZN(n4562) );
  OAI211_X1 U5094 ( .C1(n4586), .C2(n4649), .A(n4563), .B(n4562), .ZN(U3256)
         );
  AOI221_X1 U5095 ( .B1(n4566), .B2(n4565), .C1(n4564), .C2(n4565), .A(n4574), 
        .ZN(n4567) );
  AOI211_X1 U5096 ( .C1(n4578), .C2(ADDR_REG_17__SCAN_IN), .A(n4568), .B(n4567), .ZN(n4572) );
  OAI221_X1 U5097 ( .B1(n4570), .B2(n2240), .C1(n4570), .C2(n4569), .A(n4580), 
        .ZN(n4571) );
  OAI211_X1 U5098 ( .C1(n4586), .C2(n4648), .A(n4572), .B(n4571), .ZN(U3257)
         );
  INV_X1 U5099 ( .A(n4573), .ZN(n4577) );
  OAI211_X1 U5100 ( .C1(n4582), .C2(n4581), .A(n4580), .B(n4579), .ZN(n4583)
         );
  OAI211_X1 U5101 ( .C1(n4586), .C2(n4585), .A(n4584), .B(n4583), .ZN(U3258)
         );
  XNOR2_X1 U5102 ( .A(n4587), .B(n4588), .ZN(n4703) );
  XNOR2_X1 U5103 ( .A(n4589), .B(n4588), .ZN(n4599) );
  OAI22_X1 U5104 ( .A1(n4593), .A2(n4592), .B1(n4591), .B2(n4590), .ZN(n4594)
         );
  AOI21_X1 U5105 ( .B1(n4596), .B2(n4595), .A(n4594), .ZN(n4597) );
  OAI21_X1 U5106 ( .B1(n4599), .B2(n4598), .A(n4597), .ZN(n4600) );
  AOI21_X1 U5107 ( .B1(n4601), .B2(n4703), .A(n4600), .ZN(n4705) );
  AOI22_X1 U5108 ( .A1(n4602), .A2(n4622), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4634), .ZN(n4607) );
  AOI21_X1 U5109 ( .B1(n4605), .B2(n4604), .A(n4603), .ZN(n4700) );
  AOI22_X1 U5110 ( .A1(n4703), .A2(n4631), .B1(n4629), .B2(n4700), .ZN(n4606)
         );
  OAI211_X1 U5111 ( .C1(n4634), .C2(n4705), .A(n4607), .B(n4606), .ZN(U3279)
         );
  OAI21_X1 U5112 ( .B1(n2307), .B2(n2306), .A(n4608), .ZN(n4620) );
  AOI22_X1 U5113 ( .A1(n4611), .A2(n4610), .B1(n4625), .B2(n4609), .ZN(n4612)
         );
  OAI21_X1 U5114 ( .B1(n2516), .B2(n4613), .A(n4612), .ZN(n4619) );
  OR2_X1 U5115 ( .A1(n2789), .A2(n4614), .ZN(n4615) );
  NAND2_X1 U5116 ( .A1(n4616), .A2(n4615), .ZN(n4670) );
  NOR2_X1 U5117 ( .A1(n4670), .A2(n4617), .ZN(n4618) );
  AOI211_X1 U5118 ( .C1(n4621), .C2(n4620), .A(n4619), .B(n4618), .ZN(n4667)
         );
  AOI22_X1 U5119 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4622), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4634), .ZN(n4633) );
  INV_X1 U5120 ( .A(n4670), .ZN(n4630) );
  INV_X1 U5121 ( .A(n4623), .ZN(n4627) );
  NAND2_X1 U5122 ( .A1(n4625), .A2(n4624), .ZN(n4626) );
  NAND2_X1 U5123 ( .A1(n4627), .A2(n4626), .ZN(n4668) );
  INV_X1 U5124 ( .A(n4668), .ZN(n4628) );
  AOI22_X1 U5125 ( .A1(n4631), .A2(n4630), .B1(n4629), .B2(n4628), .ZN(n4632)
         );
  OAI211_X1 U5126 ( .C1(n4634), .C2(n4667), .A(n4633), .B(n4632), .ZN(U3289)
         );
  INV_X1 U5127 ( .A(D_REG_31__SCAN_IN), .ZN(n4891) );
  NOR2_X1 U5128 ( .A1(n4643), .A2(n4891), .ZN(U3291) );
  INV_X1 U5129 ( .A(D_REG_30__SCAN_IN), .ZN(n4758) );
  NOR2_X1 U5130 ( .A1(n4643), .A2(n4758), .ZN(U3292) );
  INV_X1 U5131 ( .A(D_REG_29__SCAN_IN), .ZN(n4840) );
  NOR2_X1 U5132 ( .A1(n4643), .A2(n4840), .ZN(U3293) );
  INV_X1 U5133 ( .A(D_REG_28__SCAN_IN), .ZN(n5037) );
  NOR2_X1 U5134 ( .A1(n4643), .A2(n5037), .ZN(U3294) );
  INV_X1 U5135 ( .A(D_REG_27__SCAN_IN), .ZN(n4635) );
  NOR2_X1 U5136 ( .A1(n4643), .A2(n4635), .ZN(U3295) );
  INV_X1 U5137 ( .A(D_REG_26__SCAN_IN), .ZN(n4636) );
  NOR2_X1 U5138 ( .A1(n4643), .A2(n4636), .ZN(U3296) );
  INV_X1 U5139 ( .A(D_REG_25__SCAN_IN), .ZN(n5024) );
  NOR2_X1 U5140 ( .A1(n4643), .A2(n5024), .ZN(U3297) );
  INV_X1 U5141 ( .A(D_REG_24__SCAN_IN), .ZN(n4637) );
  NOR2_X1 U5142 ( .A1(n4643), .A2(n4637), .ZN(U3298) );
  INV_X1 U5143 ( .A(D_REG_23__SCAN_IN), .ZN(n5021) );
  NOR2_X1 U5144 ( .A1(n4643), .A2(n5021), .ZN(U3299) );
  INV_X1 U5145 ( .A(D_REG_22__SCAN_IN), .ZN(n4868) );
  NOR2_X1 U5146 ( .A1(n4643), .A2(n4868), .ZN(U3300) );
  INV_X1 U5147 ( .A(D_REG_21__SCAN_IN), .ZN(n5019) );
  NOR2_X1 U5148 ( .A1(n4643), .A2(n5019), .ZN(U3301) );
  INV_X1 U5149 ( .A(D_REG_20__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U5150 ( .A1(n4643), .A2(n4638), .ZN(U3302) );
  INV_X1 U5151 ( .A(D_REG_19__SCAN_IN), .ZN(n4639) );
  NOR2_X1 U5152 ( .A1(n4643), .A2(n4639), .ZN(U3303) );
  INV_X1 U5153 ( .A(D_REG_18__SCAN_IN), .ZN(n5041) );
  NOR2_X1 U5154 ( .A1(n4643), .A2(n5041), .ZN(U3304) );
  INV_X1 U5155 ( .A(D_REG_17__SCAN_IN), .ZN(n5018) );
  NOR2_X1 U5156 ( .A1(n4643), .A2(n5018), .ZN(U3305) );
  INV_X1 U5157 ( .A(D_REG_16__SCAN_IN), .ZN(n4887) );
  NOR2_X1 U5158 ( .A1(n4643), .A2(n4887), .ZN(U3306) );
  INV_X1 U5159 ( .A(D_REG_15__SCAN_IN), .ZN(n4855) );
  NOR2_X1 U5160 ( .A1(n4643), .A2(n4855), .ZN(U3307) );
  INV_X1 U5161 ( .A(D_REG_14__SCAN_IN), .ZN(n5040) );
  NOR2_X1 U5162 ( .A1(n4643), .A2(n5040), .ZN(U3308) );
  INV_X1 U5163 ( .A(D_REG_13__SCAN_IN), .ZN(n5022) );
  NOR2_X1 U5164 ( .A1(n4643), .A2(n5022), .ZN(U3309) );
  INV_X1 U5165 ( .A(D_REG_12__SCAN_IN), .ZN(n4640) );
  NOR2_X1 U5166 ( .A1(n4643), .A2(n4640), .ZN(U3310) );
  INV_X1 U5167 ( .A(D_REG_11__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U5168 ( .A1(n4643), .A2(n4844), .ZN(U3311) );
  INV_X1 U5169 ( .A(D_REG_10__SCAN_IN), .ZN(n4879) );
  NOR2_X1 U5170 ( .A1(n4643), .A2(n4879), .ZN(U3312) );
  INV_X1 U5171 ( .A(D_REG_9__SCAN_IN), .ZN(n4829) );
  NOR2_X1 U5172 ( .A1(n4643), .A2(n4829), .ZN(U3313) );
  INV_X1 U5173 ( .A(D_REG_8__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U5174 ( .A1(n4643), .A2(n4641), .ZN(U3314) );
  INV_X1 U5175 ( .A(D_REG_7__SCAN_IN), .ZN(n4642) );
  NOR2_X1 U5176 ( .A1(n4643), .A2(n4642), .ZN(U3315) );
  INV_X1 U5177 ( .A(D_REG_6__SCAN_IN), .ZN(n5043) );
  NOR2_X1 U5178 ( .A1(n4643), .A2(n5043), .ZN(U3316) );
  INV_X1 U5179 ( .A(D_REG_5__SCAN_IN), .ZN(n5044) );
  NOR2_X1 U5180 ( .A1(n4643), .A2(n5044), .ZN(U3317) );
  INV_X1 U5181 ( .A(D_REG_4__SCAN_IN), .ZN(n4818) );
  NOR2_X1 U5182 ( .A1(n4643), .A2(n4818), .ZN(U3318) );
  INV_X1 U5183 ( .A(D_REG_3__SCAN_IN), .ZN(n5038) );
  NOR2_X1 U5184 ( .A1(n4643), .A2(n5038), .ZN(U3319) );
  INV_X1 U5185 ( .A(D_REG_2__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U5186 ( .A1(n4643), .A2(n5025), .ZN(U3320) );
  INV_X1 U5187 ( .A(DATAI_23_), .ZN(n5046) );
  AOI21_X1 U5188 ( .B1(U3149), .B2(n5046), .A(n4644), .ZN(U3329) );
  OAI22_X1 U5189 ( .A1(U3149), .A2(n4645), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4646) );
  INV_X1 U5190 ( .A(n4646), .ZN(U3334) );
  INV_X1 U5191 ( .A(DATAI_17_), .ZN(n4647) );
  AOI22_X1 U5192 ( .A1(STATE_REG_SCAN_IN), .A2(n4648), .B1(n4647), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5193 ( .A(DATAI_16_), .ZN(n4843) );
  AOI22_X1 U5194 ( .A1(STATE_REG_SCAN_IN), .A2(n4649), .B1(n4843), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5195 ( .A(DATAI_15_), .ZN(n4828) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n4650), .B1(n4828), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5197 ( .A(DATAI_14_), .ZN(n4651) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4652), .B1(n4651), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5199 ( .A1(STATE_REG_SCAN_IN), .A2(n4653), .B1(n2637), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5200 ( .A1(STATE_REG_SCAN_IN), .A2(n4654), .B1(n5082), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5201 ( .A(DATAI_11_), .ZN(n4805) );
  AOI22_X1 U5202 ( .A1(STATE_REG_SCAN_IN), .A2(n4655), .B1(n4805), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5203 ( .A(DATAI_10_), .ZN(n4656) );
  AOI22_X1 U5204 ( .A1(STATE_REG_SCAN_IN), .A2(n2377), .B1(n4656), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5205 ( .A(DATAI_9_), .ZN(n4876) );
  AOI22_X1 U5206 ( .A1(STATE_REG_SCAN_IN), .A2(n4657), .B1(n4876), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5207 ( .A(DATAI_8_), .ZN(n4867) );
  AOI22_X1 U5208 ( .A1(STATE_REG_SCAN_IN), .A2(n2378), .B1(n4867), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5209 ( .A(DATAI_7_), .ZN(n4658) );
  AOI22_X1 U5210 ( .A1(STATE_REG_SCAN_IN), .A2(n4659), .B1(n4658), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5211 ( .A(DATAI_6_), .ZN(n4660) );
  AOI22_X1 U5212 ( .A1(STATE_REG_SCAN_IN), .A2(n4661), .B1(n4660), .B2(U3149), 
        .ZN(U3346) );
  INV_X1 U5213 ( .A(DATAI_5_), .ZN(n5081) );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(n4662), .B1(n5081), .B2(U3149), 
        .ZN(U3347) );
  OAI211_X1 U5215 ( .C1(n4665), .C2(n4669), .A(n4664), .B(n4663), .ZN(n4666)
         );
  INV_X1 U5216 ( .A(n4666), .ZN(n4710) );
  INV_X1 U5217 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U5218 ( .A1(n4708), .A2(n4710), .B1(n4996), .B2(n4706), .ZN(U3467)
         );
  INV_X1 U5219 ( .A(n4667), .ZN(n4672) );
  OAI22_X1 U5220 ( .A1(n4670), .A2(n4669), .B1(n4693), .B2(n4668), .ZN(n4671)
         );
  NOR2_X1 U5221 ( .A1(n4672), .A2(n4671), .ZN(n4712) );
  INV_X1 U5222 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5223 ( .A1(n4708), .A2(n4712), .B1(n4673), .B2(n4706), .ZN(U3469)
         );
  AOI21_X1 U5224 ( .B1(n4702), .B2(n4675), .A(n4674), .ZN(n4717) );
  INV_X1 U5225 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4676) );
  OAI22_X1 U5226 ( .A1(n4677), .A2(n4713), .B1(n4708), .B2(n4676), .ZN(n4678)
         );
  INV_X1 U5227 ( .A(n4678), .ZN(n4679) );
  OAI21_X1 U5228 ( .B1(n4717), .B2(n4706), .A(n4679), .ZN(U3471) );
  INV_X1 U5229 ( .A(n4680), .ZN(n4682) );
  AOI211_X1 U5230 ( .C1(n4683), .C2(n4702), .A(n4682), .B(n4681), .ZN(n4719)
         );
  INV_X1 U5231 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4998) );
  AOI22_X1 U5232 ( .A1(n4708), .A2(n4719), .B1(n4998), .B2(n4706), .ZN(U3475)
         );
  AOI211_X1 U5233 ( .C1(n4687), .C2(n4686), .A(n4685), .B(n4684), .ZN(n4721)
         );
  INV_X1 U5234 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5235 ( .A1(n4708), .A2(n4721), .B1(n4781), .B2(n4706), .ZN(U3481)
         );
  NOR3_X1 U5236 ( .A1(n4689), .A2(n4688), .A3(n4693), .ZN(n4691) );
  AOI211_X1 U5237 ( .C1(n4692), .C2(n4702), .A(n4691), .B(n4690), .ZN(n4723)
         );
  INV_X1 U5238 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5005) );
  AOI22_X1 U5239 ( .A1(n4708), .A2(n4723), .B1(n5005), .B2(n4706), .ZN(U3483)
         );
  NOR3_X1 U5240 ( .A1(n4695), .A2(n4694), .A3(n4693), .ZN(n4697) );
  AOI211_X1 U5241 ( .C1(n4698), .C2(n4702), .A(n4697), .B(n4696), .ZN(n4725)
         );
  INV_X1 U5242 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U5243 ( .A1(n4708), .A2(n4725), .B1(n4699), .B2(n4706), .ZN(U3487)
         );
  AOI22_X1 U5244 ( .A1(n4703), .A2(n4702), .B1(n4701), .B2(n4700), .ZN(n4704)
         );
  AND2_X1 U5245 ( .A1(n4705), .A2(n4704), .ZN(n4728) );
  INV_X1 U5246 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5247 ( .A1(n4708), .A2(n4728), .B1(n4707), .B2(n4706), .ZN(U3489)
         );
  AOI22_X1 U5248 ( .A1(n4729), .A2(n4710), .B1(n4709), .B2(n4726), .ZN(U3518)
         );
  INV_X1 U5249 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5250 ( .A1(n4729), .A2(n4712), .B1(n4711), .B2(n4726), .ZN(U3519)
         );
  OAI22_X1 U5251 ( .A1(n4714), .A2(n4713), .B1(n4729), .B2(n2893), .ZN(n4715)
         );
  INV_X1 U5252 ( .A(n4715), .ZN(n4716) );
  OAI21_X1 U5253 ( .B1(n4717), .B2(n4726), .A(n4716), .ZN(U3520) );
  AOI22_X1 U5254 ( .A1(n4729), .A2(n4719), .B1(n4718), .B2(n4726), .ZN(U3522)
         );
  INV_X1 U5255 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4720) );
  AOI22_X1 U5256 ( .A1(n4729), .A2(n4721), .B1(n4720), .B2(n4726), .ZN(U3525)
         );
  INV_X1 U5257 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5258 ( .A1(n4729), .A2(n4723), .B1(n4722), .B2(n4726), .ZN(U3526)
         );
  INV_X1 U5259 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4724) );
  AOI22_X1 U5260 ( .A1(n4729), .A2(n4725), .B1(n4724), .B2(n4726), .ZN(U3528)
         );
  AOI22_X1 U5261 ( .A1(n4729), .A2(n4728), .B1(n4727), .B2(n4726), .ZN(U3529)
         );
  OAI22_X1 U5262 ( .A1(IR_REG_10__SCAN_IN), .A2(keyinput_g65), .B1(
        keyinput_g120), .B2(REG0_REG_1__SCAN_IN), .ZN(n4730) );
  AOI221_X1 U5263 ( .B1(IR_REG_10__SCAN_IN), .B2(keyinput_g65), .C1(
        REG0_REG_1__SCAN_IN), .C2(keyinput_g120), .A(n4730), .ZN(n4737) );
  OAI22_X1 U5264 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_g57), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .ZN(n4731) );
  AOI221_X1 U5265 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g50), .C2(REG3_REG_4__SCAN_IN), .A(n4731), .ZN(n4736) );
  OAI22_X1 U5266 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_g82), .B1(
        keyinput_g54), .B2(REG3_REG_13__SCAN_IN), .ZN(n4732) );
  AOI221_X1 U5267 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_g82), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_g54), .A(n4732), .ZN(n4735) );
  OAI22_X1 U5268 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput_g90), .B1(
        D_REG_18__SCAN_IN), .B2(keyinput_g105), .ZN(n4733) );
  AOI221_X1 U5269 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput_g90), .C1(
        keyinput_g105), .C2(D_REG_18__SCAN_IN), .A(n4733), .ZN(n4734) );
  NAND4_X1 U5270 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4766)
         );
  OAI22_X1 U5271 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput_g106), .B1(
        keyinput_g40), .B2(REG3_REG_28__SCAN_IN), .ZN(n4738) );
  AOI221_X1 U5272 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput_g106), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_g40), .A(n4738), .ZN(n4745) );
  OAI22_X1 U5273 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput_g99), .B1(DATAI_6_), 
        .B2(keyinput_g25), .ZN(n4739) );
  AOI221_X1 U5274 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput_g99), .C1(
        keyinput_g25), .C2(DATAI_6_), .A(n4739), .ZN(n4744) );
  OAI22_X1 U5275 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_g89), .B1(keyinput_g51), 
        .B2(REG3_REG_9__SCAN_IN), .ZN(n4740) );
  AOI221_X1 U5276 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_g89), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_g51), .A(n4740), .ZN(n4743) );
  OAI22_X1 U5277 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_g112), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput_g100), .ZN(n4741) );
  AOI221_X1 U5278 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g100), .C2(D_REG_13__SCAN_IN), .A(n4741), .ZN(n4742) );
  NAND4_X1 U5279 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4765)
         );
  OAI22_X1 U5280 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(keyinput_g7), .B2(
        DATAI_24_), .ZN(n4746) );
  AOI221_X1 U5281 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_24_), .C2(
        keyinput_g7), .A(n4746), .ZN(n4753) );
  OAI22_X1 U5282 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput_g94), .B1(
        REG0_REG_0__SCAN_IN), .B2(keyinput_g119), .ZN(n4747) );
  AOI221_X1 U5283 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g119), .C2(REG0_REG_0__SCAN_IN), .A(n4747), .ZN(n4752) );
  OAI22_X1 U5284 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_g66), .B1(
        keyinput_g61), .B2(IR_REG_6__SCAN_IN), .ZN(n4748) );
  AOI221_X1 U5285 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput_g66), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n4748), .ZN(n4751) );
  OAI22_X1 U5286 ( .A1(IR_REG_29__SCAN_IN), .A2(keyinput_g84), .B1(DATAI_3_), 
        .B2(keyinput_g28), .ZN(n4749) );
  AOI221_X1 U5287 ( .B1(IR_REG_29__SCAN_IN), .B2(keyinput_g84), .C1(
        keyinput_g28), .C2(DATAI_3_), .A(n4749), .ZN(n4750) );
  NAND4_X1 U5288 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4764)
         );
  OAI22_X1 U5289 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput_g113), .B1(
        keyinput_g47), .B2(REG3_REG_5__SCAN_IN), .ZN(n4754) );
  AOI221_X1 U5290 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput_g113), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_g47), .A(n4754), .ZN(n4762) );
  OAI22_X1 U5291 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_g86), .B1(DATAI_10_), 
        .B2(keyinput_g21), .ZN(n4755) );
  AOI221_X1 U5292 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g21), .C2(DATAI_10_), .A(n4755), .ZN(n4761) );
  OAI22_X1 U5293 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g124), .B2(REG0_REG_5__SCAN_IN), .ZN(n4756) );
  AOI221_X1 U5294 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput_g110), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput_g124), .A(n4756), .ZN(n4760) );
  OAI22_X1 U5295 ( .A1(n4758), .A2(keyinput_g117), .B1(keyinput_g87), .B2(
        D_REG_0__SCAN_IN), .ZN(n4757) );
  AOI221_X1 U5296 ( .B1(n4758), .B2(keyinput_g117), .C1(D_REG_0__SCAN_IN), 
        .C2(keyinput_g87), .A(n4757), .ZN(n4759) );
  NAND4_X1 U5297 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4763)
         );
  NOR4_X1 U5298 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n5107)
         );
  OAI22_X1 U5299 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g75), .B2(IR_REG_20__SCAN_IN), .ZN(n4767) );
  AOI221_X1 U5300 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_g79), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_g75), .A(n4767), .ZN(n4774) );
  OAI22_X1 U5301 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_g52), .B1(DATAI_30_), 
        .B2(keyinput_g1), .ZN(n4768) );
  AOI221_X1 U5302 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g1), .C2(DATAI_30_), .A(n4768), .ZN(n4773) );
  OAI22_X1 U5303 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_g35), .B1(
        keyinput_g13), .B2(DATAI_18_), .ZN(n4769) );
  AOI221_X1 U5304 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_g35), .C1(
        DATAI_18_), .C2(keyinput_g13), .A(n4769), .ZN(n4772) );
  OAI22_X1 U5305 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput_g114), .B1(
        D_REG_24__SCAN_IN), .B2(keyinput_g111), .ZN(n4770) );
  AOI221_X1 U5306 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g111), .C2(D_REG_24__SCAN_IN), .A(n4770), .ZN(n4771) );
  NAND4_X1 U5307 ( .A1(n4774), .A2(n4773), .A3(n4772), .A4(n4771), .ZN(n4905)
         );
  OAI22_X1 U5308 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(DATAI_17_), .B2(
        keyinput_g14), .ZN(n4775) );
  AOI221_X1 U5309 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(keyinput_g14), .C2(
        DATAI_17_), .A(n4775), .ZN(n4801) );
  OAI22_X1 U5310 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(keyinput_g24), .B2(
        DATAI_7_), .ZN(n4776) );
  AOI221_X1 U5311 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(DATAI_7_), .C2(
        keyinput_g24), .A(n4776), .ZN(n4779) );
  OAI22_X1 U5312 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_g48), .B1(DATAI_14_), .B2(keyinput_g17), .ZN(n4777) );
  AOI221_X1 U5313 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .C1(
        keyinput_g17), .C2(DATAI_14_), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5314 ( .C1(n4781), .C2(keyinput_g126), .A(n4779), .B(n4778), .ZN(
        n4780) );
  AOI21_X1 U5315 ( .B1(n4781), .B2(keyinput_g126), .A(n4780), .ZN(n4800) );
  AOI22_X1 U5316 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput_g95), .B1(
        D_REG_20__SCAN_IN), .B2(keyinput_g107), .ZN(n4782) );
  OAI221_X1 U5317 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput_g95), .C1(
        D_REG_20__SCAN_IN), .C2(keyinput_g107), .A(n4782), .ZN(n4789) );
  AOI22_X1 U5318 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput_g56), .ZN(n4783) );
  OAI221_X1 U5319 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput_g56), .A(n4783), .ZN(n4788) );
  AOI22_X1 U5320 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_g58), .ZN(n4784) );
  OAI221_X1 U5321 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_g58), .A(n4784), .ZN(n4787) );
  AOI22_X1 U5322 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput_g83), .B1(
        D_REG_1__SCAN_IN), .B2(keyinput_g88), .ZN(n4785) );
  OAI221_X1 U5323 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput_g83), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput_g88), .A(n4785), .ZN(n4786) );
  NOR4_X1 U5324 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4799)
         );
  AOI22_X1 U5325 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_g104), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput_g93), .ZN(n4790) );
  OAI221_X1 U5326 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_g104), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput_g93), .A(n4790), .ZN(n4797) );
  AOI22_X1 U5327 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(DATAI_23_), .B2(
        keyinput_g8), .ZN(n4791) );
  OAI221_X1 U5328 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(DATAI_23_), .C2(
        keyinput_g8), .A(n4791), .ZN(n4796) );
  AOI22_X1 U5329 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(REG3_REG_12__SCAN_IN), 
        .B2(keyinput_g44), .ZN(n4792) );
  OAI221_X1 U5330 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(REG3_REG_12__SCAN_IN), .C2(keyinput_g44), .A(n4792), .ZN(n4795) );
  AOI22_X1 U5331 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput_g76), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput_g78), .ZN(n4793) );
  OAI221_X1 U5332 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput_g76), .C1(
        IR_REG_23__SCAN_IN), .C2(keyinput_g78), .A(n4793), .ZN(n4794) );
  NOR4_X1 U5333 ( .A1(n4797), .A2(n4796), .A3(n4795), .A4(n4794), .ZN(n4798)
         );
  NAND4_X1 U5334 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4904)
         );
  INV_X1 U5335 ( .A(DATAI_25_), .ZN(n4956) );
  AOI22_X1 U5336 ( .A1(n4803), .A2(keyinput_g46), .B1(keyinput_g6), .B2(n4956), 
        .ZN(n4802) );
  OAI221_X1 U5337 ( .B1(n4803), .B2(keyinput_g46), .C1(n4956), .C2(keyinput_g6), .A(n4802), .ZN(n4814) );
  AOI22_X1 U5338 ( .A1(n5044), .A2(keyinput_g92), .B1(keyinput_g20), .B2(n4805), .ZN(n4804) );
  OAI221_X1 U5339 ( .B1(n5044), .B2(keyinput_g92), .C1(n4805), .C2(
        keyinput_g20), .A(n4804), .ZN(n4813) );
  INV_X1 U5340 ( .A(DATAI_4_), .ZN(n4807) );
  AOI22_X1 U5341 ( .A1(n4808), .A2(keyinput_g49), .B1(keyinput_g27), .B2(n4807), .ZN(n4806) );
  OAI221_X1 U5342 ( .B1(n4808), .B2(keyinput_g49), .C1(n4807), .C2(
        keyinput_g27), .A(n4806), .ZN(n4812) );
  XOR2_X1 U5343 ( .A(n2781), .B(keyinput_g74), .Z(n4810) );
  XNOR2_X1 U5344 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_g60), .ZN(n4809) );
  NAND2_X1 U5345 ( .A1(n4810), .A2(n4809), .ZN(n4811) );
  NOR4_X1 U5346 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4853)
         );
  AOI22_X1 U5347 ( .A1(n2277), .A2(keyinput_g55), .B1(keyinput_g36), .B2(n4816), .ZN(n4815) );
  OAI221_X1 U5348 ( .B1(n2277), .B2(keyinput_g55), .C1(n4816), .C2(
        keyinput_g36), .A(n4815), .ZN(n4826) );
  AOI22_X1 U5349 ( .A1(n4985), .A2(keyinput_g2), .B1(n4818), .B2(keyinput_g91), 
        .ZN(n4817) );
  OAI221_X1 U5350 ( .B1(n4985), .B2(keyinput_g2), .C1(n4818), .C2(keyinput_g91), .A(n4817), .ZN(n4825) );
  AOI22_X1 U5351 ( .A1(n4820), .A2(keyinput_g37), .B1(keyinput_g19), .B2(n5082), .ZN(n4819) );
  OAI221_X1 U5352 ( .B1(n4820), .B2(keyinput_g37), .C1(n5082), .C2(
        keyinput_g19), .A(n4819), .ZN(n4824) );
  XNOR2_X1 U5353 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_g62), .ZN(n4822) );
  XNOR2_X1 U5354 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_g41), .ZN(n4821) );
  NAND2_X1 U5355 ( .A1(n4822), .A2(n4821), .ZN(n4823) );
  NOR4_X1 U5356 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n4852)
         );
  AOI22_X1 U5357 ( .A1(n4829), .A2(keyinput_g96), .B1(keyinput_g16), .B2(n4828), .ZN(n4827) );
  OAI221_X1 U5358 ( .B1(n4829), .B2(keyinput_g96), .C1(n4828), .C2(
        keyinput_g16), .A(n4827), .ZN(n4838) );
  INV_X1 U5359 ( .A(IR_REG_16__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U5360 ( .A1(n2519), .A2(keyinput_g38), .B1(n4831), .B2(keyinput_g71), .ZN(n4830) );
  OAI221_X1 U5361 ( .B1(n2519), .B2(keyinput_g38), .C1(n4831), .C2(
        keyinput_g71), .A(n4830), .ZN(n4837) );
  INV_X1 U5362 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4999) );
  XOR2_X1 U5363 ( .A(n4999), .B(keyinput_g122), .Z(n4835) );
  XNOR2_X1 U5364 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_g63), .ZN(n4834) );
  XNOR2_X1 U5365 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_g53), .ZN(n4833) );
  XNOR2_X1 U5366 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_g59), .ZN(n4832) );
  NAND4_X1 U5367 ( .A1(n4835), .A2(n4834), .A3(n4833), .A4(n4832), .ZN(n4836)
         );
  NOR3_X1 U5368 ( .A1(n4838), .A2(n4837), .A3(n4836), .ZN(n4851) );
  AOI22_X1 U5369 ( .A1(n3580), .A2(keyinput_g43), .B1(n4840), .B2(
        keyinput_g116), .ZN(n4839) );
  OAI221_X1 U5370 ( .B1(n3580), .B2(keyinput_g43), .C1(n4840), .C2(
        keyinput_g116), .A(n4839), .ZN(n4849) );
  INV_X1 U5371 ( .A(DATAI_0_), .ZN(n5070) );
  AOI22_X1 U5372 ( .A1(n4676), .A2(keyinput_g121), .B1(keyinput_g31), .B2(
        n5070), .ZN(n4841) );
  OAI221_X1 U5373 ( .B1(n4676), .B2(keyinput_g121), .C1(n5070), .C2(
        keyinput_g31), .A(n4841), .ZN(n4848) );
  AOI22_X1 U5374 ( .A1(n4844), .A2(keyinput_g98), .B1(keyinput_g15), .B2(n4843), .ZN(n4842) );
  OAI221_X1 U5375 ( .B1(n4844), .B2(keyinput_g98), .C1(n4843), .C2(
        keyinput_g15), .A(n4842), .ZN(n4847) );
  INV_X1 U5376 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5008) );
  AOI22_X1 U5377 ( .A1(n5008), .A2(keyinput_g125), .B1(n5019), .B2(
        keyinput_g108), .ZN(n4845) );
  OAI221_X1 U5378 ( .B1(n5008), .B2(keyinput_g125), .C1(n5019), .C2(
        keyinput_g108), .A(n4845), .ZN(n4846) );
  NOR4_X1 U5379 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4850)
         );
  NAND4_X1 U5380 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4903)
         );
  AOI22_X1 U5381 ( .A1(n2455), .A2(keyinput_g69), .B1(keyinput_g102), .B2(
        n4855), .ZN(n4854) );
  OAI221_X1 U5382 ( .B1(n2455), .B2(keyinput_g69), .C1(n4855), .C2(
        keyinput_g102), .A(n4854), .ZN(n4863) );
  INV_X1 U5383 ( .A(REG3_REG_19__SCAN_IN), .ZN(n5068) );
  AOI22_X1 U5384 ( .A1(n2971), .A2(keyinput_g42), .B1(n5068), .B2(keyinput_g39), .ZN(n4856) );
  OAI221_X1 U5385 ( .B1(n2971), .B2(keyinput_g42), .C1(n5068), .C2(
        keyinput_g39), .A(n4856), .ZN(n4862) );
  XOR2_X1 U5386 ( .A(n5005), .B(keyinput_g127), .Z(n4860) );
  XNOR2_X1 U5387 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_g77), .ZN(n4859) );
  XNOR2_X1 U5388 ( .A(DATAI_2_), .B(keyinput_g29), .ZN(n4858) );
  XNOR2_X1 U5389 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_g68), .ZN(n4857) );
  NAND4_X1 U5390 ( .A1(n4860), .A2(n4859), .A3(n4858), .A4(n4857), .ZN(n4861)
         );
  NOR3_X1 U5391 ( .A1(n4863), .A2(n4862), .A3(n4861), .ZN(n4901) );
  AOI22_X1 U5392 ( .A1(U3149), .A2(keyinput_g32), .B1(n2689), .B2(keyinput_g72), .ZN(n4864) );
  OAI221_X1 U5393 ( .B1(U3149), .B2(keyinput_g32), .C1(n2689), .C2(
        keyinput_g72), .A(n4864), .ZN(n4874) );
  INV_X1 U5394 ( .A(DATAI_26_), .ZN(n5058) );
  AOI22_X1 U5395 ( .A1(n4986), .A2(keyinput_g0), .B1(n5058), .B2(keyinput_g5), 
        .ZN(n4865) );
  OAI221_X1 U5396 ( .B1(n4986), .B2(keyinput_g0), .C1(n5058), .C2(keyinput_g5), 
        .A(n4865), .ZN(n4873) );
  AOI22_X1 U5397 ( .A1(n4868), .A2(keyinput_g109), .B1(keyinput_g23), .B2(
        n4867), .ZN(n4866) );
  OAI221_X1 U5398 ( .B1(n4868), .B2(keyinput_g109), .C1(n4867), .C2(
        keyinput_g23), .A(n4866), .ZN(n4872) );
  XOR2_X1 U5399 ( .A(n2637), .B(keyinput_g18), .Z(n4870) );
  XNOR2_X1 U5400 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_g67), .ZN(n4869) );
  NAND2_X1 U5401 ( .A1(n4870), .A2(n4869), .ZN(n4871) );
  NOR4_X1 U5402 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(n4900)
         );
  INV_X1 U5403 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4980) );
  AOI22_X1 U5404 ( .A1(n4980), .A2(keyinput_g34), .B1(keyinput_g22), .B2(n4876), .ZN(n4875) );
  OAI221_X1 U5405 ( .B1(n4980), .B2(keyinput_g34), .C1(n4876), .C2(
        keyinput_g22), .A(n4875), .ZN(n4885) );
  AOI22_X1 U5406 ( .A1(n5037), .A2(keyinput_g115), .B1(keyinput_g10), .B2(
        n5055), .ZN(n4877) );
  OAI221_X1 U5407 ( .B1(n5037), .B2(keyinput_g115), .C1(n5055), .C2(
        keyinput_g10), .A(n4877), .ZN(n4884) );
  AOI22_X1 U5408 ( .A1(n4998), .A2(keyinput_g123), .B1(n4879), .B2(
        keyinput_g97), .ZN(n4878) );
  OAI221_X1 U5409 ( .B1(n4998), .B2(keyinput_g123), .C1(n4879), .C2(
        keyinput_g97), .A(n4878), .ZN(n4883) );
  XOR2_X1 U5410 ( .A(n2467), .B(keyinput_g64), .Z(n4881) );
  XNOR2_X1 U5411 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_g80), .ZN(n4880) );
  NAND2_X1 U5412 ( .A1(n4881), .A2(n4880), .ZN(n4882) );
  NOR4_X1 U5413 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n4899)
         );
  AOI22_X1 U5414 ( .A1(n2665), .A2(keyinput_g70), .B1(keyinput_g103), .B2(
        n4887), .ZN(n4886) );
  OAI221_X1 U5415 ( .B1(n2665), .B2(keyinput_g70), .C1(n4887), .C2(
        keyinput_g103), .A(n4886), .ZN(n4897) );
  INV_X1 U5416 ( .A(DATAI_22_), .ZN(n4889) );
  AOI22_X1 U5417 ( .A1(n4889), .A2(keyinput_g9), .B1(n5052), .B2(keyinput_g4), 
        .ZN(n4888) );
  OAI221_X1 U5418 ( .B1(n4889), .B2(keyinput_g9), .C1(n5052), .C2(keyinput_g4), 
        .A(n4888), .ZN(n4896) );
  AOI22_X1 U5419 ( .A1(n5040), .A2(keyinput_g101), .B1(n4891), .B2(
        keyinput_g118), .ZN(n4890) );
  OAI221_X1 U5420 ( .B1(n5040), .B2(keyinput_g101), .C1(n4891), .C2(
        keyinput_g118), .A(n4890), .ZN(n4895) );
  XNOR2_X1 U5421 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_g81), .ZN(n4893) );
  XNOR2_X1 U5422 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4892) );
  NAND2_X1 U5423 ( .A1(n4893), .A2(n4892), .ZN(n4894) );
  NOR4_X1 U5424 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4898)
         );
  NAND4_X1 U5425 ( .A1(n4901), .A2(n4900), .A3(n4899), .A4(n4898), .ZN(n4902)
         );
  NOR4_X1 U5426 ( .A1(n4905), .A2(n4904), .A3(n4903), .A4(n4902), .ZN(n5106)
         );
  OAI22_X1 U5427 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(keyinput_f57), .B2(IR_REG_2__SCAN_IN), .ZN(n4906) );
  AOI221_X1 U5428 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_f57), .A(n4906), .ZN(n4913) );
  OAI22_X1 U5429 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f126), .B2(REG0_REG_7__SCAN_IN), .ZN(n4907) );
  AOI221_X1 U5430 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_f62), .C1(
        REG0_REG_7__SCAN_IN), .C2(keyinput_f126), .A(n4907), .ZN(n4912) );
  OAI22_X1 U5431 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(keyinput_f22), .B2(
        DATAI_9_), .ZN(n4908) );
  AOI221_X1 U5432 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(DATAI_9_), .C2(
        keyinput_f22), .A(n4908), .ZN(n4911) );
  OAI22_X1 U5433 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_f88), .B1(keyinput_f82), 
        .B2(IR_REG_27__SCAN_IN), .ZN(n4909) );
  AOI221_X1 U5434 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_f88), .C1(
        IR_REG_27__SCAN_IN), .C2(keyinput_f82), .A(n4909), .ZN(n4910) );
  NAND4_X1 U5435 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4941)
         );
  OAI22_X1 U5436 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_f73), .B1(
        D_REG_15__SCAN_IN), .B2(keyinput_f102), .ZN(n4914) );
  AOI221_X1 U5437 ( .B1(IR_REG_18__SCAN_IN), .B2(keyinput_f73), .C1(
        keyinput_f102), .C2(D_REG_15__SCAN_IN), .A(n4914), .ZN(n4921) );
  OAI22_X1 U5438 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_f91), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n4915) );
  AOI221_X1 U5439 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_f91), .C1(
        keyinput_f117), .C2(D_REG_30__SCAN_IN), .A(n4915), .ZN(n4920) );
  OAI22_X1 U5440 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput_f98), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput_f116), .ZN(n4916) );
  AOI221_X1 U5441 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput_f98), .C1(
        keyinput_f116), .C2(D_REG_29__SCAN_IN), .A(n4916), .ZN(n4919) );
  OAI22_X1 U5442 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_f96), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput_f103), .ZN(n4917) );
  AOI221_X1 U5443 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput_f96), .C1(
        keyinput_f103), .C2(D_REG_16__SCAN_IN), .A(n4917), .ZN(n4918) );
  NAND4_X1 U5444 ( .A1(n4921), .A2(n4920), .A3(n4919), .A4(n4918), .ZN(n4940)
         );
  OAI22_X1 U5445 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_f109), .B1(
        D_REG_10__SCAN_IN), .B2(keyinput_f97), .ZN(n4922) );
  AOI221_X1 U5446 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_f109), .C1(
        keyinput_f97), .C2(D_REG_10__SCAN_IN), .A(n4922), .ZN(n4929) );
  OAI22_X1 U5447 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput_f118), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput_f87), .ZN(n4923) );
  AOI221_X1 U5448 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput_f118), .C1(
        keyinput_f87), .C2(D_REG_0__SCAN_IN), .A(n4923), .ZN(n4928) );
  OAI22_X1 U5449 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput_f76), .B1(
        keyinput_f15), .B2(DATAI_16_), .ZN(n4924) );
  AOI221_X1 U5450 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput_f76), .C1(DATAI_16_), 
        .C2(keyinput_f15), .A(n4924), .ZN(n4927) );
  OAI22_X1 U5451 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_f36), .B1(
        keyinput_f16), .B2(DATAI_15_), .ZN(n4925) );
  AOI221_X1 U5452 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .C1(
        DATAI_15_), .C2(keyinput_f16), .A(n4925), .ZN(n4926) );
  NAND4_X1 U5453 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .ZN(n4939)
         );
  OAI22_X1 U5454 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(DATAI_11_), .B2(keyinput_f20), .ZN(n4930) );
  AOI221_X1 U5455 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(
        keyinput_f20), .C2(DATAI_11_), .A(n4930), .ZN(n4937) );
  OAI22_X1 U5456 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_f79), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_f37), .ZN(n4931) );
  AOI221_X1 U5457 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_f79), .C1(
        keyinput_f37), .C2(REG3_REG_10__SCAN_IN), .A(n4931), .ZN(n4936) );
  OAI22_X1 U5458 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput_f68), .B1(
        keyinput_f60), .B2(IR_REG_5__SCAN_IN), .ZN(n4932) );
  AOI221_X1 U5459 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput_f68), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_f60), .A(n4932), .ZN(n4935) );
  OAI22_X1 U5460 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_f67), .B1(DATAI_8_), 
        .B2(keyinput_f23), .ZN(n4933) );
  AOI221_X1 U5461 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_f67), .C1(
        keyinput_f23), .C2(DATAI_8_), .A(n4933), .ZN(n4934) );
  NAND4_X1 U5462 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(n4938)
         );
  NOR4_X1 U5463 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n5100)
         );
  OAI22_X1 U5464 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(DATAI_18_), .B2(
        keyinput_f13), .ZN(n4942) );
  AOI221_X1 U5465 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(keyinput_f13), .C2(
        DATAI_18_), .A(n4942), .ZN(n4949) );
  OAI22_X1 U5466 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(REG3_REG_1__SCAN_IN), 
        .B2(keyinput_f42), .ZN(n4943) );
  AOI221_X1 U5467 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(keyinput_f42), .C2(
        REG3_REG_1__SCAN_IN), .A(n4943), .ZN(n4948) );
  OAI22_X1 U5468 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_f48), .B1(
        keyinput_f47), .B2(REG3_REG_5__SCAN_IN), .ZN(n4944) );
  AOI221_X1 U5469 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_f48), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_f47), .A(n4944), .ZN(n4947) );
  OAI22_X1 U5470 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput_f114), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput_f113), .ZN(n4945) );
  AOI221_X1 U5471 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput_f114), .C1(
        keyinput_f113), .C2(D_REG_26__SCAN_IN), .A(n4945), .ZN(n4946) );
  NAND4_X1 U5472 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n5098)
         );
  OAI22_X1 U5473 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_f32), .B1(DATAI_19_), 
        .B2(keyinput_f12), .ZN(n4950) );
  AOI221_X1 U5474 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        keyinput_f12), .C2(DATAI_19_), .A(n4950), .ZN(n4976) );
  OAI22_X1 U5475 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_f49), .B1(DATAI_30_), .B2(keyinput_f1), .ZN(n4951) );
  AOI221_X1 U5476 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_f49), .C1(
        keyinput_f1), .C2(DATAI_30_), .A(n4951), .ZN(n4954) );
  OAI22_X1 U5477 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_f40), .B1(
        keyinput_f11), .B2(DATAI_20_), .ZN(n4952) );
  AOI221_X1 U5478 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .C1(
        DATAI_20_), .C2(keyinput_f11), .A(n4952), .ZN(n4953) );
  OAI211_X1 U5479 ( .C1(n4956), .C2(keyinput_f6), .A(n4954), .B(n4953), .ZN(
        n4955) );
  AOI21_X1 U5480 ( .B1(n4956), .B2(keyinput_f6), .A(n4955), .ZN(n4975) );
  AOI22_X1 U5481 ( .A1(D_REG_20__SCAN_IN), .A2(keyinput_f107), .B1(
        D_REG_24__SCAN_IN), .B2(keyinput_f111), .ZN(n4957) );
  OAI221_X1 U5482 ( .B1(D_REG_20__SCAN_IN), .B2(keyinput_f107), .C1(
        D_REG_24__SCAN_IN), .C2(keyinput_f111), .A(n4957), .ZN(n4964) );
  AOI22_X1 U5483 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput_f99), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput_f106), .ZN(n4958) );
  OAI221_X1 U5484 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput_f99), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput_f106), .A(n4958), .ZN(n4963) );
  AOI22_X1 U5485 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput_f94), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput_f95), .ZN(n4959) );
  OAI221_X1 U5486 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput_f94), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput_f95), .A(n4959), .ZN(n4962) );
  AOI22_X1 U5487 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput_f69), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput_f86), .ZN(n4960) );
  OAI221_X1 U5488 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput_f69), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput_f86), .A(n4960), .ZN(n4961) );
  NOR4_X1 U5489 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n4974)
         );
  AOI22_X1 U5490 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_f70), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput_f71), .ZN(n4965) );
  OAI221_X1 U5491 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_f70), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput_f71), .A(n4965), .ZN(n4972) );
  AOI22_X1 U5492 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n4966) );
  OAI221_X1 U5493 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n4966), .ZN(n4971) );
  AOI22_X1 U5494 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_6_), .B2(
        keyinput_f25), .ZN(n4967) );
  OAI221_X1 U5495 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(DATAI_6_), .C2(
        keyinput_f25), .A(n4967), .ZN(n4970) );
  AOI22_X1 U5496 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput_f120), .B1(
        IR_REG_10__SCAN_IN), .B2(keyinput_f65), .ZN(n4968) );
  OAI221_X1 U5497 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput_f120), .C1(
        IR_REG_10__SCAN_IN), .C2(keyinput_f65), .A(n4968), .ZN(n4969) );
  NOR4_X1 U5498 ( .A1(n4972), .A2(n4971), .A3(n4970), .A4(n4969), .ZN(n4973)
         );
  NAND4_X1 U5499 ( .A1(n4976), .A2(n4975), .A3(n4974), .A4(n4973), .ZN(n5097)
         );
  INV_X1 U5500 ( .A(DATAI_24_), .ZN(n4978) );
  AOI22_X1 U5501 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput_f64), .B1(n4978), .B2(
        keyinput_f7), .ZN(n4977) );
  OAI221_X1 U5502 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput_f64), .C1(n4978), 
        .C2(keyinput_f7), .A(n4977), .ZN(n4990) );
  INV_X1 U5503 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U5504 ( .A1(n4981), .A2(keyinput_f52), .B1(n4980), .B2(keyinput_f34), .ZN(n4979) );
  OAI221_X1 U5505 ( .B1(n4981), .B2(keyinput_f52), .C1(n4980), .C2(
        keyinput_f34), .A(n4979), .ZN(n4989) );
  AOI22_X1 U5506 ( .A1(n3580), .A2(keyinput_f43), .B1(keyinput_f53), .B2(n4983), .ZN(n4982) );
  OAI221_X1 U5507 ( .B1(n3580), .B2(keyinput_f43), .C1(n4983), .C2(
        keyinput_f53), .A(n4982), .ZN(n4988) );
  AOI22_X1 U5508 ( .A1(n4986), .A2(keyinput_f0), .B1(n4985), .B2(keyinput_f2), 
        .ZN(n4984) );
  OAI221_X1 U5509 ( .B1(n4986), .B2(keyinput_f0), .C1(n4985), .C2(keyinput_f2), 
        .A(n4984), .ZN(n4987) );
  NOR4_X1 U5510 ( .A1(n4990), .A2(n4989), .A3(n4988), .A4(n4987), .ZN(n5035)
         );
  AOI22_X1 U5511 ( .A1(n2519), .A2(keyinput_f38), .B1(n2277), .B2(keyinput_f55), .ZN(n4991) );
  OAI221_X1 U5512 ( .B1(n2519), .B2(keyinput_f38), .C1(n2277), .C2(
        keyinput_f55), .A(n4991), .ZN(n5003) );
  AOI22_X1 U5513 ( .A1(n4993), .A2(keyinput_f35), .B1(n3444), .B2(keyinput_f85), .ZN(n4992) );
  OAI221_X1 U5514 ( .B1(n4993), .B2(keyinput_f35), .C1(n3444), .C2(
        keyinput_f85), .A(n4992), .ZN(n5002) );
  INV_X1 U5515 ( .A(IR_REG_1__SCAN_IN), .ZN(n4995) );
  AOI22_X1 U5516 ( .A1(n4996), .A2(keyinput_f119), .B1(n4995), .B2(
        keyinput_f56), .ZN(n4994) );
  OAI221_X1 U5517 ( .B1(n4996), .B2(keyinput_f119), .C1(n4995), .C2(
        keyinput_f56), .A(n4994), .ZN(n5001) );
  AOI22_X1 U5518 ( .A1(n4999), .A2(keyinput_f122), .B1(keyinput_f123), .B2(
        n4998), .ZN(n4997) );
  OAI221_X1 U5519 ( .B1(n4999), .B2(keyinput_f122), .C1(n4998), .C2(
        keyinput_f123), .A(n4997), .ZN(n5000) );
  NOR4_X1 U5520 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n5034)
         );
  AOI22_X1 U5521 ( .A1(n5006), .A2(keyinput_f33), .B1(keyinput_f127), .B2(
        n5005), .ZN(n5004) );
  OAI221_X1 U5522 ( .B1(n5006), .B2(keyinput_f33), .C1(n5005), .C2(
        keyinput_f127), .A(n5004), .ZN(n5016) );
  INV_X1 U5523 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5009) );
  AOI22_X1 U5524 ( .A1(n5009), .A2(keyinput_f124), .B1(n5008), .B2(
        keyinput_f125), .ZN(n5007) );
  OAI221_X1 U5525 ( .B1(n5009), .B2(keyinput_f124), .C1(n5008), .C2(
        keyinput_f125), .A(n5007), .ZN(n5015) );
  XOR2_X1 U5526 ( .A(n2527), .B(keyinput_f50), .Z(n5013) );
  XOR2_X1 U5527 ( .A(n2585), .B(keyinput_f51), .Z(n5012) );
  XNOR2_X1 U5528 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n5011) );
  XNOR2_X1 U5529 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_f66), .ZN(n5010) );
  NAND4_X1 U5530 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n5014)
         );
  NOR3_X1 U5531 ( .A1(n5016), .A2(n5015), .A3(n5014), .ZN(n5033) );
  AOI22_X1 U5532 ( .A1(n5019), .A2(keyinput_f108), .B1(keyinput_f104), .B2(
        n5018), .ZN(n5017) );
  OAI221_X1 U5533 ( .B1(n5019), .B2(keyinput_f108), .C1(n5018), .C2(
        keyinput_f104), .A(n5017), .ZN(n5031) );
  AOI22_X1 U5534 ( .A1(n5022), .A2(keyinput_f100), .B1(keyinput_f110), .B2(
        n5021), .ZN(n5020) );
  OAI221_X1 U5535 ( .B1(n5022), .B2(keyinput_f100), .C1(n5021), .C2(
        keyinput_f110), .A(n5020), .ZN(n5030) );
  AOI22_X1 U5536 ( .A1(n5025), .A2(keyinput_f89), .B1(keyinput_f112), .B2(
        n5024), .ZN(n5023) );
  OAI221_X1 U5537 ( .B1(n5025), .B2(keyinput_f89), .C1(n5024), .C2(
        keyinput_f112), .A(n5023), .ZN(n5029) );
  XOR2_X1 U5538 ( .A(n2628), .B(keyinput_f54), .Z(n5027) );
  XNOR2_X1 U5539 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_f83), .ZN(n5026) );
  NAND2_X1 U5540 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  NOR4_X1 U5541 ( .A1(n5031), .A2(n5030), .A3(n5029), .A4(n5028), .ZN(n5032)
         );
  NAND4_X1 U5542 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5032), .ZN(n5096)
         );
  AOI22_X1 U5543 ( .A1(n5038), .A2(keyinput_f90), .B1(keyinput_f115), .B2(
        n5037), .ZN(n5036) );
  OAI221_X1 U5544 ( .B1(n5038), .B2(keyinput_f90), .C1(n5037), .C2(
        keyinput_f115), .A(n5036), .ZN(n5050) );
  AOI22_X1 U5545 ( .A1(n5041), .A2(keyinput_f105), .B1(keyinput_f101), .B2(
        n5040), .ZN(n5039) );
  OAI221_X1 U5546 ( .B1(n5041), .B2(keyinput_f105), .C1(n5040), .C2(
        keyinput_f101), .A(n5039), .ZN(n5049) );
  AOI22_X1 U5547 ( .A1(n5044), .A2(keyinput_f92), .B1(keyinput_f93), .B2(n5043), .ZN(n5042) );
  OAI221_X1 U5548 ( .B1(n5044), .B2(keyinput_f92), .C1(n5043), .C2(
        keyinput_f93), .A(n5042), .ZN(n5048) );
  AOI22_X1 U5549 ( .A1(n2314), .A2(keyinput_f84), .B1(keyinput_f8), .B2(n5046), 
        .ZN(n5045) );
  OAI221_X1 U5550 ( .B1(n2314), .B2(keyinput_f84), .C1(n5046), .C2(keyinput_f8), .A(n5045), .ZN(n5047) );
  NOR4_X1 U5551 ( .A1(n5050), .A2(n5049), .A3(n5048), .A4(n5047), .ZN(n5094)
         );
  INV_X1 U5552 ( .A(DATAI_1_), .ZN(n5053) );
  AOI22_X1 U5553 ( .A1(n5053), .A2(keyinput_f30), .B1(n5052), .B2(keyinput_f4), 
        .ZN(n5051) );
  OAI221_X1 U5554 ( .B1(n5053), .B2(keyinput_f30), .C1(n5052), .C2(keyinput_f4), .A(n5051), .ZN(n5064) );
  AOI22_X1 U5555 ( .A1(n5055), .A2(keyinput_f10), .B1(n2689), .B2(keyinput_f72), .ZN(n5054) );
  OAI221_X1 U5556 ( .B1(n5055), .B2(keyinput_f10), .C1(n2689), .C2(
        keyinput_f72), .A(n5054), .ZN(n5063) );
  INV_X1 U5557 ( .A(DATAI_2_), .ZN(n5057) );
  AOI22_X1 U5558 ( .A1(n5058), .A2(keyinput_f5), .B1(n5057), .B2(keyinput_f29), 
        .ZN(n5056) );
  OAI221_X1 U5559 ( .B1(n5058), .B2(keyinput_f5), .C1(n5057), .C2(keyinput_f29), .A(n5056), .ZN(n5062) );
  XOR2_X1 U5560 ( .A(n2846), .B(keyinput_f78), .Z(n5060) );
  XNOR2_X1 U5561 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_f80), .ZN(n5059) );
  NAND2_X1 U5562 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  NOR4_X1 U5563 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n5093)
         );
  AOI22_X1 U5564 ( .A1(n5066), .A2(keyinput_f3), .B1(keyinput_f121), .B2(n4676), .ZN(n5065) );
  OAI221_X1 U5565 ( .B1(n5066), .B2(keyinput_f3), .C1(n4676), .C2(
        keyinput_f121), .A(n5065), .ZN(n5077) );
  INV_X1 U5566 ( .A(DATAI_3_), .ZN(n5069) );
  AOI22_X1 U5567 ( .A1(n5069), .A2(keyinput_f28), .B1(n5068), .B2(keyinput_f39), .ZN(n5067) );
  OAI221_X1 U5568 ( .B1(n5069), .B2(keyinput_f28), .C1(n5068), .C2(
        keyinput_f39), .A(n5067), .ZN(n5076) );
  XOR2_X1 U5569 ( .A(n5070), .B(keyinput_f31), .Z(n5074) );
  XNOR2_X1 U5570 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_f77), .ZN(n5073) );
  XNOR2_X1 U5571 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n5072) );
  XNOR2_X1 U5572 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_f63), .ZN(n5071) );
  NAND4_X1 U5573 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n5075)
         );
  NOR3_X1 U5574 ( .A1(n5077), .A2(n5076), .A3(n5075), .ZN(n5092) );
  INV_X1 U5575 ( .A(REG3_REG_12__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U5576 ( .A1(n2781), .A2(keyinput_f74), .B1(keyinput_f44), .B2(n5079), .ZN(n5078) );
  OAI221_X1 U5577 ( .B1(n2781), .B2(keyinput_f74), .C1(n5079), .C2(
        keyinput_f44), .A(n5078), .ZN(n5090) );
  AOI22_X1 U5578 ( .A1(n5082), .A2(keyinput_f19), .B1(keyinput_f26), .B2(n5081), .ZN(n5080) );
  OAI221_X1 U5579 ( .B1(n5082), .B2(keyinput_f19), .C1(n5081), .C2(
        keyinput_f26), .A(n5080), .ZN(n5089) );
  AOI22_X1 U5580 ( .A1(n2782), .A2(keyinput_f75), .B1(keyinput_f41), .B2(n5084), .ZN(n5083) );
  OAI221_X1 U5581 ( .B1(n2782), .B2(keyinput_f75), .C1(n5084), .C2(
        keyinput_f41), .A(n5083), .ZN(n5088) );
  XNOR2_X1 U5582 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_f81), .ZN(n5086) );
  XNOR2_X1 U5583 ( .A(DATAI_4_), .B(keyinput_f27), .ZN(n5085) );
  NAND2_X1 U5584 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  NOR4_X1 U5585 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n5087), .ZN(n5091)
         );
  NAND4_X1 U5586 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n5095)
         );
  NOR4_X1 U5587 ( .A1(n5098), .A2(n5097), .A3(n5096), .A4(n5095), .ZN(n5099)
         );
  NAND2_X1 U5588 ( .A1(n5100), .A2(n5099), .ZN(n5102) );
  AOI21_X1 U5589 ( .B1(keyinput_f45), .B2(n5102), .A(keyinput_g45), .ZN(n5104)
         );
  INV_X1 U5590 ( .A(keyinput_f45), .ZN(n5101) );
  AOI21_X1 U5591 ( .B1(n5102), .B2(n5101), .A(n2736), .ZN(n5103) );
  AOI22_X1 U5592 ( .A1(n2736), .A2(n5104), .B1(keyinput_g45), .B2(n5103), .ZN(
        n5105) );
  AOI21_X1 U5593 ( .B1(n5107), .B2(n5106), .A(n5105), .ZN(n5109) );
  AOI22_X1 U5594 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5108) );
  XNOR2_X1 U5595 ( .A(n5109), .B(n5108), .ZN(U3352) );
  AND2_X1 U2471 ( .A1(n3225), .A2(n3224), .ZN(n3326) );
  CLKBUF_X1 U2475 ( .A(n2508), .Z(n2606) );
  INV_X1 U2477 ( .A(n4206), .ZN(n4209) );
  NAND2_X1 U2478 ( .A1(n4206), .A2(n3401), .ZN(n4402) );
endmodule

