

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045;

  CLKBUF_X2 U3531 ( .A(n3444), .Z(n4343) );
  CLKBUF_X2 U3533 ( .A(n3379), .Z(n4352) );
  CLKBUF_X2 U3534 ( .A(n3512), .Z(n4347) );
  CLKBUF_X2 U3535 ( .A(n3431), .Z(n4086) );
  AND3_X1 U3536 ( .A1(n3223), .A2(n3224), .A3(n4728), .ZN(n3744) );
  AND2_X1 U3537 ( .A1(n4372), .A2(n3771), .ZN(n3398) );
  CLKBUF_X2 U3539 ( .A(n3378), .Z(n4353) );
  INV_X1 U3540 ( .A(n4367), .ZN(n4408) );
  INV_X2 U3541 ( .A(n5354), .ZN(n3791) );
  NOR2_X1 U3542 ( .A1(n4169), .A2(n3131), .ZN(n3130) );
  NAND2_X1 U3543 ( .A1(n3915), .A2(n3914), .ZN(n4679) );
  INV_X2 U3545 ( .A(n5586), .ZN(n6396) );
  NAND2_X1 U3546 ( .A1(n4901), .A2(n4902), .ZN(n4900) );
  AND2_X1 U3547 ( .A1(n6292), .A2(n6291), .ZN(n6359) );
  NAND2_X1 U3548 ( .A1(n4847), .A2(n4910), .ZN(n6597) );
  AND4_X1 U3549 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3083)
         );
  NOR3_X2 U3550 ( .A1(n4297), .A2(n4296), .A3(n4334), .ZN(n4335) );
  NOR2_X2 U3551 ( .A1(n5262), .A2(n5264), .ZN(n5249) );
  INV_X2 U3552 ( .A(n5366), .ZN(n3084) );
  NAND2_X1 U3553 ( .A1(n3769), .A2(n3768), .ZN(n3882) );
  NAND3_X1 U3555 ( .A1(n3408), .A2(n3407), .A3(n3409), .ZN(n3504) );
  CLKBUF_X1 U3556 ( .A(n3775), .Z(n4785) );
  INV_X2 U3557 ( .A(n4736), .ZN(n4630) );
  INV_X2 U3558 ( .A(n3392), .ZN(n3147) );
  INV_X2 U3559 ( .A(n3552), .ZN(n3149) );
  AND2_X2 U3560 ( .A1(n3780), .A2(n3280), .ZN(n3723) );
  INV_X1 U3561 ( .A(n4628), .ZN(n3399) );
  NOR2_X1 U3563 ( .A1(n3290), .A2(n3289), .ZN(n3151) );
  AOI22_X1 U3564 ( .A1(n3444), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3288) );
  CLKBUF_X2 U3565 ( .A(n3449), .Z(n4344) );
  CLKBUF_X2 U3566 ( .A(n3464), .Z(n4345) );
  BUF_X2 U3567 ( .A(n4346), .Z(n4279) );
  BUF_X2 U3568 ( .A(n3430), .Z(n4355) );
  AND2_X2 U3569 ( .A1(n4763), .A2(n4790), .ZN(n3430) );
  AND2_X1 U3570 ( .A1(n3169), .A2(n3118), .ZN(n5735) );
  AND2_X1 U3571 ( .A1(n4504), .A2(n4503), .ZN(n4505) );
  XNOR2_X1 U3572 ( .A(n5230), .B(n3268), .ZN(n5689) );
  XNOR2_X1 U3573 ( .A(n3267), .B(n4410), .ZN(n5213) );
  OR2_X1 U3574 ( .A1(n5629), .A2(n5885), .ZN(n4504) );
  AND2_X1 U3575 ( .A1(n5231), .A2(n5232), .ZN(n3171) );
  AOI21_X1 U3576 ( .B1(n5251), .B2(n5250), .A(n4499), .ZN(n5706) );
  AND2_X1 U3577 ( .A1(n3143), .A2(n3139), .ZN(n3138) );
  NAND2_X1 U3578 ( .A1(n5814), .A2(n3669), .ZN(n5775) );
  NAND2_X1 U3579 ( .A1(n3225), .A2(n3194), .ZN(n3193) );
  OR2_X1 U3580 ( .A1(n5777), .A2(n3666), .ZN(n5850) );
  NOR2_X1 U3581 ( .A1(n6073), .A2(n3871), .ZN(n6043) );
  XNOR2_X1 U3582 ( .A(n3619), .B(n6974), .ZN(n4951) );
  XNOR2_X1 U3583 ( .A(n3574), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4754)
         );
  INV_X2 U3584 ( .A(n3671), .ZN(n5777) );
  NAND2_X1 U3585 ( .A1(n5513), .A2(n4484), .ZN(n6387) );
  NAND2_X1 U3586 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  NAND2_X1 U3587 ( .A1(n3933), .A2(n3932), .ZN(n4686) );
  NAND2_X1 U3588 ( .A1(n3160), .A2(n3591), .ZN(n3592) );
  XNOR2_X1 U3589 ( .A(n3643), .B(n3642), .ZN(n3949) );
  NAND2_X1 U3590 ( .A1(n3632), .A2(n3631), .ZN(n3934) );
  OR2_X1 U3591 ( .A1(n3922), .A2(n3724), .ZN(n3160) );
  NAND2_X1 U3592 ( .A1(n3156), .A2(n3109), .ZN(n3643) );
  NAND2_X1 U3593 ( .A1(n3882), .A2(n3868), .ZN(n6061) );
  AND2_X1 U3594 ( .A1(n3569), .A2(n3609), .ZN(n4798) );
  OR2_X2 U3595 ( .A1(n6424), .A2(n4672), .ZN(n6436) );
  INV_X1 U3596 ( .A(n3609), .ZN(n3156) );
  OAI21_X1 U3597 ( .B1(n4630), .B2(n4465), .A(n4627), .ZN(n6421) );
  NAND2_X2 U3598 ( .A1(n5618), .A2(n3422), .ZN(n5623) );
  NAND2_X1 U3599 ( .A1(n4631), .A2(n4507), .ZN(n5210) );
  NAND2_X1 U3600 ( .A1(n3565), .A2(n3564), .ZN(n4699) );
  OR2_X1 U3601 ( .A1(n4804), .A2(n4515), .ZN(n4631) );
  OR2_X2 U3602 ( .A1(n4804), .A2(n6617), .ZN(n5892) );
  AOI21_X1 U3603 ( .B1(n3892), .B2(n3893), .A(n6326), .ZN(n4611) );
  NAND2_X1 U3604 ( .A1(n3530), .A2(n3529), .ZN(n3567) );
  NAND2_X1 U3605 ( .A1(n3550), .A2(n3549), .ZN(n6199) );
  NOR2_X1 U3606 ( .A1(n4931), .A2(n3220), .ZN(n3219) );
  AND2_X1 U3607 ( .A1(n3390), .A2(n3270), .ZN(n4518) );
  OR2_X1 U3608 ( .A1(n4807), .A2(n4814), .ZN(n3778) );
  CLKBUF_X1 U3609 ( .A(n3770), .Z(n5523) );
  INV_X1 U3610 ( .A(n3399), .ZN(n4736) );
  OR2_X1 U3612 ( .A1(n3455), .A2(n3454), .ZN(n3656) );
  AND2_X2 U3613 ( .A1(n3389), .A2(n4628), .ZN(n3483) );
  NAND2_X2 U3614 ( .A1(n3098), .A2(n3274), .ZN(n4728) );
  NAND2_X1 U3615 ( .A1(n3151), .A2(n3296), .ZN(n3384) );
  INV_X1 U3616 ( .A(n3389), .ZN(n3391) );
  NAND2_X2 U3617 ( .A1(n3318), .A2(n3317), .ZN(n4724) );
  AND2_X1 U3618 ( .A1(n3337), .A2(n3336), .ZN(n3274) );
  NAND2_X2 U3619 ( .A1(n3328), .A2(n3327), .ZN(n3401) );
  AND4_X1 U3620 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3296)
         );
  AND3_X1 U3621 ( .A1(n3335), .A2(n3334), .A3(n3333), .ZN(n3336) );
  AND4_X1 U3622 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3306)
         );
  AND4_X1 U3623 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3367)
         );
  AND4_X1 U3624 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  AND2_X1 U3625 ( .A1(n3939), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3950)
         );
  AND4_X1 U3626 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3327)
         );
  AND2_X1 U3627 ( .A1(n3312), .A2(n3311), .ZN(n3313) );
  AOI22_X1 U3628 ( .A1(n3517), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3292) );
  BUF_X2 U3629 ( .A(n3369), .Z(n4306) );
  BUF_X2 U3630 ( .A(n3517), .Z(n3085) );
  BUF_X2 U3631 ( .A(n3377), .Z(n4354) );
  NAND2_X1 U3632 ( .A1(n6725), .A2(n6326), .ZN(n6284) );
  BUF_X2 U3633 ( .A(n3577), .Z(n3086) );
  AND2_X2 U3634 ( .A1(n3281), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5178)
         );
  AND2_X2 U3635 ( .A1(n3283), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5179)
         );
  AND2_X2 U3636 ( .A1(n3282), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3291)
         );
  NAND2_X1 U3637 ( .A1(n3202), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4768) );
  INV_X2 U3638 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6326) );
  INV_X1 U3639 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3282) );
  NOR2_X2 U3640 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4762) );
  OAI211_X1 U3641 ( .C1(n3388), .C2(n3896), .A(n3423), .B(n3387), .ZN(n3395)
         );
  NOR2_X2 U3642 ( .A1(n5291), .A2(n5292), .ZN(n5276) );
  AND2_X2 U3643 ( .A1(n4499), .A2(n3265), .ZN(n5230) );
  AOI21_X2 U3644 ( .B1(n5523), .B2(n5545), .A(n6397), .ZN(n5596) );
  AND2_X2 U3645 ( .A1(n5249), .A2(n5248), .ZN(n4499) );
  XNOR2_X1 U3646 ( .A(n4783), .B(n6199), .ZN(n4701) );
  NOR2_X1 U3647 ( .A1(n5252), .A2(n5253), .ZN(n4446) );
  NAND2_X1 U3648 ( .A1(n4584), .A2(n6640), .ZN(n4804) );
  NAND2_X1 U3649 ( .A1(n3155), .A2(n3195), .ZN(n4419) );
  AOI21_X1 U3650 ( .B1(n3199), .B2(n3196), .A(n3115), .ZN(n3195) );
  OAI211_X1 U3651 ( .C1(n3230), .C2(n3154), .A(n3198), .B(n3153), .ZN(n3155)
         );
  NAND2_X1 U3652 ( .A1(n4458), .A2(n3402), .ZN(n3394) );
  OR2_X1 U3653 ( .A1(n3728), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3727)
         );
  NOR2_X1 U3654 ( .A1(n5232), .A2(n3266), .ZN(n3265) );
  INV_X1 U3655 ( .A(n4500), .ZN(n3266) );
  INV_X1 U3656 ( .A(n4369), .ZN(n4332) );
  AND2_X1 U3657 ( .A1(n3090), .A2(n5377), .ZN(n3253) );
  NOR2_X1 U3658 ( .A1(n5180), .A2(n6642), .ZN(n4369) );
  INV_X1 U3659 ( .A(n5617), .ZN(n3251) );
  INV_X1 U3660 ( .A(n5217), .ZN(n4390) );
  NAND2_X1 U3661 ( .A1(n3668), .A2(n5850), .ZN(n3237) );
  NOR2_X2 U3662 ( .A1(n4750), .A2(n4934), .ZN(n4933) );
  OAI21_X1 U3663 ( .B1(n3946), .B2(n3724), .A(n3618), .ZN(n3619) );
  NAND2_X1 U3664 ( .A1(n3149), .A2(n3656), .ZN(n3653) );
  INV_X1 U3665 ( .A(n3723), .ZN(n3714) );
  INV_X1 U3666 ( .A(n4518), .ZN(n4459) );
  OR3_X1 U3667 ( .A1(n4631), .A2(n4630), .A3(READY_N), .ZN(n4813) );
  XNOR2_X1 U3668 ( .A(n4427), .B(n5228), .ZN(n4492) );
  NAND2_X1 U3669 ( .A1(n4426), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4427)
         );
  INV_X1 U3670 ( .A(n4425), .ZN(n4426) );
  NAND2_X1 U3671 ( .A1(n4335), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4425)
         );
  NAND2_X1 U3672 ( .A1(n3130), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4199)
         );
  NAND2_X1 U3673 ( .A1(n4446), .A2(n4394), .ZN(n4395) );
  AND2_X2 U3674 ( .A1(n4628), .A2(n4728), .ZN(n5354) );
  NAND2_X1 U3675 ( .A1(n4421), .A2(n4420), .ZN(n4439) );
  AND2_X1 U3676 ( .A1(n3244), .A2(n3242), .ZN(n3241) );
  INV_X1 U3677 ( .A(n5754), .ZN(n3242) );
  INV_X1 U3678 ( .A(n3239), .ZN(n3238) );
  AOI21_X1 U3679 ( .B1(n3244), .B2(n3240), .A(n5741), .ZN(n3239) );
  NOR2_X1 U3680 ( .A1(n5754), .A2(n3247), .ZN(n3240) );
  XNOR2_X1 U3681 ( .A(n3671), .B(n6902), .ZN(n5822) );
  OR2_X1 U3682 ( .A1(n6039), .A2(n6042), .ZN(n6070) );
  INV_X1 U3683 ( .A(n6061), .ZN(n6464) );
  OR2_X1 U3684 ( .A1(n3773), .A2(n3772), .ZN(n6617) );
  NAND2_X1 U3685 ( .A1(n3799), .A2(n3791), .ZN(n5215) );
  INV_X1 U3686 ( .A(n3739), .ZN(n3740) );
  BUF_X1 U3687 ( .A(n3907), .Z(n6099) );
  INV_X1 U3688 ( .A(n3146), .ZN(n3696) );
  OAI211_X1 U3689 ( .C1(n3551), .C2(n4630), .A(n3148), .B(n3147), .ZN(n3146)
         );
  NAND2_X1 U3690 ( .A1(n3149), .A2(n4736), .ZN(n3148) );
  AOI22_X1 U3691 ( .A1(n3577), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U3692 ( .A1(n3369), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U3693 ( .A1(n3182), .A2(n3698), .ZN(n3181) );
  INV_X1 U3694 ( .A(n3704), .ZN(n3182) );
  NAND2_X1 U3695 ( .A1(n3156), .A2(n3271), .ZN(n3632) );
  NAND2_X1 U3696 ( .A1(n3422), .A2(n3896), .ZN(n3743) );
  OR2_X1 U3697 ( .A1(n3563), .A2(n3562), .ZN(n3571) );
  NOR2_X1 U3698 ( .A1(n3727), .A2(n6614), .ZN(n3754) );
  NAND2_X1 U3699 ( .A1(n6390), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3141)
         );
  NOR2_X1 U3700 ( .A1(n5481), .A2(n3144), .ZN(n5467) );
  NAND2_X1 U3701 ( .A1(n3145), .A2(REIP_REG_11__SCAN_IN), .ZN(n3144) );
  AND2_X1 U3702 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3411), .ZN(n3412) );
  OR2_X1 U3703 ( .A1(n4785), .A2(n4579), .ZN(n4808) );
  AND2_X1 U3704 ( .A1(n3371), .A2(n3370), .ZN(n3375) );
  NOR2_X1 U3705 ( .A1(n3257), .A2(n5367), .ZN(n3168) );
  NAND2_X1 U3706 ( .A1(n3258), .A2(n3259), .ZN(n3257) );
  INV_X1 U3707 ( .A(n5315), .ZN(n3258) );
  AND2_X1 U3708 ( .A1(n4082), .A2(n3256), .ZN(n3255) );
  INV_X1 U3709 ( .A(n5449), .ZN(n3256) );
  INV_X1 U3710 ( .A(n4615), .ZN(n3912) );
  INV_X1 U3711 ( .A(n3231), .ZN(n3152) );
  NAND2_X1 U3712 ( .A1(n5327), .A2(n5317), .ZN(n3217) );
  NOR2_X1 U3713 ( .A1(n3096), .A2(n3206), .ZN(n3205) );
  INV_X1 U3714 ( .A(n5426), .ZN(n3206) );
  NAND2_X1 U3715 ( .A1(n3193), .A2(n3111), .ZN(n5830) );
  NAND2_X1 U3716 ( .A1(n4466), .A2(n3791), .ZN(n4389) );
  INV_X1 U3717 ( .A(n4804), .ZN(n3188) );
  NOR2_X1 U3718 ( .A1(n3767), .A2(n3401), .ZN(n3187) );
  XNOR2_X1 U3719 ( .A(n3531), .B(n3532), .ZN(n3482) );
  NAND2_X1 U3720 ( .A1(n4587), .A2(n6642), .ZN(n3530) );
  OR2_X1 U3721 ( .A1(n5051), .A2(n6099), .ZN(n6239) );
  NAND2_X1 U3722 ( .A1(n3369), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U3723 ( .A1(n3518), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3312)
         );
  AOI22_X1 U3724 ( .A1(n3369), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3337) );
  AND2_X1 U3725 ( .A1(n4707), .A2(n6642), .ZN(n6113) );
  AND2_X1 U3726 ( .A1(n5014), .A2(n3509), .ZN(n4835) );
  INV_X1 U3727 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6610) );
  INV_X1 U3728 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U3729 ( .A1(n3730), .A2(n3729), .ZN(n3759) );
  AND2_X1 U3730 ( .A1(n5349), .A2(n4488), .ZN(n5316) );
  INV_X1 U3731 ( .A(n4098), .ZN(n4407) );
  INV_X1 U3732 ( .A(n4340), .ZN(n5232) );
  AND2_X1 U3733 ( .A1(n4500), .A2(n5248), .ZN(n3170) );
  NAND2_X1 U3734 ( .A1(n3128), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4294)
         );
  INV_X1 U3735 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3131) );
  AND3_X1 U3736 ( .A1(n3947), .A2(n4925), .A3(n4906), .ZN(n3948) );
  NAND2_X1 U3737 ( .A1(n5710), .A2(n5681), .ZN(n5692) );
  AND2_X1 U3738 ( .A1(n4393), .A2(n4392), .ZN(n4447) );
  INV_X1 U3739 ( .A(n4395), .ZN(n4448) );
  INV_X1 U3740 ( .A(n4446), .ZN(n5255) );
  NAND2_X1 U3741 ( .A1(n5777), .A2(n4437), .ZN(n4438) );
  NAND2_X1 U3742 ( .A1(n4439), .A2(n4438), .ZN(n5710) );
  AND2_X1 U3743 ( .A1(n3117), .A2(n3245), .ZN(n3244) );
  NAND2_X1 U3744 ( .A1(n3247), .A2(n3246), .ZN(n3245) );
  NOR2_X1 U3745 ( .A1(n5353), .A2(n5357), .ZN(n3836) );
  AND2_X1 U3746 ( .A1(n3882), .A2(n3870), .ZN(n6042) );
  INV_X1 U3747 ( .A(n5830), .ZN(n3236) );
  INV_X1 U3748 ( .A(n3237), .ZN(n3233) );
  INV_X1 U3749 ( .A(n5822), .ZN(n3158) );
  OR2_X1 U3750 ( .A1(n6734), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5207) );
  INV_X1 U3751 ( .A(n5484), .ZN(n3218) );
  OR2_X1 U3752 ( .A1(n4951), .A2(n3094), .ZN(n3162) );
  INV_X1 U3753 ( .A(n3094), .ZN(n3165) );
  INV_X1 U3754 ( .A(n6021), .ZN(n6074) );
  NAND2_X1 U3755 ( .A1(n3574), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3576)
         );
  OAI21_X1 U3756 ( .B1(n6430), .B2(n6426), .A(n6427), .ZN(n4753) );
  OR2_X1 U3757 ( .A1(n3773), .A2(n5198), .ZN(n4803) );
  AND2_X1 U3758 ( .A1(n3882), .A2(n6601), .ZN(n6039) );
  OAI21_X1 U3759 ( .B1(n3892), .B2(n3724), .A(n3499), .ZN(n4624) );
  OAI211_X1 U3760 ( .C1(n3714), .C2(n3480), .A(n3479), .B(n3478), .ZN(n3491)
         );
  AND2_X1 U3761 ( .A1(n6316), .A2(n6484), .ZN(n6323) );
  AND2_X1 U3762 ( .A1(n3275), .A2(n3087), .ZN(n6320) );
  AND2_X1 U3763 ( .A1(n4835), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6487) );
  AND2_X1 U3764 ( .A1(n4700), .A2(n6099), .ZN(n4709) );
  NOR3_X1 U3765 ( .A1(n6839), .A2(n6610), .A3(n7013), .ZN(n4829) );
  AOI21_X1 U3766 ( .B1(n6281), .B2(STATE2_REG_3__SCAN_IN), .A(n5077), .ZN(
        n6286) );
  INV_X1 U3767 ( .A(n5523), .ZN(n5198) );
  NOR2_X1 U3768 ( .A1(n3134), .A2(n3132), .ZN(n3139) );
  NOR2_X1 U3769 ( .A1(n3142), .A2(n3133), .ZN(n3132) );
  NAND2_X1 U3770 ( .A1(n3136), .A2(n3135), .ZN(n3134) );
  AND2_X1 U3771 ( .A1(n5271), .A2(n4481), .ZN(n5244) );
  NOR2_X2 U3772 ( .A1(n4468), .A2(n4467), .ZN(n6393) );
  INV_X1 U3773 ( .A(n4491), .ZN(n3127) );
  NAND2_X1 U3774 ( .A1(n4379), .A2(n4378), .ZN(n5618) );
  OR2_X1 U3775 ( .A1(n4377), .A2(n4376), .ZN(n4378) );
  OR3_X1 U3776 ( .A1(n4584), .A2(n6638), .A3(n4593), .ZN(n4379) );
  AND2_X1 U3777 ( .A1(n5678), .A2(n4816), .ZN(n5660) );
  AND2_X1 U3778 ( .A1(n5678), .A2(n4818), .ZN(n5661) );
  INV_X1 U3779 ( .A(n5678), .ZN(n5673) );
  OR3_X1 U3780 ( .A1(n4804), .A2(n4525), .A3(n6664), .ZN(n4553) );
  OAI22_X1 U3781 ( .A1(n4439), .A2(n3114), .B1(n4423), .B2(n5691), .ZN(n3157)
         );
  OR2_X1 U3782 ( .A1(n6651), .A2(n6284), .ZN(n5885) );
  XNOR2_X1 U3783 ( .A(n3215), .B(n3214), .ZN(n5899) );
  INV_X1 U3784 ( .A(n5222), .ZN(n3214) );
  NAND2_X1 U3785 ( .A1(n3112), .A2(n4444), .ZN(n3186) );
  XNOR2_X1 U3786 ( .A(n4399), .B(n5219), .ZN(n5904) );
  NOR2_X1 U3787 ( .A1(n5970), .A2(n3885), .ZN(n5949) );
  INV_X1 U3788 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6281) );
  INV_X1 U3789 ( .A(n6284), .ZN(n6484) );
  CLKBUF_X1 U3790 ( .A(n4587), .Z(n6101) );
  INV_X1 U3791 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6839) );
  OR2_X1 U3792 ( .A1(n5019), .A2(n6099), .ZN(n6206) );
  AND2_X1 U3793 ( .A1(n6626), .A2(n6625), .ZN(n6639) );
  NAND2_X1 U3794 ( .A1(n3697), .A2(n3739), .ZN(n3178) );
  NAND2_X1 U3795 ( .A1(n3696), .A2(n3695), .ZN(n3692) );
  AND2_X1 U3796 ( .A1(n3483), .A2(n3771), .ZN(n3418) );
  NOR2_X1 U3797 ( .A1(n3395), .A2(n4736), .ZN(n3419) );
  OR2_X2 U3798 ( .A1(n3780), .A2(n6642), .ZN(n3551) );
  NAND2_X1 U3799 ( .A1(n3400), .A2(n4728), .ZN(n3423) );
  NAND2_X1 U3800 ( .A1(n3771), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3552) );
  INV_X1 U3801 ( .A(n5448), .ZN(n3254) );
  OR2_X1 U3802 ( .A1(n3604), .A2(n3603), .ZN(n3616) );
  OR2_X1 U3803 ( .A1(n3587), .A2(n3586), .ZN(n3613) );
  INV_X1 U3804 ( .A(n3401), .ZN(n3859) );
  OR2_X1 U3805 ( .A1(n3442), .A2(n3441), .ZN(n3484) );
  CLKBUF_X1 U3806 ( .A(n3485), .Z(n3857) );
  OR2_X1 U3807 ( .A1(n3524), .A2(n3523), .ZN(n3526) );
  NAND2_X1 U3808 ( .A1(n3747), .A2(n3771), .ZN(n3224) );
  AND2_X1 U3809 ( .A1(n4372), .A2(n3422), .ZN(n3223) );
  NAND2_X1 U3810 ( .A1(n3746), .A2(n4469), .ZN(n3222) );
  INV_X1 U3811 ( .A(n3418), .ZN(n3221) );
  AOI21_X1 U3812 ( .B1(n3402), .B2(n3392), .A(n3401), .ZN(n3403) );
  AND2_X1 U3813 ( .A1(n3711), .A2(n3712), .ZN(n3179) );
  AOI21_X1 U3814 ( .B1(n3754), .B2(n3723), .A(n3722), .ZN(n3733) );
  AND2_X1 U3815 ( .A1(n6642), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3722)
         );
  OR2_X1 U3816 ( .A1(n4274), .A2(n4273), .ZN(n4290) );
  OR2_X1 U3817 ( .A1(n4240), .A2(n4239), .ZN(n4254) );
  AND2_X1 U3818 ( .A1(n5326), .A2(n3260), .ZN(n3259) );
  INV_X1 U3819 ( .A(n3261), .ZN(n3260) );
  NAND2_X1 U3820 ( .A1(n5335), .A2(n3262), .ZN(n3261) );
  NAND2_X1 U3821 ( .A1(n4137), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4138)
         );
  INV_X1 U3822 ( .A(n4136), .ZN(n4137) );
  NOR2_X1 U3823 ( .A1(n4084), .A2(n4083), .ZN(n3129) );
  AND2_X1 U3824 ( .A1(n4043), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4047)
         );
  INV_X1 U3825 ( .A(n4900), .ZN(n3971) );
  AND2_X1 U3826 ( .A1(n4816), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3908) );
  NOR2_X1 U3827 ( .A1(n3200), .A2(n4416), .ZN(n3198) );
  INV_X1 U3828 ( .A(n3669), .ZN(n3154) );
  AND2_X1 U3829 ( .A1(n3197), .A2(n3095), .ZN(n3196) );
  INV_X1 U3830 ( .A(n4416), .ZN(n3197) );
  INV_X1 U3831 ( .A(n3674), .ZN(n3246) );
  INV_X1 U3832 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5787) );
  AOI21_X1 U3833 ( .B1(n3234), .B2(n3232), .A(n3102), .ZN(n3231) );
  INV_X1 U3834 ( .A(n3276), .ZN(n3232) );
  INV_X1 U3835 ( .A(n5439), .ZN(n3207) );
  NOR2_X1 U3836 ( .A1(n4588), .A2(n3866), .ZN(n3869) );
  NOR2_X1 U3837 ( .A1(n5470), .A2(n3209), .ZN(n3208) );
  INV_X1 U3838 ( .A(n5450), .ZN(n3209) );
  OR2_X1 U3839 ( .A1(n6078), .A2(n6079), .ZN(n3871) );
  INV_X1 U3840 ( .A(n4973), .ZN(n3220) );
  NAND2_X1 U3841 ( .A1(n4798), .A2(n3483), .ZN(n3573) );
  OR2_X1 U3842 ( .A1(n3474), .A2(n3473), .ZN(n3497) );
  OR2_X1 U3843 ( .A1(n3743), .A2(n3742), .ZN(n5180) );
  NOR2_X1 U3844 ( .A1(n4728), .A2(n3401), .ZN(n4375) );
  AND2_X1 U3845 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U3846 ( .A1(n3436), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3310) );
  AND2_X1 U3847 ( .A1(n4797), .A2(n6099), .ZN(n4975) );
  AND2_X1 U3848 ( .A1(n3761), .A2(n3760), .ZN(n4517) );
  NAND2_X1 U3849 ( .A1(n5899), .A2(n6393), .ZN(n3136) );
  AOI21_X1 U3850 ( .B1(n5224), .B2(REIP_REG_31__SCAN_IN), .A(n3140), .ZN(n3135) );
  NAND2_X1 U3851 ( .A1(n5227), .A2(n3141), .ZN(n3140) );
  INV_X1 U3852 ( .A(n5225), .ZN(n3133) );
  NAND2_X1 U3853 ( .A1(n5467), .A2(REIP_REG_12__SCAN_IN), .ZN(n5437) );
  INV_X1 U3854 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U3855 ( .A1(n5577), .A2(n4477), .ZN(n5481) );
  INV_X1 U3856 ( .A(n3503), .ZN(n3250) );
  NAND2_X1 U3857 ( .A1(n3504), .A2(n3502), .ZN(n3249) );
  MUX2_X1 U3858 ( .A(n4316), .B(n5240), .S(n4460), .Z(n4500) );
  NOR2_X1 U3859 ( .A1(n3264), .A2(n3268), .ZN(n3263) );
  INV_X1 U3860 ( .A(n3265), .ZN(n3264) );
  NAND2_X1 U3861 ( .A1(n4295), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4297)
         );
  INV_X1 U3862 ( .A(n4294), .ZN(n4295) );
  CLKBUF_X1 U3863 ( .A(n5262), .Z(n5263) );
  NAND2_X1 U3864 ( .A1(n4200), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4202)
         );
  INV_X1 U3865 ( .A(n4199), .ZN(n4200) );
  INV_X1 U3866 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4201) );
  AND2_X1 U3867 ( .A1(n3168), .A2(n4227), .ZN(n3167) );
  NAND2_X1 U3868 ( .A1(n3129), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4136)
         );
  INV_X1 U3869 ( .A(n3129), .ZN(n4104) );
  NAND2_X1 U3870 ( .A1(n4047), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4084)
         );
  AND2_X1 U3871 ( .A1(n4031), .A2(n4030), .ZN(n5449) );
  AND3_X1 U3872 ( .A1(n4029), .A2(n4028), .A3(n4027), .ZN(n4030) );
  NAND2_X1 U3873 ( .A1(n4015), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4016)
         );
  NOR2_X1 U3874 ( .A1(n6878), .A2(n4016), .ZN(n4043) );
  AND3_X1 U3875 ( .A1(n4001), .A2(n4000), .A3(n3999), .ZN(n5617) );
  CLKBUF_X1 U3876 ( .A(n5459), .Z(n5460) );
  NAND2_X1 U3877 ( .A1(n3982), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3983)
         );
  NOR2_X1 U3878 ( .A1(n6919), .A2(n3983), .ZN(n4012) );
  AND3_X1 U3879 ( .A1(n3969), .A2(n3968), .A3(n3967), .ZN(n4965) );
  AND2_X1 U3880 ( .A1(n3950), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3982)
         );
  NAND2_X1 U3881 ( .A1(n3159), .A2(n3937), .ZN(n4925) );
  NOR2_X1 U3882 ( .A1(n3938), .A2(n3942), .ZN(n3939) );
  OR2_X1 U3883 ( .A1(n4747), .A2(n4746), .ZN(n4907) );
  AND2_X1 U3884 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3918), .ZN(n3923)
         );
  NAND2_X1 U3885 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3924) );
  NAND2_X1 U3886 ( .A1(n3913), .A2(n3912), .ZN(n3914) );
  INV_X1 U3887 ( .A(n3911), .ZN(n3913) );
  NAND2_X1 U3888 ( .A1(n4616), .A2(n4614), .ZN(n4615) );
  AND2_X1 U3889 ( .A1(n4385), .A2(n4384), .ZN(n5266) );
  INV_X1 U3890 ( .A(n5265), .ZN(n5283) );
  OR2_X1 U3891 ( .A1(n3217), .A2(n5305), .ZN(n3216) );
  AND2_X1 U3892 ( .A1(n3835), .A2(n3834), .ZN(n5357) );
  INV_X1 U3893 ( .A(n6469), .ZN(n5983) );
  NOR2_X1 U3894 ( .A1(n5615), .A2(n5470), .ZN(n5469) );
  NAND2_X1 U3895 ( .A1(n4933), .A2(n3099), .ZN(n5483) );
  NAND2_X1 U3896 ( .A1(n3172), .A2(n3126), .ZN(n6073) );
  NAND2_X1 U3897 ( .A1(n4933), .A2(n4973), .ZN(n4971) );
  NOR2_X1 U3898 ( .A1(n6061), .A2(n3173), .ZN(n3172) );
  INV_X1 U3899 ( .A(n6077), .ZN(n3173) );
  CLKBUF_X1 U3900 ( .A(n4933), .Z(n4972) );
  NOR2_X1 U3901 ( .A1(n4690), .A2(n3210), .ZN(n3211) );
  NOR2_X1 U3902 ( .A1(n4690), .A2(n3213), .ZN(n3212) );
  INV_X1 U3903 ( .A(n4682), .ZN(n3213) );
  OR2_X1 U3904 ( .A1(n3500), .A2(n6470), .ZN(n3501) );
  NAND2_X1 U3905 ( .A1(n4683), .A2(n4682), .ZN(n4689) );
  NAND2_X1 U3906 ( .A1(n3188), .A2(n3187), .ZN(n3768) );
  AND2_X1 U3907 ( .A1(n3786), .A2(n3785), .ZN(n4608) );
  NAND2_X1 U3908 ( .A1(n3481), .A2(n3491), .ZN(n3495) );
  INV_X1 U3909 ( .A(n4698), .ZN(n5127) );
  XNOR2_X1 U3910 ( .A(n3544), .B(n3545), .ZN(n4587) );
  CLKBUF_X1 U3911 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n6980) );
  NOR2_X1 U3912 ( .A1(n4459), .A2(n4630), .ZN(n6601) );
  INV_X1 U3913 ( .A(n5058), .ZN(n5053) );
  AND2_X1 U3914 ( .A1(n6099), .A2(n4796), .ZN(n5128) );
  NOR2_X1 U3915 ( .A1(n6239), .A2(n6238), .ZN(n6292) );
  INV_X1 U3916 ( .A(n3892), .ZN(n6291) );
  INV_X1 U3917 ( .A(n6239), .ZN(n4847) );
  AND2_X1 U3918 ( .A1(n6238), .A2(n6291), .ZN(n4920) );
  AND2_X1 U3919 ( .A1(n6113), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4737) );
  AND2_X1 U3920 ( .A1(n4975), .A2(n6291), .ZN(n4834) );
  NAND2_X1 U3921 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4792) );
  AND2_X1 U3922 ( .A1(n4786), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3764) );
  AND2_X1 U3923 ( .A1(n6642), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4461) );
  INV_X1 U3924 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U3925 ( .A1(n6713), .A2(REIP_REG_31__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3926 ( .A1(n5259), .A2(n3092), .ZN(n5237) );
  NAND2_X1 U3927 ( .A1(n3150), .A2(n5501), .ZN(n5271) );
  NAND2_X1 U3928 ( .A1(n5316), .A2(n3125), .ZN(n3150) );
  INV_X1 U3929 ( .A(n5522), .ZN(n6397) );
  CLKBUF_X1 U3930 ( .A(n4702), .Z(n4703) );
  INV_X1 U3931 ( .A(n5618), .ZN(n5621) );
  OAI21_X1 U3932 ( .B1(n4499), .B2(n4500), .A(n5231), .ZN(n5629) );
  INV_X1 U3933 ( .A(n5827), .ZN(n5668) );
  NAND2_X1 U3934 ( .A1(n4820), .A2(n4819), .ZN(n5674) );
  AND2_X1 U3935 ( .A1(n4811), .A2(n4810), .ZN(n4812) );
  OR2_X1 U3936 ( .A1(n4804), .A2(n4803), .ZN(n4811) );
  INV_X1 U3937 ( .A(n5674), .ZN(n5679) );
  AND2_X1 U3938 ( .A1(n4553), .A2(n5208), .ZN(n6746) );
  INV_X1 U3939 ( .A(n4553), .ZN(n6745) );
  CLKBUF_X1 U3940 ( .A(n6421), .Z(n4693) );
  INV_X1 U3941 ( .A(n4813), .ZN(n6415) );
  NOR2_X1 U3942 ( .A1(n5230), .A2(n3171), .ZN(n5697) );
  INV_X1 U3943 ( .A(n3128), .ZN(n4260) );
  INV_X1 U3944 ( .A(n3130), .ZN(n4171) );
  OAI21_X1 U3945 ( .B1(n3262), .B2(n5348), .A(n3103), .ZN(n5774) );
  AND2_X1 U3946 ( .A1(n5366), .A2(n5378), .ZN(n5792) );
  OR2_X1 U3947 ( .A1(n3097), .A2(n5394), .ZN(n5798) );
  INV_X1 U3948 ( .A(n6436), .ZN(n5889) );
  AND2_X2 U3949 ( .A1(n5892), .A2(n4429), .ZN(n6424) );
  NAND2_X1 U3950 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  NAND2_X1 U3951 ( .A1(n5692), .A2(n5915), .ZN(n5683) );
  OR2_X1 U3952 ( .A1(n4449), .A2(n4448), .ZN(n5600) );
  AOI21_X1 U3953 ( .B1(n4441), .B2(n5699), .A(n4440), .ZN(n4443) );
  NAND2_X1 U3954 ( .A1(n4439), .A2(n3089), .ZN(n4441) );
  OR2_X1 U3955 ( .A1(n5943), .A2(n4445), .ZN(n5926) );
  NAND2_X1 U3956 ( .A1(n4439), .A2(n3088), .ZN(n5700) );
  INV_X1 U3957 ( .A(n4439), .ZN(n5717) );
  NAND2_X1 U3958 ( .A1(n3243), .A2(n3108), .ZN(n3169) );
  NOR3_X1 U3959 ( .A1(n5337), .A2(n3843), .A3(n3845), .ZN(n5318) );
  XNOR2_X1 U3960 ( .A(n5745), .B(n5744), .ZN(n5963) );
  AOI21_X1 U3961 ( .B1(n5732), .B2(n3241), .A(n3238), .ZN(n5745) );
  OAI21_X1 U3962 ( .B1(n3192), .B2(n3191), .A(n3190), .ZN(n5970) );
  NOR2_X1 U3963 ( .A1(n5979), .A2(n3110), .ZN(n3190) );
  NOR2_X1 U3964 ( .A1(n5980), .A2(n3884), .ZN(n3192) );
  AND2_X1 U3965 ( .A1(n3875), .A2(n6006), .ZN(n5965) );
  NOR2_X1 U3966 ( .A1(n5337), .A2(n3843), .ZN(n5328) );
  NAND2_X1 U3967 ( .A1(n3243), .A2(n3244), .ZN(n5753) );
  NAND2_X1 U3968 ( .A1(n3235), .A2(n3234), .ZN(n5821) );
  AND2_X1 U3969 ( .A1(n3235), .A2(n3233), .ZN(n5823) );
  NAND2_X1 U3970 ( .A1(n3236), .A2(n3276), .ZN(n3235) );
  INV_X1 U3971 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U3972 ( .A1(n5875), .A2(n5876), .ZN(n3229) );
  NAND2_X1 U3973 ( .A1(n4951), .A2(n3166), .ZN(n3161) );
  INV_X1 U3974 ( .A(n3172), .ZN(n4957) );
  NAND2_X1 U3975 ( .A1(n6070), .A2(n4641), .ZN(n6469) );
  OR2_X1 U3976 ( .A1(n6070), .A2(n6464), .ZN(n6021) );
  OR2_X1 U3977 ( .A1(n6039), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4641)
         );
  INV_X1 U3978 ( .A(n5127), .ZN(n6238) );
  INV_X1 U3979 ( .A(n4798), .ZN(n5051) );
  INV_X1 U3980 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U3981 ( .A1(n4791), .A2(n5077), .ZN(n6475) );
  INV_X1 U3982 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3283) );
  OAI21_X1 U3983 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6725), .A(n6367), .ZN(
        n6732) );
  NAND2_X1 U3984 ( .A1(n4709), .A2(n6291), .ZN(n6152) );
  OAI21_X1 U3985 ( .B1(n6205), .B2(n6204), .A(n6203), .ZN(n6230) );
  OR2_X1 U3986 ( .A1(n6247), .A2(n6246), .ZN(n6275) );
  AOI22_X1 U3987 ( .A1(n6323), .A2(n6320), .B1(n6477), .B2(n6318), .ZN(n6362)
         );
  OAI21_X1 U3988 ( .B1(n4846), .B2(n4845), .A(n4844), .ZN(n6594) );
  NOR2_X1 U3989 ( .A1(n4828), .A2(n5077), .ZN(n6562) );
  AND2_X1 U3990 ( .A1(n4737), .A2(n4724), .ZN(n6542) );
  NAND2_X1 U3991 ( .A1(n6431), .A2(DATAI_22_), .ZN(n6515) );
  NAND2_X1 U3992 ( .A1(n6431), .A2(DATAI_23_), .ZN(n6589) );
  INV_X1 U3993 ( .A(n5073), .ZN(n5115) );
  NOR2_X1 U3994 ( .A1(n4824), .A2(n5077), .ZN(n6569) );
  NOR2_X1 U3995 ( .A1(n4826), .A2(n5077), .ZN(n6534) );
  AND2_X1 U3996 ( .A1(n4737), .A2(n3401), .ZN(n6532) );
  NOR2_X1 U3997 ( .A1(n4821), .A2(n5077), .ZN(n6576) );
  AND2_X1 U3998 ( .A1(n4737), .A2(n4728), .ZN(n6538) );
  NOR2_X1 U3999 ( .A1(n4909), .A2(n5077), .ZN(n6583) );
  AND2_X1 U4000 ( .A1(n4737), .A2(n3147), .ZN(n6508) );
  NOR2_X1 U4001 ( .A1(n7023), .A2(n5077), .ZN(n6553) );
  NOR2_X1 U4002 ( .A1(n4905), .A2(n5077), .ZN(n6593) );
  AND2_X1 U4003 ( .A1(n4737), .A2(n3422), .ZN(n6517) );
  INV_X1 U4004 ( .A(n4834), .ZN(n5010) );
  INV_X1 U4005 ( .A(n6562), .ZN(n6330) );
  INV_X1 U4006 ( .A(n6569), .ZN(n6334) );
  INV_X1 U4007 ( .A(n6528), .ZN(n6566) );
  INV_X1 U4008 ( .A(n6534), .ZN(n6338) );
  INV_X1 U4009 ( .A(n6576), .ZN(n6342) );
  INV_X1 U4010 ( .A(n6538), .ZN(n6573) );
  INV_X1 U4011 ( .A(n6544), .ZN(n6346) );
  INV_X1 U4012 ( .A(n6542), .ZN(n6264) );
  INV_X1 U4013 ( .A(n6508), .ZN(n6580) );
  INV_X1 U4014 ( .A(n6581), .ZN(n6303) );
  INV_X1 U4015 ( .A(n6548), .ZN(n6271) );
  NAND2_X1 U4016 ( .A1(n6431), .A2(DATAI_30_), .ZN(n6558) );
  NAND2_X1 U4017 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4829), .ZN(n4738) );
  INV_X1 U4018 ( .A(n6593), .ZN(n6361) );
  INV_X1 U4019 ( .A(n6517), .ZN(n6588) );
  INV_X1 U4020 ( .A(n6152), .ZN(n4741) );
  OAI211_X1 U4021 ( .C1(n4829), .C2(n6484), .A(n4708), .B(n6286), .ZN(n4735)
         );
  INV_X1 U4022 ( .A(n4894), .ZN(n4744) );
  NAND2_X1 U4023 ( .A1(n4584), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6635) );
  INV_X1 U4024 ( .A(n6640), .ZN(n6638) );
  AND2_X1 U4025 ( .A1(n6632), .A2(n6631), .ZN(n6648) );
  NAND2_X1 U4026 ( .A1(n6725), .A2(n4786), .ZN(n6734) );
  INV_X1 U4027 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U4028 ( .A1(n4786), .A2(n6326), .ZN(n6650) );
  INV_X1 U4029 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6725) );
  INV_X1 U4030 ( .A(n6648), .ZN(n6724) );
  INV_X1 U4031 ( .A(n6654), .ZN(n6722) );
  NAND2_X1 U4032 ( .A1(n3753), .A2(n3752), .ZN(n6664) );
  AND2_X1 U4033 ( .A1(n3752), .A2(STATE_REG_1__SCAN_IN), .ZN(n6719) );
  INV_X2 U4034 ( .A(n6719), .ZN(n6743) );
  NAND2_X1 U4035 ( .A1(n5259), .A2(n3093), .ZN(n3143) );
  NOR2_X1 U4036 ( .A1(n5586), .A2(n5727), .ZN(n5296) );
  AOI21_X1 U4037 ( .B1(n4403), .B2(n4402), .A(n4401), .ZN(n4404) );
  NOR2_X1 U4038 ( .A1(n5618), .A2(n4400), .ZN(n4401) );
  NAND2_X1 U4039 ( .A1(n3112), .A2(n4424), .ZN(n4435) );
  NAND2_X1 U4040 ( .A1(n5898), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3184) );
  AOI21_X1 U4041 ( .B1(n5899), .B2(n6463), .A(n5897), .ZN(n3185) );
  NAND2_X1 U4042 ( .A1(n5348), .A2(n3259), .ZN(n5313) );
  NAND2_X1 U4043 ( .A1(n3971), .A2(n3121), .ZN(n5479) );
  NOR2_X1 U4045 ( .A1(n5347), .A2(n3261), .ZN(n5325) );
  AND2_X1 U4046 ( .A1(n4438), .A2(n3122), .ZN(n3088) );
  AND2_X1 U4047 ( .A1(n4438), .A2(n3113), .ZN(n3089) );
  NAND2_X1 U4048 ( .A1(n3084), .A2(n4135), .ZN(n5347) );
  AND2_X1 U4049 ( .A1(n3255), .A2(n5393), .ZN(n3090) );
  OR2_X1 U4050 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3091) );
  NAND2_X1 U4051 ( .A1(n3204), .A2(n3208), .ZN(n5438) );
  NAND2_X1 U4052 ( .A1(n5577), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5585) );
  INV_X1 U4053 ( .A(n5585), .ZN(n6390) );
  AND2_X1 U4054 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n3092) );
  AND3_X1 U4055 ( .A1(n3137), .A2(n3092), .A3(REIP_REG_30__SCAN_IN), .ZN(n3093) );
  NOR2_X1 U4056 ( .A1(n5448), .A2(n5449), .ZN(n5406) );
  AND2_X1 U4057 ( .A1(n3619), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3094)
         );
  INV_X1 U4058 ( .A(n3422), .ZN(n5191) );
  NAND2_X1 U4059 ( .A1(n3252), .A2(n3255), .ZN(n5391) );
  AND2_X1 U4060 ( .A1(n3084), .A2(n3168), .ZN(n5300) );
  NAND2_X1 U4061 ( .A1(n3971), .A2(n3970), .ZN(n4964) );
  AND2_X1 U4062 ( .A1(n5832), .A2(n3672), .ZN(n3095) );
  NAND2_X1 U4063 ( .A1(n3208), .A2(n3207), .ZN(n3096) );
  AND2_X1 U4064 ( .A1(n3252), .A2(n3090), .ZN(n3097) );
  AND4_X1 U4065 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3098)
         );
  AND2_X1 U4066 ( .A1(n3219), .A2(n4967), .ZN(n3099) );
  AND4_X1 U4067 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3100)
         );
  NAND2_X1 U4068 ( .A1(n3084), .A2(n3167), .ZN(n5291) );
  NAND2_X1 U4069 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3500)
         );
  NAND2_X1 U4070 ( .A1(n3193), .A2(n3662), .ZN(n5853) );
  AND2_X1 U4071 ( .A1(n5732), .A2(n3674), .ZN(n3101) );
  AND2_X1 U4072 ( .A1(n5777), .A2(n6902), .ZN(n3102) );
  AND2_X1 U4073 ( .A1(n4589), .A2(n3780), .ZN(n4458) );
  AOI21_X1 U4074 ( .B1(n5685), .B2(n4460), .A(n4371), .ZN(n4406) );
  INV_X1 U4075 ( .A(n4406), .ZN(n3268) );
  OR2_X1 U4076 ( .A1(n5347), .A2(n5346), .ZN(n3103) );
  NOR3_X1 U4077 ( .A1(n5437), .A2(n6690), .A3(n6688), .ZN(n3104) );
  INV_X1 U4078 ( .A(n5867), .ZN(n3228) );
  INV_X1 U4079 ( .A(n3227), .ZN(n3226) );
  OAI21_X1 U4080 ( .B1(n3652), .B2(n3228), .A(n3661), .ZN(n3227) );
  NAND2_X1 U4081 ( .A1(n3495), .A2(n3653), .ZN(n3533) );
  OR2_X1 U4082 ( .A1(n4297), .A2(n4296), .ZN(n3105) );
  AND2_X1 U4083 ( .A1(n3224), .A2(n3223), .ZN(n3106) );
  NAND2_X1 U4084 ( .A1(n3221), .A2(n3222), .ZN(n3107) );
  AND2_X1 U4085 ( .A1(n3241), .A2(n5742), .ZN(n3108) );
  INV_X1 U4086 ( .A(n6072), .ZN(n3191) );
  AND2_X1 U4087 ( .A1(n3271), .A2(n3630), .ZN(n3109) );
  AND2_X1 U4088 ( .A1(n6070), .A2(n3884), .ZN(n3110) );
  NOR2_X1 U4089 ( .A1(n5281), .A2(n5280), .ZN(n5265) );
  INV_X1 U4090 ( .A(n3200), .ZN(n3199) );
  OAI21_X1 U4091 ( .B1(n3670), .B2(n3095), .A(n3673), .ZN(n3200) );
  AND2_X1 U4092 ( .A1(n3664), .A2(n3662), .ZN(n3111) );
  XOR2_X1 U4093 ( .A(n3157), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n3112) );
  AND2_X1 U4094 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3113)
         );
  NAND2_X1 U4095 ( .A1(n5681), .A2(n4422), .ZN(n3114) );
  NOR2_X1 U4096 ( .A1(n5777), .A2(n4415), .ZN(n3115) );
  AND2_X1 U4097 ( .A1(n5876), .A2(n5867), .ZN(n3116) );
  NAND2_X1 U4098 ( .A1(n5459), .A2(n5461), .ZN(n5448) );
  XNOR2_X1 U4099 ( .A(n3482), .B(n3533), .ZN(n4698) );
  OR2_X1 U4100 ( .A1(n5777), .A2(n3675), .ZN(n3117) );
  NOR2_X1 U4101 ( .A1(n3237), .A2(n3158), .ZN(n3234) );
  NAND2_X1 U4102 ( .A1(n5733), .A2(n5734), .ZN(n3118) );
  INV_X1 U4103 ( .A(n3593), .ZN(n3166) );
  XNOR2_X1 U4104 ( .A(n3250), .B(n3249), .ZN(n4702) );
  AND2_X1 U4105 ( .A1(n3099), .A2(n3218), .ZN(n3119) );
  NOR2_X1 U4106 ( .A1(n5411), .A2(n5412), .ZN(n5381) );
  INV_X1 U4107 ( .A(n3789), .ZN(n4683) );
  AND2_X1 U4108 ( .A1(n4933), .A2(n3119), .ZN(n5482) );
  AND2_X1 U4109 ( .A1(n4933), .A2(n3219), .ZN(n4930) );
  AND2_X1 U4110 ( .A1(n3212), .A2(n4683), .ZN(n4688) );
  OR3_X1 U4111 ( .A1(n5337), .A2(n3843), .A3(n3217), .ZN(n3120) );
  AND2_X1 U4112 ( .A1(n3124), .A2(n3970), .ZN(n3121) );
  OAI211_X1 U4113 ( .C1(n3163), .C2(n3594), .A(n3161), .B(n3165), .ZN(n5119)
         );
  NAND2_X1 U4114 ( .A1(n3594), .A2(n3593), .ZN(n4950) );
  NAND2_X1 U4115 ( .A1(n3229), .A2(n3652), .ZN(n5866) );
  NAND3_X1 U4116 ( .A1(n3505), .A2(n3545), .A3(n3504), .ZN(n4783) );
  OAI21_X1 U4117 ( .B1(n3922), .B2(n3945), .A(n3921), .ZN(n4745) );
  NOR2_X1 U4118 ( .A1(n5615), .A2(n3096), .ZN(n5425) );
  NAND2_X1 U4119 ( .A1(n3896), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3945) );
  INV_X1 U4120 ( .A(n3945), .ZN(n4073) );
  NAND2_X1 U4121 ( .A1(n4615), .A2(n3911), .ZN(n4678) );
  AND2_X1 U4122 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3122)
         );
  AND2_X1 U4123 ( .A1(n4679), .A2(n3948), .ZN(n4901) );
  NAND2_X1 U4124 ( .A1(n3121), .A2(n3251), .ZN(n3123) );
  OAI21_X1 U4125 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n4906) );
  NAND2_X1 U4126 ( .A1(n3906), .A2(n3905), .ZN(n4614) );
  OR2_X1 U4127 ( .A1(n5207), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6075) );
  INV_X2 U4128 ( .A(n5885), .ZN(n6431) );
  INV_X1 U4129 ( .A(n5346), .ZN(n3262) );
  INV_X1 U4130 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4170) );
  NAND3_X1 U4131 ( .A1(n3988), .A2(n3987), .A3(n3986), .ZN(n3124) );
  NAND2_X1 U4132 ( .A1(n3393), .A2(n3391), .ZN(n4372) );
  INV_X1 U4133 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6902) );
  AND2_X1 U4134 ( .A1(n4479), .A2(n5278), .ZN(n3125) );
  INV_X1 U4135 ( .A(n5464), .ZN(n3145) );
  INV_X1 U4136 ( .A(REIP_REG_31__SCAN_IN), .ZN(n3142) );
  AND2_X1 U4137 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3126) );
  NAND2_X2 U4138 ( .A1(n4492), .A2(n3127), .ZN(n5586) );
  NOR2_X2 U4139 ( .A1(n4258), .A2(n4228), .ZN(n3128) );
  OAI21_X1 U4140 ( .B1(n5229), .B2(n5522), .A(n3138), .ZN(U2796) );
  NAND2_X2 U4141 ( .A1(n3551), .A2(n3552), .ZN(n3731) );
  AND2_X4 U4142 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4574) );
  NAND2_X2 U4143 ( .A1(n3189), .A2(n3741), .ZN(n4584) );
  NAND2_X1 U4145 ( .A1(n3896), .A2(n3389), .ZN(n3400) );
  NAND2_X1 U4146 ( .A1(n3152), .A2(n3669), .ZN(n3153) );
  NAND2_X1 U4147 ( .A1(n3230), .A2(n3231), .ZN(n5814) );
  NAND2_X1 U4148 ( .A1(n3505), .A2(n3504), .ZN(n3544) );
  NAND2_X1 U4149 ( .A1(n3934), .A2(n4073), .ZN(n3159) );
  XNOR2_X1 U4150 ( .A(n3592), .B(n3795), .ZN(n4860) );
  NAND2_X1 U4151 ( .A1(n3589), .A2(n3608), .ZN(n3922) );
  INV_X1 U4152 ( .A(n4951), .ZN(n3163) );
  NAND3_X1 U4153 ( .A1(n3164), .A2(n3162), .A3(n5120), .ZN(n3639) );
  NAND3_X1 U4154 ( .A1(n3594), .A2(n3165), .A3(n3593), .ZN(n3164) );
  INV_X1 U4155 ( .A(n4768), .ZN(n3203) );
  AND2_X2 U4156 ( .A1(n3203), .A2(n4790), .ZN(n3512) );
  INV_X1 U4157 ( .A(n4768), .ZN(n3201) );
  NOR2_X2 U4158 ( .A1(n4900), .A2(n3123), .ZN(n5459) );
  AND2_X2 U4159 ( .A1(n3243), .A2(n3241), .ZN(n5752) );
  OR2_X2 U4160 ( .A1(n5732), .A2(n3676), .ZN(n3243) );
  NAND2_X1 U4161 ( .A1(n5249), .A2(n3170), .ZN(n5231) );
  AND2_X2 U4162 ( .A1(n3348), .A2(n3398), .ZN(n4589) );
  INV_X2 U4163 ( .A(n4724), .ZN(n3771) );
  NAND2_X1 U4164 ( .A1(n3176), .A2(n3174), .ZN(n3177) );
  INV_X1 U4165 ( .A(n3175), .ZN(n3174) );
  OAI22_X1 U4166 ( .A1(n3696), .A2(n3695), .B1(n3739), .B2(n3757), .ZN(n3175)
         );
  NAND3_X1 U4167 ( .A1(n3691), .A2(n3692), .A3(n3178), .ZN(n3176) );
  NAND2_X1 U4168 ( .A1(n3177), .A2(n3181), .ZN(n3180) );
  NAND2_X1 U4169 ( .A1(n3180), .A2(n3179), .ZN(n3716) );
  NAND4_X1 U4170 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(U2987)
         );
  NAND3_X1 U4171 ( .A1(n5901), .A2(n5893), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3183) );
  NAND3_X1 U4172 ( .A1(n3738), .A2(n3736), .A3(n3737), .ZN(n3189) );
  NAND2_X1 U4173 ( .A1(n3225), .A2(n3226), .ZN(n5859) );
  NOR2_X1 U4174 ( .A1(n3227), .A2(n3663), .ZN(n3194) );
  OAI21_X1 U4175 ( .B1(n5775), .B2(n3095), .A(n3199), .ZN(n5767) );
  NAND2_X2 U4176 ( .A1(n3495), .A2(n3494), .ZN(n3892) );
  AND2_X2 U4177 ( .A1(n3203), .A2(n4574), .ZN(n3436) );
  INV_X2 U4178 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3202) );
  AND2_X2 U4179 ( .A1(n3201), .A2(n5179), .ZN(n3517) );
  AND2_X2 U4180 ( .A1(n3201), .A2(n5178), .ZN(n3431) );
  INV_X1 U4181 ( .A(n5615), .ZN(n3204) );
  NAND2_X1 U4182 ( .A1(n3204), .A2(n3205), .ZN(n5411) );
  NAND2_X1 U4183 ( .A1(n4749), .A2(n4682), .ZN(n3210) );
  NAND2_X1 U4184 ( .A1(n4683), .A2(n3211), .ZN(n4750) );
  OAI22_X1 U4185 ( .A1(n5221), .A2(n5354), .B1(n4395), .B2(n5220), .ZN(n3215)
         );
  NOR2_X2 U4186 ( .A1(n4395), .A2(n5218), .ZN(n5221) );
  NOR3_X4 U4187 ( .A1(n5337), .A2(n3216), .A3(n3843), .ZN(n3853) );
  NAND4_X1 U4188 ( .A1(n3744), .A2(n3403), .A3(n3222), .A4(n3221), .ZN(n3404)
         );
  AND2_X4 U4189 ( .A1(n3399), .A2(n3780), .ZN(n4469) );
  NAND2_X1 U4190 ( .A1(n3398), .A2(n3422), .ZN(n3746) );
  NAND2_X1 U4191 ( .A1(n5875), .A2(n3116), .ZN(n3225) );
  NAND2_X1 U4192 ( .A1(n5830), .A2(n3234), .ZN(n3230) );
  INV_X1 U4193 ( .A(n3676), .ZN(n3247) );
  AND2_X4 U4194 ( .A1(n5178), .A2(n4763), .ZN(n3379) );
  AND2_X2 U4195 ( .A1(n5178), .A2(n4762), .ZN(n3444) );
  AND2_X2 U4196 ( .A1(n3291), .A2(n5178), .ZN(n3577) );
  NAND2_X2 U4197 ( .A1(n3248), .A2(n3443), .ZN(n3531) );
  NAND2_X1 U4198 ( .A1(n4702), .A2(n6642), .ZN(n3248) );
  NAND2_X1 U4199 ( .A1(n3608), .A2(n3607), .ZN(n3612) );
  NAND4_X1 U4200 ( .A1(n4699), .A2(n3568), .A3(n3588), .A4(n3567), .ZN(n3608)
         );
  NAND3_X1 U4201 ( .A1(n4699), .A2(n3568), .A3(n3567), .ZN(n3609) );
  NAND2_X1 U4202 ( .A1(n3254), .A2(n3253), .ZN(n5366) );
  CLKBUF_X1 U4203 ( .A(n3254), .Z(n3252) );
  NAND2_X1 U4204 ( .A1(n4499), .A2(n3263), .ZN(n3267) );
  INV_X1 U4205 ( .A(n5689), .ZN(n5197) );
  NAND2_X1 U4206 ( .A1(n5689), .A2(n4380), .ZN(n4405) );
  NAND2_X1 U4207 ( .A1(n5752), .A2(n3680), .ZN(n3685) );
  NAND2_X1 U4208 ( .A1(n3506), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3407) );
  NAND2_X1 U4209 ( .A1(n3882), .A2(n3779), .ZN(n6088) );
  INV_X1 U4210 ( .A(n6088), .ZN(n6463) );
  INV_X2 U4211 ( .A(n4629), .ZN(n4692) );
  INV_X1 U4212 ( .A(n5892), .ZN(n4424) );
  INV_X1 U4213 ( .A(n3655), .ZN(n3671) );
  INV_X1 U4214 ( .A(n5300), .ZN(n5314) );
  INV_X1 U4215 ( .A(n5732), .ZN(n5733) );
  NOR2_X1 U4216 ( .A1(n3950), .A2(n3935), .ZN(n3269) );
  AND3_X1 U4217 ( .A1(n3771), .A2(n4526), .A3(n3147), .ZN(n3270) );
  AND2_X1 U4218 ( .A1(n3611), .A2(n3588), .ZN(n3271) );
  NOR2_X2 U4219 ( .A1(n5018), .A2(n6099), .ZN(n3272) );
  OR2_X1 U4220 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3273)
         );
  NOR2_X1 U4221 ( .A1(n6097), .A2(n6101), .ZN(n3275) );
  NOR2_X1 U4222 ( .A1(n5840), .A2(n5831), .ZN(n3276) );
  INV_X1 U4223 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5769) );
  INV_X1 U4224 ( .A(n4227), .ZN(n5302) );
  NAND2_X1 U4225 ( .A1(n5618), .A2(n5191), .ZN(n5620) );
  INV_X1 U4226 ( .A(n5620), .ZN(n4402) );
  NOR2_X1 U4227 ( .A1(n3422), .A2(n6326), .ZN(n4097) );
  NOR2_X1 U4228 ( .A1(n6477), .A2(n6112), .ZN(n3277) );
  OR2_X1 U4229 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3278)
         );
  OR3_X1 U4230 ( .A1(n3684), .A2(n3683), .A3(n3889), .ZN(n3279) );
  INV_X1 U4231 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4437) );
  AND2_X1 U4232 ( .A1(n4724), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3280) );
  INV_X1 U4233 ( .A(n3804), .ZN(n3846) );
  OR2_X1 U4234 ( .A1(n3410), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3411)
         );
  INV_X1 U4235 ( .A(n3400), .ZN(n3747) );
  NAND2_X1 U4236 ( .A1(n3369), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3370) );
  INV_X1 U4237 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U4238 ( .A1(n3462), .A2(n3460), .ZN(n3503) );
  INV_X1 U4239 ( .A(n3415), .ZN(n3416) );
  AOI22_X1 U4240 ( .A1(n3449), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3374) );
  INV_X1 U4241 ( .A(n4081), .ZN(n4082) );
  INV_X1 U4242 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4334) );
  OR2_X1 U4243 ( .A1(n3629), .A2(n3628), .ZN(n3645) );
  INV_X1 U4244 ( .A(n3526), .ZN(n3538) );
  INV_X1 U4245 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4246 ( .A1(n3723), .A2(n3483), .ZN(n3739) );
  INV_X1 U4247 ( .A(n4447), .ZN(n4394) );
  OR2_X1 U4248 ( .A1(n4312), .A2(n4311), .ZN(n4329) );
  INV_X1 U4249 ( .A(n4965), .ZN(n3970) );
  INV_X1 U4250 ( .A(n5367), .ZN(n4135) );
  NAND2_X1 U4251 ( .A1(n4518), .A2(n4630), .ZN(n3775) );
  AND4_X1 U4252 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3365)
         );
  OR2_X1 U4253 ( .A1(n4782), .A2(n6991), .ZN(n4788) );
  OR2_X1 U4254 ( .A1(n4463), .A2(n6633), .ZN(n4464) );
  NAND2_X2 U4255 ( .A1(n3100), .A2(n3083), .ZN(n4628) );
  AND2_X1 U4256 ( .A1(n4120), .A2(n4119), .ZN(n5377) );
  INV_X1 U4257 ( .A(n5406), .ZN(n5407) );
  INV_X1 U4258 ( .A(n5896), .ZN(n5897) );
  AND2_X1 U4259 ( .A1(n5708), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4440)
         );
  INV_X1 U4260 ( .A(n5718), .ZN(n4420) );
  INV_X1 U4261 ( .A(n3483), .ZN(n3724) );
  NAND2_X1 U4262 ( .A1(n6635), .A2(n4706), .ZN(n4707) );
  INV_X1 U4263 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4776) );
  AND2_X1 U4264 ( .A1(n4911), .A2(n6484), .ZN(n4917) );
  AND2_X1 U4265 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5076), .ZN(n5005)
         );
  NAND2_X1 U4266 ( .A1(n3740), .A2(n3759), .ZN(n3741) );
  INV_X1 U4267 ( .A(n4458), .ZN(n4515) );
  AND2_X1 U4268 ( .A1(n6396), .A2(n5685), .ZN(n4493) );
  INV_X1 U4269 ( .A(n6393), .ZN(n5517) );
  INV_X1 U4270 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3942) );
  INV_X1 U4271 ( .A(n4409), .ZN(n4410) );
  INV_X1 U4272 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6878) );
  INV_X1 U4273 ( .A(n6424), .ZN(n5884) );
  NAND2_X1 U4274 ( .A1(n5691), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5682) );
  AND2_X1 U4275 ( .A1(n5777), .A2(n5964), .ZN(n5741) );
  NAND2_X1 U4276 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3674) );
  AND2_X1 U4277 ( .A1(n5830), .A2(n5850), .ZN(n5843) );
  NAND2_X1 U4278 ( .A1(n3490), .A2(n3489), .ZN(n4636) );
  OR2_X1 U4279 ( .A1(n5052), .A2(n6099), .ZN(n5058) );
  OAI21_X1 U4280 ( .B1(n5136), .B2(n6643), .A(n6484), .ZN(n6205) );
  NAND2_X1 U4281 ( .A1(n4847), .A2(n4920), .ZN(n6590) );
  INV_X1 U4282 ( .A(n4977), .ZN(n5007) );
  INV_X1 U4283 ( .A(n6524), .ZN(n6559) );
  INV_X1 U4284 ( .A(n6532), .ZN(n6257) );
  AND2_X1 U4285 ( .A1(n4781), .A2(n4780), .ZN(n6624) );
  OR2_X1 U4286 ( .A1(n4494), .A2(n4493), .ZN(n4495) );
  AND2_X1 U4287 ( .A1(n4012), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4015)
         );
  NAND2_X1 U4288 ( .A1(n5577), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4491) );
  AND2_X1 U4289 ( .A1(n5678), .A2(n5191), .ZN(n5192) );
  NOR2_X1 U4290 ( .A1(n4553), .A2(n4526), .ZN(n6409) );
  NOR2_X2 U4291 ( .A1(n4792), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6744) );
  INV_X1 U4292 ( .A(n6084), .ZN(n4444) );
  INV_X1 U4293 ( .A(n5743), .ZN(n5744) );
  XNOR2_X1 U4294 ( .A(n3500), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4638)
         );
  INV_X1 U4295 ( .A(n6113), .ZN(n5077) );
  OAI21_X1 U4296 ( .B1(n6117), .B2(n6116), .A(n6115), .ZN(n6154) );
  NOR2_X2 U4297 ( .A1(n5058), .A2(n6291), .ZN(n6159) );
  OAI21_X1 U4298 ( .B1(n6166), .B2(n6165), .A(n6325), .ZN(n6191) );
  OAI21_X1 U4299 ( .B1(n5024), .B2(n5023), .A(n5022), .ZN(n5047) );
  INV_X1 U4300 ( .A(n6206), .ZN(n6234) );
  INV_X1 U4301 ( .A(n4913), .ZN(n6549) );
  AND2_X1 U4302 ( .A1(n5128), .A2(n4920), .ZN(n6551) );
  AND2_X1 U4303 ( .A1(n4737), .A2(n4736), .ZN(n6528) );
  XNOR2_X1 U4304 ( .A(n6281), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6477)
         );
  NOR2_X1 U4305 ( .A1(n4822), .A2(n5077), .ZN(n6544) );
  AND2_X1 U4306 ( .A1(n6238), .A2(n3892), .ZN(n4910) );
  INV_X1 U4307 ( .A(n6565), .ZN(n6491) );
  INV_X1 U4308 ( .A(n6579), .ZN(n6501) );
  INV_X1 U4309 ( .A(n6598), .ZN(n6520) );
  OAI211_X1 U4310 ( .C1(n4893), .C2(n6725), .A(n4833), .B(n4832), .ZN(n4898)
         );
  INV_X1 U4311 ( .A(n6574), .ZN(n6539) );
  INV_X1 U4312 ( .A(n6515), .ZN(n6550) );
  AND2_X1 U4313 ( .A1(n3764), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6640) );
  INV_X1 U4314 ( .A(STATE_REG_0__SCAN_IN), .ZN(n3752) );
  INV_X1 U4315 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6673) );
  INV_X1 U4316 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6643) );
  NOR2_X1 U4317 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  INV_X1 U4318 ( .A(n5792), .ZN(n5659) );
  NAND2_X1 U4319 ( .A1(n4813), .A2(n4812), .ZN(n5678) );
  NAND2_X2 U4320 ( .A1(n5678), .A2(n4815), .ZN(n5680) );
  INV_X1 U4321 ( .A(n6409), .ZN(n4572) );
  INV_X1 U4322 ( .A(n6744), .ZN(n5208) );
  INV_X1 U4323 ( .A(n6746), .ZN(n6408) );
  INV_X1 U4324 ( .A(n4433), .ZN(n4434) );
  INV_X1 U4325 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6932) );
  AND2_X1 U4326 ( .A1(n6019), .A2(n6018), .ZN(n6444) );
  NAND2_X1 U4327 ( .A1(n3882), .A2(n3777), .ZN(n6084) );
  NAND2_X1 U4328 ( .A1(n5053), .A2(n6291), .ZN(n6197) );
  AOI22_X1 U4329 ( .A1(n5021), .A2(n5023), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5017), .ZN(n5050) );
  OR2_X1 U4330 ( .A1(n5136), .A2(n6291), .ZN(n6237) );
  AOI211_X2 U4331 ( .C1(n6201), .C2(n6284), .A(n5133), .B(n5132), .ZN(n5170)
         );
  NAND2_X1 U4332 ( .A1(n5128), .A2(n4910), .ZN(n6557) );
  NAND2_X1 U4333 ( .A1(n6292), .A2(n3892), .ZN(n6314) );
  INV_X1 U4334 ( .A(n6583), .ZN(n6350) );
  INV_X1 U4335 ( .A(n6553), .ZN(n6354) );
  NOR2_X1 U4336 ( .A1(n5079), .A2(n5078), .ZN(n5118) );
  NAND2_X1 U4337 ( .A1(n6431), .A2(DATAI_21_), .ZN(n6581) );
  NAND2_X1 U4338 ( .A1(n6431), .A2(DATAI_24_), .ZN(n6565) );
  NAND2_X1 U4339 ( .A1(n6431), .A2(DATAI_27_), .ZN(n6579) );
  NAND2_X1 U4340 ( .A1(n6431), .A2(DATAI_31_), .ZN(n6598) );
  OAI221_X1 U4341 ( .B1(n6673), .B2(n3752), .C1(STATE_REG_1__SCAN_IN), .C2(
        n3752), .A(n6743), .ZN(n6654) );
  INV_X1 U4342 ( .A(n6722), .ZN(n6655) );
  INV_X1 U4343 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6690) );
  CLKBUF_X1 U4344 ( .A(n6716), .Z(n6705) );
  INV_X1 U4345 ( .A(n6709), .ZN(n6716) );
  OAI21_X1 U4346 ( .B1(n5197), .B2(n5522), .A(n4497), .ZN(U2797) );
  INV_X1 U4347 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3281) );
  AND2_X2 U4348 ( .A1(n5179), .A2(n4762), .ZN(n3377) );
  AOI22_X1 U4349 ( .A1(n3577), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3285) );
  AND2_X4 U4350 ( .A1(n3291), .A2(n4574), .ZN(n3369) );
  AND2_X4 U4351 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4763) );
  NOR2_X4 U4352 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U4353 ( .A1(n3369), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4354 ( .A1(n3285), .A2(n3284), .ZN(n3290) );
  AND2_X4 U4355 ( .A1(n4763), .A2(n4574), .ZN(n3372) );
  NAND2_X1 U4356 ( .A1(n3372), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3287)
         );
  NAND2_X1 U4357 ( .A1(n3431), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3286)
         );
  NAND3_X1 U4358 ( .A1(n3288), .A2(n3287), .A3(n3286), .ZN(n3289) );
  AND2_X2 U4359 ( .A1(n4762), .A2(n4790), .ZN(n3378) );
  AOI22_X1 U4360 ( .A1(n3512), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3295) );
  AND2_X2 U4361 ( .A1(n3291), .A2(n4790), .ZN(n3464) );
  AND2_X4 U4362 ( .A1(n5179), .A2(n4763), .ZN(n3518) );
  AOI22_X1 U4363 ( .A1(n3464), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3294) );
  AND2_X4 U4364 ( .A1(n4574), .A2(n4762), .ZN(n4346) );
  AOI22_X1 U4365 ( .A1(n3436), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3293) );
  AND2_X4 U4366 ( .A1(n5179), .A2(n3291), .ZN(n3449) );
  AOI22_X1 U4367 ( .A1(n3436), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4368 ( .A1(n3444), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4369 ( .A1(n3379), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4370 ( .A1(n3517), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4371 ( .A1(n3449), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4372 ( .A1(n3431), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3301) );
  NAND2_X2 U4373 ( .A1(n3306), .A2(n3305), .ZN(n3389) );
  AOI22_X1 U4374 ( .A1(n3577), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4375 ( .A1(n3444), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4376 ( .A1(n3379), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4378 ( .A1(n3517), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4379 ( .A1(n3449), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4380 ( .A1(n3431), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3314) );
  AND4_X2 U4381 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3317)
         );
  AOI22_X1 U4382 ( .A1(n3449), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4383 ( .A1(n3436), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4384 ( .A1(n3431), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4385 ( .A1(n3444), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3319) );
  AND4_X2 U4386 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3328)
         );
  AOI22_X1 U4387 ( .A1(n3577), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4388 ( .A1(n3517), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4389 ( .A1(n3379), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4390 ( .A1(n3369), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4391 ( .A1(n3436), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4392 ( .A1(n3577), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4393 ( .A1(n3444), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4394 ( .A1(n3379), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4395 ( .A1(n3517), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4396 ( .A1(n3449), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4397 ( .A1(n3431), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4398 ( .A1(n3859), .A2(n4728), .ZN(n3485) );
  AOI22_X1 U4399 ( .A1(n3436), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4400 ( .A1(n3577), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4401 ( .A1(n3444), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4402 ( .A1(n3379), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4403 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3347)
         );
  AOI22_X1 U4404 ( .A1(n3369), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4405 ( .A1(n3517), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4406 ( .A1(n3449), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4407 ( .A1(n3431), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4408 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  OR2_X2 U4409 ( .A1(n3347), .A2(n3346), .ZN(n3422) );
  NAND2_X1 U4410 ( .A1(n3391), .A2(n3422), .ZN(n4817) );
  NOR2_X1 U4411 ( .A1(n3485), .A2(n4817), .ZN(n3348) );
  NAND2_X1 U4412 ( .A1(n3444), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4413 ( .A1(n3430), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3350)
         );
  NAND2_X1 U4414 ( .A1(n3436), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3349)
         );
  NAND3_X1 U4415 ( .A1(n3351), .A2(n3350), .A3(n3349), .ZN(n3352) );
  AOI21_X2 U4416 ( .B1(n3577), .B2(INSTQUEUE_REG_6__0__SCAN_IN), .A(n3352), 
        .ZN(n3368) );
  NAND2_X1 U4417 ( .A1(n3449), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4418 ( .A1(n3431), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3355)
         );
  NAND2_X1 U4419 ( .A1(n3379), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3354)
         );
  NAND2_X1 U4420 ( .A1(n3518), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3353)
         );
  NAND2_X1 U4421 ( .A1(n3464), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3360) );
  NAND2_X1 U4422 ( .A1(n3517), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4423 ( .A1(n3369), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3358) );
  BUF_X4 U4424 ( .A(n3372), .Z(n4317) );
  NAND2_X1 U4425 ( .A1(n4317), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3357)
         );
  AND4_X2 U4426 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3366)
         );
  NAND2_X1 U4427 ( .A1(n3512), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4428 ( .A1(n3377), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4429 ( .A1(n3378), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U4430 ( .A1(n4346), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3361) );
  NAND4_X4 U4431 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3780)
         );
  AOI22_X1 U4432 ( .A1(n3517), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4433 ( .A1(n3518), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3371)
         );
  AOI22_X1 U4434 ( .A1(n3431), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4435 ( .A1(n3436), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3512), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4436 ( .A1(n3577), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4437 ( .A1(n3444), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4438 ( .A1(n3379), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3380) );
  XNOR2_X1 U4439 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3751) );
  NAND2_X1 U4440 ( .A1(n3399), .A2(n3751), .ZN(n3402) );
  XNOR2_X1 U4441 ( .A(n3389), .B(n3401), .ZN(n3388) );
  NAND2_X1 U4442 ( .A1(n3401), .A2(n4724), .ZN(n3385) );
  OAI211_X1 U4443 ( .C1(n3393), .C2(n4724), .A(n3385), .B(n3422), .ZN(n3386)
         );
  INV_X1 U4444 ( .A(n3386), .ZN(n3387) );
  INV_X1 U4445 ( .A(n3395), .ZN(n3390) );
  INV_X2 U4446 ( .A(n3780), .ZN(n4526) );
  NOR2_X1 U4447 ( .A1(n4628), .A2(n3780), .ZN(n3770) );
  BUF_X1 U4448 ( .A(n3391), .Z(n3392) );
  NAND3_X1 U4449 ( .A1(n3770), .A2(n4375), .A3(n3392), .ZN(n4807) );
  NAND2_X1 U4450 ( .A1(n3393), .A2(n3422), .ZN(n4814) );
  NAND3_X1 U4451 ( .A1(n3394), .A2(n3775), .A3(n3778), .ZN(n3413) );
  NAND2_X1 U4452 ( .A1(n3413), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4453 ( .A1(n3723), .A2(n3400), .ZN(n3396) );
  OAI21_X1 U4454 ( .B1(n3419), .B2(n3551), .A(n3396), .ZN(n3397) );
  INV_X1 U4455 ( .A(n3397), .ZN(n3406) );
  NAND2_X1 U4456 ( .A1(n3404), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3405) );
  NAND2_X2 U4457 ( .A1(n3406), .A2(n3405), .ZN(n3506) );
  INV_X1 U4458 ( .A(n5207), .ZN(n3414) );
  INV_X1 U4459 ( .A(n3764), .ZN(n4373) );
  AOI22_X1 U4460 ( .A1(n3414), .A2(n6477), .B1(n4373), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3409) );
  INV_X1 U4461 ( .A(n3409), .ZN(n3410) );
  NAND2_X1 U4462 ( .A1(n3413), .A2(n3412), .ZN(n3502) );
  NAND2_X1 U4463 ( .A1(n3506), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3417) );
  MUX2_X1 U4464 ( .A(n4373), .B(n3414), .S(n6281), .Z(n3415) );
  NAND2_X1 U4465 ( .A1(n3417), .A2(n3416), .ZN(n3462) );
  NOR2_X1 U4466 ( .A1(n3419), .A2(n3418), .ZN(n3421) );
  NAND2_X1 U4467 ( .A1(n3780), .A2(n3859), .ZN(n3420) );
  NAND2_X1 U4468 ( .A1(n3421), .A2(n3420), .ZN(n3865) );
  INV_X1 U4469 ( .A(n3743), .ZN(n3893) );
  NAND4_X1 U4470 ( .A1(n3893), .A2(n4526), .A3(n4375), .A4(n4724), .ZN(n4770)
         );
  INV_X1 U4471 ( .A(n6734), .ZN(n6364) );
  NAND2_X1 U4472 ( .A1(n3423), .A2(n4469), .ZN(n3424) );
  NAND4_X1 U4473 ( .A1(n4770), .A2(n6364), .A3(STATE2_REG_0__SCAN_IN), .A4(
        n3424), .ZN(n3425) );
  NOR2_X1 U4474 ( .A1(n3107), .A2(n3425), .ZN(n3429) );
  INV_X1 U4475 ( .A(n3744), .ZN(n3427) );
  AND2_X1 U4476 ( .A1(n3400), .A2(n4724), .ZN(n3426) );
  OAI21_X1 U4477 ( .B1(n3427), .B2(n3426), .A(n4736), .ZN(n3428) );
  NAND3_X1 U4478 ( .A1(n3865), .A2(n3429), .A3(n3428), .ZN(n3460) );
  AOI22_X1 U4479 ( .A1(n4347), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4480 ( .A1(n3449), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4481 ( .A1(n3557), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4482 ( .A1(n4086), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4483 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3442)
         );
  AOI22_X1 U4484 ( .A1(n3577), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4485 ( .A1(n4345), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4486 ( .A1(n4322), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4487 ( .A1(n3085), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4488 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3441)
         );
  NAND2_X1 U4489 ( .A1(n3149), .A2(n3484), .ZN(n3443) );
  AOI22_X1 U4490 ( .A1(n4322), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4491 ( .A1(n3086), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4492 ( .A1(n3444), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4493 ( .A1(n4352), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3445) );
  NAND4_X1 U4494 ( .A1(n3448), .A2(n3447), .A3(n3446), .A4(n3445), .ZN(n3455)
         );
  AOI22_X1 U4495 ( .A1(n3085), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4496 ( .A1(n4306), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4497 ( .A1(n3449), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3430), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4498 ( .A1(n4086), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3450) );
  NAND4_X1 U4499 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3454)
         );
  INV_X1 U4500 ( .A(n3656), .ZN(n3456) );
  NAND2_X1 U4501 ( .A1(n3149), .A2(n3456), .ZN(n3476) );
  INV_X1 U4502 ( .A(n3551), .ZN(n3457) );
  NAND2_X1 U4503 ( .A1(n3457), .A2(n3484), .ZN(n3458) );
  OAI211_X1 U4504 ( .C1(n3459), .C2(n3714), .A(n3476), .B(n3458), .ZN(n3532)
         );
  INV_X1 U4505 ( .A(n3460), .ZN(n3461) );
  XNOR2_X1 U4506 ( .A(n3462), .B(n3461), .ZN(n3894) );
  NAND2_X1 U4507 ( .A1(n3894), .A2(n6642), .ZN(n3477) );
  INV_X1 U4508 ( .A(n3436), .ZN(n3463) );
  INV_X2 U4509 ( .A(n3463), .ZN(n4322) );
  AOI22_X1 U4510 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4322), .B1(n3085), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4511 ( .A1(n3464), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4512 ( .A1(n3444), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4513 ( .A1(n4086), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3465) );
  NAND4_X1 U4514 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3474)
         );
  AOI22_X1 U4515 ( .A1(n3086), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4516 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3449), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4517 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4347), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4518 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3557), .B1(n3430), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3469) );
  NAND4_X1 U4519 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), .ZN(n3473)
         );
  INV_X1 U4520 ( .A(n3497), .ZN(n3475) );
  MUX2_X1 U4521 ( .A(n3476), .B(n3653), .S(n3475), .Z(n3493) );
  NAND2_X1 U4522 ( .A1(n3477), .A2(n3493), .ZN(n3481) );
  AOI21_X1 U4523 ( .B1(n3771), .B2(n3656), .A(n6642), .ZN(n3479) );
  NAND2_X1 U4524 ( .A1(n4526), .A2(n3497), .ZN(n3478) );
  NAND2_X1 U4525 ( .A1(n4698), .A2(n3483), .ZN(n3490) );
  NAND2_X1 U4526 ( .A1(n3484), .A2(n3497), .ZN(n3537) );
  OAI21_X1 U4527 ( .B1(n3497), .B2(n3484), .A(n3537), .ZN(n3487) );
  INV_X1 U4528 ( .A(n4469), .ZN(n5201) );
  INV_X1 U4529 ( .A(n3857), .ZN(n3486) );
  OAI211_X1 U4530 ( .C1(n3487), .C2(n5201), .A(n3486), .B(n3147), .ZN(n3488)
         );
  INV_X1 U4531 ( .A(n3488), .ZN(n3489) );
  INV_X1 U4532 ( .A(n3491), .ZN(n3492) );
  NAND2_X1 U4533 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  AND2_X1 U4534 ( .A1(n4526), .A2(n4728), .ZN(n3539) );
  INV_X1 U4535 ( .A(n3539), .ZN(n3496) );
  OAI21_X1 U4536 ( .B1(n5201), .B2(n3497), .A(n3496), .ZN(n3498) );
  INV_X1 U4537 ( .A(n3498), .ZN(n3499) );
  NAND2_X1 U4538 ( .A1(n4636), .A2(n4638), .ZN(n4637) );
  NAND2_X1 U4539 ( .A1(n4637), .A2(n3501), .ZN(n6430) );
  NAND2_X1 U4540 ( .A1(n3503), .A2(n3502), .ZN(n3505) );
  NAND2_X1 U4541 ( .A1(n3507), .A2(n6610), .ZN(n5014) );
  INV_X1 U4542 ( .A(n3507), .ZN(n3508) );
  NAND2_X1 U4543 ( .A1(n3508), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3509) );
  OAI22_X1 U4544 ( .A1(n4835), .A2(n5207), .B1(n3764), .B2(n6610), .ZN(n3510)
         );
  AOI21_X1 U4545 ( .B1(n3506), .B2(n6980), .A(n3510), .ZN(n3511) );
  INV_X1 U4546 ( .A(n3511), .ZN(n3545) );
  INV_X1 U4547 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4548 ( .A1(n4322), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4549 ( .A1(n3577), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3515) );
  INV_X1 U4550 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6887) );
  AOI22_X1 U4551 ( .A1(n4343), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4552 ( .A1(n4352), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4553 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3524)
         );
  AOI22_X1 U4554 ( .A1(n3085), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4555 ( .A1(n4306), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4556 ( .A1(n3449), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4557 ( .A1(n4086), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4558 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3523)
         );
  OAI22_X1 U4559 ( .A1(n3714), .A2(n3525), .B1(n3538), .B2(n3551), .ZN(n3528)
         );
  AND2_X1 U4560 ( .A1(n3149), .A2(n3526), .ZN(n3527) );
  XNOR2_X1 U4561 ( .A(n3528), .B(n3527), .ZN(n3529) );
  INV_X1 U4562 ( .A(n3567), .ZN(n3536) );
  OAI21_X2 U4563 ( .B1(n3533), .B2(n3532), .A(n3531), .ZN(n3535) );
  NAND2_X1 U4564 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  NAND2_X2 U4565 ( .A1(n3535), .A2(n3534), .ZN(n3568) );
  XNOR2_X1 U4566 ( .A(n3536), .B(n3568), .ZN(n3907) );
  NAND2_X1 U4567 ( .A1(n3907), .A2(n3483), .ZN(n3542) );
  NAND2_X1 U4568 ( .A1(n3537), .A2(n3538), .ZN(n3570) );
  OAI21_X1 U4569 ( .B1(n3538), .B2(n3537), .A(n3570), .ZN(n3540) );
  AOI21_X1 U4570 ( .B1(n3540), .B2(n4469), .A(n3539), .ZN(n3541) );
  NAND2_X1 U4571 ( .A1(n3542), .A2(n3541), .ZN(n3543) );
  AND2_X1 U4572 ( .A1(n3543), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6426)
         );
  OR2_X1 U4573 ( .A1(n3543), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6427)
         );
  NAND2_X1 U4574 ( .A1(n3568), .A2(n3567), .ZN(n3566) );
  NAND2_X1 U4575 ( .A1(n3506), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3550) );
  NAND3_X1 U4576 ( .A1(n6839), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6481) );
  INV_X1 U4577 ( .A(n6481), .ZN(n3546) );
  NAND2_X1 U4578 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3546), .ZN(n4913) );
  NAND2_X1 U4579 ( .A1(n6839), .A2(n4913), .ZN(n3547) );
  NAND2_X1 U4580 ( .A1(n3547), .A2(n4738), .ZN(n6111) );
  OAI22_X1 U4581 ( .A1(n5207), .A2(n6111), .B1(n3764), .B2(n6839), .ZN(n3548)
         );
  INV_X1 U4582 ( .A(n3548), .ZN(n3549) );
  NAND2_X1 U4583 ( .A1(n4701), .A2(n6642), .ZN(n3565) );
  AOI22_X1 U4584 ( .A1(n4322), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4585 ( .A1(n3086), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4586 ( .A1(n4343), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4587 ( .A1(n4352), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3553) );
  NAND4_X1 U4588 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3563)
         );
  AOI22_X1 U4589 ( .A1(n3085), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4590 ( .A1(n4306), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4591 ( .A1(n3449), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4592 ( .A1(n4086), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4593 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3562)
         );
  AOI22_X1 U4594 ( .A1(n3731), .A2(n3571), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3723), .ZN(n3564) );
  INV_X1 U4595 ( .A(n4699), .ZN(n4796) );
  NAND2_X1 U4596 ( .A1(n3566), .A2(n4796), .ZN(n3569) );
  NAND2_X1 U4597 ( .A1(n3570), .A2(n3571), .ZN(n3615) );
  OAI211_X1 U4598 ( .C1(n3571), .C2(n3570), .A(n3615), .B(n4469), .ZN(n3572)
         );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3575) );
  OAI21_X2 U4600 ( .B1(n4753), .B2(n4754), .A(n3576), .ZN(n4859) );
  AOI22_X1 U4601 ( .A1(n4322), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4602 ( .A1(n4344), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4603 ( .A1(n4306), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4604 ( .A1(n4345), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4605 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3587)
         );
  AOI22_X1 U4606 ( .A1(n4343), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4607 ( .A1(n4347), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4608 ( .A1(n3085), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4609 ( .A1(n4086), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4610 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  AOI22_X1 U4611 ( .A1(n3731), .A2(n3613), .B1(n3723), .B2(
        INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3610) );
  INV_X1 U4612 ( .A(n3610), .ZN(n3588) );
  NAND2_X1 U4613 ( .A1(n3609), .A2(n3610), .ZN(n3589) );
  XNOR2_X1 U4614 ( .A(n3615), .B(n3613), .ZN(n3590) );
  NAND2_X1 U4615 ( .A1(n3590), .A2(n4469), .ZN(n3591) );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4617 ( .A1(n4859), .A2(n4860), .ZN(n3594) );
  NAND2_X1 U4618 ( .A1(n3592), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3593)
         );
  AOI22_X1 U4619 ( .A1(n4322), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4620 ( .A1(n3577), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4621 ( .A1(n4343), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4622 ( .A1(n4352), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4623 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3604)
         );
  INV_X1 U4624 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6888) );
  AOI22_X1 U4625 ( .A1(n3085), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4626 ( .A1(n4306), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4627 ( .A1(n4344), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4628 ( .A1(n4086), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4629 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  NAND2_X1 U4630 ( .A1(n3731), .A2(n3616), .ZN(n3606) );
  NAND2_X1 U4631 ( .A1(n3723), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4632 ( .A1(n3606), .A2(n3605), .ZN(n3611) );
  INV_X1 U4633 ( .A(n3611), .ZN(n3607) );
  NAND2_X1 U4634 ( .A1(n3612), .A2(n3632), .ZN(n3946) );
  INV_X1 U4635 ( .A(n3613), .ZN(n3614) );
  NOR2_X1 U4636 ( .A1(n3615), .A2(n3614), .ZN(n3617) );
  NAND2_X1 U4637 ( .A1(n3617), .A2(n3616), .ZN(n3644) );
  OAI211_X1 U4638 ( .C1(n3617), .C2(n3616), .A(n3644), .B(n4469), .ZN(n3618)
         );
  AOI22_X1 U4639 ( .A1(n4322), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4640 ( .A1(n4343), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4641 ( .A1(n4352), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4642 ( .A1(n3557), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3620) );
  NAND4_X1 U4643 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3629)
         );
  AOI22_X1 U4644 ( .A1(n3085), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4645 ( .A1(n4345), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4646 ( .A1(n3086), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4647 ( .A1(n4086), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4648 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3628)
         );
  AOI22_X1 U4649 ( .A1(n3731), .A2(n3645), .B1(n3723), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3631) );
  INV_X1 U4650 ( .A(n3631), .ZN(n3630) );
  NAND3_X1 U4651 ( .A1(n3643), .A2(n3483), .A3(n3934), .ZN(n3635) );
  XNOR2_X1 U4652 ( .A(n3644), .B(n3645), .ZN(n3633) );
  NAND2_X1 U4653 ( .A1(n3633), .A2(n4469), .ZN(n3634) );
  NAND2_X1 U4654 ( .A1(n3635), .A2(n3634), .ZN(n3637) );
  INV_X1 U4655 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3636) );
  XNOR2_X1 U4656 ( .A(n3637), .B(n3636), .ZN(n5120) );
  NAND2_X1 U4657 ( .A1(n3637), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3638)
         );
  NAND2_X1 U4658 ( .A1(n3639), .A2(n3638), .ZN(n5875) );
  INV_X1 U4659 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U4660 ( .A1(n3731), .A2(n3656), .ZN(n3640) );
  OAI21_X1 U4661 ( .B1(n3641), .B2(n3714), .A(n3640), .ZN(n3642) );
  NAND2_X1 U4662 ( .A1(n3949), .A2(n3483), .ZN(n3649) );
  INV_X1 U4663 ( .A(n3644), .ZN(n3646) );
  NAND2_X1 U4664 ( .A1(n3646), .A2(n3645), .ZN(n3658) );
  XNOR2_X1 U4665 ( .A(n3658), .B(n3656), .ZN(n3647) );
  NAND2_X1 U4666 ( .A1(n3647), .A2(n4469), .ZN(n3648) );
  NAND2_X1 U4667 ( .A1(n3649), .A2(n3648), .ZN(n3651) );
  INV_X1 U4668 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3650) );
  XNOR2_X1 U4669 ( .A(n3651), .B(n3650), .ZN(n5876) );
  NAND2_X1 U4670 ( .A1(n3651), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3652)
         );
  NOR2_X1 U4671 ( .A1(n3653), .A2(n3724), .ZN(n3654) );
  NAND2_X1 U4672 ( .A1(n3643), .A2(n3654), .ZN(n3655) );
  NAND2_X1 U4673 ( .A1(n4469), .A2(n3656), .ZN(n3657) );
  OR2_X1 U4674 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  NAND2_X1 U4675 ( .A1(n3655), .A2(n3659), .ZN(n3660) );
  INV_X1 U4676 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3805) );
  XNOR2_X1 U4677 ( .A(n3660), .B(n3805), .ZN(n5867) );
  NAND2_X1 U4678 ( .A1(n3660), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3661)
         );
  NOR2_X1 U4679 ( .A1(n5777), .A2(n6801), .ZN(n3663) );
  NAND2_X1 U4680 ( .A1(n5777), .A2(n6801), .ZN(n3662) );
  INV_X1 U4681 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3666) );
  AND2_X1 U4682 ( .A1(n5777), .A2(n3666), .ZN(n5851) );
  INV_X1 U4683 ( .A(n5851), .ZN(n3664) );
  INV_X1 U4684 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6443) );
  AND2_X1 U4685 ( .A1(n5777), .A2(n6443), .ZN(n5840) );
  INV_X1 U4686 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3665) );
  AND2_X1 U4687 ( .A1(n5777), .A2(n3665), .ZN(n5831) );
  NOR2_X1 U4688 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3667) );
  OR2_X1 U4689 ( .A1(n5777), .A2(n3667), .ZN(n3668) );
  INV_X1 U4690 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6044) );
  OR2_X1 U4691 ( .A1(n5777), .A2(n6044), .ZN(n3669) );
  NAND2_X1 U4692 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U4693 ( .A1(n5777), .A2(n6014), .ZN(n3670) );
  INV_X1 U4694 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6005) );
  INV_X1 U4695 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6003) );
  INV_X1 U4696 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5776) );
  NAND4_X1 U4697 ( .A1(n5787), .A2(n6005), .A3(n6003), .A4(n5776), .ZN(n3672)
         );
  NAND2_X1 U4698 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3856) );
  OAI21_X1 U4699 ( .B1(n5787), .B2(n3856), .A(n5777), .ZN(n3673) );
  XNOR2_X1 U4700 ( .A(n5777), .B(n6932), .ZN(n5768) );
  OR2_X2 U4701 ( .A1(n5767), .A2(n5768), .ZN(n5732) );
  NOR2_X1 U4702 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3676)
         );
  INV_X1 U4703 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3675) );
  XNOR2_X1 U4704 ( .A(n5832), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5754)
         );
  INV_X1 U4705 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5948) );
  INV_X1 U4706 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U4707 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3681) );
  NOR4_X1 U4708 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n3682), 
        .A4(n3681), .ZN(n3677) );
  AOI21_X1 U4709 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n5948), .A(n3677), 
        .ZN(n3678) );
  NOR2_X1 U4710 ( .A1(n5752), .A2(n3678), .ZN(n3687) );
  NOR2_X1 U4711 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5742)
         );
  AND2_X1 U4712 ( .A1(n5742), .A2(n5948), .ZN(n3684) );
  INV_X1 U4713 ( .A(n3684), .ZN(n3679) );
  AND2_X1 U4714 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4412) );
  INV_X1 U4715 ( .A(n4412), .ZN(n4450) );
  OAI21_X1 U4716 ( .B1(n3679), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n4450), 
        .ZN(n3680) );
  NOR3_X1 U4717 ( .A1(n5832), .A2(n3682), .A3(n3681), .ZN(n3683) );
  INV_X1 U4718 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3889) );
  NAND2_X1 U4719 ( .A1(n3685), .A2(n3279), .ZN(n3686) );
  NOR2_X1 U4720 ( .A1(n3687), .A2(n3686), .ZN(n5731) );
  XNOR2_X1 U4721 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4722 ( .A1(n6281), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3699) );
  XNOR2_X1 U4723 ( .A(n3700), .B(n3699), .ZN(n3757) );
  NAND2_X1 U4724 ( .A1(n3757), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3695) );
  INV_X1 U4725 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U4726 ( .A1(n6727), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U4727 ( .A1(n3699), .A2(n3688), .ZN(n3693) );
  AOI21_X1 U4728 ( .B1(n3149), .B2(n3147), .A(n3693), .ZN(n3690) );
  NAND2_X1 U4729 ( .A1(n3392), .A2(n3780), .ZN(n3689) );
  NAND2_X1 U4730 ( .A1(n3689), .A2(n4630), .ZN(n3698) );
  OAI21_X1 U4731 ( .B1(n3690), .B2(n4526), .A(n3698), .ZN(n3691) );
  INV_X1 U4732 ( .A(n3693), .ZN(n3694) );
  NAND2_X1 U4733 ( .A1(n3731), .A2(n3694), .ZN(n3697) );
  INV_X1 U4734 ( .A(n3698), .ZN(n3710) );
  INV_X1 U4735 ( .A(n3699), .ZN(n3701) );
  NAND2_X1 U4736 ( .A1(n3701), .A2(n3700), .ZN(n3703) );
  NAND2_X1 U4737 ( .A1(n7013), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4738 ( .A1(n3703), .A2(n3702), .ZN(n3707) );
  XNOR2_X1 U4739 ( .A(n3202), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3705)
         );
  XNOR2_X1 U4740 ( .A(n3707), .B(n3705), .ZN(n3756) );
  MUX2_X1 U4741 ( .A(n3723), .B(n3731), .S(n3756), .Z(n3704) );
  INV_X1 U4742 ( .A(n3705), .ZN(n3706) );
  NAND2_X1 U4743 ( .A1(n3707), .A2(n3706), .ZN(n3709) );
  NAND2_X1 U4744 ( .A1(n6610), .A2(n6980), .ZN(n3708) );
  NAND2_X1 U4745 ( .A1(n3709), .A2(n3708), .ZN(n3719) );
  XNOR2_X1 U4746 ( .A(n4776), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3717)
         );
  XNOR2_X1 U4747 ( .A(n3719), .B(n3717), .ZN(n3755) );
  INV_X1 U4748 ( .A(n3755), .ZN(n3713) );
  NAND2_X1 U4749 ( .A1(n3483), .A2(n3713), .ZN(n3712) );
  NAND3_X1 U4750 ( .A1(n3710), .A2(n3731), .A3(n3756), .ZN(n3711) );
  NAND2_X1 U4751 ( .A1(n3714), .A2(n3713), .ZN(n3715) );
  NAND2_X1 U4752 ( .A1(n3716), .A2(n3715), .ZN(n3732) );
  INV_X1 U4753 ( .A(n3717), .ZN(n3718) );
  NAND2_X1 U4754 ( .A1(n3719), .A2(n3718), .ZN(n3721) );
  NAND2_X1 U4755 ( .A1(n6839), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4756 ( .A1(n3721), .A2(n3720), .ZN(n3728) );
  NAND2_X1 U4757 ( .A1(n3732), .A2(n3733), .ZN(n3726) );
  OAI21_X1 U4758 ( .B1(n3731), .B2(n3724), .A(n3754), .ZN(n3725) );
  NAND2_X1 U4759 ( .A1(n3726), .A2(n3725), .ZN(n3738) );
  NAND2_X1 U4760 ( .A1(n3727), .A2(n6614), .ZN(n3730) );
  NAND2_X1 U4761 ( .A1(n3728), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U4762 ( .A1(n3731), .A2(n3759), .ZN(n3737) );
  INV_X1 U4763 ( .A(n3732), .ZN(n3735) );
  INV_X1 U4764 ( .A(n3733), .ZN(n3734) );
  NAND2_X1 U4765 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  NAND2_X1 U4766 ( .A1(n4724), .A2(n3147), .ZN(n3742) );
  NOR2_X1 U4767 ( .A1(n5180), .A2(n4630), .ZN(n3867) );
  INV_X1 U4768 ( .A(n3867), .ZN(n3763) );
  AOI21_X1 U4769 ( .B1(n5180), .B2(n4526), .A(n3401), .ZN(n3745) );
  NAND2_X1 U4770 ( .A1(n3744), .A2(n3745), .ZN(n3773) );
  OAI21_X1 U4771 ( .B1(n3747), .B2(n4526), .A(n5201), .ZN(n3748) );
  OAI21_X1 U4772 ( .B1(n3746), .B2(n3747), .A(n3748), .ZN(n3862) );
  INV_X1 U4773 ( .A(n3862), .ZN(n3749) );
  OR2_X1 U4774 ( .A1(n3773), .A2(n3749), .ZN(n3750) );
  NAND2_X1 U4775 ( .A1(n3750), .A2(n4459), .ZN(n4581) );
  INV_X1 U4776 ( .A(n3751), .ZN(n3753) );
  NAND2_X1 U4777 ( .A1(n4628), .A2(n6664), .ZN(n5203) );
  INV_X1 U4778 ( .A(n3754), .ZN(n3761) );
  AND3_X1 U4779 ( .A1(n3757), .A2(n3756), .A3(n3755), .ZN(n3758) );
  OR2_X1 U4780 ( .A1(n3759), .A2(n3758), .ZN(n3760) );
  NOR2_X1 U4781 ( .A1(n4517), .A2(READY_N), .ZN(n4578) );
  NAND3_X1 U4782 ( .A1(n5203), .A2(n4578), .A3(n3401), .ZN(n3762) );
  OAI211_X1 U4783 ( .C1(n4584), .C2(n3763), .A(n4581), .B(n3762), .ZN(n3765)
         );
  NAND2_X1 U4784 ( .A1(n3765), .A2(n6640), .ZN(n3769) );
  AOI21_X1 U4785 ( .B1(n4630), .B2(n6664), .A(READY_N), .ZN(n4576) );
  NAND2_X1 U4786 ( .A1(n4814), .A2(n3780), .ZN(n3766) );
  AOI21_X1 U4787 ( .B1(n4589), .B2(n4576), .A(n3766), .ZN(n3767) );
  NAND2_X1 U4788 ( .A1(n3771), .A2(n3147), .ZN(n3772) );
  INV_X1 U4789 ( .A(n3778), .ZN(n3774) );
  INV_X4 U4790 ( .A(n3787), .ZN(n4466) );
  AOI22_X1 U4791 ( .A1(n3774), .A2(n4724), .B1(n4589), .B2(n4466), .ZN(n3776)
         );
  NAND4_X1 U4792 ( .A1(n4803), .A2(n6617), .A3(n3776), .A4(n4785), .ZN(n3777)
         );
  NAND2_X1 U4793 ( .A1(n4589), .A2(n4469), .ZN(n6630) );
  OAI21_X1 U4794 ( .B1(n3778), .B2(n4724), .A(n6630), .ZN(n3779) );
  NAND2_X2 U4795 ( .A1(n5354), .A2(n4466), .ZN(n5217) );
  INV_X1 U4796 ( .A(n4728), .ZN(n3781) );
  NAND2_X1 U4797 ( .A1(n3781), .A2(n3780), .ZN(n3799) );
  INV_X1 U4798 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4799 ( .A1(n4466), .A2(n3782), .ZN(n3783) );
  OAI211_X1 U4800 ( .C1(n3804), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n3783), 
        .B(n3791), .ZN(n3784) );
  OAI21_X2 U4801 ( .B1(EBX_REG_1__SCAN_IN), .B2(n5217), .A(n3784), .ZN(n3788)
         );
  INV_X1 U4802 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U4803 ( .A1(n3791), .A2(n4612), .ZN(n3786) );
  NAND2_X1 U4804 ( .A1(n3799), .A2(EBX_REG_0__SCAN_IN), .ZN(n3785) );
  XNOR2_X1 U4805 ( .A(n3788), .B(n4608), .ZN(n4617) );
  OAI21_X1 U4806 ( .B1(n4617), .B2(n3787), .A(n3788), .ZN(n3789) );
  INV_X1 U4807 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4808 ( .A1(n3799), .A2(n3790), .ZN(n3792) );
  OAI211_X1 U4809 ( .C1(n3787), .C2(EBX_REG_2__SCAN_IN), .A(n3792), .B(n3791), 
        .ZN(n3793) );
  OAI21_X1 U4810 ( .B1(n5217), .B2(EBX_REG_2__SCAN_IN), .A(n3793), .ZN(n4682)
         );
  MUX2_X1 U4811 ( .A(n4389), .B(n3791), .S(EBX_REG_3__SCAN_IN), .Z(n3794) );
  NAND2_X1 U4812 ( .A1(n3278), .A2(n3794), .ZN(n4690) );
  NAND2_X1 U4813 ( .A1(n3799), .A2(n3795), .ZN(n3796) );
  OAI211_X1 U4814 ( .C1(n3787), .C2(EBX_REG_4__SCAN_IN), .A(n3796), .B(n3791), 
        .ZN(n3797) );
  OAI21_X1 U4815 ( .B1(n5217), .B2(EBX_REG_4__SCAN_IN), .A(n3797), .ZN(n4749)
         );
  MUX2_X1 U4816 ( .A(n4389), .B(n3791), .S(EBX_REG_5__SCAN_IN), .Z(n3798) );
  OAI21_X1 U4817 ( .B1(n5215), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n3798), 
        .ZN(n4934) );
  INV_X1 U4818 ( .A(n3799), .ZN(n3804) );
  MUX2_X1 U4819 ( .A(n5217), .B(n3846), .S(EBX_REG_6__SCAN_IN), .Z(n3802) );
  NAND2_X1 U4820 ( .A1(n3787), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3800)
         );
  OR2_X1 U4821 ( .A1(n4466), .A2(n3846), .ZN(n3815) );
  AND2_X1 U4822 ( .A1(n3800), .A2(n3815), .ZN(n3801) );
  NAND2_X1 U4823 ( .A1(n3802), .A2(n3801), .ZN(n4973) );
  MUX2_X1 U4824 ( .A(n4389), .B(n3791), .S(EBX_REG_7__SCAN_IN), .Z(n3803) );
  NAND2_X1 U4825 ( .A1(n3273), .A2(n3803), .ZN(n4931) );
  NAND2_X1 U4826 ( .A1(n3846), .A2(n3805), .ZN(n3806) );
  OAI211_X1 U4827 ( .C1(n5214), .C2(EBX_REG_8__SCAN_IN), .A(n3806), .B(n3791), 
        .ZN(n3807) );
  OAI21_X1 U4828 ( .B1(n5217), .B2(EBX_REG_8__SCAN_IN), .A(n3807), .ZN(n4967)
         );
  MUX2_X1 U4829 ( .A(n4389), .B(n3791), .S(EBX_REG_9__SCAN_IN), .Z(n3808) );
  OAI21_X1 U4830 ( .B1(n5215), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n3808), 
        .ZN(n5484) );
  MUX2_X1 U4831 ( .A(n5217), .B(n3846), .S(EBX_REG_10__SCAN_IN), .Z(n3811) );
  NAND2_X1 U4832 ( .A1(n3787), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3809) );
  AND2_X1 U4833 ( .A1(n3809), .A2(n3815), .ZN(n3810) );
  NAND2_X1 U4834 ( .A1(n3811), .A2(n3810), .ZN(n5616) );
  NAND2_X1 U4835 ( .A1(n5482), .A2(n5616), .ZN(n5615) );
  INV_X1 U4836 ( .A(EBX_REG_11__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4837 ( .A1(n4466), .A2(n3812), .ZN(n3813) );
  OAI211_X1 U4838 ( .C1(n5354), .C2(n6443), .A(n3813), .B(n3846), .ZN(n3814)
         );
  OAI21_X1 U4839 ( .B1(n4389), .B2(EBX_REG_11__SCAN_IN), .A(n3814), .ZN(n5470)
         );
  MUX2_X1 U4840 ( .A(n5217), .B(n3846), .S(EBX_REG_12__SCAN_IN), .Z(n3818) );
  NAND2_X1 U4841 ( .A1(n5214), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3816) );
  AND2_X1 U4842 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  NAND2_X1 U4843 ( .A1(n3818), .A2(n3817), .ZN(n5450) );
  INV_X1 U4844 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6979) );
  NAND2_X1 U4845 ( .A1(n4466), .A2(n6979), .ZN(n3819) );
  OAI211_X1 U4846 ( .C1(n5354), .C2(n6902), .A(n3819), .B(n3846), .ZN(n3820)
         );
  OAI21_X1 U4847 ( .B1(n4389), .B2(EBX_REG_13__SCAN_IN), .A(n3820), .ZN(n5439)
         );
  MUX2_X1 U4848 ( .A(n5217), .B(n3846), .S(EBX_REG_14__SCAN_IN), .Z(n3822) );
  NAND2_X1 U4849 ( .A1(n5214), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3821) );
  NAND2_X1 U4850 ( .A1(n3822), .A2(n3821), .ZN(n5426) );
  NAND2_X1 U4851 ( .A1(n3791), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3823) );
  OAI211_X1 U4852 ( .C1(n5214), .C2(EBX_REG_15__SCAN_IN), .A(n3846), .B(n3823), 
        .ZN(n3824) );
  OAI21_X1 U4853 ( .B1(n4389), .B2(EBX_REG_15__SCAN_IN), .A(n3824), .ZN(n5412)
         );
  MUX2_X1 U4854 ( .A(n5217), .B(n3799), .S(EBX_REG_16__SCAN_IN), .Z(n3826) );
  NAND2_X1 U4855 ( .A1(n5214), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4856 ( .A1(n3826), .A2(n3825), .ZN(n5397) );
  INV_X1 U4857 ( .A(n4389), .ZN(n3827) );
  INV_X1 U4858 ( .A(EBX_REG_17__SCAN_IN), .ZN(n7012) );
  NAND2_X1 U4859 ( .A1(n3827), .A2(n7012), .ZN(n3830) );
  NAND2_X1 U4860 ( .A1(n3791), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3828) );
  OAI211_X1 U4861 ( .C1(n5214), .C2(EBX_REG_17__SCAN_IN), .A(n3846), .B(n3828), 
        .ZN(n3829) );
  AND2_X1 U4862 ( .A1(n3830), .A2(n3829), .ZN(n5382) );
  AND2_X1 U4863 ( .A1(n5397), .A2(n5382), .ZN(n3831) );
  NAND2_X1 U4864 ( .A1(n5381), .A2(n3831), .ZN(n5353) );
  INV_X1 U4865 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4866 ( .A1(n4390), .A2(n3832), .ZN(n3835) );
  NAND2_X1 U4867 ( .A1(n3846), .A2(n6932), .ZN(n3833) );
  OAI211_X1 U4868 ( .C1(EBX_REG_19__SCAN_IN), .C2(n5214), .A(n3833), .B(n3791), 
        .ZN(n3834) );
  INV_X1 U4869 ( .A(n3836), .ZN(n5337) );
  OR2_X1 U4870 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3838)
         );
  INV_X1 U4871 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U4872 ( .A1(n4466), .A2(n7019), .ZN(n3837) );
  AND2_X1 U4873 ( .A1(n3838), .A2(n3837), .ZN(n5338) );
  OR2_X1 U4874 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3840)
         );
  INV_X1 U4875 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4876 ( .A1(n4466), .A2(n3839), .ZN(n5355) );
  NAND2_X1 U4877 ( .A1(n3840), .A2(n5355), .ZN(n5356) );
  NAND2_X1 U4878 ( .A1(n5354), .A2(EBX_REG_20__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4879 ( .A1(n5356), .A2(n3791), .ZN(n3841) );
  OAI211_X1 U4880 ( .C1(n5338), .C2(n5356), .A(n3842), .B(n3841), .ZN(n3843)
         );
  MUX2_X1 U4881 ( .A(n4389), .B(n3791), .S(EBX_REG_21__SCAN_IN), .Z(n3844) );
  OAI21_X1 U4882 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5215), .A(n3844), 
        .ZN(n3845) );
  INV_X1 U4883 ( .A(n3845), .ZN(n5327) );
  MUX2_X1 U4884 ( .A(n5217), .B(n3846), .S(EBX_REG_22__SCAN_IN), .Z(n3848) );
  NAND2_X1 U4885 ( .A1(n5214), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3847) );
  NAND2_X1 U4886 ( .A1(n3848), .A2(n3847), .ZN(n5317) );
  NAND2_X1 U4887 ( .A1(n3791), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3849) );
  OAI211_X1 U4888 ( .C1(n5214), .C2(EBX_REG_23__SCAN_IN), .A(n3846), .B(n3849), 
        .ZN(n3850) );
  OAI21_X1 U4889 ( .B1(n4389), .B2(EBX_REG_23__SCAN_IN), .A(n3850), .ZN(n5305)
         );
  MUX2_X1 U4890 ( .A(n5217), .B(n3799), .S(EBX_REG_24__SCAN_IN), .Z(n3852) );
  NAND2_X1 U4891 ( .A1(n5214), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3851) );
  NAND2_X1 U4892 ( .A1(n3852), .A2(n3851), .ZN(n3854) );
  NAND2_X1 U4893 ( .A1(n3853), .A2(n3854), .ZN(n5281) );
  OR2_X1 U4894 ( .A1(n3853), .A2(n3854), .ZN(n3855) );
  AND2_X1 U4895 ( .A1(n5281), .A2(n3855), .ZN(n5602) );
  AND2_X1 U4896 ( .A1(n5868), .A2(REIP_REG_24__SCAN_IN), .ZN(n5725) );
  INV_X1 U4897 ( .A(n3856), .ZN(n5973) );
  AND2_X1 U4898 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U4899 ( .A1(n5973), .A2(n5975), .ZN(n3884) );
  INV_X1 U4900 ( .A(n3884), .ZN(n3875) );
  NAND2_X1 U4901 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6041) );
  NOR2_X1 U4902 ( .A1(n6902), .A2(n6041), .ZN(n6020) );
  INV_X1 U4903 ( .A(n4814), .ZN(n4816) );
  NAND2_X1 U4904 ( .A1(n5215), .A2(n3857), .ZN(n3858) );
  NAND2_X1 U4905 ( .A1(n4526), .A2(n4736), .ZN(n5543) );
  OR2_X1 U4906 ( .A1(n5543), .A2(n3401), .ZN(n4580) );
  OAI211_X1 U4907 ( .C1(n3859), .C2(n4816), .A(n3858), .B(n4580), .ZN(n3860)
         );
  INV_X1 U4908 ( .A(n3860), .ZN(n3861) );
  OAI211_X1 U4909 ( .C1(n3106), .C2(n3791), .A(n3862), .B(n3861), .ZN(n3863)
         );
  INV_X1 U4910 ( .A(n3863), .ZN(n3864) );
  NAND2_X1 U4911 ( .A1(n3865), .A2(n3864), .ZN(n4588) );
  INV_X1 U4912 ( .A(n4770), .ZN(n3866) );
  NAND2_X1 U4913 ( .A1(n3869), .A2(n3867), .ZN(n4593) );
  INV_X1 U4914 ( .A(n4593), .ZN(n3868) );
  AOI21_X1 U4915 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4758) );
  NAND2_X1 U4916 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4864) );
  NOR2_X1 U4917 ( .A1(n4758), .A2(n4864), .ZN(n6077) );
  NOR2_X1 U4918 ( .A1(n3650), .A2(n3805), .ZN(n6089) );
  INV_X1 U4919 ( .A(n6089), .ZN(n6078) );
  NAND2_X1 U4920 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6079) );
  INV_X1 U4921 ( .A(n6043), .ZN(n3872) );
  INV_X1 U4922 ( .A(n3869), .ZN(n3870) );
  NAND2_X1 U4923 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4756) );
  NOR2_X1 U4924 ( .A1(n4864), .A2(n4756), .ZN(n4956) );
  NAND3_X1 U4925 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4956), .ZN(n6071) );
  NOR2_X1 U4926 ( .A1(n3871), .A2(n6071), .ZN(n3876) );
  NAND2_X1 U4927 ( .A1(n5983), .A2(n3876), .ZN(n6060) );
  NAND2_X1 U4928 ( .A1(n3872), .A2(n6060), .ZN(n6439) );
  NAND2_X1 U4929 ( .A1(n6020), .A2(n6439), .ZN(n6036) );
  INV_X1 U4930 ( .A(n6036), .ZN(n3873) );
  NAND2_X1 U4931 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n3873), .ZN(n3874) );
  NOR2_X2 U4932 ( .A1(n6014), .A2(n3874), .ZN(n6006) );
  AND2_X1 U4933 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U4934 ( .A1(n5965), .A2(n4411), .ZN(n5947) );
  NOR2_X1 U4935 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4414) );
  INV_X1 U4936 ( .A(n3876), .ZN(n3877) );
  NAND2_X1 U4937 ( .A1(n6070), .A2(n3877), .ZN(n6018) );
  NOR2_X1 U4938 ( .A1(n6014), .A2(n5787), .ZN(n3878) );
  AND2_X1 U4939 ( .A1(n6020), .A2(n3878), .ZN(n3881) );
  INV_X1 U4940 ( .A(n3881), .ZN(n3879) );
  NAND2_X1 U4941 ( .A1(n6070), .A2(n3879), .ZN(n3880) );
  NAND2_X1 U4942 ( .A1(n6018), .A2(n3880), .ZN(n5979) );
  NAND2_X1 U4943 ( .A1(n6043), .A2(n3881), .ZN(n5980) );
  OR2_X1 U4944 ( .A1(n3882), .A2(n5868), .ZN(n4620) );
  INV_X1 U4945 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6726) );
  INV_X1 U4946 ( .A(n6042), .ZN(n3883) );
  NAND2_X1 U4947 ( .A1(n3883), .A2(n6061), .ZN(n6037) );
  NAND2_X1 U4948 ( .A1(n6726), .A2(n6037), .ZN(n4619) );
  NAND2_X1 U4949 ( .A1(n4620), .A2(n4619), .ZN(n4755) );
  INV_X1 U4950 ( .A(n4755), .ZN(n4639) );
  NAND2_X1 U4951 ( .A1(n6061), .A2(n4639), .ZN(n6072) );
  INV_X1 U4952 ( .A(n4411), .ZN(n5957) );
  AND2_X1 U4953 ( .A1(n6021), .A2(n5957), .ZN(n3885) );
  NAND2_X1 U4954 ( .A1(n6469), .A2(n6061), .ZN(n3886) );
  NAND2_X1 U4955 ( .A1(n3886), .A2(n4450), .ZN(n3887) );
  NAND2_X1 U4956 ( .A1(n5949), .A2(n3887), .ZN(n5943) );
  INV_X1 U4957 ( .A(n5943), .ZN(n3888) );
  AOI211_X1 U4958 ( .C1(n3889), .C2(n5947), .A(n4414), .B(n3888), .ZN(n3890)
         );
  AOI211_X1 U4959 ( .C1(n6463), .C2(n5602), .A(n5725), .B(n3890), .ZN(n3891)
         );
  OAI21_X1 U4960 ( .B1(n5731), .B2(n6084), .A(n3891), .ZN(U2994) );
  NAND2_X1 U4962 ( .A1(n3895), .A2(n4073), .ZN(n3900) );
  AOI22_X1 U4963 ( .A1(n4408), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6326), .ZN(n3898) );
  NAND2_X1 U4964 ( .A1(n3908), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3897) );
  AND2_X1 U4965 ( .A1(n3898), .A2(n3897), .ZN(n3899) );
  NAND2_X1 U4966 ( .A1(n3900), .A2(n3899), .ZN(n4610) );
  NAND2_X1 U4967 ( .A1(n4611), .A2(n4610), .ZN(n4609) );
  INV_X1 U4968 ( .A(n4610), .ZN(n3901) );
  NAND2_X1 U4969 ( .A1(n3901), .A2(n4460), .ZN(n3902) );
  NAND2_X1 U4970 ( .A1(n4609), .A2(n3902), .ZN(n4616) );
  NAND2_X1 U4971 ( .A1(n4698), .A2(n4073), .ZN(n3906) );
  AOI22_X1 U4972 ( .A1(n4408), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6326), .ZN(n3904) );
  NAND2_X1 U4973 ( .A1(n3908), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3903) );
  AND2_X1 U4974 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  NAND2_X1 U4975 ( .A1(n6326), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4098) );
  AOI21_X1 U4976 ( .B1(n3907), .B2(n4073), .A(n4407), .ZN(n3911) );
  INV_X1 U4977 ( .A(n3908), .ZN(n3930) );
  INV_X2 U4978 ( .A(n3091), .ZN(n4460) );
  OAI21_X1 U4979 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3924), .ZN(n6435) );
  AOI22_X1 U4980 ( .A1(n4407), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4460), 
        .B2(n6435), .ZN(n3910) );
  NAND2_X1 U4981 ( .A1(n4097), .A2(EAX_REG_2__SCAN_IN), .ZN(n3909) );
  OAI211_X1 U4982 ( .C1(n3930), .C2(n3202), .A(n3910), .B(n3909), .ZN(n4681)
         );
  NAND2_X1 U4983 ( .A1(n4678), .A2(n4681), .ZN(n3915) );
  INV_X1 U4984 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U4985 ( .A1(n6326), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3917)
         );
  NAND2_X1 U4986 ( .A1(n4408), .A2(EAX_REG_4__SCAN_IN), .ZN(n3916) );
  OAI211_X1 U4987 ( .C1(n3930), .C2(n6991), .A(n3917), .B(n3916), .ZN(n3919)
         );
  INV_X1 U4988 ( .A(n3924), .ZN(n3918) );
  NAND2_X1 U4989 ( .A1(n3923), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3938)
         );
  OAI21_X1 U4990 ( .B1(n3923), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3938), 
        .ZN(n5537) );
  MUX2_X1 U4991 ( .A(n3919), .B(n5537), .S(n4460), .Z(n3920) );
  INV_X1 U4992 ( .A(n3920), .ZN(n3921) );
  NAND2_X1 U4993 ( .A1(n4798), .A2(n4073), .ZN(n3933) );
  INV_X1 U4994 ( .A(n3923), .ZN(n3927) );
  INV_X1 U4995 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3925) );
  NAND2_X1 U4996 ( .A1(n3925), .A2(n3924), .ZN(n3926) );
  NAND2_X1 U4997 ( .A1(n3927), .A2(n3926), .ZN(n5559) );
  AOI22_X1 U4998 ( .A1(n5559), .A2(n4460), .B1(n4407), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4999 ( .A1(n4097), .A2(EAX_REG_3__SCAN_IN), .ZN(n3928) );
  OAI211_X1 U5000 ( .C1(n3930), .C2(n4776), .A(n3929), .B(n3928), .ZN(n3931)
         );
  INV_X1 U5001 ( .A(n3931), .ZN(n3932) );
  AND2_X1 U5002 ( .A1(n4745), .A2(n4686), .ZN(n3947) );
  NOR2_X1 U5003 ( .A1(n3939), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3935)
         );
  AOI22_X1 U5004 ( .A1(n4408), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6326), .ZN(n3936) );
  MUX2_X1 U5005 ( .A(n3269), .B(n3936), .S(n3091), .Z(n3937) );
  AND2_X1 U5006 ( .A1(n3938), .A2(n3942), .ZN(n3940) );
  OR2_X1 U5007 ( .A1(n3940), .A2(n3939), .ZN(n5536) );
  NAND2_X1 U5008 ( .A1(n5536), .A2(n4460), .ZN(n3941) );
  OAI21_X1 U5009 ( .B1(n3942), .B2(n4098), .A(n3941), .ZN(n3943) );
  AOI21_X1 U5010 ( .B1(n4097), .B2(EAX_REG_5__SCAN_IN), .A(n3943), .ZN(n3944)
         );
  NAND2_X1 U5011 ( .A1(n3949), .A2(n4073), .ZN(n3955) );
  NAND2_X1 U5012 ( .A1(n4408), .A2(EAX_REG_7__SCAN_IN), .ZN(n3953) );
  NOR2_X1 U5013 ( .A1(n3950), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3951)
         );
  OR2_X1 U5014 ( .A1(n3982), .A2(n3951), .ZN(n5878) );
  AOI22_X1 U5015 ( .A1(n5878), .A2(n4460), .B1(n4407), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3952) );
  AND2_X1 U5016 ( .A1(n3953), .A2(n3952), .ZN(n3954) );
  NAND2_X1 U5017 ( .A1(n3955), .A2(n3954), .ZN(n4902) );
  AOI22_X1 U5018 ( .A1(n4322), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U5019 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4086), .B1(n4345), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U5020 ( .A1(n4354), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U5021 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3085), .B1(n4355), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U5022 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3965)
         );
  AOI22_X1 U5023 ( .A1(n3086), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U5024 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4344), .B1(n4306), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U5025 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4352), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U5026 ( .A1(n3557), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U5027 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  OAI21_X1 U5028 ( .B1(n3965), .B2(n3964), .A(n4073), .ZN(n3969) );
  XOR2_X1 U5029 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3982), .Z(n5873) );
  INV_X1 U5030 ( .A(n5873), .ZN(n3966) );
  AOI22_X1 U5031 ( .A1(n4407), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4460), 
        .B2(n3966), .ZN(n3968) );
  NAND2_X1 U5032 ( .A1(n4097), .A2(EAX_REG_8__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U5033 ( .A1(n4347), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U5034 ( .A1(n4352), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U5035 ( .A1(n4345), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5036 ( .A1(n3557), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U5037 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3981)
         );
  AOI22_X1 U5038 ( .A1(n3577), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U5039 ( .A1(n3085), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5040 ( .A1(n4086), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5041 ( .A1(n4322), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U5042 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  OAI21_X1 U5043 ( .B1(n3981), .B2(n3980), .A(n4073), .ZN(n3988) );
  INV_X1 U5044 ( .A(n3983), .ZN(n3985) );
  INV_X1 U5045 ( .A(n4012), .ZN(n3984) );
  OAI21_X1 U5046 ( .B1(PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n3985), .A(n3984), 
        .ZN(n5861) );
  AOI22_X1 U5047 ( .A1(n4460), .A2(n5861), .B1(n4407), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U5048 ( .A1(n4097), .A2(EAX_REG_9__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U5049 ( .A1(n4322), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U5050 ( .A1(n4344), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U5051 ( .A1(n4343), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U5052 ( .A1(n4345), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U5053 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3998)
         );
  AOI22_X1 U5054 ( .A1(n3086), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U5055 ( .A1(n4306), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5056 ( .A1(n3085), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U5057 ( .A1(n4086), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U5058 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3997)
         );
  OAI21_X1 U5059 ( .B1(n3998), .B2(n3997), .A(n4073), .ZN(n4001) );
  XOR2_X1 U5060 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4012), .Z(n6395) );
  INV_X1 U5061 ( .A(n6395), .ZN(n5856) );
  AOI22_X1 U5062 ( .A1(n4407), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n4460), 
        .B2(n5856), .ZN(n4000) );
  NAND2_X1 U5063 ( .A1(n4097), .A2(EAX_REG_10__SCAN_IN), .ZN(n3999) );
  INV_X1 U5064 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5671) );
  AOI22_X1 U5065 ( .A1(n3086), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U5066 ( .A1(n4347), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5067 ( .A1(n4344), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5068 ( .A1(n4355), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U5069 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4011)
         );
  AOI22_X1 U5070 ( .A1(n4322), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5071 ( .A1(n3085), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5072 ( .A1(n4345), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5073 ( .A1(n4086), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U5074 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  OAI21_X1 U5075 ( .B1(n4011), .B2(n4010), .A(n4073), .ZN(n4014) );
  XNOR2_X1 U5076 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4015), .ZN(n5845)
         );
  AOI22_X1 U5077 ( .A1(n4460), .A2(n5845), .B1(n4407), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4013) );
  OAI211_X1 U5078 ( .C1(n4367), .C2(n5671), .A(n4014), .B(n4013), .ZN(n5461)
         );
  AOI21_X1 U5079 ( .B1(n6878), .B2(n4016), .A(n4043), .ZN(n5836) );
  OR2_X1 U5080 ( .A1(n5836), .A2(n3091), .ZN(n4031) );
  AOI22_X1 U5081 ( .A1(n3086), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5082 ( .A1(n3085), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5083 ( .A1(n4322), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5084 ( .A1(n4352), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4017) );
  NAND4_X1 U5085 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4026)
         );
  AOI22_X1 U5086 ( .A1(n4347), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5087 ( .A1(n4345), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5088 ( .A1(n4343), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5089 ( .A1(n4086), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4021) );
  NAND4_X1 U5090 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4025)
         );
  OAI21_X1 U5091 ( .B1(n4026), .B2(n4025), .A(n4073), .ZN(n4029) );
  NAND2_X1 U5092 ( .A1(n4097), .A2(EAX_REG_12__SCAN_IN), .ZN(n4028) );
  NAND2_X1 U5093 ( .A1(n4407), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4027)
         );
  AOI22_X1 U5094 ( .A1(n4322), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5095 ( .A1(n3086), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5096 ( .A1(n4343), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5097 ( .A1(n4352), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U5098 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4041)
         );
  AOI22_X1 U5099 ( .A1(n3085), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5100 ( .A1(n4306), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5101 ( .A1(n4344), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5102 ( .A1(n4086), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U5103 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4040)
         );
  OR2_X1 U5104 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  AND2_X1 U5105 ( .A1(n4073), .A2(n4042), .ZN(n5435) );
  INV_X1 U5106 ( .A(n4047), .ZN(n4064) );
  OR2_X1 U5107 ( .A1(n4043), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4044)
         );
  NAND2_X1 U5108 ( .A1(n4064), .A2(n4044), .ZN(n5825) );
  NAND2_X1 U5109 ( .A1(n5825), .A2(n4460), .ZN(n4046) );
  AOI22_X1 U5110 ( .A1(n4408), .A2(EAX_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4407), .ZN(n4045) );
  NAND2_X1 U5111 ( .A1(n4046), .A2(n4045), .ZN(n5408) );
  INV_X1 U5112 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U5113 ( .A(n4084), .B(n5414), .ZN(n5809) );
  NAND2_X1 U5114 ( .A1(n5809), .A2(n4460), .ZN(n4062) );
  AOI22_X1 U5115 ( .A1(n4322), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5116 ( .A1(n4344), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5117 ( .A1(n4086), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5118 ( .A1(n4352), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U5119 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4057)
         );
  AOI22_X1 U5120 ( .A1(n3086), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5121 ( .A1(n4347), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5122 ( .A1(n3085), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5123 ( .A1(n4306), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U5124 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4056)
         );
  OAI21_X1 U5125 ( .B1(n4057), .B2(n4056), .A(n4073), .ZN(n4060) );
  NAND2_X1 U5126 ( .A1(n4097), .A2(EAX_REG_15__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U5127 ( .A1(n4407), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4058)
         );
  AND3_X1 U5128 ( .A1(n4060), .A2(n4059), .A3(n4058), .ZN(n4061) );
  NAND2_X1 U5129 ( .A1(n4062), .A2(n4061), .ZN(n5410) );
  INV_X1 U5130 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4063) );
  XNOR2_X1 U5131 ( .A(n4064), .B(n4063), .ZN(n5817) );
  NAND2_X1 U5132 ( .A1(n5817), .A2(n4460), .ZN(n4080) );
  AOI22_X1 U5133 ( .A1(n3085), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5134 ( .A1(n4345), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5135 ( .A1(n4086), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5136 ( .A1(n4354), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4065) );
  NAND4_X1 U5137 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4075)
         );
  AOI22_X1 U5138 ( .A1(n3086), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5139 ( .A1(n4322), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5140 ( .A1(n4347), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5141 ( .A1(n4355), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4069) );
  NAND4_X1 U5142 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4074)
         );
  OAI21_X1 U5143 ( .B1(n4075), .B2(n4074), .A(n4073), .ZN(n4078) );
  NAND2_X1 U5144 ( .A1(n4097), .A2(EAX_REG_14__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U5145 ( .A1(n4407), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4076)
         );
  AND3_X1 U5146 ( .A1(n4078), .A2(n4077), .A3(n4076), .ZN(n4079) );
  NAND2_X1 U5147 ( .A1(n4080), .A2(n4079), .ZN(n5409) );
  OAI211_X1 U5148 ( .C1(n5435), .C2(n5408), .A(n5410), .B(n5409), .ZN(n4081)
         );
  INV_X1 U5149 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6814) );
  OAI21_X1 U5150 ( .B1(n4084), .B2(n5414), .A(n6814), .ZN(n4085) );
  NAND2_X1 U5151 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4083) );
  NAND2_X1 U5152 ( .A1(n4085), .A2(n4104), .ZN(n5800) );
  NAND2_X1 U5153 ( .A1(n5800), .A2(n4460), .ZN(n4103) );
  AOI22_X1 U5154 ( .A1(n4322), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5155 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3085), .B1(n4345), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5156 ( .A1(n4086), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5157 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4352), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U5158 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4096)
         );
  AOI22_X1 U5159 ( .A1(n3086), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5160 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4347), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5161 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n4344), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5162 ( .A1(n4306), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4091) );
  NAND4_X1 U5163 ( .A1(n4094), .A2(n4093), .A3(n4092), .A4(n4091), .ZN(n4095)
         );
  OR2_X1 U5164 ( .A1(n4096), .A2(n4095), .ZN(n4101) );
  INV_X1 U5165 ( .A(n4097), .ZN(n4367) );
  INV_X1 U5166 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4099) );
  OAI22_X1 U5167 ( .A1(n4367), .A2(n4099), .B1(n6814), .B2(n4098), .ZN(n4100)
         );
  AOI21_X1 U5168 ( .B1(n4369), .B2(n4101), .A(n4100), .ZN(n4102) );
  NAND2_X1 U5169 ( .A1(n4103), .A2(n4102), .ZN(n5393) );
  INV_X1 U5170 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U5171 ( .A1(n4104), .A2(n6837), .ZN(n4105) );
  NAND2_X1 U5172 ( .A1(n4136), .A2(n4105), .ZN(n5790) );
  OR2_X1 U5173 ( .A1(n5790), .A2(n3091), .ZN(n4120) );
  AOI22_X1 U5174 ( .A1(n4322), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5175 ( .A1(n3085), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5176 ( .A1(n4086), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5177 ( .A1(n4344), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5178 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4115)
         );
  AOI22_X1 U5179 ( .A1(n3086), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5180 ( .A1(n4347), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5181 ( .A1(n4352), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5182 ( .A1(n4306), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4110) );
  NAND4_X1 U5183 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4114)
         );
  NOR2_X1 U5184 ( .A1(n4115), .A2(n4114), .ZN(n4118) );
  OAI21_X1 U5185 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6643), .A(n6326), 
        .ZN(n4117) );
  NAND2_X1 U5186 ( .A1(n4408), .A2(EAX_REG_17__SCAN_IN), .ZN(n4116) );
  OAI211_X1 U5187 ( .C1(n4332), .C2(n4118), .A(n4117), .B(n4116), .ZN(n4119)
         );
  AOI22_X1 U5188 ( .A1(n4343), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5189 ( .A1(n3085), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5190 ( .A1(n4306), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5191 ( .A1(n4322), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5192 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4130)
         );
  AOI22_X1 U5193 ( .A1(n4347), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5194 ( .A1(n3086), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5195 ( .A1(n4345), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5196 ( .A1(n4086), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4125) );
  NAND4_X1 U5197 ( .A1(n4128), .A2(n4127), .A3(n4126), .A4(n4125), .ZN(n4129)
         );
  OR2_X1 U5198 ( .A1(n4130), .A2(n4129), .ZN(n4133) );
  INV_X1 U5199 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4131) );
  INV_X1 U5200 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5781) );
  OAI22_X1 U5201 ( .A1(n4367), .A2(n4131), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5781), .ZN(n4132) );
  AOI21_X1 U5202 ( .B1(n4369), .B2(n4133), .A(n4132), .ZN(n4134) );
  XNOR2_X1 U5203 ( .A(n4136), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5783)
         );
  MUX2_X1 U5204 ( .A(n4134), .B(n5783), .S(n4460), .Z(n5367) );
  OR2_X2 U5205 ( .A1(n4138), .A2(n5769), .ZN(n4169) );
  NAND2_X1 U5206 ( .A1(n4138), .A2(n5769), .ZN(n4139) );
  NAND2_X1 U5207 ( .A1(n4169), .A2(n4139), .ZN(n5363) );
  AOI22_X1 U5208 ( .A1(n4343), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5209 ( .A1(n3085), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5210 ( .A1(n4344), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5211 ( .A1(n4086), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4140) );
  NAND4_X1 U5212 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4149)
         );
  AOI22_X1 U5213 ( .A1(n4322), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5214 ( .A1(n4345), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5215 ( .A1(n3086), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5216 ( .A1(n4352), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4144) );
  NAND4_X1 U5217 ( .A1(n4147), .A2(n4146), .A3(n4145), .A4(n4144), .ZN(n4148)
         );
  NOR2_X1 U5218 ( .A1(n4149), .A2(n4148), .ZN(n4152) );
  OAI21_X1 U5219 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6643), .A(n6326), 
        .ZN(n4151) );
  NAND2_X1 U5220 ( .A1(n4097), .A2(EAX_REG_19__SCAN_IN), .ZN(n4150) );
  OAI211_X1 U5221 ( .C1(n4332), .C2(n4152), .A(n4151), .B(n4150), .ZN(n4153)
         );
  OAI21_X1 U5222 ( .B1(n5363), .B2(n3091), .A(n4153), .ZN(n5346) );
  XNOR2_X1 U5223 ( .A(n4169), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5761)
         );
  AOI22_X1 U5224 ( .A1(n4322), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5225 ( .A1(n3086), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5226 ( .A1(n4343), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5227 ( .A1(n4352), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4154) );
  NAND4_X1 U5228 ( .A1(n4157), .A2(n4156), .A3(n4155), .A4(n4154), .ZN(n4163)
         );
  AOI22_X1 U5229 ( .A1(n3085), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5230 ( .A1(n4306), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5231 ( .A1(n4344), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5232 ( .A1(n4086), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U5233 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4162)
         );
  OR2_X1 U5234 ( .A1(n4163), .A2(n4162), .ZN(n4167) );
  INV_X1 U5235 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4165) );
  OAI21_X1 U5236 ( .B1(n6643), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n6326), 
        .ZN(n4164) );
  OAI21_X1 U5237 ( .B1(n4367), .B2(n4165), .A(n4164), .ZN(n4166) );
  AOI21_X1 U5238 ( .B1(n4369), .B2(n4167), .A(n4166), .ZN(n4168) );
  AOI21_X1 U5239 ( .B1(n5761), .B2(n4460), .A(n4168), .ZN(n5335) );
  NAND2_X1 U5240 ( .A1(n4171), .A2(n4170), .ZN(n4172) );
  NAND2_X1 U5241 ( .A1(n4199), .A2(n4172), .ZN(n5756) );
  AOI22_X1 U5242 ( .A1(n3086), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5243 ( .A1(n4347), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5244 ( .A1(n3085), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5245 ( .A1(n4345), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4173) );
  NAND4_X1 U5246 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4182)
         );
  AOI22_X1 U5247 ( .A1(n4354), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5248 ( .A1(n4322), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5249 ( .A1(n4306), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5250 ( .A1(n4086), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4177) );
  NAND4_X1 U5251 ( .A1(n4180), .A2(n4179), .A3(n4178), .A4(n4177), .ZN(n4181)
         );
  NOR2_X1 U5252 ( .A1(n4182), .A2(n4181), .ZN(n4184) );
  AOI22_X1 U5253 ( .A1(n4408), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6326), .ZN(n4183) );
  OAI21_X1 U5254 ( .B1(n4332), .B2(n4184), .A(n4183), .ZN(n4185) );
  MUX2_X1 U5255 ( .A(n5756), .B(n4185), .S(n3091), .Z(n5326) );
  AOI22_X1 U5256 ( .A1(n4322), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5257 ( .A1(n3085), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5258 ( .A1(n4343), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5259 ( .A1(n4352), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U5260 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4195)
         );
  AOI22_X1 U5261 ( .A1(n4345), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5262 ( .A1(n3086), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5263 ( .A1(n4344), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5264 ( .A1(n3557), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4190) );
  NAND4_X1 U5265 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4194)
         );
  OR2_X1 U5266 ( .A1(n4195), .A2(n4194), .ZN(n4197) );
  INV_X1 U5267 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4571) );
  INV_X1 U5268 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5748) );
  OAI22_X1 U5269 ( .A1(n4367), .A2(n4571), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5748), .ZN(n4196) );
  AOI21_X1 U5270 ( .B1(n4369), .B2(n4197), .A(n4196), .ZN(n4198) );
  XNOR2_X1 U5271 ( .A(n4199), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5746)
         );
  MUX2_X1 U5272 ( .A(n4198), .B(n5746), .S(n4460), .Z(n5315) );
  OR2_X2 U5273 ( .A1(n4202), .A2(n4201), .ZN(n4258) );
  NAND2_X1 U5274 ( .A1(n4202), .A2(n4201), .ZN(n4203) );
  NAND2_X1 U5275 ( .A1(n4258), .A2(n4203), .ZN(n5737) );
  AOI22_X1 U5276 ( .A1(n4343), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5277 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4344), .B1(n4345), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5278 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4347), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5279 ( .A1(n3557), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4204) );
  NAND4_X1 U5280 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4213)
         );
  AOI22_X1 U5281 ( .A1(n4322), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3086), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5282 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4086), .B1(n4306), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5283 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n4352), .B1(n4279), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5284 ( .A1(n3085), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4208) );
  NAND4_X1 U5285 ( .A1(n4211), .A2(n4210), .A3(n4209), .A4(n4208), .ZN(n4212)
         );
  NOR2_X1 U5286 ( .A1(n4213), .A2(n4212), .ZN(n4229) );
  AOI22_X1 U5287 ( .A1(n4345), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5288 ( .A1(n4347), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5289 ( .A1(n4352), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5290 ( .A1(n4086), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4214) );
  NAND4_X1 U5291 ( .A1(n4217), .A2(n4216), .A3(n4215), .A4(n4214), .ZN(n4223)
         );
  AOI22_X1 U5292 ( .A1(n3086), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5293 ( .A1(n4322), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5294 ( .A1(n3085), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5295 ( .A1(n4344), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4218) );
  NAND4_X1 U5296 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(n4222)
         );
  NOR2_X1 U5297 ( .A1(n4223), .A2(n4222), .ZN(n4230) );
  XNOR2_X1 U5298 ( .A(n4229), .B(n4230), .ZN(n4225) );
  AOI22_X1 U5299 ( .A1(n4408), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6326), .ZN(n4224) );
  OAI21_X1 U5300 ( .B1(n4332), .B2(n4225), .A(n4224), .ZN(n4226) );
  MUX2_X1 U5301 ( .A(n5737), .B(n4226), .S(n3091), .Z(n4227) );
  INV_X1 U5302 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4228) );
  XNOR2_X1 U5303 ( .A(n4258), .B(n4228), .ZN(n5727) );
  NOR2_X1 U5304 ( .A1(n4230), .A2(n4229), .ZN(n4255) );
  AOI22_X1 U5305 ( .A1(n4322), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U5306 ( .A1(n3086), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5307 ( .A1(n4343), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U5308 ( .A1(n4352), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4231) );
  NAND4_X1 U5309 ( .A1(n4234), .A2(n4233), .A3(n4232), .A4(n4231), .ZN(n4240)
         );
  AOI22_X1 U5310 ( .A1(n3085), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U5311 ( .A1(n4306), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5312 ( .A1(n4344), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5313 ( .A1(n4086), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4235) );
  NAND4_X1 U5314 ( .A1(n4238), .A2(n4237), .A3(n4236), .A4(n4235), .ZN(n4239)
         );
  XNOR2_X1 U5315 ( .A(n4255), .B(n4254), .ZN(n4242) );
  AOI22_X1 U5316 ( .A1(n4408), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4407), .ZN(n4241) );
  OAI21_X1 U5317 ( .B1(n4242), .B2(n4332), .A(n4241), .ZN(n4243) );
  AOI21_X1 U5318 ( .B1(n5727), .B2(n4460), .A(n4243), .ZN(n5292) );
  AOI22_X1 U5319 ( .A1(n4322), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U5320 ( .A1(n3086), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U5321 ( .A1(n4343), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4245) );
  AOI22_X1 U5322 ( .A1(n4352), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4244) );
  NAND4_X1 U5323 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(n4253)
         );
  AOI22_X1 U5324 ( .A1(n3085), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U5325 ( .A1(n4306), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U5326 ( .A1(n4344), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U5327 ( .A1(n4086), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4248) );
  NAND4_X1 U5328 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4252)
         );
  NOR2_X1 U5329 ( .A1(n4253), .A2(n4252), .ZN(n4264) );
  NAND2_X1 U5330 ( .A1(n4255), .A2(n4254), .ZN(n4263) );
  XNOR2_X1 U5331 ( .A(n4264), .B(n4263), .ZN(n4257) );
  AOI22_X1 U5332 ( .A1(n4408), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6326), .ZN(n4256) );
  OAI21_X1 U5333 ( .B1(n4257), .B2(n4332), .A(n4256), .ZN(n4262) );
  INV_X1 U5334 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U5335 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  NAND2_X1 U5336 ( .A1(n4294), .A2(n4261), .ZN(n5721) );
  MUX2_X1 U5337 ( .A(n4262), .B(n5721), .S(n4460), .Z(n5277) );
  NAND2_X1 U5338 ( .A1(n5276), .A2(n5277), .ZN(n5262) );
  NOR2_X1 U5339 ( .A1(n4264), .A2(n4263), .ZN(n4291) );
  AOI22_X1 U5340 ( .A1(n4322), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5341 ( .A1(n3086), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U5342 ( .A1(n4343), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U5343 ( .A1(n3379), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4265) );
  NAND4_X1 U5344 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(n4274)
         );
  AOI22_X1 U5345 ( .A1(n3085), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5346 ( .A1(n4306), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U5347 ( .A1(n4344), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U5348 ( .A1(n4086), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4269) );
  NAND4_X1 U5349 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), .ZN(n4273)
         );
  XOR2_X1 U5350 ( .A(n4291), .B(n4290), .Z(n4277) );
  INV_X1 U5351 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4275) );
  INV_X1 U5352 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5713) );
  OAI22_X1 U5353 ( .A1(n4367), .A2(n4275), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5713), .ZN(n4276) );
  AOI21_X1 U5354 ( .B1(n4277), .B2(n4369), .A(n4276), .ZN(n4278) );
  XNOR2_X1 U5355 ( .A(n4294), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5711)
         );
  MUX2_X1 U5356 ( .A(n4278), .B(n5711), .S(n4460), .Z(n5264) );
  AOI22_X1 U5357 ( .A1(n4345), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4283) );
  AOI22_X1 U5358 ( .A1(n4347), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U5359 ( .A1(n4322), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U5360 ( .A1(n4344), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4280) );
  NAND4_X1 U5361 ( .A1(n4283), .A2(n4282), .A3(n4281), .A4(n4280), .ZN(n4289)
         );
  AOI22_X1 U5362 ( .A1(n3086), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4287) );
  AOI22_X1 U5363 ( .A1(n4343), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U5364 ( .A1(n3085), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U5365 ( .A1(n4086), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4284) );
  NAND4_X1 U5366 ( .A1(n4287), .A2(n4286), .A3(n4285), .A4(n4284), .ZN(n4288)
         );
  NOR2_X1 U5367 ( .A1(n4289), .A2(n4288), .ZN(n4301) );
  NAND2_X1 U5368 ( .A1(n4291), .A2(n4290), .ZN(n4300) );
  XNOR2_X1 U5369 ( .A(n4301), .B(n4300), .ZN(n4293) );
  AOI22_X1 U5370 ( .A1(n4408), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6326), .ZN(n4292) );
  OAI21_X1 U5371 ( .B1(n4293), .B2(n4332), .A(n4292), .ZN(n4299) );
  INV_X1 U5372 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U5373 ( .A1(n4297), .A2(n4296), .ZN(n4298) );
  NAND2_X1 U5374 ( .A1(n3105), .A2(n4298), .ZN(n5704) );
  MUX2_X1 U5375 ( .A(n4299), .B(n5704), .S(n4460), .Z(n5248) );
  NOR2_X1 U5376 ( .A1(n4301), .A2(n4300), .ZN(n4330) );
  AOI22_X1 U5377 ( .A1(n4322), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U5378 ( .A1(n3086), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U5379 ( .A1(n4343), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U5380 ( .A1(n3379), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4302) );
  NAND4_X1 U5381 ( .A1(n4305), .A2(n4304), .A3(n4303), .A4(n4302), .ZN(n4312)
         );
  AOI22_X1 U5382 ( .A1(n3085), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3464), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U5383 ( .A1(n4306), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U5384 ( .A1(n4344), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U5385 ( .A1(n4086), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4307) );
  NAND4_X1 U5386 ( .A1(n4310), .A2(n4309), .A3(n4308), .A4(n4307), .ZN(n4311)
         );
  XNOR2_X1 U5387 ( .A(n4330), .B(n4329), .ZN(n4314) );
  AOI22_X1 U5388 ( .A1(n4408), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6326), .ZN(n4313) );
  OAI21_X1 U5389 ( .B1(n4314), .B2(n4332), .A(n4313), .ZN(n4316) );
  INV_X1 U5390 ( .A(n3105), .ZN(n4315) );
  XNOR2_X1 U5391 ( .A(n4315), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5240)
         );
  AOI22_X1 U5392 ( .A1(n3085), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U5393 ( .A1(n3086), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U5394 ( .A1(n4355), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U5395 ( .A1(n4086), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4318) );
  NAND4_X1 U5396 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(n4328)
         );
  AOI22_X1 U5397 ( .A1(n4343), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U5398 ( .A1(n4322), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4347), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5399 ( .A1(n4344), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5400 ( .A1(n4345), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U5401 ( .A1(n4326), .A2(n4325), .A3(n4324), .A4(n4323), .ZN(n4327)
         );
  NOR2_X1 U5402 ( .A1(n4328), .A2(n4327), .ZN(n4342) );
  NAND2_X1 U5403 ( .A1(n4330), .A2(n4329), .ZN(n4341) );
  XNOR2_X1 U5404 ( .A(n4342), .B(n4341), .ZN(n4333) );
  AOI22_X1 U5405 ( .A1(n4408), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6326), .ZN(n4331) );
  OAI21_X1 U5406 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(n4339) );
  INV_X1 U5407 ( .A(n4335), .ZN(n4337) );
  INV_X1 U5408 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4336) );
  NAND2_X1 U5409 ( .A1(n4337), .A2(n4336), .ZN(n4338) );
  NAND2_X1 U5410 ( .A1(n4425), .A2(n4338), .ZN(n5695) );
  MUX2_X1 U5411 ( .A(n4339), .B(n5695), .S(n4460), .Z(n4340) );
  XNOR2_X1 U5412 ( .A(n4425), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5685)
         );
  NOR2_X1 U5413 ( .A1(n4342), .A2(n4341), .ZN(n4364) );
  AOI22_X1 U5414 ( .A1(n3086), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4351) );
  AOI22_X1 U5415 ( .A1(n3085), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4344), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U5416 ( .A1(n4086), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U5417 ( .A1(n4347), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4348) );
  NAND4_X1 U5418 ( .A1(n4351), .A2(n4350), .A3(n4349), .A4(n4348), .ZN(n4362)
         );
  AOI22_X1 U5419 ( .A1(n4322), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U5420 ( .A1(n4354), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U5421 ( .A1(n4306), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U5422 ( .A1(n3557), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4356), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4357) );
  NAND4_X1 U5423 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), .ZN(n4361)
         );
  NOR2_X1 U5424 ( .A1(n4362), .A2(n4361), .ZN(n4363) );
  XNOR2_X1 U5425 ( .A(n4364), .B(n4363), .ZN(n4370) );
  INV_X1 U5426 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4366) );
  OAI21_X1 U5427 ( .B1(n6643), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6326), 
        .ZN(n4365) );
  OAI21_X1 U5428 ( .B1(n4367), .B2(n4366), .A(n4365), .ZN(n4368) );
  AOI21_X1 U5429 ( .B1(n4370), .B2(n4369), .A(n4368), .ZN(n4371) );
  INV_X1 U5430 ( .A(n4372), .ZN(n4374) );
  NOR2_X1 U5431 ( .A1(n3422), .A2(n4373), .ZN(n4805) );
  NAND3_X1 U5432 ( .A1(n4374), .A2(n4466), .A3(n4805), .ZN(n4377) );
  NAND2_X1 U5433 ( .A1(n3149), .A2(n4375), .ZN(n4376) );
  INV_X1 U5434 ( .A(n5623), .ZN(n4380) );
  NAND2_X1 U5435 ( .A1(n3791), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4381) );
  OAI211_X1 U5436 ( .C1(n5214), .C2(EBX_REG_25__SCAN_IN), .A(n3846), .B(n4381), 
        .ZN(n4382) );
  OAI21_X1 U5437 ( .B1(n4389), .B2(EBX_REG_25__SCAN_IN), .A(n4382), .ZN(n5280)
         );
  INV_X1 U5438 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U5439 ( .A1(n4390), .A2(n6892), .ZN(n4385) );
  INV_X1 U5440 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5441 ( .A1(n3846), .A2(n5708), .ZN(n4383) );
  OAI211_X1 U5442 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5214), .A(n4383), .B(n3791), 
        .ZN(n4384) );
  INV_X1 U5443 ( .A(n5266), .ZN(n4386) );
  NAND2_X1 U5444 ( .A1(n5265), .A2(n4386), .ZN(n5252) );
  NAND2_X1 U5445 ( .A1(n3791), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4387) );
  OAI211_X1 U5446 ( .C1(n5214), .C2(EBX_REG_27__SCAN_IN), .A(n3846), .B(n4387), 
        .ZN(n4388) );
  OAI21_X1 U5447 ( .B1(n4389), .B2(EBX_REG_27__SCAN_IN), .A(n4388), .ZN(n5253)
         );
  INV_X1 U5448 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U5449 ( .A1(n4390), .A2(n5601), .ZN(n4393) );
  INV_X1 U5450 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U5451 ( .A1(n3846), .A2(n4442), .ZN(n4391) );
  OAI211_X1 U5452 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5214), .A(n4391), .B(n3791), 
        .ZN(n4392) );
  INV_X1 U5453 ( .A(n5215), .ZN(n4397) );
  INV_X1 U5454 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U5455 ( .A1(n5214), .A2(EBX_REG_29__SCAN_IN), .ZN(n4396) );
  AOI21_X1 U5456 ( .B1(n4397), .B2(n5915), .A(n4396), .ZN(n5216) );
  AOI21_X1 U5457 ( .B1(n5354), .B2(n4395), .A(n5221), .ZN(n4399) );
  AND2_X1 U5458 ( .A1(n5214), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4398)
         );
  AOI21_X1 U5459 ( .B1(n5215), .B2(EBX_REG_30__SCAN_IN), .A(n4398), .ZN(n5219)
         );
  INV_X1 U5460 ( .A(n5904), .ZN(n4403) );
  INV_X1 U5461 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5462 ( .A1(n4405), .A2(n4404), .ZN(U2829) );
  AOI22_X1 U5463 ( .A1(n4408), .A2(EAX_REG_31__SCAN_IN), .B1(n4407), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U5464 ( .A1(n4461), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6651) );
  NAND2_X1 U5465 ( .A1(n5213), .A2(n6431), .ZN(n4436) );
  NAND2_X1 U5466 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4423) );
  AND2_X1 U5467 ( .A1(n4411), .A2(n5975), .ZN(n5734) );
  NAND2_X1 U5468 ( .A1(n5734), .A2(n4412), .ZN(n4413) );
  AND2_X1 U5469 ( .A1(n5777), .A2(n4413), .ZN(n4416) );
  NOR2_X1 U5470 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5955) );
  NOR2_X1 U5471 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5974) );
  AND3_X1 U5472 ( .A1(n5955), .A2(n4414), .A3(n5974), .ZN(n4415) );
  NAND2_X1 U5473 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U5474 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5910) );
  NOR2_X1 U5475 ( .A1(n5931), .A2(n5910), .ZN(n4417) );
  AND2_X1 U5476 ( .A1(n5777), .A2(n4417), .ZN(n4418) );
  NAND2_X1 U5477 ( .A1(n4419), .A2(n4418), .ZN(n5691) );
  INV_X1 U5478 ( .A(n4419), .ZN(n4421) );
  XOR2_X1 U5479 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n5777), .Z(n5718) );
  INV_X1 U5480 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U5481 ( .A1(n5920), .A2(n4442), .ZN(n4452) );
  NOR3_X1 U5482 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n4452), 
        .ZN(n5681) );
  INV_X1 U5483 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5900) );
  AND2_X1 U5484 ( .A1(n5900), .A2(n5915), .ZN(n4422) );
  INV_X1 U5485 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U5486 ( .A1(n5207), .A2(n6284), .ZN(n4428) );
  NAND2_X1 U5487 ( .A1(n4428), .A2(n6642), .ZN(n4429) );
  NAND2_X1 U5488 ( .A1(n6642), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5489 ( .A1(n6643), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4430) );
  AND2_X1 U5490 ( .A1(n4431), .A2(n4430), .ZN(n4672) );
  INV_X2 U5491 ( .A(n6075), .ZN(n5868) );
  NAND2_X1 U5492 ( .A1(n5868), .A2(REIP_REG_31__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U5493 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4432)
         );
  OAI211_X1 U5494 ( .C1(n4492), .C2(n6436), .A(n5896), .B(n4432), .ZN(n4433)
         );
  NAND3_X1 U5495 ( .A1(n4436), .A2(n4435), .A3(n4434), .ZN(U2955) );
  NOR2_X1 U5496 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5929) );
  NAND3_X1 U5497 ( .A1(n4421), .A2(n5832), .A3(n5929), .ZN(n5699) );
  XNOR2_X1 U5498 ( .A(n4443), .B(n4442), .ZN(n4498) );
  NAND2_X1 U5499 ( .A1(n4498), .A2(n4444), .ZN(n4457) );
  AND2_X1 U5500 ( .A1(n6021), .A2(n5931), .ZN(n4445) );
  AND2_X1 U5501 ( .A1(n5255), .A2(n4447), .ZN(n4449) );
  INV_X1 U5502 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U5503 ( .A1(n6075), .A2(n6707), .ZN(n4502) );
  INV_X1 U5504 ( .A(n4502), .ZN(n4454) );
  NOR2_X1 U5505 ( .A1(n5947), .A2(n4450), .ZN(n5939) );
  INV_X1 U5506 ( .A(n5931), .ZN(n4451) );
  NAND2_X1 U5507 ( .A1(n5939), .A2(n4451), .ZN(n5911) );
  INV_X1 U5508 ( .A(n5911), .ZN(n5921) );
  NAND3_X1 U5509 ( .A1(n5921), .A2(n4452), .A3(n5910), .ZN(n4453) );
  OAI211_X1 U5510 ( .C1(n5600), .C2(n6088), .A(n4454), .B(n4453), .ZN(n4455)
         );
  AOI21_X1 U5511 ( .B1(n5926), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n4455), 
        .ZN(n4456) );
  NAND2_X1 U5512 ( .A1(n4457), .A2(n4456), .ZN(U2990) );
  NOR2_X1 U5513 ( .A1(n4459), .A2(n4517), .ZN(n4509) );
  NAND2_X1 U5514 ( .A1(n4509), .A2(n6640), .ZN(n4507) );
  AND2_X1 U5515 ( .A1(n4461), .A2(n4460), .ZN(n4463) );
  NAND2_X1 U5516 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .ZN(n4462) );
  NOR2_X1 U5517 ( .A1(n6650), .A2(n4462), .ZN(n6633) );
  OR3_X4 U5518 ( .A1(n5210), .A2(n5868), .A3(n4464), .ZN(n5577) );
  OR2_X4 U5519 ( .A1(n4492), .A2(n4491), .ZN(n5522) );
  AND2_X2 U5520 ( .A1(n5577), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5545) );
  INV_X1 U5521 ( .A(n5545), .ZN(n4468) );
  INV_X1 U5522 ( .A(READY_N), .ZN(n4465) );
  NAND2_X1 U5523 ( .A1(n4465), .A2(n6643), .ZN(n4473) );
  NAND3_X1 U5524 ( .A1(n4466), .A2(EBX_REG_31__SCAN_IN), .A3(n4473), .ZN(n4467) );
  OR2_X1 U5525 ( .A1(n6664), .A2(n4473), .ZN(n6629) );
  AND2_X1 U5526 ( .A1(n4469), .A2(n6629), .ZN(n5226) );
  INV_X1 U5527 ( .A(n5226), .ZN(n4471) );
  INV_X1 U5528 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5597) );
  NAND3_X1 U5529 ( .A1(n3780), .A2(n5597), .A3(n4473), .ZN(n4470) );
  NAND2_X1 U5530 ( .A1(n4471), .A2(n4470), .ZN(n4472) );
  AND2_X2 U5531 ( .A1(n5545), .A2(n4472), .ZN(n6394) );
  AOI22_X1 U5532 ( .A1(n6394), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6390), .ZN(n4483) );
  INV_X1 U5533 ( .A(n6664), .ZN(n5202) );
  NAND2_X1 U5534 ( .A1(n3780), .A2(n5202), .ZN(n4474) );
  AOI21_X1 U5535 ( .B1(n5214), .B2(n4474), .A(n4473), .ZN(n4475) );
  AND2_X2 U5536 ( .A1(n5545), .A2(n4475), .ZN(n5565) );
  INV_X1 U5537 ( .A(n5565), .ZN(n5223) );
  NAND2_X1 U5538 ( .A1(n5223), .A2(n5577), .ZN(n5501) );
  AND2_X1 U5539 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4486) );
  INV_X1 U5540 ( .A(n4486), .ZN(n5395) );
  INV_X1 U5541 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6688) );
  INV_X1 U5542 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U5543 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5464) );
  NAND3_X1 U5544 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U5545 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .ZN(
        n4476) );
  NOR2_X1 U5546 ( .A1(n5539), .A2(n4476), .ZN(n5499) );
  AND3_X1 U5547 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n4484) );
  AND2_X1 U5548 ( .A1(n5499), .A2(n4484), .ZN(n4477) );
  NAND2_X1 U5549 ( .A1(REIP_REG_17__SCAN_IN), .A2(n3104), .ZN(n4478) );
  NOR2_X1 U5550 ( .A1(n5395), .A2(n4478), .ZN(n5349) );
  AND3_X1 U5551 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_20__SCAN_IN), .ZN(n4488) );
  AND2_X1 U5552 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5303) );
  NAND2_X1 U5553 ( .A1(n5303), .A2(REIP_REG_23__SCAN_IN), .ZN(n4489) );
  INV_X1 U5554 ( .A(n4489), .ZN(n5278) );
  AND2_X1 U5555 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5270) );
  NAND2_X1 U5556 ( .A1(n5270), .A2(REIP_REG_26__SCAN_IN), .ZN(n4490) );
  INV_X1 U5557 ( .A(n4490), .ZN(n4479) );
  INV_X1 U5558 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6708) );
  OR2_X1 U5559 ( .A1(n6707), .A2(n6708), .ZN(n4480) );
  NAND2_X1 U5560 ( .A1(n5565), .A2(n4480), .ZN(n4481) );
  OAI21_X1 U5561 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5223), .A(n5244), .ZN(n5225) );
  NAND2_X1 U5562 ( .A1(n5225), .A2(REIP_REG_30__SCAN_IN), .ZN(n4482) );
  OAI211_X1 U5563 ( .C1(n5904), .C2(n5517), .A(n4483), .B(n4482), .ZN(n4496)
         );
  AND2_X2 U5564 ( .A1(n5565), .A2(n5499), .ZN(n5513) );
  NAND2_X1 U5565 ( .A1(n3145), .A2(REIP_REG_11__SCAN_IN), .ZN(n4485) );
  NOR2_X2 U5566 ( .A1(n6387), .A2(n4485), .ZN(n5453) );
  NAND2_X1 U5567 ( .A1(n5453), .A2(REIP_REG_12__SCAN_IN), .ZN(n5436) );
  OR3_X2 U5568 ( .A1(n5436), .A2(n6690), .A3(n6688), .ZN(n5418) );
  NAND2_X1 U5569 ( .A1(n4486), .A2(REIP_REG_17__SCAN_IN), .ZN(n4487) );
  NOR2_X2 U5570 ( .A1(n5418), .A2(n4487), .ZN(n5362) );
  NAND2_X1 U5571 ( .A1(n5362), .A2(n4488), .ZN(n5330) );
  OR2_X2 U5572 ( .A1(n5330), .A2(n4489), .ZN(n5269) );
  NOR2_X2 U5573 ( .A1(n5269), .A2(n4490), .ZN(n5259) );
  INV_X1 U5574 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6713) );
  NOR3_X1 U5575 ( .A1(n5237), .A2(REIP_REG_30__SCAN_IN), .A3(n6713), .ZN(n4494) );
  NAND2_X1 U5576 ( .A1(n4498), .A2(n4424), .ZN(n4506) );
  NOR2_X1 U5577 ( .A1(n5240), .A2(n6436), .ZN(n4501) );
  AOI211_X1 U5578 ( .C1(n6424), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n4502), 
        .B(n4501), .ZN(n4503) );
  NAND2_X1 U5579 ( .A1(n4506), .A2(n4505), .ZN(U2958) );
  OR2_X1 U5580 ( .A1(n6284), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6370) );
  INV_X1 U5581 ( .A(n6370), .ZN(n5351) );
  INV_X1 U5582 ( .A(n4631), .ZN(n4627) );
  AOI211_X1 U5583 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4507), .A(n5351), .B(
        n4627), .ZN(n4508) );
  INV_X1 U5584 ( .A(n4508), .ZN(U2788) );
  OR2_X1 U5585 ( .A1(n4584), .A2(n5523), .ZN(n4511) );
  OR2_X1 U5586 ( .A1(n4509), .A2(n4458), .ZN(n4510) );
  NAND2_X1 U5587 ( .A1(n4511), .A2(n4510), .ZN(n6368) );
  NOR2_X1 U5588 ( .A1(n5523), .A2(n5202), .ZN(n4512) );
  AOI21_X1 U5589 ( .B1(n4512), .B2(n5214), .A(READY_N), .ZN(n4513) );
  OR2_X1 U5590 ( .A1(n6368), .A2(n4513), .ZN(n6619) );
  NAND2_X1 U5591 ( .A1(n6619), .A2(n6640), .ZN(n4521) );
  INV_X1 U5592 ( .A(n4521), .ZN(n4514) );
  INV_X1 U5593 ( .A(FLUSH_REG_SCAN_IN), .ZN(n4778) );
  OAI21_X1 U5594 ( .B1(n4514), .B2(n4778), .A(n5892), .ZN(U2793) );
  AND3_X1 U5595 ( .A1(n4803), .A2(n6617), .A3(n4515), .ZN(n4516) );
  MUX2_X1 U5596 ( .A(n4516), .B(n4593), .S(n4584), .Z(n4520) );
  NAND2_X1 U5597 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  AND2_X1 U5598 ( .A1(n4520), .A2(n4519), .ZN(n6618) );
  INV_X1 U5599 ( .A(MORE_REG_SCAN_IN), .ZN(n4522) );
  MUX2_X1 U5600 ( .A(n6618), .B(n4522), .S(n4521), .Z(n4523) );
  INV_X1 U5601 ( .A(n4523), .ZN(U3471) );
  INV_X1 U5602 ( .A(n6630), .ZN(n4524) );
  NOR2_X1 U5603 ( .A1(n6601), .A2(n4524), .ZN(n4525) );
  AOI222_X1 U5604 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6409), .B1(n6746), .B2(
        DATAO_REG_18__SCAN_IN), .C1(n6744), .C2(UWORD_REG_2__SCAN_IN), .ZN(
        n4527) );
  INV_X1 U5605 ( .A(n4527), .ZN(U2905) );
  AOI222_X1 U5606 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_15__SCAN_IN), .C1(n6744), .C2(LWORD_REG_15__SCAN_IN), .ZN(
        n4528) );
  INV_X1 U5607 ( .A(n4528), .ZN(U2908) );
  AOI222_X1 U5608 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_12__SCAN_IN), .C1(n6744), .C2(LWORD_REG_12__SCAN_IN), .ZN(
        n4529) );
  INV_X1 U5609 ( .A(n4529), .ZN(U2911) );
  AOI222_X1 U5610 ( .A1(EAX_REG_3__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_3__SCAN_IN), .C1(n6744), .C2(LWORD_REG_3__SCAN_IN), .ZN(
        n4530) );
  INV_X1 U5611 ( .A(n4530), .ZN(U2920) );
  AOI222_X1 U5612 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_4__SCAN_IN), .C1(n6744), .C2(LWORD_REG_4__SCAN_IN), .ZN(
        n4531) );
  INV_X1 U5613 ( .A(n4531), .ZN(U2919) );
  AOI222_X1 U5614 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_9__SCAN_IN), .C1(n6744), .C2(LWORD_REG_9__SCAN_IN), .ZN(
        n4532) );
  INV_X1 U5615 ( .A(n4532), .ZN(U2914) );
  AOI222_X1 U5616 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6409), .B1(n6746), .B2(
        DATAO_REG_21__SCAN_IN), .C1(n6744), .C2(UWORD_REG_5__SCAN_IN), .ZN(
        n4533) );
  INV_X1 U5617 ( .A(n4533), .ZN(U2902) );
  AOI222_X1 U5618 ( .A1(EAX_REG_1__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_1__SCAN_IN), .C1(n6744), .C2(LWORD_REG_1__SCAN_IN), .ZN(
        n4534) );
  INV_X1 U5619 ( .A(n4534), .ZN(U2922) );
  AOI222_X1 U5620 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_8__SCAN_IN), .C1(n6744), .C2(LWORD_REG_8__SCAN_IN), .ZN(
        n4535) );
  INV_X1 U5621 ( .A(n4535), .ZN(U2915) );
  INV_X1 U5622 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4827) );
  AOI222_X1 U5623 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6745), .B1(n6746), .B2(
        DATAO_REG_0__SCAN_IN), .C1(n6744), .C2(LWORD_REG_0__SCAN_IN), .ZN(
        n4536) );
  INV_X1 U5624 ( .A(n4536), .ZN(U2923) );
  INV_X1 U5625 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5626 ( .A1(n6745), .A2(EAX_REG_7__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n4537) );
  OAI21_X1 U5627 ( .B1(n6408), .B2(n4538), .A(n4537), .ZN(U2916) );
  INV_X1 U5628 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4540) );
  AOI22_X1 U5629 ( .A1(n6409), .A2(EAX_REG_19__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4539) );
  OAI21_X1 U5630 ( .B1(n6408), .B2(n4540), .A(n4539), .ZN(U2904) );
  INV_X1 U5631 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5632 ( .A1(n6745), .A2(EAX_REG_5__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n4541) );
  OAI21_X1 U5633 ( .B1(n6408), .B2(n4542), .A(n4541), .ZN(U2918) );
  INV_X1 U5634 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5635 ( .A1(n6745), .A2(EAX_REG_2__SCAN_IN), .B1(n6744), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4543) );
  OAI21_X1 U5636 ( .B1(n6408), .B2(n4544), .A(n4543), .ZN(U2921) );
  INV_X1 U5637 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4546) );
  AOI22_X1 U5638 ( .A1(n6409), .A2(EAX_REG_17__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4545) );
  OAI21_X1 U5639 ( .B1(n6408), .B2(n4546), .A(n4545), .ZN(U2906) );
  INV_X1 U5640 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4548) );
  AOI22_X1 U5641 ( .A1(n6409), .A2(EAX_REG_25__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U5642 ( .B1(n6408), .B2(n4548), .A(n4547), .ZN(U2898) );
  INV_X1 U5643 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4550) );
  INV_X1 U5644 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n4549) );
  OAI222_X1 U5645 ( .A1(n4550), .A2(n6408), .B1(n4553), .B2(n5671), .C1(n5208), 
        .C2(n4549), .ZN(U2912) );
  INV_X1 U5646 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4554) );
  INV_X1 U5647 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4552) );
  INV_X1 U5648 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4551) );
  OAI222_X1 U5649 ( .A1(n4554), .A2(n6408), .B1(n4553), .B2(n4552), .C1(n5208), 
        .C2(n4551), .ZN(U2917) );
  INV_X1 U5650 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4556) );
  INV_X1 U5651 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4555) );
  OAI222_X1 U5652 ( .A1(n4556), .A2(n6408), .B1(n4572), .B2(n4099), .C1(n5208), 
        .C2(n4555), .ZN(U2907) );
  INV_X1 U5653 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4558) );
  INV_X1 U5654 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4557) );
  OAI222_X1 U5655 ( .A1(n4558), .A2(n6408), .B1(n4572), .B2(n4165), .C1(n5208), 
        .C2(n4557), .ZN(U2903) );
  INV_X1 U5656 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4561) );
  INV_X1 U5657 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4560) );
  INV_X1 U5658 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4559) );
  OAI222_X1 U5659 ( .A1(n4561), .A2(n6408), .B1(n4572), .B2(n4560), .C1(n5208), 
        .C2(n4559), .ZN(U2899) );
  INV_X1 U5660 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4563) );
  INV_X1 U5661 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n4562) );
  OAI222_X1 U5662 ( .A1(n4563), .A2(n6408), .B1(n4572), .B2(n4366), .C1(n5208), 
        .C2(n4562), .ZN(U2893) );
  INV_X1 U5663 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4566) );
  INV_X1 U5664 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4565) );
  INV_X1 U5665 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4564) );
  OAI222_X1 U5666 ( .A1(n4566), .A2(n6408), .B1(n4572), .B2(n4565), .C1(n5208), 
        .C2(n4564), .ZN(U2896) );
  INV_X1 U5667 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4569) );
  INV_X1 U5668 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4568) );
  INV_X1 U5669 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n4567) );
  OAI222_X1 U5670 ( .A1(n4569), .A2(n6408), .B1(n4572), .B2(n4568), .C1(n5208), 
        .C2(n4567), .ZN(U2895) );
  INV_X1 U5671 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4573) );
  INV_X1 U5672 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4570) );
  OAI222_X1 U5673 ( .A1(n5208), .A2(n4573), .B1(n4572), .B2(n4571), .C1(n6408), 
        .C2(n4570), .ZN(U2901) );
  INV_X1 U5674 ( .A(n6635), .ZN(n6728) );
  INV_X1 U5675 ( .A(n4574), .ZN(n4601) );
  MUX2_X1 U5676 ( .A(n4593), .B(n4803), .S(n4584), .Z(n4586) );
  OR2_X1 U5677 ( .A1(n4458), .A2(n5202), .ZN(n4575) );
  OAI211_X1 U5678 ( .C1(n6601), .C2(n4589), .A(n4576), .B(n4575), .ZN(n4577)
         );
  INV_X1 U5679 ( .A(n4577), .ZN(n4583) );
  INV_X1 U5680 ( .A(n4578), .ZN(n4579) );
  NAND3_X1 U5681 ( .A1(n4808), .A2(n4581), .A3(n4580), .ZN(n4582) );
  AOI21_X1 U5682 ( .B1(n4584), .B2(n4583), .A(n4582), .ZN(n4585) );
  NAND2_X1 U5683 ( .A1(n4586), .A2(n4585), .ZN(n6604) );
  NOR2_X1 U5684 ( .A1(n6642), .A2(n4792), .ZN(n6649) );
  AOI22_X1 U5685 ( .A1(n6640), .A2(n6604), .B1(FLUSH_REG_SCAN_IN), .B2(n6649), 
        .ZN(n6367) );
  INV_X1 U5686 ( .A(n6732), .ZN(n4604) );
  AOI21_X1 U5687 ( .B1(n6728), .B2(n4601), .A(n4604), .ZN(n4606) );
  INV_X1 U5688 ( .A(n4588), .ZN(n4592) );
  INV_X1 U5689 ( .A(n4589), .ZN(n4590) );
  AND3_X1 U5690 ( .A1(n4785), .A2(n4807), .A3(n4590), .ZN(n4591) );
  NAND2_X1 U5691 ( .A1(n4592), .A2(n4591), .ZN(n6600) );
  NAND2_X1 U5692 ( .A1(n6101), .A2(n6600), .ZN(n4599) );
  NAND2_X1 U5693 ( .A1(n4593), .A2(n4803), .ZN(n4766) );
  XNOR2_X1 U5694 ( .A(n4574), .B(n6980), .ZN(n4597) );
  INV_X1 U5695 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U5696 ( .A(n5190), .B(n6980), .ZN(n4594) );
  NAND2_X1 U5697 ( .A1(n6601), .A2(n4594), .ZN(n4595) );
  OAI21_X1 U5698 ( .B1(n4597), .B2(n4770), .A(n4595), .ZN(n4596) );
  AOI21_X1 U5699 ( .B1(n4766), .B2(n4597), .A(n4596), .ZN(n4598) );
  NAND2_X1 U5700 ( .A1(n4599), .A2(n4598), .ZN(n4761) );
  NOR2_X1 U5701 ( .A1(n4786), .A2(n6726), .ZN(n5184) );
  INV_X1 U5702 ( .A(n5184), .ZN(n4600) );
  INV_X1 U5703 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5893) );
  INV_X1 U5704 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6470) );
  AOI22_X1 U5705 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5893), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6470), .ZN(n5185) );
  NOR2_X1 U5706 ( .A1(n4600), .A2(n5185), .ZN(n4603) );
  NOR3_X1 U5707 ( .A1(n6635), .A2(n6980), .A3(n4601), .ZN(n4602) );
  AOI211_X1 U5708 ( .C1(n6364), .C2(n4761), .A(n4603), .B(n4602), .ZN(n4605)
         );
  OAI22_X1 U5709 ( .A1(n4606), .A2(n3202), .B1(n4605), .B2(n4604), .ZN(U3459)
         );
  NOR2_X1 U5710 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4607)
         );
  NOR2_X1 U5711 ( .A1(n4608), .A2(n4607), .ZN(n5588) );
  INV_X1 U5712 ( .A(n5588), .ZN(n4613) );
  OAI21_X1 U5713 ( .B1(n4611), .B2(n4610), .A(n4609), .ZN(n5595) );
  OAI222_X1 U5714 ( .A1(n4613), .A2(n5620), .B1(n5618), .B2(n4612), .C1(n5623), 
        .C2(n5595), .ZN(U2859) );
  OAI21_X1 U5715 ( .B1(n4614), .B2(n4616), .A(n4615), .ZN(n5584) );
  XNOR2_X1 U5716 ( .A(n4617), .B(n5214), .ZN(n5576) );
  AOI22_X1 U5717 ( .A1(n4402), .A2(n5576), .B1(n5621), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4618) );
  OAI21_X1 U5718 ( .B1(n5584), .B2(n5623), .A(n4618), .ZN(U2858) );
  INV_X1 U5719 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6740) );
  OAI21_X1 U5720 ( .B1(n6075), .B2(n6740), .A(n4619), .ZN(n4623) );
  INV_X1 U5721 ( .A(n6039), .ZN(n4621) );
  AOI21_X1 U5722 ( .B1(n4621), .B2(n4620), .A(n6726), .ZN(n4622) );
  AOI211_X1 U5723 ( .C1(n5588), .C2(n6463), .A(n4623), .B(n4622), .ZN(n4626)
         );
  OR2_X1 U5724 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4674)
         );
  NAND3_X1 U5725 ( .A1(n4674), .A2(n4444), .A3(n3500), .ZN(n4625) );
  NAND2_X1 U5726 ( .A1(n4626), .A2(n4625), .ZN(U3018) );
  OR2_X1 U5727 ( .A1(n4631), .A2(n4628), .ZN(n4629) );
  AOI22_X1 U5728 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5729 ( .A1(n6415), .A2(DATAI_4_), .ZN(n4658) );
  NAND2_X1 U5730 ( .A1(n4632), .A2(n4658), .ZN(U2928) );
  AOI22_X1 U5731 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5732 ( .A1(n6415), .A2(DATAI_2_), .ZN(n4664) );
  NAND2_X1 U5733 ( .A1(n4633), .A2(n4664), .ZN(U2926) );
  AOI22_X1 U5734 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5735 ( .A1(n6415), .A2(DATAI_3_), .ZN(n4662) );
  NAND2_X1 U5736 ( .A1(n4634), .A2(n4662), .ZN(U2927) );
  AOI22_X1 U5737 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U5738 ( .A1(n6415), .A2(DATAI_1_), .ZN(n4646) );
  NAND2_X1 U5739 ( .A1(n4635), .A2(n4646), .ZN(U2925) );
  OAI21_X1 U5740 ( .B1(n4638), .B2(n4636), .A(n4637), .ZN(n4943) );
  AND2_X1 U5741 ( .A1(n5868), .A2(REIP_REG_1__SCAN_IN), .ZN(n4938) );
  NOR2_X1 U5742 ( .A1(n4639), .A2(n6470), .ZN(n4640) );
  AOI211_X1 U5743 ( .C1(n6463), .C2(n5576), .A(n4938), .B(n4640), .ZN(n4643)
         );
  NAND3_X1 U5744 ( .A1(n6021), .A2(n6470), .A3(n4641), .ZN(n4642) );
  OAI211_X1 U5745 ( .C1(n4943), .C2(n6084), .A(n4643), .B(n4642), .ZN(U3017)
         );
  AOI22_X1 U5746 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n4644) );
  INV_X1 U5747 ( .A(DATAI_12_), .ZN(n5669) );
  OR2_X1 U5748 ( .A1(n4813), .A2(n5669), .ZN(n4694) );
  NAND2_X1 U5749 ( .A1(n4644), .A2(n4694), .ZN(U2936) );
  AOI22_X1 U5750 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4645) );
  NAND2_X1 U5751 ( .A1(n6415), .A2(DATAI_9_), .ZN(n4655) );
  NAND2_X1 U5752 ( .A1(n4645), .A2(n4655), .ZN(U2948) );
  AOI22_X1 U5753 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U5754 ( .A1(n4647), .A2(n4646), .ZN(U2940) );
  AOI22_X1 U5755 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5756 ( .A1(n6415), .A2(DATAI_0_), .ZN(n4696) );
  NAND2_X1 U5757 ( .A1(n4648), .A2(n4696), .ZN(U2939) );
  AOI22_X1 U5758 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4649) );
  NAND2_X1 U5759 ( .A1(n6415), .A2(DATAI_7_), .ZN(n4651) );
  NAND2_X1 U5760 ( .A1(n4649), .A2(n4651), .ZN(U2931) );
  AOI22_X1 U5761 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4650) );
  NAND2_X1 U5762 ( .A1(n6415), .A2(DATAI_6_), .ZN(n4670) );
  NAND2_X1 U5763 ( .A1(n4650), .A2(n4670), .ZN(U2945) );
  AOI22_X1 U5764 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U5765 ( .A1(n4652), .A2(n4651), .ZN(U2946) );
  AOI22_X1 U5766 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U5767 ( .A1(n6415), .A2(DATAI_8_), .ZN(n4668) );
  NAND2_X1 U5768 ( .A1(n4653), .A2(n4668), .ZN(U2932) );
  AOI22_X1 U5769 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U5770 ( .A1(n6415), .A2(DATAI_5_), .ZN(n4666) );
  NAND2_X1 U5771 ( .A1(n4654), .A2(n4666), .ZN(U2929) );
  AOI22_X1 U5772 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n4656) );
  NAND2_X1 U5773 ( .A1(n4656), .A2(n4655), .ZN(U2933) );
  AOI22_X1 U5774 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5775 ( .A1(n6415), .A2(DATAI_13_), .ZN(n4660) );
  NAND2_X1 U5776 ( .A1(n4657), .A2(n4660), .ZN(U2937) );
  AOI22_X1 U5777 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U5778 ( .A1(n4659), .A2(n4658), .ZN(U2943) );
  AOI22_X1 U5779 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5780 ( .A1(n4661), .A2(n4660), .ZN(U2952) );
  AOI22_X1 U5781 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4663) );
  NAND2_X1 U5782 ( .A1(n4663), .A2(n4662), .ZN(U2942) );
  AOI22_X1 U5783 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5784 ( .A1(n4665), .A2(n4664), .ZN(U2941) );
  AOI22_X1 U5785 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5786 ( .A1(n4667), .A2(n4666), .ZN(U2944) );
  AOI22_X1 U5787 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5788 ( .A1(n4669), .A2(n4668), .ZN(U2947) );
  AOI22_X1 U5789 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5790 ( .A1(n4671), .A2(n4670), .ZN(U2930) );
  NAND2_X1 U5791 ( .A1(n5884), .A2(n4672), .ZN(n4673) );
  AOI22_X1 U5792 ( .A1(n4673), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n5868), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4676) );
  NAND3_X1 U5793 ( .A1(n4674), .A2(n4424), .A3(n3500), .ZN(n4675) );
  OAI211_X1 U5794 ( .C1(n5595), .C2(n5885), .A(n4676), .B(n4675), .ZN(U2986)
         );
  AOI222_X1 U5795 ( .A1(EAX_REG_15__SCAN_IN), .A2(n4692), .B1(DATAI_15_), .B2(
        n6415), .C1(n4693), .C2(LWORD_REG_15__SCAN_IN), .ZN(n4677) );
  INV_X1 U5796 ( .A(n4677), .ZN(U2954) );
  INV_X1 U5797 ( .A(n4679), .ZN(n4680) );
  OAI21_X1 U5798 ( .B1(n4681), .B2(n4678), .A(n4680), .ZN(n6425) );
  OR2_X1 U5799 ( .A1(n4683), .A2(n4682), .ZN(n4684) );
  AND2_X1 U5800 ( .A1(n4684), .A2(n4689), .ZN(n6462) );
  AOI22_X1 U5801 ( .A1(n6462), .A2(n4402), .B1(n5621), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4685) );
  OAI21_X1 U5802 ( .B1(n6425), .B2(n5623), .A(n4685), .ZN(U2857) );
  NAND2_X1 U5803 ( .A1(n4679), .A2(n4686), .ZN(n4747) );
  OR2_X1 U5804 ( .A1(n4679), .A2(n4686), .ZN(n4687) );
  NAND2_X1 U5805 ( .A1(n4747), .A2(n4687), .ZN(n5564) );
  AOI21_X1 U5806 ( .B1(n4690), .B2(n4689), .A(n4688), .ZN(n5554) );
  AOI22_X1 U5807 ( .A1(n4402), .A2(n5554), .B1(n5621), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4691) );
  OAI21_X1 U5808 ( .B1(n5564), .B2(n5623), .A(n4691), .ZN(U2856) );
  AOI22_X1 U5809 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4693), .B1(n4692), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5810 ( .A1(n4695), .A2(n4694), .ZN(U2951) );
  AOI22_X1 U5811 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U5812 ( .A1(n4697), .A2(n4696), .ZN(U2924) );
  AND2_X1 U5813 ( .A1(n4699), .A2(n6238), .ZN(n4700) );
  AND2_X1 U5814 ( .A1(n4709), .A2(n3892), .ZN(n4894) );
  NOR2_X1 U5815 ( .A1(n6284), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6200) );
  INV_X1 U5816 ( .A(n6200), .ZN(n6244) );
  OAI21_X1 U5817 ( .B1(n4709), .B2(n5885), .A(n6244), .ZN(n4705) );
  AND2_X1 U5818 ( .A1(n3087), .A2(n3895), .ZN(n6283) );
  NAND2_X1 U5819 ( .A1(n6101), .A2(n4703), .ZN(n6485) );
  INV_X1 U5820 ( .A(n6485), .ZN(n4915) );
  INV_X1 U5821 ( .A(n4738), .ZN(n4704) );
  AOI21_X1 U5822 ( .B1(n6283), .B2(n4915), .A(n4704), .ZN(n4710) );
  NAND2_X1 U5823 ( .A1(n4705), .A2(n4710), .ZN(n4708) );
  NAND2_X1 U5824 ( .A1(n6650), .A2(n4792), .ZN(n4706) );
  NAND2_X1 U5825 ( .A1(n4735), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4714)
         );
  INV_X1 U5826 ( .A(n4710), .ZN(n4711) );
  AOI22_X1 U5827 ( .A1(n4711), .A2(n6484), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4829), .ZN(n4739) );
  INV_X1 U5828 ( .A(DATAI_6_), .ZN(n7023) );
  AND2_X1 U5829 ( .A1(n4737), .A2(n3393), .ZN(n6548) );
  OAI22_X1 U5830 ( .A1(n4739), .A2(n6354), .B1(n6271), .B2(n4738), .ZN(n4712)
         );
  AOI21_X1 U5831 ( .B1(n4741), .B2(n6550), .A(n4712), .ZN(n4713) );
  OAI211_X1 U5832 ( .C1(n4744), .C2(n6558), .A(n4714), .B(n4713), .ZN(U3146)
         );
  NAND2_X1 U5833 ( .A1(n4735), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4717)
         );
  INV_X1 U5834 ( .A(n6589), .ZN(n6311) );
  INV_X1 U5835 ( .A(DATAI_7_), .ZN(n4905) );
  OAI22_X1 U5836 ( .A1(n4739), .A2(n6361), .B1(n6588), .B2(n4738), .ZN(n4715)
         );
  AOI21_X1 U5837 ( .B1(n4741), .B2(n6311), .A(n4715), .ZN(n4716) );
  OAI211_X1 U5838 ( .C1(n4744), .C2(n6598), .A(n4717), .B(n4716), .ZN(U3147)
         );
  NAND2_X1 U5839 ( .A1(n4735), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4720)
         );
  NAND2_X1 U5840 ( .A1(n6431), .A2(DATAI_16_), .ZN(n6560) );
  INV_X1 U5841 ( .A(n6560), .ZN(n6525) );
  INV_X1 U5842 ( .A(DATAI_0_), .ZN(n4828) );
  AND2_X1 U5843 ( .A1(n4737), .A2(n3780), .ZN(n6524) );
  OAI22_X1 U5844 ( .A1(n4739), .A2(n6330), .B1(n6559), .B2(n4738), .ZN(n4718)
         );
  AOI21_X1 U5845 ( .B1(n4741), .B2(n6525), .A(n4718), .ZN(n4719) );
  OAI211_X1 U5846 ( .C1(n4744), .C2(n6565), .A(n4720), .B(n4719), .ZN(U3140)
         );
  NAND2_X1 U5847 ( .A1(n6431), .A2(DATAI_29_), .ZN(n6586) );
  NAND2_X1 U5848 ( .A1(n4735), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4723)
         );
  INV_X1 U5849 ( .A(DATAI_5_), .ZN(n4909) );
  OAI22_X1 U5850 ( .A1(n4739), .A2(n6350), .B1(n6580), .B2(n4738), .ZN(n4721)
         );
  AOI21_X1 U5851 ( .B1(n4741), .B2(n6303), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5852 ( .C1(n4744), .C2(n6586), .A(n4723), .B(n4722), .ZN(U3145)
         );
  NAND2_X1 U5853 ( .A1(n6431), .A2(DATAI_28_), .ZN(n6547) );
  NAND2_X1 U5854 ( .A1(n4735), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4727)
         );
  NAND2_X1 U5855 ( .A1(n6431), .A2(DATAI_20_), .ZN(n6507) );
  INV_X1 U5856 ( .A(n6507), .ZN(n6543) );
  INV_X1 U5857 ( .A(DATAI_4_), .ZN(n4822) );
  OAI22_X1 U5858 ( .A1(n4739), .A2(n6346), .B1(n6264), .B2(n4738), .ZN(n4725)
         );
  AOI21_X1 U5859 ( .B1(n4741), .B2(n6543), .A(n4725), .ZN(n4726) );
  OAI211_X1 U5860 ( .C1(n4744), .C2(n6547), .A(n4727), .B(n4726), .ZN(U3144)
         );
  NAND2_X1 U5861 ( .A1(n4735), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4731)
         );
  NAND2_X1 U5862 ( .A1(n6431), .A2(DATAI_19_), .ZN(n6574) );
  INV_X1 U5863 ( .A(DATAI_3_), .ZN(n4821) );
  OAI22_X1 U5864 ( .A1(n4739), .A2(n6342), .B1(n6573), .B2(n4738), .ZN(n4729)
         );
  AOI21_X1 U5865 ( .B1(n4741), .B2(n6539), .A(n4729), .ZN(n4730) );
  OAI211_X1 U5866 ( .C1(n4744), .C2(n6579), .A(n4731), .B(n4730), .ZN(U3143)
         );
  NAND2_X1 U5867 ( .A1(n6431), .A2(DATAI_26_), .ZN(n6537) );
  NAND2_X1 U5868 ( .A1(n4735), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4734)
         );
  NAND2_X1 U5869 ( .A1(n6431), .A2(DATAI_18_), .ZN(n6500) );
  INV_X1 U5870 ( .A(n6500), .ZN(n6533) );
  INV_X1 U5871 ( .A(DATAI_2_), .ZN(n4826) );
  OAI22_X1 U5872 ( .A1(n4739), .A2(n6338), .B1(n6257), .B2(n4738), .ZN(n4732)
         );
  AOI21_X1 U5873 ( .B1(n4741), .B2(n6533), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5874 ( .C1(n4744), .C2(n6537), .A(n4734), .B(n4733), .ZN(U3142)
         );
  NAND2_X1 U5875 ( .A1(n6431), .A2(DATAI_25_), .ZN(n6572) );
  NAND2_X1 U5876 ( .A1(n4735), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4743)
         );
  NAND2_X1 U5877 ( .A1(n6431), .A2(DATAI_17_), .ZN(n6567) );
  INV_X1 U5878 ( .A(n6567), .ZN(n6529) );
  INV_X1 U5879 ( .A(DATAI_1_), .ZN(n4824) );
  OAI22_X1 U5880 ( .A1(n4739), .A2(n6334), .B1(n6566), .B2(n4738), .ZN(n4740)
         );
  AOI21_X1 U5881 ( .B1(n4741), .B2(n6529), .A(n4740), .ZN(n4742) );
  OAI211_X1 U5882 ( .C1(n4744), .C2(n6572), .A(n4743), .B(n4742), .ZN(U3141)
         );
  INV_X1 U5883 ( .A(n4745), .ZN(n4746) );
  NAND2_X1 U5884 ( .A1(n4747), .A2(n4746), .ZN(n4748) );
  NAND2_X1 U5885 ( .A1(n4907), .A2(n4748), .ZN(n5553) );
  OR2_X1 U5886 ( .A1(n4749), .A2(n4688), .ZN(n4751) );
  NAND2_X1 U5887 ( .A1(n4751), .A2(n4750), .ZN(n4861) );
  INV_X1 U5888 ( .A(n4861), .ZN(n5538) );
  AOI22_X1 U5889 ( .A1(n4402), .A2(n5538), .B1(n5621), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4752) );
  OAI21_X1 U5890 ( .B1(n5553), .B2(n5623), .A(n4752), .ZN(U2855) );
  XNOR2_X1 U5891 ( .A(n4754), .B(n4753), .ZN(n4949) );
  AOI22_X1 U5892 ( .A1(n6061), .A2(n4755), .B1(n6070), .B2(n4756), .ZN(n6466)
         );
  NAND2_X1 U5893 ( .A1(n6464), .A2(n4758), .ZN(n6472) );
  NAND2_X1 U5894 ( .A1(n6466), .A2(n6472), .ZN(n4863) );
  OAI21_X1 U5895 ( .B1(n6469), .B2(n4756), .A(n6061), .ZN(n6076) );
  INV_X1 U5896 ( .A(n6076), .ZN(n4757) );
  NOR2_X1 U5897 ( .A1(n4758), .A2(n4757), .ZN(n4865) );
  AOI22_X1 U5898 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4863), .B1(n4865), 
        .B2(n3575), .ZN(n4760) );
  AND2_X1 U5899 ( .A1(n5868), .A2(REIP_REG_3__SCAN_IN), .ZN(n4944) );
  AOI21_X1 U5900 ( .B1(n6463), .B2(n5554), .A(n4944), .ZN(n4759) );
  OAI211_X1 U5901 ( .C1(n4949), .C2(n6084), .A(n4760), .B(n4759), .ZN(U3015)
         );
  MUX2_X1 U5902 ( .A(n6980), .B(n4761), .S(n6604), .Z(n6609) );
  MUX2_X1 U5903 ( .A(n4762), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4574), 
        .Z(n4764) );
  NOR2_X1 U5904 ( .A1(n4764), .A2(n4763), .ZN(n4765) );
  NAND2_X1 U5905 ( .A1(n4766), .A2(n4765), .ZN(n4774) );
  NAND2_X1 U5906 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n6980), .ZN(n4767) );
  XNOR2_X1 U5907 ( .A(n4767), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4772)
         );
  OAI21_X1 U5908 ( .B1(n4574), .B2(n4776), .A(n4768), .ZN(n4769) );
  NOR2_X1 U5909 ( .A1(n4769), .A2(n4306), .ZN(n6106) );
  NOR2_X1 U5910 ( .A1(n4770), .A2(n6106), .ZN(n4771) );
  AOI21_X1 U5911 ( .B1(n6601), .B2(n4772), .A(n4771), .ZN(n4773) );
  NAND2_X1 U5912 ( .A1(n4774), .A2(n4773), .ZN(n4775) );
  AOI21_X1 U5913 ( .B1(n3087), .B2(n6600), .A(n4775), .ZN(n6107) );
  MUX2_X1 U5914 ( .A(n4776), .B(n6107), .S(n6604), .Z(n6611) );
  INV_X1 U5915 ( .A(n6611), .ZN(n4777) );
  NAND3_X1 U5916 ( .A1(n6609), .A2(n4777), .A3(n4786), .ZN(n4781) );
  AND2_X1 U5917 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4778), .ZN(n4779) );
  NAND2_X1 U5918 ( .A1(n4763), .A2(n4779), .ZN(n4780) );
  MUX2_X1 U5919 ( .A(FLUSH_REG_SCAN_IN), .B(n6604), .S(n4786), .Z(n4782) );
  INV_X1 U5920 ( .A(n6199), .ZN(n4912) );
  NOR2_X1 U5921 ( .A1(n4783), .A2(n4912), .ZN(n4784) );
  XNOR2_X1 U5922 ( .A(n4784), .B(n6991), .ZN(n6365) );
  INV_X1 U5923 ( .A(n4785), .ZN(n6363) );
  NAND3_X1 U5924 ( .A1(n6365), .A2(n6363), .A3(n4786), .ZN(n4787) );
  NAND2_X1 U5925 ( .A1(n4788), .A2(n4787), .ZN(n6622) );
  INV_X1 U5926 ( .A(n6622), .ZN(n4789) );
  OAI21_X1 U5927 ( .B1(n6624), .B2(n4790), .A(n4789), .ZN(n4793) );
  OAI21_X1 U5928 ( .B1(n4793), .B2(FLUSH_REG_SCAN_IN), .A(n6649), .ZN(n4791)
         );
  NOR2_X1 U5929 ( .A1(n4793), .A2(n4792), .ZN(n6634) );
  INV_X1 U5930 ( .A(n3895), .ZN(n5016) );
  AND2_X1 U5931 ( .A1(n6725), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6102) );
  OAI22_X1 U5932 ( .A1(n3892), .A2(n6284), .B1(n5016), .B2(n6102), .ZN(n4794)
         );
  OAI21_X1 U5933 ( .B1(n6634), .B2(n4794), .A(n6475), .ZN(n4795) );
  OAI21_X1 U5934 ( .B1(n6475), .B2(n6281), .A(n4795), .ZN(U3465) );
  NOR2_X1 U5935 ( .A1(n6238), .A2(n4796), .ZN(n4797) );
  NAND2_X1 U5936 ( .A1(n4975), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4978) );
  NAND2_X1 U5937 ( .A1(n4978), .A2(n6239), .ZN(n5012) );
  INV_X1 U5938 ( .A(n5012), .ZN(n4799) );
  NAND2_X1 U5939 ( .A1(n6238), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6095) );
  INV_X1 U5940 ( .A(n6095), .ZN(n6100) );
  NAND2_X1 U5941 ( .A1(n5128), .A2(n6100), .ZN(n4911) );
  AOI21_X1 U5942 ( .B1(n4799), .B2(n4911), .A(n6284), .ZN(n4801) );
  INV_X1 U5943 ( .A(n3087), .ZN(n6207) );
  OAI22_X1 U5944 ( .A1(n5051), .A2(n6244), .B1(n6207), .B2(n6102), .ZN(n4800)
         );
  OAI21_X1 U5945 ( .B1(n4801), .B2(n4800), .A(n6475), .ZN(n4802) );
  OAI21_X1 U5946 ( .B1(n6475), .B2(n6839), .A(n4802), .ZN(U3462) );
  NAND3_X1 U5947 ( .A1(n3149), .A2(n4805), .A3(n3393), .ZN(n4806) );
  OAI22_X1 U5948 ( .A1(n4808), .A2(n6638), .B1(n4807), .B2(n4806), .ZN(n4809)
         );
  INV_X1 U5949 ( .A(n4809), .ZN(n4810) );
  AND2_X1 U5950 ( .A1(n4817), .A2(n4814), .ZN(n4815) );
  INV_X1 U5951 ( .A(n5660), .ZN(n4820) );
  INV_X1 U5952 ( .A(n4817), .ZN(n4818) );
  INV_X1 U5953 ( .A(n5661), .ZN(n4819) );
  INV_X1 U5954 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6977) );
  OAI222_X1 U5955 ( .A1(n5564), .A2(n5680), .B1(n5679), .B2(n4821), .C1(n5678), 
        .C2(n6977), .ZN(U2888) );
  INV_X1 U5956 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6863) );
  OAI222_X1 U5957 ( .A1(n5553), .A2(n5680), .B1(n5679), .B2(n4822), .C1(n5678), 
        .C2(n6863), .ZN(U2887) );
  INV_X1 U5958 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4823) );
  OAI222_X1 U5959 ( .A1(n5584), .A2(n5680), .B1(n5679), .B2(n4824), .C1(n5678), 
        .C2(n4823), .ZN(U2890) );
  INV_X1 U5960 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4825) );
  OAI222_X1 U5961 ( .A1(n6425), .A2(n5680), .B1(n5679), .B2(n4826), .C1(n5678), 
        .C2(n4825), .ZN(U2889) );
  OAI222_X1 U5962 ( .A1(n5595), .A2(n5680), .B1(n5679), .B2(n4828), .C1(n5678), 
        .C2(n4827), .ZN(U2891) );
  INV_X1 U5963 ( .A(n4829), .ZN(n4830) );
  NOR2_X1 U5964 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4830), .ZN(n4893)
         );
  OAI21_X1 U5965 ( .B1(n6477), .B2(n6326), .A(n6113), .ZN(n6486) );
  NOR3_X1 U5966 ( .A1(n6486), .A2(n6839), .A3(n6487), .ZN(n4833) );
  OAI21_X1 U5967 ( .B1(n4834), .B2(n4894), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4831) );
  NAND3_X1 U5968 ( .A1(n6485), .A2(n6484), .A3(n4831), .ZN(n4832) );
  INV_X1 U5969 ( .A(n4898), .ZN(n4842) );
  INV_X1 U5970 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4841) );
  AND2_X1 U5971 ( .A1(n4915), .A2(n6484), .ZN(n6476) );
  NAND2_X1 U5972 ( .A1(n6476), .A2(n3087), .ZN(n4837) );
  NOR2_X1 U5973 ( .A1(n4835), .A2(n6326), .ZN(n6478) );
  NAND3_X1 U5974 ( .A1(n6478), .A2(n6477), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U5975 ( .A1(n4837), .A2(n4836), .ZN(n4892) );
  AOI22_X1 U5976 ( .A1(n6524), .A2(n4893), .B1(n6562), .B2(n4892), .ZN(n4838)
         );
  OAI21_X1 U5977 ( .B1(n5010), .B2(n6565), .A(n4838), .ZN(n4839) );
  AOI21_X1 U5978 ( .B1(n6525), .B2(n4894), .A(n4839), .ZN(n4840) );
  OAI21_X1 U5979 ( .B1(n4842), .B2(n4841), .A(n4840), .ZN(U3132) );
  OAI21_X1 U5980 ( .B1(n6239), .B2(n6095), .A(n6484), .ZN(n4846) );
  INV_X1 U5981 ( .A(n4703), .ZN(n6097) );
  NOR2_X1 U5982 ( .A1(n5014), .A2(n6839), .ZN(n4848) );
  AOI21_X1 U5983 ( .B1(n6320), .B2(n3895), .A(n4848), .ZN(n4843) );
  NAND3_X1 U5984 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6610), .ZN(n6319) );
  OAI22_X1 U5985 ( .A1(n4846), .A2(n4843), .B1(n6319), .B2(n6326), .ZN(n6592)
         );
  INV_X1 U5986 ( .A(n6592), .ZN(n4858) );
  INV_X1 U5987 ( .A(n4843), .ZN(n4845) );
  INV_X1 U5988 ( .A(n6286), .ZN(n5133) );
  AOI21_X1 U5989 ( .B1(n6284), .B2(n6319), .A(n5133), .ZN(n4844) );
  NOR2_X1 U5990 ( .A1(n6597), .A2(n6537), .ZN(n4850) );
  INV_X1 U5991 ( .A(n4848), .ZN(n6587) );
  OAI22_X1 U5992 ( .A1(n6590), .A2(n6500), .B1(n6257), .B2(n6587), .ZN(n4849)
         );
  AOI211_X1 U5993 ( .C1(n6594), .C2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4850), 
        .B(n4849), .ZN(n4851) );
  OAI21_X1 U5994 ( .B1(n4858), .B2(n6338), .A(n4851), .ZN(U3110) );
  NOR2_X1 U5995 ( .A1(n6597), .A2(n6558), .ZN(n4853) );
  OAI22_X1 U5996 ( .A1(n6590), .A2(n6515), .B1(n6271), .B2(n6587), .ZN(n4852)
         );
  AOI211_X1 U5997 ( .C1(n6594), .C2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4853), 
        .B(n4852), .ZN(n4854) );
  OAI21_X1 U5998 ( .B1(n4858), .B2(n6354), .A(n4854), .ZN(U3114) );
  NOR2_X1 U5999 ( .A1(n6597), .A2(n6547), .ZN(n4856) );
  OAI22_X1 U6000 ( .A1(n6590), .A2(n6507), .B1(n6264), .B2(n6587), .ZN(n4855)
         );
  AOI211_X1 U6001 ( .C1(n6594), .C2(INSTQUEUE_REG_11__4__SCAN_IN), .A(n4856), 
        .B(n4855), .ZN(n4857) );
  OAI21_X1 U6002 ( .B1(n4858), .B2(n6346), .A(n4857), .ZN(U3112) );
  XNOR2_X1 U6003 ( .A(n4860), .B(n4859), .ZN(n5177) );
  NAND2_X1 U6004 ( .A1(n5868), .A2(REIP_REG_4__SCAN_IN), .ZN(n5171) );
  OAI21_X1 U6005 ( .B1(n6088), .B2(n4861), .A(n5171), .ZN(n4862) );
  AOI21_X1 U6006 ( .B1(n4863), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4862), 
        .ZN(n4867) );
  OAI211_X1 U6007 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4865), .B(n4864), .ZN(n4866) );
  OAI211_X1 U6008 ( .C1(n6084), .C2(n5177), .A(n4867), .B(n4866), .ZN(U3014)
         );
  AOI22_X1 U6009 ( .A1(n6528), .A2(n4893), .B1(n6569), .B2(n4892), .ZN(n4869)
         );
  NAND2_X1 U6010 ( .A1(n4894), .A2(n6529), .ZN(n4868) );
  OAI211_X1 U6011 ( .C1(n5010), .C2(n6572), .A(n4869), .B(n4868), .ZN(n4870)
         );
  AOI21_X1 U6012 ( .B1(n4898), .B2(INSTQUEUE_REG_14__1__SCAN_IN), .A(n4870), 
        .ZN(n4871) );
  INV_X1 U6013 ( .A(n4871), .ZN(U3133) );
  AOI22_X1 U6014 ( .A1(n6517), .A2(n4893), .B1(n6593), .B2(n4892), .ZN(n4873)
         );
  NAND2_X1 U6015 ( .A1(n4894), .A2(n6311), .ZN(n4872) );
  OAI211_X1 U6016 ( .C1(n5010), .C2(n6598), .A(n4873), .B(n4872), .ZN(n4874)
         );
  AOI21_X1 U6017 ( .B1(n4898), .B2(INSTQUEUE_REG_14__7__SCAN_IN), .A(n4874), 
        .ZN(n4875) );
  INV_X1 U6018 ( .A(n4875), .ZN(U3139) );
  AOI22_X1 U6019 ( .A1(n6548), .A2(n4893), .B1(n6553), .B2(n4892), .ZN(n4877)
         );
  NAND2_X1 U6020 ( .A1(n4894), .A2(n6550), .ZN(n4876) );
  OAI211_X1 U6021 ( .C1(n5010), .C2(n6558), .A(n4877), .B(n4876), .ZN(n4878)
         );
  AOI21_X1 U6022 ( .B1(n4898), .B2(INSTQUEUE_REG_14__6__SCAN_IN), .A(n4878), 
        .ZN(n4879) );
  INV_X1 U6023 ( .A(n4879), .ZN(U3138) );
  AOI22_X1 U6024 ( .A1(n6538), .A2(n4893), .B1(n6576), .B2(n4892), .ZN(n4881)
         );
  NAND2_X1 U6025 ( .A1(n4894), .A2(n6539), .ZN(n4880) );
  OAI211_X1 U6026 ( .C1(n5010), .C2(n6579), .A(n4881), .B(n4880), .ZN(n4882)
         );
  AOI21_X1 U6027 ( .B1(n4898), .B2(INSTQUEUE_REG_14__3__SCAN_IN), .A(n4882), 
        .ZN(n4883) );
  INV_X1 U6028 ( .A(n4883), .ZN(U3135) );
  AOI22_X1 U6029 ( .A1(n6542), .A2(n4893), .B1(n6544), .B2(n4892), .ZN(n4885)
         );
  NAND2_X1 U6030 ( .A1(n4894), .A2(n6543), .ZN(n4884) );
  OAI211_X1 U6031 ( .C1(n5010), .C2(n6547), .A(n4885), .B(n4884), .ZN(n4886)
         );
  AOI21_X1 U6032 ( .B1(n4898), .B2(INSTQUEUE_REG_14__4__SCAN_IN), .A(n4886), 
        .ZN(n4887) );
  INV_X1 U6033 ( .A(n4887), .ZN(U3136) );
  AOI22_X1 U6034 ( .A1(n6532), .A2(n4893), .B1(n6534), .B2(n4892), .ZN(n4889)
         );
  NAND2_X1 U6035 ( .A1(n4894), .A2(n6533), .ZN(n4888) );
  OAI211_X1 U6036 ( .C1(n5010), .C2(n6537), .A(n4889), .B(n4888), .ZN(n4890)
         );
  AOI21_X1 U6037 ( .B1(n4898), .B2(INSTQUEUE_REG_14__2__SCAN_IN), .A(n4890), 
        .ZN(n4891) );
  INV_X1 U6038 ( .A(n4891), .ZN(U3134) );
  AOI22_X1 U6039 ( .A1(n6508), .A2(n4893), .B1(n6583), .B2(n4892), .ZN(n4896)
         );
  NAND2_X1 U6040 ( .A1(n4894), .A2(n6303), .ZN(n4895) );
  OAI211_X1 U6041 ( .C1(n5010), .C2(n6586), .A(n4896), .B(n4895), .ZN(n4897)
         );
  AOI21_X1 U6042 ( .B1(n4898), .B2(INSTQUEUE_REG_14__5__SCAN_IN), .A(n4897), 
        .ZN(n4899) );
  INV_X1 U6043 ( .A(n4899), .ZN(U3137) );
  OR2_X1 U6044 ( .A1(n4901), .A2(n4902), .ZN(n4903) );
  NAND2_X1 U6045 ( .A1(n4900), .A2(n4903), .ZN(n5882) );
  INV_X1 U6046 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4904) );
  OAI222_X1 U6047 ( .A1(n5882), .A2(n5680), .B1(n5679), .B2(n4905), .C1(n5678), 
        .C2(n4904), .ZN(U2884) );
  INV_X1 U6048 ( .A(n4906), .ZN(n4908) );
  NOR2_X1 U6049 ( .A1(n4907), .A2(n4908), .ZN(n4926) );
  AOI21_X1 U6050 ( .B1(n4908), .B2(n4907), .A(n4926), .ZN(n5524) );
  INV_X1 U6051 ( .A(n5524), .ZN(n4935) );
  INV_X1 U6052 ( .A(EAX_REG_5__SCAN_IN), .ZN(n7006) );
  OAI222_X1 U6053 ( .A1(n4935), .A2(n5680), .B1(n5679), .B2(n4909), .C1(n5678), 
        .C2(n7006), .ZN(U2886) );
  NAND2_X1 U6054 ( .A1(n3895), .A2(n4912), .ZN(n5129) );
  INV_X1 U6055 ( .A(n5129), .ZN(n4914) );
  AOI21_X1 U6056 ( .B1(n4915), .B2(n4914), .A(n6549), .ZN(n4919) );
  AOI22_X1 U6057 ( .A1(n4917), .A2(n4919), .B1(n6481), .B2(n6284), .ZN(n4916)
         );
  NAND2_X1 U6058 ( .A1(n6286), .A2(n4916), .ZN(n6554) );
  INV_X1 U6059 ( .A(n4917), .ZN(n4918) );
  OAI22_X1 U6060 ( .A1(n4919), .A2(n4918), .B1(n6326), .B2(n6481), .ZN(n6552)
         );
  AOI22_X1 U6061 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6554), .B1(n6583), 
        .B2(n6552), .ZN(n4922) );
  AOI22_X1 U6062 ( .A1(n6551), .A2(n6303), .B1(n6549), .B2(n6508), .ZN(n4921)
         );
  OAI211_X1 U6063 ( .C1(n6586), .C2(n6557), .A(n4922), .B(n4921), .ZN(U3081)
         );
  AOI22_X1 U6064 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6554), .B1(n6593), 
        .B2(n6552), .ZN(n4924) );
  AOI22_X1 U6065 ( .A1(n6551), .A2(n6311), .B1(n6549), .B2(n6517), .ZN(n4923)
         );
  OAI211_X1 U6066 ( .C1(n6598), .C2(n6557), .A(n4924), .B(n4923), .ZN(U3083)
         );
  OR2_X1 U6067 ( .A1(n4926), .A2(n4925), .ZN(n4928) );
  INV_X1 U6068 ( .A(n4901), .ZN(n4927) );
  NAND2_X1 U6069 ( .A1(n4928), .A2(n4927), .ZN(n5886) );
  AOI22_X1 U6070 ( .A1(n5674), .A2(DATAI_6_), .B1(EAX_REG_6__SCAN_IN), .B2(
        n5673), .ZN(n4929) );
  OAI21_X1 U6071 ( .B1(n5886), .B2(n5680), .A(n4929), .ZN(U2885) );
  AOI21_X1 U6072 ( .B1(n4931), .B2(n4971), .A(n4930), .ZN(n6455) );
  INV_X1 U6073 ( .A(n6455), .ZN(n5508) );
  INV_X1 U6074 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4932) );
  OAI222_X1 U6075 ( .A1(n5508), .A2(n5620), .B1(n4932), .B2(n5618), .C1(n5882), 
        .C2(n5623), .ZN(U2852) );
  AOI21_X1 U6076 ( .B1(n4934), .B2(n4750), .A(n4972), .ZN(n5533) );
  INV_X1 U6077 ( .A(n5533), .ZN(n4937) );
  INV_X1 U6078 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4936) );
  OAI222_X1 U6079 ( .A1(n4937), .A2(n5620), .B1(n5618), .B2(n4936), .C1(n5623), 
        .C2(n4935), .ZN(U2854) );
  INV_X1 U6080 ( .A(n5584), .ZN(n4941) );
  INV_X1 U6081 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n7029) );
  AOI21_X1 U6082 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4938), 
        .ZN(n4939) );
  OAI21_X1 U6083 ( .B1(n6436), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4939), 
        .ZN(n4940) );
  AOI21_X1 U6084 ( .B1(n4941), .B2(n6431), .A(n4940), .ZN(n4942) );
  OAI21_X1 U6085 ( .B1(n5892), .B2(n4943), .A(n4942), .ZN(U2985) );
  INV_X1 U6086 ( .A(n5564), .ZN(n4947) );
  AOI21_X1 U6087 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4944), 
        .ZN(n4945) );
  OAI21_X1 U6088 ( .B1(n6436), .B2(n5559), .A(n4945), .ZN(n4946) );
  AOI21_X1 U6089 ( .B1(n4947), .B2(n6431), .A(n4946), .ZN(n4948) );
  OAI21_X1 U6090 ( .B1(n4949), .B2(n5892), .A(n4948), .ZN(U2983) );
  XNOR2_X1 U6091 ( .A(n4950), .B(n4951), .ZN(n4963) );
  AND2_X1 U6092 ( .A1(n5868), .A2(REIP_REG_5__SCAN_IN), .ZN(n4960) );
  AOI21_X1 U6093 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4960), 
        .ZN(n4952) );
  OAI21_X1 U6094 ( .B1(n6436), .B2(n5536), .A(n4952), .ZN(n4953) );
  AOI21_X1 U6095 ( .B1(n5524), .B2(n6431), .A(n4953), .ZN(n4954) );
  OAI21_X1 U6096 ( .B1(n5892), .B2(n4963), .A(n4954), .ZN(U2981) );
  AND2_X1 U6097 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6077), .ZN(n4955)
         );
  OAI21_X1 U6098 ( .B1(n6074), .B2(n4955), .A(n6466), .ZN(n5124) );
  INV_X1 U6099 ( .A(n4956), .ZN(n4958) );
  INV_X1 U6100 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6974) );
  OAI211_X1 U6101 ( .C1(n4958), .C2(n6469), .A(n4957), .B(n6974), .ZN(n4959)
         );
  NAND2_X1 U6102 ( .A1(n5124), .A2(n4959), .ZN(n4962) );
  AOI21_X1 U6103 ( .B1(n6463), .B2(n5533), .A(n4960), .ZN(n4961) );
  OAI211_X1 U6104 ( .C1(n4963), .C2(n6084), .A(n4962), .B(n4961), .ZN(U3013)
         );
  NAND2_X1 U6105 ( .A1(n4900), .A2(n4965), .ZN(n4966) );
  NAND2_X1 U6106 ( .A1(n4964), .A2(n4966), .ZN(n5870) );
  OR2_X1 U6107 ( .A1(n4967), .A2(n4930), .ZN(n4968) );
  NAND2_X1 U6108 ( .A1(n4968), .A2(n5483), .ZN(n6087) );
  INV_X1 U6109 ( .A(n6087), .ZN(n4969) );
  AOI22_X1 U6110 ( .A1(n4402), .A2(n4969), .B1(n5621), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4970) );
  OAI21_X1 U6111 ( .B1(n5870), .B2(n5623), .A(n4970), .ZN(U2851) );
  OAI21_X1 U6112 ( .B1(n4973), .B2(n4972), .A(n4971), .ZN(n5518) );
  INV_X1 U6113 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4974) );
  OAI222_X1 U6114 ( .A1(n5518), .A2(n5620), .B1(n4974), .B2(n5618), .C1(n5886), 
        .C2(n5623), .ZN(U2853) );
  NAND2_X1 U6115 ( .A1(n4975), .A2(n3892), .ZN(n5073) );
  NAND2_X1 U6116 ( .A1(n6101), .A2(n6097), .ZN(n6198) );
  INV_X1 U6117 ( .A(n6198), .ZN(n5075) );
  NAND2_X1 U6118 ( .A1(n7013), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5126) );
  NOR2_X1 U6119 ( .A1(n6839), .A2(n5126), .ZN(n5076) );
  AOI21_X1 U6120 ( .B1(n6283), .B2(n5075), .A(n5005), .ZN(n4979) );
  NAND2_X1 U6121 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4976) );
  OAI22_X1 U6122 ( .A1(n4979), .A2(n6284), .B1(n4976), .B2(n5126), .ZN(n4977)
         );
  NAND2_X1 U6123 ( .A1(n4979), .A2(n4978), .ZN(n4982) );
  INV_X1 U6124 ( .A(n5076), .ZN(n4980) );
  NAND2_X1 U6125 ( .A1(n6284), .A2(n4980), .ZN(n4981) );
  OAI211_X1 U6126 ( .C1(n6284), .C2(n4982), .A(n6286), .B(n4981), .ZN(n5004)
         );
  AOI22_X1 U6127 ( .A1(n6524), .A2(n5005), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n5004), .ZN(n4983) );
  OAI21_X1 U6128 ( .B1(n5007), .B2(n6330), .A(n4983), .ZN(n4984) );
  AOI21_X1 U6129 ( .B1(n6491), .B2(n5115), .A(n4984), .ZN(n4985) );
  OAI21_X1 U6130 ( .B1(n6560), .B2(n5010), .A(n4985), .ZN(U3124) );
  AOI22_X1 U6131 ( .A1(n6517), .A2(n5005), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n5004), .ZN(n4986) );
  OAI21_X1 U6132 ( .B1(n5007), .B2(n6361), .A(n4986), .ZN(n4987) );
  AOI21_X1 U6133 ( .B1(n6520), .B2(n5115), .A(n4987), .ZN(n4988) );
  OAI21_X1 U6134 ( .B1(n6589), .B2(n5010), .A(n4988), .ZN(U3131) );
  INV_X1 U6135 ( .A(n6572), .ZN(n6494) );
  AOI22_X1 U6136 ( .A1(n6528), .A2(n5005), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n5004), .ZN(n4989) );
  OAI21_X1 U6137 ( .B1(n5007), .B2(n6334), .A(n4989), .ZN(n4990) );
  AOI21_X1 U6138 ( .B1(n6494), .B2(n5115), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6139 ( .B1(n6567), .B2(n5010), .A(n4991), .ZN(U3125) );
  INV_X1 U6140 ( .A(n6586), .ZN(n6509) );
  AOI22_X1 U6141 ( .A1(n6508), .A2(n5005), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n5004), .ZN(n4992) );
  OAI21_X1 U6142 ( .B1(n5007), .B2(n6350), .A(n4992), .ZN(n4993) );
  AOI21_X1 U6143 ( .B1(n6509), .B2(n5115), .A(n4993), .ZN(n4994) );
  OAI21_X1 U6144 ( .B1(n6581), .B2(n5010), .A(n4994), .ZN(U3129) );
  AOI22_X1 U6145 ( .A1(n6538), .A2(n5005), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n5004), .ZN(n4995) );
  OAI21_X1 U6146 ( .B1(n5007), .B2(n6342), .A(n4995), .ZN(n4996) );
  AOI21_X1 U6147 ( .B1(n6501), .B2(n5115), .A(n4996), .ZN(n4997) );
  OAI21_X1 U6148 ( .B1(n6574), .B2(n5010), .A(n4997), .ZN(U3127) );
  INV_X1 U6149 ( .A(n6537), .ZN(n6497) );
  AOI22_X1 U6150 ( .A1(n6532), .A2(n5005), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n5004), .ZN(n4998) );
  OAI21_X1 U6151 ( .B1(n5007), .B2(n6338), .A(n4998), .ZN(n4999) );
  AOI21_X1 U6152 ( .B1(n6497), .B2(n5115), .A(n4999), .ZN(n5000) );
  OAI21_X1 U6153 ( .B1(n6500), .B2(n5010), .A(n5000), .ZN(U3126) );
  INV_X1 U6154 ( .A(n6547), .ZN(n6504) );
  AOI22_X1 U6155 ( .A1(n6542), .A2(n5005), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n5004), .ZN(n5001) );
  OAI21_X1 U6156 ( .B1(n5007), .B2(n6346), .A(n5001), .ZN(n5002) );
  AOI21_X1 U6157 ( .B1(n6504), .B2(n5115), .A(n5002), .ZN(n5003) );
  OAI21_X1 U6158 ( .B1(n6507), .B2(n5010), .A(n5003), .ZN(U3128) );
  INV_X1 U6159 ( .A(n6558), .ZN(n6512) );
  AOI22_X1 U6160 ( .A1(n6548), .A2(n5005), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n5004), .ZN(n5006) );
  OAI21_X1 U6161 ( .B1(n5007), .B2(n6354), .A(n5006), .ZN(n5008) );
  AOI21_X1 U6162 ( .B1(n6512), .B2(n5115), .A(n5008), .ZN(n5009) );
  OAI21_X1 U6163 ( .B1(n6515), .B2(n5010), .A(n5009), .ZN(U3130) );
  INV_X1 U6164 ( .A(DATAI_8_), .ZN(n6978) );
  INV_X1 U6165 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5011) );
  OAI222_X1 U6166 ( .A1(n5870), .A2(n5680), .B1(n5679), .B2(n6978), .C1(n5678), 
        .C2(n5011), .ZN(U2883) );
  NOR3_X1 U6167 ( .A1(n5012), .A2(n6099), .A3(n6095), .ZN(n5013) );
  NOR2_X1 U6168 ( .A1(n5013), .A2(n6284), .ZN(n5021) );
  NAND2_X1 U6169 ( .A1(n6207), .A2(n3275), .ZN(n6167) );
  INV_X1 U6170 ( .A(n5014), .ZN(n5015) );
  NAND2_X1 U6171 ( .A1(n5015), .A2(n6839), .ZN(n5045) );
  OAI21_X1 U6172 ( .B1(n6167), .B2(n5016), .A(n5045), .ZN(n5023) );
  NAND3_X1 U6173 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6839), .A3(n6610), .ZN(n6162) );
  INV_X1 U6174 ( .A(n6162), .ZN(n5017) );
  NAND3_X1 U6175 ( .A1(n5051), .A2(n3892), .A3(n6238), .ZN(n5018) );
  NAND3_X1 U6176 ( .A1(n5051), .A2(n6238), .A3(n6291), .ZN(n5019) );
  OAI22_X1 U6177 ( .A1(n6206), .A2(n6515), .B1(n6271), .B2(n5045), .ZN(n5020)
         );
  AOI21_X1 U6178 ( .B1(n6512), .B2(n3272), .A(n5020), .ZN(n5026) );
  INV_X1 U6179 ( .A(n5021), .ZN(n5024) );
  AOI21_X1 U6180 ( .B1(n6284), .B2(n6162), .A(n5133), .ZN(n5022) );
  NAND2_X1 U6181 ( .A1(n5047), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5025) );
  OAI211_X1 U6182 ( .C1(n5050), .C2(n6354), .A(n5026), .B(n5025), .ZN(U3050)
         );
  OAI22_X1 U6183 ( .A1(n6206), .A2(n6589), .B1(n6588), .B2(n5045), .ZN(n5027)
         );
  AOI21_X1 U6184 ( .B1(n6520), .B2(n3272), .A(n5027), .ZN(n5029) );
  NAND2_X1 U6185 ( .A1(n5047), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5028) );
  OAI211_X1 U6186 ( .C1(n5050), .C2(n6361), .A(n5029), .B(n5028), .ZN(U3051)
         );
  OAI22_X1 U6187 ( .A1(n6206), .A2(n6500), .B1(n6257), .B2(n5045), .ZN(n5030)
         );
  AOI21_X1 U6188 ( .B1(n6497), .B2(n3272), .A(n5030), .ZN(n5032) );
  NAND2_X1 U6189 ( .A1(n5047), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5031) );
  OAI211_X1 U6190 ( .C1(n5050), .C2(n6338), .A(n5032), .B(n5031), .ZN(U3046)
         );
  OAI22_X1 U6191 ( .A1(n6206), .A2(n6574), .B1(n6573), .B2(n5045), .ZN(n5033)
         );
  AOI21_X1 U6192 ( .B1(n6501), .B2(n3272), .A(n5033), .ZN(n5035) );
  NAND2_X1 U6193 ( .A1(n5047), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5034) );
  OAI211_X1 U6194 ( .C1(n5050), .C2(n6342), .A(n5035), .B(n5034), .ZN(U3047)
         );
  OAI22_X1 U6195 ( .A1(n6206), .A2(n6581), .B1(n6580), .B2(n5045), .ZN(n5036)
         );
  AOI21_X1 U6196 ( .B1(n6509), .B2(n3272), .A(n5036), .ZN(n5038) );
  NAND2_X1 U6197 ( .A1(n5047), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5037) );
  OAI211_X1 U6198 ( .C1(n5050), .C2(n6350), .A(n5038), .B(n5037), .ZN(U3049)
         );
  OAI22_X1 U6199 ( .A1(n6206), .A2(n6507), .B1(n6264), .B2(n5045), .ZN(n5039)
         );
  AOI21_X1 U6200 ( .B1(n6504), .B2(n3272), .A(n5039), .ZN(n5041) );
  NAND2_X1 U6201 ( .A1(n5047), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5040) );
  OAI211_X1 U6202 ( .C1(n5050), .C2(n6346), .A(n5041), .B(n5040), .ZN(U3048)
         );
  OAI22_X1 U6203 ( .A1(n6206), .A2(n6567), .B1(n6566), .B2(n5045), .ZN(n5042)
         );
  AOI21_X1 U6204 ( .B1(n6494), .B2(n3272), .A(n5042), .ZN(n5044) );
  NAND2_X1 U6205 ( .A1(n5047), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5043) );
  OAI211_X1 U6206 ( .C1(n5050), .C2(n6334), .A(n5044), .B(n5043), .ZN(U3045)
         );
  OAI22_X1 U6207 ( .A1(n6206), .A2(n6560), .B1(n6559), .B2(n5045), .ZN(n5046)
         );
  AOI21_X1 U6208 ( .B1(n6491), .B2(n3272), .A(n5046), .ZN(n5049) );
  NAND2_X1 U6209 ( .A1(n5047), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5048) );
  OAI211_X1 U6210 ( .C1(n5050), .C2(n6330), .A(n5049), .B(n5048), .ZN(U3044)
         );
  NAND2_X1 U6211 ( .A1(n5051), .A2(n5127), .ZN(n5052) );
  OR2_X1 U6212 ( .A1(n6101), .A2(n4703), .ZN(n6243) );
  NOR2_X1 U6213 ( .A1(n3087), .A2(n6243), .ZN(n6117) );
  NAND3_X1 U6214 ( .A1(n6839), .A2(n6610), .A3(n7013), .ZN(n6110) );
  NOR2_X1 U6215 ( .A1(n6281), .A2(n6110), .ZN(n6158) );
  AOI21_X1 U6216 ( .B1(n6117), .B2(n3895), .A(n6158), .ZN(n5057) );
  AOI21_X1 U6217 ( .B1(n5053), .B2(STATEBS16_REG_SCAN_IN), .A(n6284), .ZN(
        n5055) );
  AOI22_X1 U6218 ( .A1(n5057), .A2(n5055), .B1(n6284), .B2(n6110), .ZN(n5054)
         );
  NAND2_X1 U6219 ( .A1(n6286), .A2(n5054), .ZN(n6157) );
  INV_X1 U6220 ( .A(n5055), .ZN(n5056) );
  OAI22_X1 U6221 ( .A1(n5057), .A2(n5056), .B1(n6326), .B2(n6110), .ZN(n6156)
         );
  AOI22_X1 U6222 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6157), .B1(n6583), 
        .B2(n6156), .ZN(n5060) );
  AOI22_X1 U6223 ( .A1(n6159), .A2(n6509), .B1(n6508), .B2(n6158), .ZN(n5059)
         );
  OAI211_X1 U6224 ( .C1(n6581), .C2(n6197), .A(n5060), .B(n5059), .ZN(U3033)
         );
  AOI22_X1 U6225 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6157), .B1(n6553), 
        .B2(n6156), .ZN(n5062) );
  AOI22_X1 U6226 ( .A1(n6159), .A2(n6512), .B1(n6548), .B2(n6158), .ZN(n5061)
         );
  OAI211_X1 U6227 ( .C1(n6515), .C2(n6197), .A(n5062), .B(n5061), .ZN(U3034)
         );
  AOI22_X1 U6228 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6157), .B1(n6569), 
        .B2(n6156), .ZN(n5064) );
  AOI22_X1 U6229 ( .A1(n6159), .A2(n6494), .B1(n6528), .B2(n6158), .ZN(n5063)
         );
  OAI211_X1 U6230 ( .C1(n6567), .C2(n6197), .A(n5064), .B(n5063), .ZN(U3029)
         );
  AOI22_X1 U6231 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6157), .B1(n6534), 
        .B2(n6156), .ZN(n5066) );
  AOI22_X1 U6232 ( .A1(n6159), .A2(n6497), .B1(n6532), .B2(n6158), .ZN(n5065)
         );
  OAI211_X1 U6233 ( .C1(n6500), .C2(n6197), .A(n5066), .B(n5065), .ZN(U3030)
         );
  AOI22_X1 U6234 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6157), .B1(n6593), 
        .B2(n6156), .ZN(n5068) );
  AOI22_X1 U6235 ( .A1(n6159), .A2(n6520), .B1(n6517), .B2(n6158), .ZN(n5067)
         );
  OAI211_X1 U6236 ( .C1(n6589), .C2(n6197), .A(n5068), .B(n5067), .ZN(U3035)
         );
  AOI22_X1 U6237 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6157), .B1(n6544), 
        .B2(n6156), .ZN(n5070) );
  AOI22_X1 U6238 ( .A1(n6159), .A2(n6504), .B1(n6542), .B2(n6158), .ZN(n5069)
         );
  OAI211_X1 U6239 ( .C1(n6507), .C2(n6197), .A(n5070), .B(n5069), .ZN(U3032)
         );
  AOI22_X1 U6240 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6157), .B1(n6576), 
        .B2(n6156), .ZN(n5072) );
  AOI22_X1 U6241 ( .A1(n6159), .A2(n6501), .B1(n6538), .B2(n6158), .ZN(n5071)
         );
  OAI211_X1 U6242 ( .C1(n6574), .C2(n6197), .A(n5072), .B(n5071), .ZN(U3031)
         );
  AOI21_X1 U6243 ( .B1(n6590), .B2(n5073), .A(n6643), .ZN(n5074) );
  AOI211_X1 U6244 ( .C1(n5075), .C2(n6199), .A(n6284), .B(n5074), .ZN(n5079)
         );
  AND2_X1 U6245 ( .A1(n6281), .A2(n5076), .ZN(n5112) );
  INV_X1 U6246 ( .A(n6487), .ZN(n6317) );
  OR2_X1 U6247 ( .A1(n6477), .A2(n6111), .ZN(n5080) );
  AOI21_X1 U6248 ( .B1(n5080), .B2(STATE2_REG_2__SCAN_IN), .A(n5077), .ZN(
        n6240) );
  OAI211_X1 U6249 ( .C1(n6725), .C2(n5112), .A(n6317), .B(n6240), .ZN(n5078)
         );
  INV_X1 U6250 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5086) );
  NOR2_X1 U6251 ( .A1(n6198), .A2(n6284), .ZN(n6208) );
  NAND2_X1 U6252 ( .A1(n6208), .A2(n3087), .ZN(n5082) );
  INV_X1 U6253 ( .A(n5080), .ZN(n6249) );
  NAND2_X1 U6254 ( .A1(n6478), .A2(n6249), .ZN(n5081) );
  NAND2_X1 U6255 ( .A1(n5082), .A2(n5081), .ZN(n5111) );
  AOI22_X1 U6256 ( .A1(n6532), .A2(n5112), .B1(n6534), .B2(n5111), .ZN(n5083)
         );
  OAI21_X1 U6257 ( .B1(n6590), .B2(n6537), .A(n5083), .ZN(n5084) );
  AOI21_X1 U6258 ( .B1(n6533), .B2(n5115), .A(n5084), .ZN(n5085) );
  OAI21_X1 U6259 ( .B1(n5118), .B2(n5086), .A(n5085), .ZN(U3118) );
  INV_X1 U6260 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5090) );
  AOI22_X1 U6261 ( .A1(n6538), .A2(n5112), .B1(n6576), .B2(n5111), .ZN(n5087)
         );
  OAI21_X1 U6262 ( .B1(n6590), .B2(n6579), .A(n5087), .ZN(n5088) );
  AOI21_X1 U6263 ( .B1(n6539), .B2(n5115), .A(n5088), .ZN(n5089) );
  OAI21_X1 U6264 ( .B1(n5118), .B2(n5090), .A(n5089), .ZN(U3119) );
  INV_X1 U6265 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5094) );
  AOI22_X1 U6266 ( .A1(n6508), .A2(n5112), .B1(n6583), .B2(n5111), .ZN(n5091)
         );
  OAI21_X1 U6267 ( .B1(n6590), .B2(n6586), .A(n5091), .ZN(n5092) );
  AOI21_X1 U6268 ( .B1(n6303), .B2(n5115), .A(n5092), .ZN(n5093) );
  OAI21_X1 U6269 ( .B1(n5118), .B2(n5094), .A(n5093), .ZN(U3121) );
  INV_X1 U6270 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5098) );
  AOI22_X1 U6271 ( .A1(n6548), .A2(n5112), .B1(n6553), .B2(n5111), .ZN(n5095)
         );
  OAI21_X1 U6272 ( .B1(n6590), .B2(n6558), .A(n5095), .ZN(n5096) );
  AOI21_X1 U6273 ( .B1(n6550), .B2(n5115), .A(n5096), .ZN(n5097) );
  OAI21_X1 U6274 ( .B1(n5118), .B2(n5098), .A(n5097), .ZN(U3122) );
  INV_X1 U6275 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5102) );
  AOI22_X1 U6276 ( .A1(n6517), .A2(n5112), .B1(n6593), .B2(n5111), .ZN(n5099)
         );
  OAI21_X1 U6277 ( .B1(n6590), .B2(n6598), .A(n5099), .ZN(n5100) );
  AOI21_X1 U6278 ( .B1(n6311), .B2(n5115), .A(n5100), .ZN(n5101) );
  OAI21_X1 U6279 ( .B1(n5118), .B2(n5102), .A(n5101), .ZN(U3123) );
  INV_X1 U6280 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5106) );
  AOI22_X1 U6281 ( .A1(n6524), .A2(n5112), .B1(n6562), .B2(n5111), .ZN(n5103)
         );
  OAI21_X1 U6282 ( .B1(n6590), .B2(n6565), .A(n5103), .ZN(n5104) );
  AOI21_X1 U6283 ( .B1(n6525), .B2(n5115), .A(n5104), .ZN(n5105) );
  OAI21_X1 U6284 ( .B1(n5118), .B2(n5106), .A(n5105), .ZN(U3116) );
  INV_X1 U6285 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5110) );
  AOI22_X1 U6286 ( .A1(n6528), .A2(n5112), .B1(n6569), .B2(n5111), .ZN(n5107)
         );
  OAI21_X1 U6287 ( .B1(n6590), .B2(n6572), .A(n5107), .ZN(n5108) );
  AOI21_X1 U6288 ( .B1(n6529), .B2(n5115), .A(n5108), .ZN(n5109) );
  OAI21_X1 U6289 ( .B1(n5118), .B2(n5110), .A(n5109), .ZN(U3117) );
  INV_X1 U6290 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5117) );
  AOI22_X1 U6291 ( .A1(n6542), .A2(n5112), .B1(n6544), .B2(n5111), .ZN(n5113)
         );
  OAI21_X1 U6292 ( .B1(n6590), .B2(n6547), .A(n5113), .ZN(n5114) );
  AOI21_X1 U6293 ( .B1(n6543), .B2(n5115), .A(n5114), .ZN(n5116) );
  OAI21_X1 U6294 ( .B1(n5118), .B2(n5117), .A(n5116), .ZN(U3120) );
  XNOR2_X1 U6295 ( .A(n5119), .B(n5120), .ZN(n5891) );
  NAND2_X1 U6296 ( .A1(n5868), .A2(REIP_REG_6__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U6297 ( .B1(n6088), .B2(n5518), .A(n5883), .ZN(n5123) );
  NAND3_X1 U6298 ( .A1(n6077), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6076), 
        .ZN(n5121) );
  NOR2_X1 U6299 ( .A1(n5121), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5122)
         );
  AOI211_X1 U6300 ( .C1(n5124), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5123), 
        .B(n5122), .ZN(n5125) );
  OAI21_X1 U6301 ( .B1(n6084), .B2(n5891), .A(n5125), .ZN(U3012) );
  OR2_X1 U6302 ( .A1(n5126), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6201)
         );
  NAND2_X1 U6303 ( .A1(n5128), .A2(n5127), .ZN(n5136) );
  OR2_X1 U6304 ( .A1(n6198), .A2(n5129), .ZN(n5131) );
  NOR2_X1 U6305 ( .A1(n6281), .A2(n6201), .ZN(n5164) );
  INV_X1 U6306 ( .A(n5164), .ZN(n5130) );
  NAND2_X1 U6307 ( .A1(n5131), .A2(n5130), .ZN(n5134) );
  NOR2_X1 U6308 ( .A1(n6205), .A2(n5134), .ZN(n5132) );
  INV_X1 U6309 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5140) );
  INV_X1 U6310 ( .A(n5134), .ZN(n5135) );
  OAI22_X1 U6311 ( .A1(n6205), .A2(n5135), .B1(n6201), .B2(n6326), .ZN(n5167)
         );
  NOR2_X2 U6312 ( .A1(n5136), .A2(n3892), .ZN(n6519) );
  AOI22_X1 U6313 ( .A1(n6519), .A2(n6550), .B1(n6548), .B2(n5164), .ZN(n5137)
         );
  OAI21_X1 U6314 ( .B1(n6558), .B2(n6237), .A(n5137), .ZN(n5138) );
  AOI21_X1 U6315 ( .B1(n6553), .B2(n5167), .A(n5138), .ZN(n5139) );
  OAI21_X1 U6316 ( .B1(n5170), .B2(n5140), .A(n5139), .ZN(U3066) );
  INV_X1 U6317 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5144) );
  AOI22_X1 U6318 ( .A1(n6519), .A2(n6311), .B1(n6517), .B2(n5164), .ZN(n5141)
         );
  OAI21_X1 U6319 ( .B1(n6598), .B2(n6237), .A(n5141), .ZN(n5142) );
  AOI21_X1 U6320 ( .B1(n6593), .B2(n5167), .A(n5142), .ZN(n5143) );
  OAI21_X1 U6321 ( .B1(n5170), .B2(n5144), .A(n5143), .ZN(U3067) );
  INV_X1 U6322 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5148) );
  AOI22_X1 U6323 ( .A1(n6519), .A2(n6539), .B1(n6538), .B2(n5164), .ZN(n5145)
         );
  OAI21_X1 U6324 ( .B1(n6579), .B2(n6237), .A(n5145), .ZN(n5146) );
  AOI21_X1 U6325 ( .B1(n6576), .B2(n5167), .A(n5146), .ZN(n5147) );
  OAI21_X1 U6326 ( .B1(n5170), .B2(n5148), .A(n5147), .ZN(U3063) );
  AOI22_X1 U6327 ( .A1(n6519), .A2(n6303), .B1(n6508), .B2(n5164), .ZN(n5149)
         );
  OAI21_X1 U6328 ( .B1(n6586), .B2(n6237), .A(n5149), .ZN(n5150) );
  AOI21_X1 U6329 ( .B1(n6583), .B2(n5167), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6330 ( .B1(n5170), .B2(n6888), .A(n5151), .ZN(U3065) );
  INV_X1 U6331 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5155) );
  AOI22_X1 U6332 ( .A1(n6519), .A2(n6529), .B1(n6528), .B2(n5164), .ZN(n5152)
         );
  OAI21_X1 U6333 ( .B1(n6572), .B2(n6237), .A(n5152), .ZN(n5153) );
  AOI21_X1 U6334 ( .B1(n6569), .B2(n5167), .A(n5153), .ZN(n5154) );
  OAI21_X1 U6335 ( .B1(n5170), .B2(n5155), .A(n5154), .ZN(U3061) );
  INV_X1 U6336 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5159) );
  AOI22_X1 U6337 ( .A1(n6519), .A2(n6525), .B1(n6524), .B2(n5164), .ZN(n5156)
         );
  OAI21_X1 U6338 ( .B1(n6565), .B2(n6237), .A(n5156), .ZN(n5157) );
  AOI21_X1 U6339 ( .B1(n6562), .B2(n5167), .A(n5157), .ZN(n5158) );
  OAI21_X1 U6340 ( .B1(n5170), .B2(n5159), .A(n5158), .ZN(U3060) );
  INV_X1 U6341 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5163) );
  AOI22_X1 U6342 ( .A1(n6519), .A2(n6543), .B1(n6542), .B2(n5164), .ZN(n5160)
         );
  OAI21_X1 U6343 ( .B1(n6547), .B2(n6237), .A(n5160), .ZN(n5161) );
  AOI21_X1 U6344 ( .B1(n6544), .B2(n5167), .A(n5161), .ZN(n5162) );
  OAI21_X1 U6345 ( .B1(n5170), .B2(n5163), .A(n5162), .ZN(U3064) );
  INV_X1 U6346 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5169) );
  AOI22_X1 U6347 ( .A1(n6519), .A2(n6533), .B1(n6532), .B2(n5164), .ZN(n5165)
         );
  OAI21_X1 U6348 ( .B1(n6537), .B2(n6237), .A(n5165), .ZN(n5166) );
  AOI21_X1 U6349 ( .B1(n6534), .B2(n5167), .A(n5166), .ZN(n5168) );
  OAI21_X1 U6350 ( .B1(n5170), .B2(n5169), .A(n5168), .ZN(U3062) );
  INV_X1 U6351 ( .A(n5553), .ZN(n5175) );
  INV_X1 U6352 ( .A(n5171), .ZN(n5172) );
  AOI21_X1 U6353 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5172), 
        .ZN(n5173) );
  OAI21_X1 U6354 ( .B1(n6436), .B2(n5537), .A(n5173), .ZN(n5174) );
  AOI21_X1 U6355 ( .B1(n5175), .B2(n6431), .A(n5174), .ZN(n5176) );
  OAI21_X1 U6356 ( .B1(n5177), .B2(n5892), .A(n5176), .ZN(U2982) );
  NAND2_X1 U6357 ( .A1(n6601), .A2(n5190), .ZN(n5182) );
  CLKBUF_X1 U6358 ( .A(n5178), .Z(n5187) );
  INV_X1 U6359 ( .A(n5180), .ZN(n6599) );
  OAI21_X1 U6360 ( .B1(n5187), .B2(n5179), .A(n6599), .ZN(n5181) );
  NAND2_X1 U6361 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  AOI21_X1 U6362 ( .B1(n4703), .B2(n6600), .A(n5183), .ZN(n6602) );
  AOI22_X1 U6363 ( .A1(n6728), .A2(n5179), .B1(n5185), .B2(n5184), .ZN(n5186)
         );
  OAI21_X1 U6364 ( .B1(n6602), .B2(n6734), .A(n5186), .ZN(n5188) );
  AOI22_X1 U6365 ( .A1(n6732), .A2(n5188), .B1(n5187), .B2(n6728), .ZN(n5189)
         );
  OAI21_X1 U6366 ( .B1(n6732), .B2(n5190), .A(n5189), .ZN(U3460) );
  NAND2_X1 U6367 ( .A1(n5213), .A2(n5192), .ZN(n5194) );
  AOI22_X1 U6368 ( .A1(n5660), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5673), .ZN(n5193) );
  NAND2_X1 U6369 ( .A1(n5194), .A2(n5193), .ZN(U2860) );
  AOI22_X1 U6370 ( .A1(n5660), .A2(DATAI_30_), .B1(n5673), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6371 ( .A1(n5661), .A2(DATAI_14_), .ZN(n5195) );
  OAI211_X1 U6372 ( .C1(n5197), .C2(n5680), .A(n5196), .B(n5195), .ZN(U2861)
         );
  INV_X1 U6373 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6803) );
  NAND2_X1 U6374 ( .A1(n6370), .A2(n6803), .ZN(n5200) );
  NAND2_X1 U6375 ( .A1(n5198), .A2(n5214), .ZN(n5199) );
  MUX2_X1 U6376 ( .A(n5200), .B(n5199), .S(n5210), .Z(U3474) );
  AOI21_X1 U6377 ( .B1(n5202), .B2(STATEBS16_REG_SCAN_IN), .A(n5201), .ZN(
        n5205) );
  OAI211_X1 U6378 ( .C1(n5203), .C2(n3780), .A(STATE2_REG_2__SCAN_IN), .B(
        n4465), .ZN(n5204) );
  OAI21_X1 U6379 ( .B1(n5205), .B2(n5204), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n5206) );
  NAND2_X1 U6380 ( .A1(n5206), .A2(n6650), .ZN(n5212) );
  OAI211_X1 U6381 ( .C1(READY_N), .C2(n5208), .A(n5207), .B(n6284), .ZN(n5209)
         );
  NOR2_X1 U6382 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  MUX2_X1 U6383 ( .A(n5212), .B(REQUESTPENDING_REG_SCAN_IN), .S(n5211), .Z(
        U3472) );
  INV_X1 U6384 ( .A(n5213), .ZN(n5229) );
  AOI22_X1 U6385 ( .A1(n5215), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5214), .ZN(n5222) );
  INV_X1 U6386 ( .A(n5216), .ZN(n5218) );
  OAI22_X1 U6387 ( .A1(n5218), .A2(n5354), .B1(EBX_REG_29__SCAN_IN), .B2(n5217), .ZN(n5233) );
  NAND2_X1 U6388 ( .A1(n5233), .A2(n5219), .ZN(n5220) );
  NOR2_X1 U6389 ( .A1(n5223), .A2(REIP_REG_30__SCAN_IN), .ZN(n5224) );
  NAND3_X1 U6390 ( .A1(n5545), .A2(EBX_REG_31__SCAN_IN), .A3(n5226), .ZN(n5227) );
  INV_X1 U6391 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6717) );
  INV_X1 U6392 ( .A(n5697), .ZN(n5626) );
  INV_X1 U6393 ( .A(n5695), .ZN(n5236) );
  XNOR2_X1 U6394 ( .A(n4448), .B(n5233), .ZN(n5909) );
  AOI22_X1 U6395 ( .A1(n6394), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6390), .ZN(n5234) );
  OAI21_X1 U6396 ( .B1(n5909), .B2(n5517), .A(n5234), .ZN(n5235) );
  AOI21_X1 U6397 ( .B1(n6396), .B2(n5236), .A(n5235), .ZN(n5239) );
  MUX2_X1 U6398 ( .A(n5237), .B(n5244), .S(REIP_REG_29__SCAN_IN), .Z(n5238) );
  OAI211_X1 U6399 ( .C1(n5626), .C2(n5522), .A(n5239), .B(n5238), .ZN(U2798)
         );
  INV_X1 U6400 ( .A(n5240), .ZN(n5243) );
  AOI22_X1 U6401 ( .A1(n6394), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6390), .ZN(n5241) );
  OAI21_X1 U6402 ( .B1(n5600), .B2(n5517), .A(n5241), .ZN(n5242) );
  AOI21_X1 U6403 ( .B1(n6396), .B2(n5243), .A(n5242), .ZN(n5247) );
  NAND2_X1 U6404 ( .A1(n5259), .A2(REIP_REG_27__SCAN_IN), .ZN(n5245) );
  MUX2_X1 U6405 ( .A(n5245), .B(n5244), .S(REIP_REG_28__SCAN_IN), .Z(n5246) );
  OAI211_X1 U6406 ( .C1(n5629), .C2(n5522), .A(n5247), .B(n5246), .ZN(U2799)
         );
  INV_X1 U6407 ( .A(n5248), .ZN(n5251) );
  INV_X1 U6408 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6409 ( .A1(n5706), .A2(n6397), .ZN(n5261) );
  NOR2_X1 U6410 ( .A1(n5271), .A2(n6708), .ZN(n5258) );
  NAND2_X1 U6411 ( .A1(n5252), .A2(n5253), .ZN(n5254) );
  NAND2_X1 U6412 ( .A1(n5255), .A2(n5254), .ZN(n5924) );
  AOI22_X1 U6413 ( .A1(n6394), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6390), .ZN(n5256) );
  OAI21_X1 U6414 ( .B1(n5924), .B2(n5517), .A(n5256), .ZN(n5257) );
  AOI211_X1 U6415 ( .C1(n5259), .C2(n6708), .A(n5258), .B(n5257), .ZN(n5260)
         );
  OAI211_X1 U6416 ( .C1(n5586), .C2(n5704), .A(n5261), .B(n5260), .ZN(U2800)
         );
  AOI21_X1 U6417 ( .B1(n5264), .B2(n5263), .A(n5249), .ZN(n5715) );
  INV_X1 U6418 ( .A(n5715), .ZN(n5635) );
  NAND2_X1 U6419 ( .A1(n5283), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U6420 ( .A1(n5252), .A2(n5267), .ZN(n5934) );
  AOI22_X1 U6421 ( .A1(n6394), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6390), .ZN(n5268) );
  OAI21_X1 U6422 ( .B1(n5934), .B2(n5517), .A(n5268), .ZN(n5274) );
  INV_X1 U6423 ( .A(n5269), .ZN(n5298) );
  AOI21_X1 U6424 ( .B1(n5298), .B2(n5270), .A(REIP_REG_26__SCAN_IN), .ZN(n5272) );
  NOR2_X1 U6425 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  AOI211_X1 U6426 ( .C1(n6396), .C2(n5711), .A(n5274), .B(n5273), .ZN(n5275)
         );
  OAI21_X1 U6427 ( .B1(n5635), .B2(n5522), .A(n5275), .ZN(U2801) );
  OAI21_X1 U6428 ( .B1(n5276), .B2(n5277), .A(n5263), .ZN(n5719) );
  XOR2_X1 U6429 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .Z(n5289) );
  NAND2_X1 U6430 ( .A1(n5316), .A2(n5278), .ZN(n5279) );
  NAND2_X1 U6431 ( .A1(n5501), .A2(n5279), .ZN(n5308) );
  INV_X1 U6432 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U6433 ( .A1(n6394), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6390), .ZN(n5286) );
  NAND2_X1 U6434 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6435 ( .A1(n5283), .A2(n5282), .ZN(n5941) );
  INV_X1 U6436 ( .A(n5941), .ZN(n5284) );
  NAND2_X1 U6437 ( .A1(n6393), .A2(n5284), .ZN(n5285) );
  OAI211_X1 U6438 ( .C1(n5308), .C2(n6936), .A(n5286), .B(n5285), .ZN(n5288)
         );
  NOR2_X1 U6439 ( .A1(n5586), .A2(n5721), .ZN(n5287) );
  AOI211_X1 U6440 ( .C1(n5298), .C2(n5289), .A(n5288), .B(n5287), .ZN(n5290)
         );
  OAI21_X1 U6441 ( .B1(n5719), .B2(n5522), .A(n5290), .ZN(U2802) );
  AND2_X1 U6442 ( .A1(n5291), .A2(n5292), .ZN(n5293) );
  NOR2_X1 U6443 ( .A1(n5276), .A2(n5293), .ZN(n5729) );
  INV_X1 U6444 ( .A(n5729), .ZN(n5640) );
  INV_X1 U6445 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6701) );
  AOI22_X1 U6446 ( .A1(n6394), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6390), .ZN(n5295) );
  NAND2_X1 U6447 ( .A1(n6393), .A2(n5602), .ZN(n5294) );
  OAI211_X1 U6448 ( .C1(n5308), .C2(n6701), .A(n5295), .B(n5294), .ZN(n5297)
         );
  AOI211_X1 U6449 ( .C1(n5298), .C2(n6701), .A(n5297), .B(n5296), .ZN(n5299)
         );
  OAI21_X1 U6450 ( .B1(n5640), .B2(n5522), .A(n5299), .ZN(U2803) );
  INV_X1 U6451 ( .A(n5291), .ZN(n5301) );
  AOI21_X1 U6452 ( .B1(n5302), .B2(n5314), .A(n5301), .ZN(n5739) );
  INV_X1 U6453 ( .A(n5739), .ZN(n5643) );
  INV_X1 U6454 ( .A(n5737), .ZN(n5311) );
  INV_X1 U6455 ( .A(n5330), .ZN(n5304) );
  AOI21_X1 U6456 ( .B1(n5304), .B2(n5303), .A(REIP_REG_23__SCAN_IN), .ZN(n5309) );
  AOI22_X1 U6457 ( .A1(n6394), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6390), .ZN(n5307) );
  AOI21_X1 U6458 ( .B1(n5305), .B2(n3120), .A(n3853), .ZN(n5952) );
  NAND2_X1 U6459 ( .A1(n6393), .A2(n5952), .ZN(n5306) );
  OAI211_X1 U6460 ( .C1(n5309), .C2(n5308), .A(n5307), .B(n5306), .ZN(n5310)
         );
  AOI21_X1 U6461 ( .B1(n5311), .B2(n6396), .A(n5310), .ZN(n5312) );
  OAI21_X1 U6462 ( .B1(n5643), .B2(n5522), .A(n5312), .ZN(U2804) );
  AOI21_X1 U6463 ( .B1(n5315), .B2(n5313), .A(n5300), .ZN(n5750) );
  INV_X1 U6464 ( .A(n5750), .ZN(n5646) );
  XNOR2_X1 U6465 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .ZN(
        n5322) );
  INV_X1 U6466 ( .A(n5501), .ZN(n5591) );
  NOR2_X1 U6467 ( .A1(n5591), .A2(n5316), .ZN(n5340) );
  OAI21_X1 U6468 ( .B1(n5318), .B2(n5317), .A(n3120), .ZN(n5960) );
  AOI22_X1 U6469 ( .A1(n6394), .A2(EBX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6390), .ZN(n5319) );
  OAI21_X1 U6470 ( .B1(n5960), .B2(n5517), .A(n5319), .ZN(n5320) );
  AOI21_X1 U6471 ( .B1(n5340), .B2(REIP_REG_22__SCAN_IN), .A(n5320), .ZN(n5321) );
  OAI21_X1 U6472 ( .B1(n5330), .B2(n5322), .A(n5321), .ZN(n5323) );
  AOI21_X1 U6473 ( .B1(n6396), .B2(n5746), .A(n5323), .ZN(n5324) );
  OAI21_X1 U6474 ( .B1(n5646), .B2(n5522), .A(n5324), .ZN(U2805) );
  OAI21_X1 U6475 ( .B1(n5325), .B2(n5326), .A(n5313), .ZN(n5649) );
  INV_X1 U6476 ( .A(n5649), .ZN(n5758) );
  NAND2_X1 U6477 ( .A1(n5758), .A2(n6397), .ZN(n5334) );
  XNOR2_X1 U6478 ( .A(n5328), .B(n5327), .ZN(n5968) );
  AOI22_X1 U6479 ( .A1(n6394), .A2(EBX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6390), .ZN(n5329) );
  OAI21_X1 U6480 ( .B1(n5517), .B2(n5968), .A(n5329), .ZN(n5332) );
  NOR2_X1 U6481 ( .A1(n5330), .A2(REIP_REG_21__SCAN_IN), .ZN(n5331) );
  AOI211_X1 U6482 ( .C1(n5340), .C2(REIP_REG_21__SCAN_IN), .A(n5332), .B(n5331), .ZN(n5333) );
  OAI211_X1 U6483 ( .C1(n5586), .C2(n5756), .A(n5334), .B(n5333), .ZN(U2806)
         );
  INV_X1 U6484 ( .A(n5335), .ZN(n5336) );
  AOI21_X1 U6485 ( .B1(n5336), .B2(n3103), .A(n5325), .ZN(n5765) );
  INV_X1 U6486 ( .A(n5765), .ZN(n5652) );
  MUX2_X1 U6487 ( .A(n5356), .B(n3791), .S(n5337), .Z(n5339) );
  XNOR2_X1 U6488 ( .A(n5339), .B(n5338), .ZN(n5978) );
  INV_X1 U6489 ( .A(n5978), .ZN(n5606) );
  INV_X1 U6490 ( .A(n5362), .ZN(n5374) );
  INV_X1 U6491 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6694) );
  INV_X1 U6492 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6998) );
  NOR3_X1 U6493 ( .A1(n5374), .A2(n6694), .A3(n6998), .ZN(n5341) );
  OAI21_X1 U6494 ( .B1(n5341), .B2(REIP_REG_20__SCAN_IN), .A(n5340), .ZN(n5343) );
  AOI22_X1 U6495 ( .A1(n6394), .A2(EBX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6390), .ZN(n5342) );
  OAI211_X1 U6496 ( .C1(n5606), .C2(n5517), .A(n5343), .B(n5342), .ZN(n5344)
         );
  AOI21_X1 U6497 ( .B1(n5761), .B2(n6396), .A(n5344), .ZN(n5345) );
  OAI21_X1 U6498 ( .B1(n5652), .B2(n5522), .A(n5345), .ZN(U2807) );
  INV_X1 U6499 ( .A(n5347), .ZN(n5348) );
  XNOR2_X1 U6500 ( .A(n6998), .B(REIP_REG_19__SCAN_IN), .ZN(n5361) );
  INV_X1 U6501 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6502 ( .A1(n5501), .A2(n5350), .ZN(n5379) );
  NAND2_X1 U6503 ( .A1(n5577), .A2(n5351), .ZN(n5540) );
  OAI21_X1 U6504 ( .B1(n5585), .B2(n5769), .A(n5540), .ZN(n5352) );
  AOI21_X1 U6505 ( .B1(n6394), .B2(EBX_REG_19__SCAN_IN), .A(n5352), .ZN(n5359)
         );
  MUX2_X1 U6506 ( .A(n5356), .B(n5355), .S(n5354), .Z(n5369) );
  NOR2_X1 U6507 ( .A1(n5353), .A2(n5369), .ZN(n5368) );
  XNOR2_X1 U6508 ( .A(n5368), .B(n5357), .ZN(n5992) );
  NAND2_X1 U6509 ( .A1(n6393), .A2(n5992), .ZN(n5358) );
  OAI211_X1 U6510 ( .C1(n5379), .C2(n6694), .A(n5359), .B(n5358), .ZN(n5360)
         );
  AOI21_X1 U6511 ( .B1(n5362), .B2(n5361), .A(n5360), .ZN(n5365) );
  INV_X1 U6512 ( .A(n5363), .ZN(n5771) );
  NAND2_X1 U6513 ( .A1(n6396), .A2(n5771), .ZN(n5364) );
  OAI211_X1 U6514 ( .C1(n5774), .C2(n5522), .A(n5365), .B(n5364), .ZN(U2808)
         );
  OAI21_X1 U6515 ( .B1(n3084), .B2(n4135), .A(n5347), .ZN(n5786) );
  AOI21_X1 U6516 ( .B1(n5353), .B2(n5369), .A(n5368), .ZN(n6000) );
  INV_X1 U6517 ( .A(n6394), .ZN(n5493) );
  NAND2_X1 U6518 ( .A1(n6394), .A2(EBX_REG_18__SCAN_IN), .ZN(n5370) );
  OAI211_X1 U6519 ( .C1(n5585), .C2(n5781), .A(n5370), .B(n5540), .ZN(n5372)
         );
  NOR2_X1 U6520 ( .A1(n5379), .A2(n6998), .ZN(n5371) );
  AOI211_X1 U6521 ( .C1(n6000), .C2(n6393), .A(n5372), .B(n5371), .ZN(n5373)
         );
  OAI21_X1 U6522 ( .B1(n5374), .B2(REIP_REG_18__SCAN_IN), .A(n5373), .ZN(n5375) );
  AOI21_X1 U6523 ( .B1(n6396), .B2(n5783), .A(n5375), .ZN(n5376) );
  OAI21_X1 U6524 ( .B1(n5786), .B2(n5522), .A(n5376), .ZN(U2809) );
  OR2_X1 U6525 ( .A1(n3097), .A2(n5377), .ZN(n5378) );
  INV_X1 U6526 ( .A(n5379), .ZN(n5389) );
  INV_X1 U6527 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5380) );
  OAI21_X1 U6528 ( .B1(n5418), .B2(n5395), .A(n5380), .ZN(n5388) );
  AND2_X1 U6529 ( .A1(n5381), .A2(n5397), .ZN(n5383) );
  OAI21_X1 U6530 ( .B1(n5383), .B2(n5382), .A(n5353), .ZN(n6009) );
  OAI21_X1 U6531 ( .B1(n5585), .B2(n6837), .A(n5540), .ZN(n5384) );
  AOI21_X1 U6532 ( .B1(n6394), .B2(EBX_REG_17__SCAN_IN), .A(n5384), .ZN(n5385)
         );
  OAI21_X1 U6533 ( .B1(n5517), .B2(n6009), .A(n5385), .ZN(n5387) );
  NOR2_X1 U6534 ( .A1(n5586), .A2(n5790), .ZN(n5386) );
  AOI211_X1 U6535 ( .C1(n5389), .C2(n5388), .A(n5387), .B(n5386), .ZN(n5390)
         );
  OAI21_X1 U6536 ( .B1(n5659), .B2(n5522), .A(n5390), .ZN(U2810) );
  INV_X1 U6537 ( .A(n5391), .ZN(n5392) );
  NOR2_X1 U6538 ( .A1(n5392), .A2(n5393), .ZN(n5394) );
  INV_X1 U6539 ( .A(n5800), .ZN(n5404) );
  NOR2_X1 U6540 ( .A1(n5591), .A2(n3104), .ZN(n5430) );
  INV_X1 U6541 ( .A(n5430), .ZN(n5402) );
  INV_X1 U6542 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7004) );
  INV_X1 U6543 ( .A(n5418), .ZN(n5396) );
  OAI211_X1 U6544 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n5396), .B(n5395), .ZN(n5401) );
  XOR2_X1 U6545 ( .A(n5397), .B(n5381), .Z(n6017) );
  NAND2_X1 U6546 ( .A1(n6394), .A2(EBX_REG_16__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6547 ( .C1(n5585), .C2(n6814), .A(n5398), .B(n5540), .ZN(n5399)
         );
  AOI21_X1 U6548 ( .B1(n6393), .B2(n6017), .A(n5399), .ZN(n5400) );
  OAI211_X1 U6549 ( .C1(n5402), .C2(n7004), .A(n5401), .B(n5400), .ZN(n5403)
         );
  AOI21_X1 U6550 ( .B1(n6396), .B2(n5404), .A(n5403), .ZN(n5405) );
  OAI21_X1 U6551 ( .B1(n5798), .B2(n5522), .A(n5405), .ZN(U2811) );
  XNOR2_X1 U6552 ( .A(n5407), .B(n5408), .ZN(n5434) );
  AOI22_X1 U6553 ( .A1(n5434), .A2(n5435), .B1(n5406), .B2(n5408), .ZN(n5424)
         );
  INV_X1 U6554 ( .A(n5409), .ZN(n5423) );
  NOR2_X1 U6555 ( .A1(n5424), .A2(n5423), .ZN(n5422) );
  OAI21_X1 U6556 ( .B1(n5422), .B2(n5410), .A(n5391), .ZN(n5813) );
  INV_X1 U6557 ( .A(n5809), .ZN(n5420) );
  AOI21_X1 U6558 ( .B1(n5412), .B2(n5411), .A(n5381), .ZN(n6029) );
  NAND2_X1 U6559 ( .A1(n6394), .A2(EBX_REG_15__SCAN_IN), .ZN(n5413) );
  OAI211_X1 U6560 ( .C1(n5585), .C2(n5414), .A(n5413), .B(n5540), .ZN(n5415)
         );
  AOI21_X1 U6561 ( .B1(n6393), .B2(n6029), .A(n5415), .ZN(n5417) );
  NAND2_X1 U6562 ( .A1(n5430), .A2(REIP_REG_15__SCAN_IN), .ZN(n5416) );
  OAI211_X1 U6563 ( .C1(n5418), .C2(REIP_REG_15__SCAN_IN), .A(n5417), .B(n5416), .ZN(n5419) );
  AOI21_X1 U6564 ( .B1(n6396), .B2(n5420), .A(n5419), .ZN(n5421) );
  OAI21_X1 U6565 ( .B1(n5813), .B2(n5522), .A(n5421), .ZN(U2812) );
  AOI21_X1 U6566 ( .B1(n5424), .B2(n5423), .A(n5422), .ZN(n5819) );
  NAND2_X1 U6567 ( .A1(n5819), .A2(n6397), .ZN(n5433) );
  OAI21_X1 U6568 ( .B1(n5436), .B2(n6688), .A(n6690), .ZN(n5431) );
  OAI21_X1 U6569 ( .B1(n5426), .B2(n5425), .A(n5411), .ZN(n6034) );
  INV_X1 U6570 ( .A(n5540), .ZN(n6389) );
  AOI21_X1 U6571 ( .B1(n6390), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6389), 
        .ZN(n5428) );
  NAND2_X1 U6572 ( .A1(n6394), .A2(EBX_REG_14__SCAN_IN), .ZN(n5427) );
  OAI211_X1 U6573 ( .C1(n5517), .C2(n6034), .A(n5428), .B(n5427), .ZN(n5429)
         );
  AOI21_X1 U6574 ( .B1(n5431), .B2(n5430), .A(n5429), .ZN(n5432) );
  OAI211_X1 U6575 ( .C1(n5586), .C2(n5817), .A(n5433), .B(n5432), .ZN(U2813)
         );
  XOR2_X1 U6576 ( .A(n5435), .B(n5434), .Z(n5827) );
  INV_X1 U6577 ( .A(n5436), .ZN(n5446) );
  NAND2_X1 U6578 ( .A1(n5501), .A2(n5437), .ZN(n5451) );
  AOI21_X1 U6579 ( .B1(n5439), .B2(n5438), .A(n5425), .ZN(n6055) );
  INV_X1 U6580 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6581 ( .A1(n6394), .A2(EBX_REG_13__SCAN_IN), .ZN(n5440) );
  OAI211_X1 U6582 ( .C1(n5585), .C2(n5441), .A(n5440), .B(n5540), .ZN(n5442)
         );
  AOI21_X1 U6583 ( .B1(n6393), .B2(n6055), .A(n5442), .ZN(n5443) );
  OAI21_X1 U6584 ( .B1(n6688), .B2(n5451), .A(n5443), .ZN(n5445) );
  NOR2_X1 U6585 ( .A1(n5586), .A2(n5825), .ZN(n5444) );
  AOI211_X1 U6586 ( .C1(n5446), .C2(n6688), .A(n5445), .B(n5444), .ZN(n5447)
         );
  OAI21_X1 U6587 ( .B1(n5668), .B2(n5522), .A(n5447), .ZN(U2814) );
  AOI21_X1 U6588 ( .B1(n5449), .B2(n5448), .A(n5406), .ZN(n5837) );
  INV_X1 U6589 ( .A(n5837), .ZN(n5670) );
  OAI21_X1 U6590 ( .B1(n5450), .B2(n5469), .A(n5438), .ZN(n6065) );
  INV_X1 U6591 ( .A(n5451), .ZN(n5452) );
  OAI21_X1 U6592 ( .B1(n5453), .B2(REIP_REG_12__SCAN_IN), .A(n5452), .ZN(n5456) );
  OAI21_X1 U6593 ( .B1(n5585), .B2(n6878), .A(n5540), .ZN(n5454) );
  AOI21_X1 U6594 ( .B1(n6394), .B2(EBX_REG_12__SCAN_IN), .A(n5454), .ZN(n5455)
         );
  OAI211_X1 U6595 ( .C1(n6065), .C2(n5517), .A(n5456), .B(n5455), .ZN(n5457)
         );
  AOI21_X1 U6596 ( .B1(n6396), .B2(n5836), .A(n5457), .ZN(n5458) );
  OAI21_X1 U6597 ( .B1(n5670), .B2(n5522), .A(n5458), .ZN(U2815) );
  OR2_X1 U6598 ( .A1(n5460), .A2(n5461), .ZN(n5462) );
  NAND2_X1 U6599 ( .A1(n5448), .A2(n5462), .ZN(n5849) );
  INV_X1 U6600 ( .A(n5849), .ZN(n5463) );
  NAND2_X1 U6601 ( .A1(n5463), .A2(n6397), .ZN(n5478) );
  INV_X1 U6602 ( .A(n6387), .ZN(n5476) );
  NOR2_X1 U6603 ( .A1(n5464), .A2(REIP_REG_11__SCAN_IN), .ZN(n5475) );
  INV_X1 U6604 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5465) );
  OAI21_X1 U6605 ( .B1(n5585), .B2(n5465), .A(n5540), .ZN(n5466) );
  AOI21_X1 U6606 ( .B1(n6394), .B2(EBX_REG_11__SCAN_IN), .A(n5466), .ZN(n5473)
         );
  INV_X1 U6607 ( .A(n5467), .ZN(n5468) );
  NAND3_X1 U6608 ( .A1(n5501), .A2(REIP_REG_11__SCAN_IN), .A3(n5468), .ZN(
        n5472) );
  AOI21_X1 U6609 ( .B1(n5470), .B2(n5615), .A(n5469), .ZN(n6438) );
  NAND2_X1 U6610 ( .A1(n6393), .A2(n6438), .ZN(n5471) );
  NAND3_X1 U6611 ( .A1(n5473), .A2(n5472), .A3(n5471), .ZN(n5474) );
  AOI21_X1 U6612 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5477) );
  OAI211_X1 U6613 ( .C1(n5586), .C2(n5845), .A(n5478), .B(n5477), .ZN(U2816)
         );
  INV_X1 U6614 ( .A(n4964), .ZN(n5480) );
  OAI21_X1 U6615 ( .B1(n5480), .B2(n3124), .A(n5479), .ZN(n5865) );
  INV_X1 U6616 ( .A(n5861), .ZN(n5490) );
  NOR2_X1 U6617 ( .A1(n6387), .A2(REIP_REG_9__SCAN_IN), .ZN(n6401) );
  INV_X1 U6618 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6619 ( .A1(n5501), .A2(n5481), .ZN(n6399) );
  AOI21_X1 U6620 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n6447) );
  NAND2_X1 U6621 ( .A1(n6394), .A2(EBX_REG_9__SCAN_IN), .ZN(n5485) );
  OAI211_X1 U6622 ( .C1(n5585), .C2(n6919), .A(n5485), .B(n5540), .ZN(n5486)
         );
  AOI21_X1 U6623 ( .B1(n6393), .B2(n6447), .A(n5486), .ZN(n5487) );
  OAI21_X1 U6624 ( .B1(n5488), .B2(n6399), .A(n5487), .ZN(n5489) );
  AOI211_X1 U6625 ( .C1(n6396), .C2(n5490), .A(n6401), .B(n5489), .ZN(n5491)
         );
  OAI21_X1 U6626 ( .B1(n5522), .B2(n5865), .A(n5491), .ZN(U2818) );
  NAND3_X1 U6627 ( .A1(n5513), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n5492) );
  INV_X1 U6628 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6683) );
  AOI21_X1 U6629 ( .B1(n5492), .B2(n6683), .A(n6399), .ZN(n5497) );
  INV_X1 U6630 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U6631 ( .A1(n5493), .A2(n6844), .ZN(n5494) );
  AOI211_X1 U6632 ( .C1(n6390), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6389), 
        .B(n5494), .ZN(n5495) );
  OAI21_X1 U6633 ( .B1(n5517), .B2(n6087), .A(n5495), .ZN(n5496) );
  AOI211_X1 U6634 ( .C1(n6396), .C2(n5873), .A(n5497), .B(n5496), .ZN(n5498)
         );
  OAI21_X1 U6635 ( .B1(n5522), .B2(n5870), .A(n5498), .ZN(U2819) );
  INV_X1 U6636 ( .A(n5878), .ZN(n5511) );
  NAND2_X1 U6637 ( .A1(n5577), .A2(n5499), .ZN(n5500) );
  NAND2_X1 U6638 ( .A1(n5501), .A2(n5500), .ZN(n5528) );
  INV_X1 U6639 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U6640 ( .A1(n5528), .A2(n6682), .ZN(n5510) );
  INV_X1 U6641 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5502) );
  OAI22_X1 U6642 ( .A1(n5502), .A2(REIP_REG_7__SCAN_IN), .B1(n6682), .B2(
        REIP_REG_6__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6643 ( .A1(n5513), .A2(n5503), .ZN(n5507) );
  INV_X1 U6644 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5504) );
  OAI21_X1 U6645 ( .B1(n5585), .B2(n5504), .A(n5540), .ZN(n5505) );
  AOI21_X1 U6646 ( .B1(n6394), .B2(EBX_REG_7__SCAN_IN), .A(n5505), .ZN(n5506)
         );
  OAI211_X1 U6647 ( .C1(n5508), .C2(n5517), .A(n5507), .B(n5506), .ZN(n5509)
         );
  AOI211_X1 U6648 ( .C1(n6396), .C2(n5511), .A(n5510), .B(n5509), .ZN(n5512)
         );
  OAI21_X1 U6649 ( .B1(n5522), .B2(n5882), .A(n5512), .ZN(U2820) );
  NOR2_X1 U6650 ( .A1(n5528), .A2(n5502), .ZN(n5520) );
  NAND2_X1 U6651 ( .A1(n5513), .A2(n5502), .ZN(n5516) );
  INV_X1 U6652 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U6653 ( .B1(n5585), .B2(n6899), .A(n5540), .ZN(n5514) );
  AOI21_X1 U6654 ( .B1(n6394), .B2(EBX_REG_6__SCAN_IN), .A(n5514), .ZN(n5515)
         );
  OAI211_X1 U6655 ( .C1(n5518), .C2(n5517), .A(n5516), .B(n5515), .ZN(n5519)
         );
  AOI211_X1 U6656 ( .C1(n6396), .C2(n3269), .A(n5520), .B(n5519), .ZN(n5521)
         );
  OAI21_X1 U6657 ( .B1(n5522), .B2(n5886), .A(n5521), .ZN(U2821) );
  INV_X1 U6658 ( .A(n5596), .ZN(n5525) );
  NAND2_X1 U6659 ( .A1(n5525), .A2(n5524), .ZN(n5535) );
  NAND2_X1 U6660 ( .A1(n6394), .A2(EBX_REG_5__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U6661 ( .C1(n3942), .C2(n5585), .A(n5526), .B(n5540), .ZN(n5532)
         );
  INV_X1 U6662 ( .A(REIP_REG_5__SCAN_IN), .ZN(n5530) );
  INV_X1 U6663 ( .A(n5539), .ZN(n5527) );
  NAND3_X1 U6664 ( .A1(n5565), .A2(REIP_REG_4__SCAN_IN), .A3(n5527), .ZN(n5529) );
  AOI21_X1 U6665 ( .B1(n5530), .B2(n5529), .A(n5528), .ZN(n5531) );
  AOI211_X1 U6666 ( .C1(n5533), .C2(n6393), .A(n5532), .B(n5531), .ZN(n5534)
         );
  OAI211_X1 U6667 ( .C1(n5586), .C2(n5536), .A(n5535), .B(n5534), .ZN(U2822)
         );
  INV_X1 U6668 ( .A(n5537), .ZN(n5551) );
  NAND2_X1 U6669 ( .A1(n5565), .A2(n5539), .ZN(n5558) );
  NAND2_X1 U6670 ( .A1(n5558), .A2(n5577), .ZN(n5562) );
  NAND2_X1 U6671 ( .A1(n5562), .A2(REIP_REG_4__SCAN_IN), .ZN(n5549) );
  AOI22_X1 U6672 ( .A1(n6393), .A2(n5538), .B1(n6394), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5548) );
  NOR2_X1 U6673 ( .A1(n5539), .A2(REIP_REG_4__SCAN_IN), .ZN(n5542) );
  INV_X1 U6674 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6824) );
  OAI21_X1 U6675 ( .B1(n5585), .B2(n6824), .A(n5540), .ZN(n5541) );
  AOI21_X1 U6676 ( .B1(n5565), .B2(n5542), .A(n5541), .ZN(n5547) );
  INV_X1 U6677 ( .A(n5543), .ZN(n5544) );
  AND2_X1 U6678 ( .A1(n5545), .A2(n5544), .ZN(n5587) );
  NAND2_X1 U6679 ( .A1(n5587), .A2(n6365), .ZN(n5546) );
  NAND4_X1 U6680 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n5550)
         );
  AOI21_X1 U6681 ( .B1(n6396), .B2(n5551), .A(n5550), .ZN(n5552) );
  OAI21_X1 U6682 ( .B1(n5596), .B2(n5553), .A(n5552), .ZN(U2823) );
  NAND2_X1 U6683 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5557) );
  AOI22_X1 U6684 ( .A1(n5554), .A2(n6393), .B1(n5587), .B2(n3087), .ZN(n5556)
         );
  AOI22_X1 U6685 ( .A1(n6394), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6390), .ZN(n5555) );
  OAI211_X1 U6686 ( .C1(n5558), .C2(n5557), .A(n5556), .B(n5555), .ZN(n5561)
         );
  NOR2_X1 U6687 ( .A1(n5586), .A2(n5559), .ZN(n5560) );
  AOI211_X1 U6688 ( .C1(REIP_REG_3__SCAN_IN), .C2(n5562), .A(n5561), .B(n5560), 
        .ZN(n5563) );
  OAI21_X1 U6689 ( .B1(n5596), .B2(n5564), .A(n5563), .ZN(U2824) );
  INV_X1 U6690 ( .A(n6435), .ZN(n5574) );
  INV_X1 U6691 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U6692 ( .A1(n5565), .A2(n6944), .ZN(n5579) );
  NAND3_X1 U6693 ( .A1(n5579), .A2(n5577), .A3(REIP_REG_2__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6694 ( .A1(n5565), .A2(REIP_REG_1__SCAN_IN), .ZN(n5567) );
  INV_X1 U6695 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U6696 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND2_X1 U6697 ( .A1(n5569), .A2(n5568), .ZN(n5572) );
  AOI22_X1 U6698 ( .A1(n6462), .A2(n6393), .B1(n5587), .B2(n6101), .ZN(n5571)
         );
  AOI22_X1 U6699 ( .A1(n6394), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6390), .ZN(n5570) );
  NAND3_X1 U6700 ( .A1(n5572), .A2(n5571), .A3(n5570), .ZN(n5573) );
  AOI21_X1 U6701 ( .B1(n6396), .B2(n5574), .A(n5573), .ZN(n5575) );
  OAI21_X1 U6702 ( .B1(n5596), .B2(n6425), .A(n5575), .ZN(U2825) );
  AOI22_X1 U6703 ( .A1(n6394), .A2(EBX_REG_1__SCAN_IN), .B1(n6393), .B2(n5576), 
        .ZN(n5581) );
  INV_X1 U6704 ( .A(n5577), .ZN(n5578) );
  AOI22_X1 U6705 ( .A1(n5587), .A2(n4703), .B1(n5578), .B2(REIP_REG_1__SCAN_IN), .ZN(n5580) );
  AND3_X1 U6706 ( .A1(n5581), .A2(n5580), .A3(n5579), .ZN(n5583) );
  MUX2_X1 U6707 ( .A(n5586), .B(n5585), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n5582) );
  OAI211_X1 U6708 ( .C1(n5596), .C2(n5584), .A(n5583), .B(n5582), .ZN(U2826)
         );
  NAND2_X1 U6709 ( .A1(n5586), .A2(n5585), .ZN(n5593) );
  AOI22_X1 U6710 ( .A1(n3895), .A2(n5587), .B1(n6394), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5590) );
  NAND2_X1 U6711 ( .A1(n6393), .A2(n5588), .ZN(n5589) );
  OAI211_X1 U6712 ( .C1(n5591), .C2(n6740), .A(n5590), .B(n5589), .ZN(n5592)
         );
  AOI21_X1 U6713 ( .B1(n5593), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5592), 
        .ZN(n5594) );
  OAI21_X1 U6714 ( .B1(n5596), .B2(n5595), .A(n5594), .ZN(U2827) );
  INV_X1 U6715 ( .A(n5899), .ZN(n5598) );
  OAI22_X1 U6716 ( .A1(n5598), .A2(n5620), .B1(n5597), .B2(n5618), .ZN(U2828)
         );
  INV_X1 U6717 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5599) );
  OAI222_X1 U6718 ( .A1(n5599), .A2(n5618), .B1(n5620), .B2(n5909), .C1(n5623), 
        .C2(n5626), .ZN(U2830) );
  OAI222_X1 U6719 ( .A1(n5601), .A2(n5618), .B1(n5620), .B2(n5600), .C1(n5629), 
        .C2(n5623), .ZN(U2831) );
  INV_X1 U6720 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6855) );
  INV_X1 U6721 ( .A(n5706), .ZN(n5632) );
  OAI222_X1 U6722 ( .A1(n6855), .A2(n5618), .B1(n5620), .B2(n5924), .C1(n5632), 
        .C2(n5623), .ZN(U2832) );
  OAI222_X1 U6723 ( .A1(n6892), .A2(n5618), .B1(n5620), .B2(n5934), .C1(n5635), 
        .C2(n5623), .ZN(U2833) );
  INV_X1 U6724 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U6725 ( .A1(n5941), .A2(n5620), .B1(n6823), .B2(n5618), .C1(n5719), 
        .C2(n5623), .ZN(U2834) );
  AOI22_X1 U6726 ( .A1(n5602), .A2(n4402), .B1(n5621), .B2(EBX_REG_24__SCAN_IN), .ZN(n5603) );
  OAI21_X1 U6727 ( .B1(n5640), .B2(n5623), .A(n5603), .ZN(U2835) );
  AOI22_X1 U6728 ( .A1(n5952), .A2(n4402), .B1(n5621), .B2(EBX_REG_23__SCAN_IN), .ZN(n5604) );
  OAI21_X1 U6729 ( .B1(n5643), .B2(n5623), .A(n5604), .ZN(U2836) );
  INV_X1 U6730 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6975) );
  OAI222_X1 U6731 ( .A1(n6975), .A2(n5618), .B1(n5620), .B2(n5960), .C1(n5646), 
        .C2(n5623), .ZN(U2837) );
  INV_X1 U6732 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5605) );
  OAI222_X1 U6733 ( .A1(n5605), .A2(n5618), .B1(n5620), .B2(n5968), .C1(n5649), 
        .C2(n5623), .ZN(U2838) );
  OAI222_X1 U6734 ( .A1(n5623), .A2(n5652), .B1(n5618), .B2(n7019), .C1(n5606), 
        .C2(n5620), .ZN(U2839) );
  AOI22_X1 U6735 ( .A1(n4402), .A2(n5992), .B1(n5621), .B2(EBX_REG_19__SCAN_IN), .ZN(n5607) );
  OAI21_X1 U6736 ( .B1(n5774), .B2(n5623), .A(n5607), .ZN(U2840) );
  AOI22_X1 U6737 ( .A1(n4402), .A2(n6000), .B1(n5621), .B2(EBX_REG_18__SCAN_IN), .ZN(n5608) );
  OAI21_X1 U6738 ( .B1(n5786), .B2(n5623), .A(n5608), .ZN(U2841) );
  OAI222_X1 U6739 ( .A1(n7012), .A2(n5618), .B1(n5620), .B2(n6009), .C1(n5659), 
        .C2(n5623), .ZN(U2842) );
  AOI22_X1 U6740 ( .A1(n4402), .A2(n6017), .B1(n5621), .B2(EBX_REG_16__SCAN_IN), .ZN(n5609) );
  OAI21_X1 U6741 ( .B1(n5798), .B2(n5623), .A(n5609), .ZN(U2843) );
  AOI22_X1 U6742 ( .A1(n4402), .A2(n6029), .B1(n5621), .B2(EBX_REG_15__SCAN_IN), .ZN(n5610) );
  OAI21_X1 U6743 ( .B1(n5813), .B2(n5623), .A(n5610), .ZN(U2844) );
  INV_X1 U6744 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5611) );
  INV_X1 U6745 ( .A(n5819), .ZN(n5666) );
  OAI222_X1 U6746 ( .A1(n6034), .A2(n5620), .B1(n5618), .B2(n5611), .C1(n5623), 
        .C2(n5666), .ZN(U2845) );
  AOI22_X1 U6747 ( .A1(n4402), .A2(n6055), .B1(n5621), .B2(EBX_REG_13__SCAN_IN), .ZN(n5612) );
  OAI21_X1 U6748 ( .B1(n5668), .B2(n5623), .A(n5612), .ZN(U2846) );
  INV_X1 U6749 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5613) );
  OAI222_X1 U6750 ( .A1(n6065), .A2(n5620), .B1(n5618), .B2(n5613), .C1(n5623), 
        .C2(n5670), .ZN(U2847) );
  AOI22_X1 U6751 ( .A1(n4402), .A2(n6438), .B1(n5621), .B2(EBX_REG_11__SCAN_IN), .ZN(n5614) );
  OAI21_X1 U6752 ( .B1(n5849), .B2(n5623), .A(n5614), .ZN(U2848) );
  OAI21_X1 U6753 ( .B1(n5616), .B2(n5482), .A(n5615), .ZN(n6391) );
  INV_X1 U6754 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5619) );
  AOI21_X1 U6755 ( .B1(n5617), .B2(n5479), .A(n5460), .ZN(n6398) );
  INV_X1 U6756 ( .A(n6398), .ZN(n5676) );
  OAI222_X1 U6757 ( .A1(n6391), .A2(n5620), .B1(n5619), .B2(n5618), .C1(n5676), 
        .C2(n5623), .ZN(U2849) );
  AOI22_X1 U6758 ( .A1(n4402), .A2(n6447), .B1(n5621), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5622) );
  OAI21_X1 U6759 ( .B1(n5865), .B2(n5623), .A(n5622), .ZN(U2850) );
  AOI22_X1 U6760 ( .A1(n5660), .A2(DATAI_29_), .B1(n5673), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U6761 ( .A1(n5661), .A2(DATAI_13_), .ZN(n5624) );
  OAI211_X1 U6762 ( .C1(n5626), .C2(n5680), .A(n5625), .B(n5624), .ZN(U2862)
         );
  AOI22_X1 U6763 ( .A1(n5660), .A2(DATAI_28_), .B1(n5673), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U6764 ( .A1(n5661), .A2(DATAI_12_), .ZN(n5627) );
  OAI211_X1 U6765 ( .C1(n5629), .C2(n5680), .A(n5628), .B(n5627), .ZN(U2863)
         );
  AOI22_X1 U6766 ( .A1(n5660), .A2(DATAI_27_), .B1(n5673), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U6767 ( .A1(n5661), .A2(DATAI_11_), .ZN(n5630) );
  OAI211_X1 U6768 ( .C1(n5632), .C2(n5680), .A(n5631), .B(n5630), .ZN(U2864)
         );
  AOI22_X1 U6769 ( .A1(n5660), .A2(DATAI_26_), .B1(n5673), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U6770 ( .A1(n5661), .A2(DATAI_10_), .ZN(n5633) );
  OAI211_X1 U6771 ( .C1(n5635), .C2(n5680), .A(n5634), .B(n5633), .ZN(U2865)
         );
  AOI22_X1 U6772 ( .A1(n5660), .A2(DATAI_25_), .B1(n5673), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U6773 ( .A1(n5661), .A2(DATAI_9_), .ZN(n5636) );
  OAI211_X1 U6774 ( .C1(n5719), .C2(n5680), .A(n5637), .B(n5636), .ZN(U2866)
         );
  AOI22_X1 U6775 ( .A1(n5660), .A2(DATAI_24_), .B1(n5673), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6776 ( .A1(n5661), .A2(DATAI_8_), .ZN(n5638) );
  OAI211_X1 U6777 ( .C1(n5640), .C2(n5680), .A(n5639), .B(n5638), .ZN(U2867)
         );
  AOI22_X1 U6778 ( .A1(n5660), .A2(DATAI_23_), .B1(n5673), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U6779 ( .A1(n5661), .A2(DATAI_7_), .ZN(n5641) );
  OAI211_X1 U6780 ( .C1(n5643), .C2(n5680), .A(n5642), .B(n5641), .ZN(U2868)
         );
  AOI22_X1 U6781 ( .A1(n5660), .A2(DATAI_22_), .B1(n5673), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6782 ( .A1(n5661), .A2(DATAI_6_), .ZN(n5644) );
  OAI211_X1 U6783 ( .C1(n5646), .C2(n5680), .A(n5645), .B(n5644), .ZN(U2869)
         );
  AOI22_X1 U6784 ( .A1(n5660), .A2(DATAI_21_), .B1(n5673), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6785 ( .A1(n5661), .A2(DATAI_5_), .ZN(n5647) );
  OAI211_X1 U6786 ( .C1(n5649), .C2(n5680), .A(n5648), .B(n5647), .ZN(U2870)
         );
  AOI22_X1 U6787 ( .A1(n5660), .A2(DATAI_20_), .B1(n5673), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U6788 ( .A1(n5661), .A2(DATAI_4_), .ZN(n5650) );
  OAI211_X1 U6789 ( .C1(n5652), .C2(n5680), .A(n5651), .B(n5650), .ZN(U2871)
         );
  AOI22_X1 U6790 ( .A1(n5660), .A2(DATAI_19_), .B1(n5673), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6791 ( .A1(n5661), .A2(DATAI_3_), .ZN(n5653) );
  OAI211_X1 U6792 ( .C1(n5774), .C2(n5680), .A(n5654), .B(n5653), .ZN(U2872)
         );
  AOI22_X1 U6793 ( .A1(n5660), .A2(DATAI_18_), .B1(n5673), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U6794 ( .A1(n5661), .A2(DATAI_2_), .ZN(n5655) );
  OAI211_X1 U6795 ( .C1(n5786), .C2(n5680), .A(n5656), .B(n5655), .ZN(U2873)
         );
  AOI22_X1 U6796 ( .A1(n5660), .A2(DATAI_17_), .B1(n5673), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U6797 ( .A1(n5661), .A2(DATAI_1_), .ZN(n5657) );
  OAI211_X1 U6798 ( .C1(n5659), .C2(n5680), .A(n5658), .B(n5657), .ZN(U2874)
         );
  AOI22_X1 U6799 ( .A1(n5660), .A2(DATAI_16_), .B1(n5673), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6800 ( .A1(n5661), .A2(DATAI_0_), .ZN(n5662) );
  OAI211_X1 U6801 ( .C1(n5798), .C2(n5680), .A(n5663), .B(n5662), .ZN(U2875)
         );
  AOI22_X1 U6802 ( .A1(n5674), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5673), .ZN(n5664) );
  OAI21_X1 U6803 ( .B1(n5813), .B2(n5680), .A(n5664), .ZN(U2876) );
  AOI22_X1 U6804 ( .A1(n5674), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5673), .ZN(n5665) );
  OAI21_X1 U6805 ( .B1(n5666), .B2(n5680), .A(n5665), .ZN(U2877) );
  AOI22_X1 U6806 ( .A1(n5674), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5673), .ZN(n5667) );
  OAI21_X1 U6807 ( .B1(n5668), .B2(n5680), .A(n5667), .ZN(U2878) );
  INV_X1 U6808 ( .A(EAX_REG_12__SCAN_IN), .ZN(n7028) );
  OAI222_X1 U6809 ( .A1(n5670), .A2(n5680), .B1(n5679), .B2(n5669), .C1(n5678), 
        .C2(n7028), .ZN(U2879) );
  INV_X1 U6810 ( .A(DATAI_11_), .ZN(n5672) );
  OAI222_X1 U6811 ( .A1(n5849), .A2(n5680), .B1(n5672), .B2(n5679), .C1(n5671), 
        .C2(n5678), .ZN(U2880) );
  AOI22_X1 U6812 ( .A1(n5674), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5673), .ZN(n5675) );
  OAI21_X1 U6813 ( .B1(n5676), .B2(n5680), .A(n5675), .ZN(U2881) );
  INV_X1 U6814 ( .A(DATAI_9_), .ZN(n6959) );
  INV_X1 U6815 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5677) );
  OAI222_X1 U6816 ( .A1(n5865), .A2(n5680), .B1(n5679), .B2(n6959), .C1(n5678), 
        .C2(n5677), .ZN(U2882) );
  XNOR2_X1 U6817 ( .A(n5684), .B(n5900), .ZN(n5908) );
  INV_X1 U6818 ( .A(n5685), .ZN(n5687) );
  NAND2_X1 U6819 ( .A1(n5868), .A2(REIP_REG_30__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U6820 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5686)
         );
  OAI211_X1 U6821 ( .C1(n5687), .C2(n6436), .A(n5903), .B(n5686), .ZN(n5688)
         );
  AOI21_X1 U6822 ( .B1(n5689), .B2(n6431), .A(n5688), .ZN(n5690) );
  OAI21_X1 U6823 ( .B1(n5908), .B2(n5892), .A(n5690), .ZN(U2956) );
  NAND2_X1 U6824 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  XNOR2_X1 U6825 ( .A(n5693), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5919)
         );
  AND2_X1 U6826 ( .A1(n5868), .A2(REIP_REG_29__SCAN_IN), .ZN(n5913) );
  AOI21_X1 U6827 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5913), 
        .ZN(n5694) );
  OAI21_X1 U6828 ( .B1(n5695), .B2(n6436), .A(n5694), .ZN(n5696) );
  AOI21_X1 U6829 ( .B1(n5697), .B2(n6431), .A(n5696), .ZN(n5698) );
  OAI21_X1 U6830 ( .B1(n5919), .B2(n5892), .A(n5698), .ZN(U2957) );
  NAND2_X1 U6831 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  XNOR2_X1 U6832 ( .A(n5701), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5928)
         );
  NAND2_X1 U6833 ( .A1(n5868), .A2(REIP_REG_27__SCAN_IN), .ZN(n5923) );
  INV_X1 U6834 ( .A(n5923), .ZN(n5702) );
  AOI21_X1 U6835 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5702), 
        .ZN(n5703) );
  OAI21_X1 U6836 ( .B1(n5704), .B2(n6436), .A(n5703), .ZN(n5705) );
  AOI21_X1 U6837 ( .B1(n5706), .B2(n6431), .A(n5705), .ZN(n5707) );
  OAI21_X1 U6838 ( .B1(n5928), .B2(n5892), .A(n5707), .ZN(U2959) );
  XNOR2_X1 U6839 ( .A(n5777), .B(n5708), .ZN(n5709) );
  XNOR2_X1 U6840 ( .A(n5710), .B(n5709), .ZN(n5937) );
  NAND2_X1 U6841 ( .A1(n5711), .A2(n5889), .ZN(n5712) );
  NAND2_X1 U6842 ( .A1(n5868), .A2(REIP_REG_26__SCAN_IN), .ZN(n5933) );
  OAI211_X1 U6843 ( .C1(n5884), .C2(n5713), .A(n5712), .B(n5933), .ZN(n5714)
         );
  AOI21_X1 U6844 ( .B1(n5715), .B2(n6431), .A(n5714), .ZN(n5716) );
  OAI21_X1 U6845 ( .B1(n5892), .B2(n5937), .A(n5716), .ZN(U2960) );
  AOI21_X1 U6846 ( .B1(n4419), .B2(n5718), .A(n5717), .ZN(n5945) );
  INV_X1 U6847 ( .A(n5719), .ZN(n5723) );
  AND2_X1 U6848 ( .A1(n5868), .A2(REIP_REG_25__SCAN_IN), .ZN(n5938) );
  AOI21_X1 U6849 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5938), 
        .ZN(n5720) );
  OAI21_X1 U6850 ( .B1(n5721), .B2(n6436), .A(n5720), .ZN(n5722) );
  AOI21_X1 U6851 ( .B1(n5723), .B2(n6431), .A(n5722), .ZN(n5724) );
  OAI21_X1 U6852 ( .B1(n5945), .B2(n5892), .A(n5724), .ZN(U2961) );
  AOI21_X1 U6853 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5725), 
        .ZN(n5726) );
  OAI21_X1 U6854 ( .B1(n5727), .B2(n6436), .A(n5726), .ZN(n5728) );
  AOI21_X1 U6855 ( .B1(n5729), .B2(n6431), .A(n5728), .ZN(n5730) );
  OAI21_X1 U6856 ( .B1(n5731), .B2(n5892), .A(n5730), .ZN(U2962) );
  XNOR2_X1 U6857 ( .A(n5735), .B(n5948), .ZN(n5954) );
  NAND2_X1 U6858 ( .A1(n5868), .A2(REIP_REG_23__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U6859 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5736)
         );
  OAI211_X1 U6860 ( .C1(n5737), .C2(n6436), .A(n5946), .B(n5736), .ZN(n5738)
         );
  AOI21_X1 U6861 ( .B1(n5739), .B2(n6431), .A(n5738), .ZN(n5740) );
  OAI21_X1 U6862 ( .B1(n5954), .B2(n5892), .A(n5740), .ZN(U2963) );
  INV_X1 U6863 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5964) );
  AOI21_X1 U6864 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5777), .A(n5742), 
        .ZN(n5743) );
  NAND2_X1 U6865 ( .A1(n5746), .A2(n5889), .ZN(n5747) );
  NAND2_X1 U6866 ( .A1(n5868), .A2(REIP_REG_22__SCAN_IN), .ZN(n5959) );
  OAI211_X1 U6867 ( .C1(n5884), .C2(n5748), .A(n5747), .B(n5959), .ZN(n5749)
         );
  AOI21_X1 U6868 ( .B1(n5750), .B2(n6431), .A(n5749), .ZN(n5751) );
  OAI21_X1 U6869 ( .B1(n5963), .B2(n5892), .A(n5751), .ZN(U2964) );
  AOI21_X1 U6870 ( .B1(n5754), .B2(n5753), .A(n5752), .ZN(n5972) );
  NAND2_X1 U6871 ( .A1(n5868), .A2(REIP_REG_21__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U6872 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5755)
         );
  OAI211_X1 U6873 ( .C1(n6436), .C2(n5756), .A(n5967), .B(n5755), .ZN(n5757)
         );
  AOI21_X1 U6874 ( .B1(n5758), .B2(n6431), .A(n5757), .ZN(n5759) );
  OAI21_X1 U6875 ( .B1(n5972), .B2(n5892), .A(n5759), .ZN(U2965) );
  XNOR2_X1 U6876 ( .A(n5832), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5760)
         );
  XNOR2_X1 U6877 ( .A(n3101), .B(n5760), .ZN(n5986) );
  INV_X1 U6878 ( .A(n5761), .ZN(n5763) );
  AND2_X1 U6879 ( .A1(n5868), .A2(REIP_REG_20__SCAN_IN), .ZN(n5977) );
  AOI21_X1 U6880 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5977), 
        .ZN(n5762) );
  OAI21_X1 U6881 ( .B1(n6436), .B2(n5763), .A(n5762), .ZN(n5764) );
  AOI21_X1 U6882 ( .B1(n5765), .B2(n6431), .A(n5764), .ZN(n5766) );
  OAI21_X1 U6883 ( .B1(n5986), .B2(n5892), .A(n5766), .ZN(U2966) );
  NAND2_X1 U6884 ( .A1(n5767), .A2(n5768), .ZN(n5988) );
  NAND3_X1 U6885 ( .A1(n5732), .A2(n4424), .A3(n5988), .ZN(n5773) );
  NAND2_X1 U6886 ( .A1(n5868), .A2(REIP_REG_19__SCAN_IN), .ZN(n5989) );
  OAI21_X1 U6887 ( .B1(n5884), .B2(n5769), .A(n5989), .ZN(n5770) );
  AOI21_X1 U6888 ( .B1(n5771), .B2(n5889), .A(n5770), .ZN(n5772) );
  OAI211_X1 U6889 ( .C1(n5885), .C2(n5774), .A(n5773), .B(n5772), .ZN(U2967)
         );
  OAI21_X1 U6890 ( .B1(n5832), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5775), 
        .ZN(n5808) );
  AND2_X1 U6891 ( .A1(n5777), .A2(n5776), .ZN(n5805) );
  NAND2_X1 U6892 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5804) );
  OAI21_X2 U6893 ( .B1(n5808), .B2(n5805), .A(n5804), .ZN(n5796) );
  NOR2_X1 U6894 ( .A1(n5777), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5794)
         );
  NAND2_X1 U6895 ( .A1(n5794), .A2(n6005), .ZN(n5779) );
  NAND4_X1 U6896 ( .A1(n5796), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A4(n5777), .ZN(n5778) );
  OAI21_X1 U6897 ( .B1(n5796), .B2(n5779), .A(n5778), .ZN(n5780) );
  XNOR2_X1 U6898 ( .A(n5780), .B(n6003), .ZN(n5996) );
  NAND2_X1 U6899 ( .A1(n5996), .A2(n4424), .ZN(n5785) );
  AND2_X1 U6900 ( .A1(n5868), .A2(REIP_REG_18__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U6901 ( .A1(n5884), .A2(n5781), .ZN(n5782) );
  AOI211_X1 U6902 ( .C1(n5889), .C2(n5783), .A(n5999), .B(n5782), .ZN(n5784)
         );
  OAI211_X1 U6903 ( .C1(n5885), .C2(n5786), .A(n5785), .B(n5784), .ZN(U2968)
         );
  NOR2_X1 U6904 ( .A1(n5832), .A2(n5787), .ZN(n5795) );
  MUX2_X1 U6905 ( .A(n5794), .B(n5795), .S(n5796), .Z(n5788) );
  XNOR2_X1 U6906 ( .A(n5788), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6013)
         );
  NAND2_X1 U6907 ( .A1(n5868), .A2(REIP_REG_17__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U6908 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5789)
         );
  OAI211_X1 U6909 ( .C1(n6436), .C2(n5790), .A(n6008), .B(n5789), .ZN(n5791)
         );
  AOI21_X1 U6910 ( .B1(n5792), .B2(n6431), .A(n5791), .ZN(n5793) );
  OAI21_X1 U6911 ( .B1(n6013), .B2(n5892), .A(n5793), .ZN(U2969) );
  NOR2_X1 U6912 ( .A1(n5795), .A2(n5794), .ZN(n5797) );
  XOR2_X1 U6913 ( .A(n5797), .B(n5796), .Z(n6025) );
  INV_X1 U6914 ( .A(n5798), .ZN(n5802) );
  AND2_X1 U6915 ( .A1(n5868), .A2(REIP_REG_16__SCAN_IN), .ZN(n6016) );
  AOI21_X1 U6916 ( .B1(n6424), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6016), 
        .ZN(n5799) );
  OAI21_X1 U6917 ( .B1(n6436), .B2(n5800), .A(n5799), .ZN(n5801) );
  AOI21_X1 U6918 ( .B1(n5802), .B2(n6431), .A(n5801), .ZN(n5803) );
  OAI21_X1 U6919 ( .B1(n6025), .B2(n5892), .A(n5803), .ZN(U2970) );
  INV_X1 U6920 ( .A(n5804), .ZN(n5806) );
  NOR2_X1 U6921 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  XNOR2_X1 U6922 ( .A(n5808), .B(n5807), .ZN(n6026) );
  NAND2_X1 U6923 ( .A1(n6026), .A2(n4424), .ZN(n5812) );
  INV_X1 U6924 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6691) );
  NOR2_X1 U6925 ( .A1(n6075), .A2(n6691), .ZN(n6028) );
  NOR2_X1 U6926 ( .A1(n6436), .A2(n5809), .ZN(n5810) );
  AOI211_X1 U6927 ( .C1(n6424), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6028), 
        .B(n5810), .ZN(n5811) );
  OAI211_X1 U6928 ( .C1(n5885), .C2(n5813), .A(n5812), .B(n5811), .ZN(U2971)
         );
  XNOR2_X1 U6929 ( .A(n5832), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5815)
         );
  XNOR2_X1 U6930 ( .A(n5814), .B(n5815), .ZN(n6051) );
  NAND2_X1 U6931 ( .A1(n5868), .A2(REIP_REG_14__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U6932 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5816)
         );
  OAI211_X1 U6933 ( .C1(n6436), .C2(n5817), .A(n6035), .B(n5816), .ZN(n5818)
         );
  AOI21_X1 U6934 ( .B1(n5819), .B2(n6431), .A(n5818), .ZN(n5820) );
  OAI21_X1 U6935 ( .B1(n5892), .B2(n6051), .A(n5820), .ZN(U2972) );
  OAI21_X1 U6936 ( .B1(n5823), .B2(n5822), .A(n5821), .ZN(n6052) );
  INV_X1 U6937 ( .A(n6052), .ZN(n5829) );
  NAND2_X1 U6938 ( .A1(n5868), .A2(REIP_REG_13__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U6939 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5824)
         );
  OAI211_X1 U6940 ( .C1(n6436), .C2(n5825), .A(n6056), .B(n5824), .ZN(n5826)
         );
  AOI21_X1 U6941 ( .B1(n5827), .B2(n6431), .A(n5826), .ZN(n5828) );
  OAI21_X1 U6942 ( .B1(n5829), .B2(n5892), .A(n5828), .ZN(U2973) );
  NAND2_X1 U6943 ( .A1(n5832), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5841) );
  OAI21_X1 U6944 ( .B1(n5843), .B2(n5840), .A(n5841), .ZN(n5834) );
  AOI21_X1 U6945 ( .B1(n5832), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5831), 
        .ZN(n5833) );
  XNOR2_X1 U6946 ( .A(n5834), .B(n5833), .ZN(n6069) );
  INV_X1 U6947 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6809) );
  NOR2_X1 U6948 ( .A1(n6075), .A2(n6809), .ZN(n6062) );
  AND2_X1 U6949 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5835)
         );
  AOI211_X1 U6950 ( .C1(n5836), .C2(n5889), .A(n6062), .B(n5835), .ZN(n5839)
         );
  NAND2_X1 U6951 ( .A1(n5837), .A2(n6431), .ZN(n5838) );
  OAI211_X1 U6952 ( .C1(n6069), .C2(n5892), .A(n5839), .B(n5838), .ZN(U2974)
         );
  INV_X1 U6953 ( .A(n5840), .ZN(n5842) );
  NAND2_X1 U6954 ( .A1(n5842), .A2(n5841), .ZN(n5844) );
  XOR2_X1 U6955 ( .A(n5844), .B(n5843), .Z(n6440) );
  NAND2_X1 U6956 ( .A1(n6440), .A2(n4424), .ZN(n5848) );
  NOR2_X1 U6957 ( .A1(n6075), .A2(n6686), .ZN(n6437) );
  NOR2_X1 U6958 ( .A1(n6436), .A2(n5845), .ZN(n5846) );
  AOI211_X1 U6959 ( .C1(n6424), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6437), 
        .B(n5846), .ZN(n5847) );
  OAI211_X1 U6960 ( .C1(n5885), .C2(n5849), .A(n5848), .B(n5847), .ZN(U2975)
         );
  INV_X1 U6961 ( .A(n5850), .ZN(n5852) );
  NOR2_X1 U6962 ( .A1(n5852), .A2(n5851), .ZN(n5854) );
  XOR2_X1 U6963 ( .A(n5854), .B(n5853), .Z(n6085) );
  AOI22_X1 U6964 ( .A1(n6424), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n5868), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5855) );
  OAI21_X1 U6965 ( .B1(n6436), .B2(n5856), .A(n5855), .ZN(n5857) );
  AOI21_X1 U6966 ( .B1(n6398), .B2(n6431), .A(n5857), .ZN(n5858) );
  OAI21_X1 U6967 ( .B1(n6085), .B2(n5892), .A(n5858), .ZN(U2976) );
  XNOR2_X1 U6968 ( .A(n5777), .B(n6801), .ZN(n5860) );
  XNOR2_X1 U6969 ( .A(n5859), .B(n5860), .ZN(n6449) );
  NAND2_X1 U6970 ( .A1(n6449), .A2(n4424), .ZN(n5864) );
  AND2_X1 U6971 ( .A1(n5868), .A2(REIP_REG_9__SCAN_IN), .ZN(n6446) );
  NOR2_X1 U6972 ( .A1(n6436), .A2(n5861), .ZN(n5862) );
  AOI211_X1 U6973 ( .C1(n6424), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6446), 
        .B(n5862), .ZN(n5863) );
  OAI211_X1 U6974 ( .C1(n5885), .C2(n5865), .A(n5864), .B(n5863), .ZN(U2977)
         );
  XNOR2_X1 U6975 ( .A(n5866), .B(n5867), .ZN(n6094) );
  INV_X1 U6976 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U6977 ( .A1(n5868), .A2(REIP_REG_8__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U6978 ( .B1(n5884), .B2(n5869), .A(n6086), .ZN(n5872) );
  NOR2_X1 U6979 ( .A1(n5870), .A2(n5885), .ZN(n5871) );
  AOI211_X1 U6980 ( .C1(n5889), .C2(n5873), .A(n5872), .B(n5871), .ZN(n5874)
         );
  OAI21_X1 U6981 ( .B1(n6094), .B2(n5892), .A(n5874), .ZN(U2978) );
  INV_X1 U6982 ( .A(n5876), .ZN(n5877) );
  XNOR2_X1 U6983 ( .A(n5875), .B(n5877), .ZN(n6453) );
  NAND2_X1 U6984 ( .A1(n6453), .A2(n4424), .ZN(n5881) );
  AND2_X1 U6985 ( .A1(n5868), .A2(REIP_REG_7__SCAN_IN), .ZN(n6454) );
  NOR2_X1 U6986 ( .A1(n6436), .A2(n5878), .ZN(n5879) );
  AOI211_X1 U6987 ( .C1(n6424), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6454), 
        .B(n5879), .ZN(n5880) );
  OAI211_X1 U6988 ( .C1(n5885), .C2(n5882), .A(n5881), .B(n5880), .ZN(U2979)
         );
  OAI21_X1 U6989 ( .B1(n5884), .B2(n6899), .A(n5883), .ZN(n5888) );
  NOR2_X1 U6990 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  AOI211_X1 U6991 ( .C1(n5889), .C2(n3269), .A(n5888), .B(n5887), .ZN(n5890)
         );
  OAI21_X1 U6992 ( .B1(n5892), .B2(n5891), .A(n5890), .ZN(U2980) );
  NOR3_X1 U6993 ( .A1(n5911), .A2(n5915), .A3(n5910), .ZN(n5901) );
  AND2_X1 U6994 ( .A1(n6021), .A2(n5910), .ZN(n5894) );
  NOR2_X1 U6995 ( .A1(n5926), .A2(n5894), .ZN(n5916) );
  OAI21_X1 U6996 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n6074), .A(n5916), 
        .ZN(n5906) );
  INV_X1 U6997 ( .A(n5906), .ZN(n5895) );
  OAI21_X1 U6998 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n6074), .A(n5895), 
        .ZN(n5898) );
  NAND2_X1 U6999 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  OAI211_X1 U7000 ( .C1(n5904), .C2(n6088), .A(n5903), .B(n5902), .ZN(n5905)
         );
  AOI21_X1 U7001 ( .B1(n5906), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5905), 
        .ZN(n5907) );
  OAI21_X1 U7002 ( .B1(n5908), .B2(n6084), .A(n5907), .ZN(U2988) );
  INV_X1 U7003 ( .A(n5909), .ZN(n5914) );
  NOR3_X1 U7004 ( .A1(n5911), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5910), 
        .ZN(n5912) );
  AOI211_X1 U7005 ( .C1(n5914), .C2(n6463), .A(n5913), .B(n5912), .ZN(n5918)
         );
  OR2_X1 U7006 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  OAI211_X1 U7007 ( .C1(n5919), .C2(n6084), .A(n5918), .B(n5917), .ZN(U2989)
         );
  NAND2_X1 U7008 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  OAI211_X1 U7009 ( .C1(n5924), .C2(n6088), .A(n5923), .B(n5922), .ZN(n5925)
         );
  AOI21_X1 U7010 ( .B1(n5926), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5925), 
        .ZN(n5927) );
  OAI21_X1 U7011 ( .B1(n5928), .B2(n6084), .A(n5927), .ZN(U2991) );
  INV_X1 U7012 ( .A(n5929), .ZN(n5930) );
  NAND3_X1 U7013 ( .A1(n5939), .A2(n5931), .A3(n5930), .ZN(n5932) );
  OAI211_X1 U7014 ( .C1(n5934), .C2(n6088), .A(n5933), .B(n5932), .ZN(n5935)
         );
  AOI21_X1 U7015 ( .B1(n5943), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5935), 
        .ZN(n5936) );
  OAI21_X1 U7016 ( .B1(n5937), .B2(n6084), .A(n5936), .ZN(U2992) );
  AOI21_X1 U7017 ( .B1(n5939), .B2(n4437), .A(n5938), .ZN(n5940) );
  OAI21_X1 U7018 ( .B1(n5941), .B2(n6088), .A(n5940), .ZN(n5942) );
  AOI21_X1 U7019 ( .B1(n5943), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5942), 
        .ZN(n5944) );
  OAI21_X1 U7020 ( .B1(n5945), .B2(n6084), .A(n5944), .ZN(U2993) );
  OAI21_X1 U7021 ( .B1(n5947), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5946), 
        .ZN(n5951) );
  NOR2_X1 U7022 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  AOI211_X1 U7023 ( .C1(n6463), .C2(n5952), .A(n5951), .B(n5950), .ZN(n5953)
         );
  OAI21_X1 U7024 ( .B1(n5954), .B2(n6084), .A(n5953), .ZN(U2995) );
  INV_X1 U7025 ( .A(n5955), .ZN(n5956) );
  NAND3_X1 U7026 ( .A1(n5965), .A2(n5957), .A3(n5956), .ZN(n5958) );
  OAI211_X1 U7027 ( .C1(n6088), .C2(n5960), .A(n5959), .B(n5958), .ZN(n5961)
         );
  AOI21_X1 U7028 ( .B1(n5970), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5961), 
        .ZN(n5962) );
  OAI21_X1 U7029 ( .B1(n5963), .B2(n6084), .A(n5962), .ZN(U2996) );
  NAND2_X1 U7030 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  OAI211_X1 U7031 ( .C1(n6088), .C2(n5968), .A(n5967), .B(n5966), .ZN(n5969)
         );
  AOI21_X1 U7032 ( .B1(n5970), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5969), 
        .ZN(n5971) );
  OAI21_X1 U7033 ( .B1(n5972), .B2(n6084), .A(n5971), .ZN(U2997) );
  NAND2_X1 U7034 ( .A1(n6006), .A2(n5973), .ZN(n5990) );
  NOR3_X1 U7035 ( .A1(n5990), .A2(n5975), .A3(n5974), .ZN(n5976) );
  AOI211_X1 U7036 ( .C1(n6463), .C2(n5978), .A(n5977), .B(n5976), .ZN(n5985)
         );
  INV_X1 U7037 ( .A(n5979), .ZN(n5982) );
  OAI21_X1 U7038 ( .B1(n5980), .B2(n6005), .A(n6072), .ZN(n5981) );
  NAND2_X1 U7039 ( .A1(n5982), .A2(n5981), .ZN(n6011) );
  AOI21_X1 U7040 ( .B1(n5983), .B2(n6005), .A(n6011), .ZN(n6004) );
  OAI21_X1 U7041 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6074), .A(n6004), 
        .ZN(n5987) );
  NAND2_X1 U7042 ( .A1(n5987), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5984) );
  OAI211_X1 U7043 ( .C1(n5986), .C2(n6084), .A(n5985), .B(n5984), .ZN(U2998)
         );
  INV_X1 U7044 ( .A(n5987), .ZN(n5995) );
  NAND3_X1 U7045 ( .A1(n5732), .A2(n4444), .A3(n5988), .ZN(n5994) );
  OAI21_X1 U7046 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5990), .A(n5989), 
        .ZN(n5991) );
  AOI21_X1 U7047 ( .B1(n6463), .B2(n5992), .A(n5991), .ZN(n5993) );
  OAI211_X1 U7048 ( .C1(n5995), .C2(n6932), .A(n5994), .B(n5993), .ZN(U2999)
         );
  NAND2_X1 U7049 ( .A1(n5996), .A2(n4444), .ZN(n6002) );
  INV_X1 U7050 ( .A(n6006), .ZN(n5997) );
  NOR3_X1 U7051 ( .A1(n5997), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6005), 
        .ZN(n5998) );
  AOI211_X1 U7052 ( .C1(n6463), .C2(n6000), .A(n5999), .B(n5998), .ZN(n6001)
         );
  OAI211_X1 U7053 ( .C1(n6004), .C2(n6003), .A(n6002), .B(n6001), .ZN(U3000)
         );
  NAND2_X1 U7054 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  OAI211_X1 U7055 ( .C1(n6088), .C2(n6009), .A(n6008), .B(n6007), .ZN(n6010)
         );
  AOI21_X1 U7056 ( .B1(n6011), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6010), 
        .ZN(n6012) );
  OAI21_X1 U7057 ( .B1(n6013), .B2(n6084), .A(n6012), .ZN(U3001) );
  NOR3_X1 U7058 ( .A1(n6014), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6036), 
        .ZN(n6015) );
  AOI211_X1 U7059 ( .C1(n6463), .C2(n6017), .A(n6016), .B(n6015), .ZN(n6024)
         );
  OR2_X1 U7060 ( .A1(n6043), .A2(n3191), .ZN(n6019) );
  INV_X1 U7061 ( .A(n6020), .ZN(n6038) );
  OAI21_X1 U7062 ( .B1(n6044), .B2(n6038), .A(n6021), .ZN(n6022) );
  NAND2_X1 U7063 ( .A1(n6444), .A2(n6022), .ZN(n6030) );
  NOR3_X1 U7064 ( .A1(n6044), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6036), 
        .ZN(n6027) );
  OAI21_X1 U7065 ( .B1(n6030), .B2(n6027), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n6023) );
  OAI211_X1 U7066 ( .C1(n6025), .C2(n6084), .A(n6024), .B(n6023), .ZN(U3002)
         );
  INV_X1 U7067 ( .A(n6026), .ZN(n6033) );
  AOI211_X1 U7068 ( .C1(n6463), .C2(n6029), .A(n6028), .B(n6027), .ZN(n6032)
         );
  NAND2_X1 U7069 ( .A1(n6030), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6031) );
  OAI211_X1 U7070 ( .C1(n6033), .C2(n6084), .A(n6032), .B(n6031), .ZN(U3003)
         );
  INV_X1 U7071 ( .A(n6034), .ZN(n6049) );
  OAI21_X1 U7072 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6036), .A(n6035), 
        .ZN(n6048) );
  AOI22_X1 U7073 ( .A1(n6039), .A2(n6038), .B1(n6041), .B2(n6037), .ZN(n6040)
         );
  NAND2_X1 U7074 ( .A1(n6444), .A2(n6040), .ZN(n6054) );
  INV_X1 U7075 ( .A(n6054), .ZN(n6046) );
  NOR2_X1 U7076 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6041), .ZN(n6053)
         );
  OAI21_X1 U7077 ( .B1(n6043), .B2(n6042), .A(n6053), .ZN(n6045) );
  AOI21_X1 U7078 ( .B1(n6046), .B2(n6045), .A(n6044), .ZN(n6047) );
  AOI211_X1 U7079 ( .C1(n6463), .C2(n6049), .A(n6048), .B(n6047), .ZN(n6050)
         );
  OAI21_X1 U7080 ( .B1(n6051), .B2(n6084), .A(n6050), .ZN(U3004) );
  NAND2_X1 U7081 ( .A1(n6052), .A2(n4444), .ZN(n6059) );
  AOI22_X1 U7082 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6054), .B1(n6053), .B2(n6439), .ZN(n6058) );
  NAND2_X1 U7083 ( .A1(n6463), .A2(n6055), .ZN(n6057) );
  NAND4_X1 U7084 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(U3005)
         );
  OAI221_X1 U7085 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6061), .C1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6060), .A(n6444), .ZN(n6067) );
  NAND3_X1 U7086 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n3665), .A3(n6439), .ZN(n6064) );
  INV_X1 U7087 ( .A(n6062), .ZN(n6063) );
  OAI211_X1 U7088 ( .C1(n6088), .C2(n6065), .A(n6064), .B(n6063), .ZN(n6066)
         );
  AOI21_X1 U7089 ( .B1(n6067), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n6066), 
        .ZN(n6068) );
  OAI21_X1 U7090 ( .B1(n6069), .B2(n6084), .A(n6068), .ZN(U3006) );
  AOI22_X1 U7091 ( .A1(n6073), .A2(n6072), .B1(n6071), .B2(n6070), .ZN(n6461)
         );
  OAI21_X1 U7092 ( .B1(n6089), .B2(n6074), .A(n6461), .ZN(n6445) );
  INV_X1 U7093 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6830) );
  OAI22_X1 U7094 ( .A1(n6088), .A2(n6391), .B1(n6830), .B2(n6075), .ZN(n6082)
         );
  NAND3_X1 U7095 ( .A1(n3126), .A2(n6077), .A3(n6076), .ZN(n6458) );
  NOR2_X1 U7096 ( .A1(n6078), .A2(n6458), .ZN(n6448) );
  OAI211_X1 U7097 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6448), .B(n6079), .ZN(n6080) );
  INV_X1 U7098 ( .A(n6080), .ZN(n6081) );
  AOI211_X1 U7099 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6445), .A(n6082), .B(n6081), .ZN(n6083) );
  OAI21_X1 U7100 ( .B1(n6085), .B2(n6084), .A(n6083), .ZN(U3008) );
  INV_X1 U7101 ( .A(n6461), .ZN(n6092) );
  OAI21_X1 U7102 ( .B1(n6088), .B2(n6087), .A(n6086), .ZN(n6091) );
  AOI211_X1 U7103 ( .C1(n3650), .C2(n3805), .A(n6089), .B(n6458), .ZN(n6090)
         );
  AOI211_X1 U7104 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6092), .A(n6091), 
        .B(n6090), .ZN(n6093) );
  OAI21_X1 U7105 ( .B1(n6084), .B2(n6094), .A(n6093), .ZN(U3010) );
  OAI211_X1 U7106 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6238), .A(n6095), .B(
        n6484), .ZN(n6096) );
  OAI21_X1 U7107 ( .B1(n6102), .B2(n6097), .A(n6096), .ZN(n6098) );
  MUX2_X1 U7108 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6098), .S(n6475), 
        .Z(U3464) );
  XNOR2_X1 U7109 ( .A(n6100), .B(n6099), .ZN(n6104) );
  INV_X1 U7110 ( .A(n6101), .ZN(n6103) );
  OAI22_X1 U7111 ( .A1(n6104), .A2(n6284), .B1(n6103), .B2(n6102), .ZN(n6105)
         );
  MUX2_X1 U7112 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6105), .S(n6475), 
        .Z(U3463) );
  OAI22_X1 U7113 ( .A1(n6107), .A2(n6734), .B1(n6106), .B2(n6635), .ZN(n6108)
         );
  MUX2_X1 U7114 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6108), .S(n6732), 
        .Z(U3456) );
  NOR2_X1 U7115 ( .A1(n6159), .A2(n6284), .ZN(n6109) );
  AOI21_X1 U7116 ( .B1(n6109), .B2(n6152), .A(n6200), .ZN(n6116) );
  NOR2_X1 U7117 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6110), .ZN(n6149)
         );
  INV_X1 U7118 ( .A(n6149), .ZN(n6114) );
  INV_X1 U7119 ( .A(n6111), .ZN(n6112) );
  OAI21_X1 U7120 ( .B1(n3277), .B2(n6326), .A(n6113), .ZN(n6202) );
  AOI211_X1 U7121 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6114), .A(n6478), .B(
        n6202), .ZN(n6115) );
  NAND2_X1 U7122 ( .A1(n6159), .A2(n6525), .ZN(n6121) );
  NAND2_X1 U7123 ( .A1(n6117), .A2(n6484), .ZN(n6119) );
  NAND2_X1 U7124 ( .A1(n3277), .A2(n6487), .ZN(n6118) );
  NAND2_X1 U7125 ( .A1(n6119), .A2(n6118), .ZN(n6148) );
  AOI22_X1 U7126 ( .A1(n6524), .A2(n6149), .B1(n6148), .B2(n6562), .ZN(n6120)
         );
  OAI211_X1 U7127 ( .C1(n6152), .C2(n6565), .A(n6121), .B(n6120), .ZN(n6122)
         );
  AOI21_X1 U7128 ( .B1(n6154), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n6122), 
        .ZN(n6123) );
  INV_X1 U7129 ( .A(n6123), .ZN(U3020) );
  NAND2_X1 U7130 ( .A1(n6159), .A2(n6529), .ZN(n6125) );
  AOI22_X1 U7131 ( .A1(n6528), .A2(n6149), .B1(n6148), .B2(n6569), .ZN(n6124)
         );
  OAI211_X1 U7132 ( .C1(n6152), .C2(n6572), .A(n6125), .B(n6124), .ZN(n6126)
         );
  AOI21_X1 U7133 ( .B1(n6154), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n6126), 
        .ZN(n6127) );
  INV_X1 U7134 ( .A(n6127), .ZN(U3021) );
  NAND2_X1 U7135 ( .A1(n6159), .A2(n6533), .ZN(n6129) );
  AOI22_X1 U7136 ( .A1(n6532), .A2(n6149), .B1(n6148), .B2(n6534), .ZN(n6128)
         );
  OAI211_X1 U7137 ( .C1(n6152), .C2(n6537), .A(n6129), .B(n6128), .ZN(n6130)
         );
  AOI21_X1 U7138 ( .B1(n6154), .B2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n6130), 
        .ZN(n6131) );
  INV_X1 U7139 ( .A(n6131), .ZN(U3022) );
  NAND2_X1 U7140 ( .A1(n6159), .A2(n6539), .ZN(n6133) );
  AOI22_X1 U7141 ( .A1(n6538), .A2(n6149), .B1(n6148), .B2(n6576), .ZN(n6132)
         );
  OAI211_X1 U7142 ( .C1(n6152), .C2(n6579), .A(n6133), .B(n6132), .ZN(n6134)
         );
  AOI21_X1 U7143 ( .B1(n6154), .B2(INSTQUEUE_REG_0__3__SCAN_IN), .A(n6134), 
        .ZN(n6135) );
  INV_X1 U7144 ( .A(n6135), .ZN(U3023) );
  NAND2_X1 U7145 ( .A1(n6159), .A2(n6543), .ZN(n6137) );
  AOI22_X1 U7146 ( .A1(n6542), .A2(n6149), .B1(n6148), .B2(n6544), .ZN(n6136)
         );
  OAI211_X1 U7147 ( .C1(n6152), .C2(n6547), .A(n6137), .B(n6136), .ZN(n6138)
         );
  AOI21_X1 U7148 ( .B1(n6154), .B2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n6138), 
        .ZN(n6139) );
  INV_X1 U7149 ( .A(n6139), .ZN(U3024) );
  NAND2_X1 U7150 ( .A1(n6159), .A2(n6303), .ZN(n6141) );
  AOI22_X1 U7151 ( .A1(n6508), .A2(n6149), .B1(n6148), .B2(n6583), .ZN(n6140)
         );
  OAI211_X1 U7152 ( .C1(n6152), .C2(n6586), .A(n6141), .B(n6140), .ZN(n6142)
         );
  AOI21_X1 U7153 ( .B1(n6154), .B2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n6142), 
        .ZN(n6143) );
  INV_X1 U7154 ( .A(n6143), .ZN(U3025) );
  NAND2_X1 U7155 ( .A1(n6159), .A2(n6550), .ZN(n6145) );
  AOI22_X1 U7156 ( .A1(n6548), .A2(n6149), .B1(n6148), .B2(n6553), .ZN(n6144)
         );
  OAI211_X1 U7157 ( .C1(n6152), .C2(n6558), .A(n6145), .B(n6144), .ZN(n6146)
         );
  AOI21_X1 U7158 ( .B1(n6154), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n6146), 
        .ZN(n6147) );
  INV_X1 U7159 ( .A(n6147), .ZN(U3026) );
  NAND2_X1 U7160 ( .A1(n6159), .A2(n6311), .ZN(n6151) );
  AOI22_X1 U7161 ( .A1(n6517), .A2(n6149), .B1(n6148), .B2(n6593), .ZN(n6150)
         );
  OAI211_X1 U7162 ( .C1(n6152), .C2(n6598), .A(n6151), .B(n6150), .ZN(n6153)
         );
  AOI21_X1 U7163 ( .B1(n6154), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n6153), 
        .ZN(n6155) );
  INV_X1 U7164 ( .A(n6155), .ZN(U3027) );
  AOI22_X1 U7165 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6157), .B1(n6562), 
        .B2(n6156), .ZN(n6161) );
  AOI22_X1 U7166 ( .A1(n6159), .A2(n6491), .B1(n6524), .B2(n6158), .ZN(n6160)
         );
  OAI211_X1 U7167 ( .C1(n6560), .C2(n6197), .A(n6161), .B(n6160), .ZN(U3028)
         );
  NOR2_X1 U7168 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6162), .ZN(n6166)
         );
  INV_X1 U7169 ( .A(n6197), .ZN(n6163) );
  OAI21_X1 U7170 ( .B1(n6163), .B2(n3272), .A(n6244), .ZN(n6164) );
  AOI21_X1 U7171 ( .B1(n6164), .B2(n6167), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6165) );
  NOR2_X1 U7172 ( .A1(n6478), .A2(n6486), .ZN(n6325) );
  NAND2_X1 U7173 ( .A1(n6191), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6172) );
  INV_X1 U7174 ( .A(n6166), .ZN(n6193) );
  INV_X1 U7175 ( .A(n6167), .ZN(n6169) );
  NOR2_X1 U7176 ( .A1(n6317), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6168)
         );
  AOI22_X1 U7177 ( .A1(n6169), .A2(n6484), .B1(n6477), .B2(n6168), .ZN(n6192)
         );
  OAI22_X1 U7178 ( .A1(n6559), .A2(n6193), .B1(n6192), .B2(n6330), .ZN(n6170)
         );
  AOI21_X1 U7179 ( .B1(n6525), .B2(n3272), .A(n6170), .ZN(n6171) );
  OAI211_X1 U7180 ( .C1(n6197), .C2(n6565), .A(n6172), .B(n6171), .ZN(U3036)
         );
  NAND2_X1 U7181 ( .A1(n6191), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6175) );
  OAI22_X1 U7182 ( .A1(n6566), .A2(n6193), .B1(n6192), .B2(n6334), .ZN(n6173)
         );
  AOI21_X1 U7183 ( .B1(n6529), .B2(n3272), .A(n6173), .ZN(n6174) );
  OAI211_X1 U7184 ( .C1(n6197), .C2(n6572), .A(n6175), .B(n6174), .ZN(U3037)
         );
  NAND2_X1 U7185 ( .A1(n6191), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6178) );
  OAI22_X1 U7186 ( .A1(n6257), .A2(n6193), .B1(n6192), .B2(n6338), .ZN(n6176)
         );
  AOI21_X1 U7187 ( .B1(n6533), .B2(n3272), .A(n6176), .ZN(n6177) );
  OAI211_X1 U7188 ( .C1(n6197), .C2(n6537), .A(n6178), .B(n6177), .ZN(U3038)
         );
  NAND2_X1 U7189 ( .A1(n6191), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6181) );
  OAI22_X1 U7190 ( .A1(n6573), .A2(n6193), .B1(n6192), .B2(n6342), .ZN(n6179)
         );
  AOI21_X1 U7191 ( .B1(n6539), .B2(n3272), .A(n6179), .ZN(n6180) );
  OAI211_X1 U7192 ( .C1(n6197), .C2(n6579), .A(n6181), .B(n6180), .ZN(U3039)
         );
  NAND2_X1 U7193 ( .A1(n6191), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6184) );
  OAI22_X1 U7194 ( .A1(n6264), .A2(n6193), .B1(n6192), .B2(n6346), .ZN(n6182)
         );
  AOI21_X1 U7195 ( .B1(n6543), .B2(n3272), .A(n6182), .ZN(n6183) );
  OAI211_X1 U7196 ( .C1(n6197), .C2(n6547), .A(n6184), .B(n6183), .ZN(U3040)
         );
  NAND2_X1 U7197 ( .A1(n6191), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6187) );
  OAI22_X1 U7198 ( .A1(n6580), .A2(n6193), .B1(n6192), .B2(n6350), .ZN(n6185)
         );
  AOI21_X1 U7199 ( .B1(n6303), .B2(n3272), .A(n6185), .ZN(n6186) );
  OAI211_X1 U7200 ( .C1(n6197), .C2(n6586), .A(n6187), .B(n6186), .ZN(U3041)
         );
  NAND2_X1 U7201 ( .A1(n6191), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6190) );
  OAI22_X1 U7202 ( .A1(n6271), .A2(n6193), .B1(n6192), .B2(n6354), .ZN(n6188)
         );
  AOI21_X1 U7203 ( .B1(n6550), .B2(n3272), .A(n6188), .ZN(n6189) );
  OAI211_X1 U7204 ( .C1(n6197), .C2(n6558), .A(n6190), .B(n6189), .ZN(U3042)
         );
  NAND2_X1 U7205 ( .A1(n6191), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6196) );
  OAI22_X1 U7206 ( .A1(n6588), .A2(n6193), .B1(n6192), .B2(n6361), .ZN(n6194)
         );
  AOI21_X1 U7207 ( .B1(n6311), .B2(n3272), .A(n6194), .ZN(n6195) );
  OAI211_X1 U7208 ( .C1(n6197), .C2(n6598), .A(n6196), .B(n6195), .ZN(U3043)
         );
  OAI22_X1 U7209 ( .A1(n6206), .A2(n6200), .B1(n6199), .B2(n6198), .ZN(n6204)
         );
  OR2_X1 U7210 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6201), .ZN(n6232)
         );
  AOI211_X1 U7211 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6232), .A(n6487), .B(
        n6202), .ZN(n6203) );
  NAND2_X1 U7212 ( .A1(n6230), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6211) );
  AOI22_X1 U7213 ( .A1(n6208), .A2(n6207), .B1(n6478), .B2(n3277), .ZN(n6231)
         );
  OAI22_X1 U7214 ( .A1(n6559), .A2(n6232), .B1(n6231), .B2(n6330), .ZN(n6209)
         );
  AOI21_X1 U7215 ( .B1(n6491), .B2(n6234), .A(n6209), .ZN(n6210) );
  OAI211_X1 U7216 ( .C1(n6560), .C2(n6237), .A(n6211), .B(n6210), .ZN(U3052)
         );
  NAND2_X1 U7217 ( .A1(n6230), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6214) );
  OAI22_X1 U7218 ( .A1(n6566), .A2(n6232), .B1(n6231), .B2(n6334), .ZN(n6212)
         );
  AOI21_X1 U7219 ( .B1(n6494), .B2(n6234), .A(n6212), .ZN(n6213) );
  OAI211_X1 U7220 ( .C1(n6237), .C2(n6567), .A(n6214), .B(n6213), .ZN(U3053)
         );
  NAND2_X1 U7221 ( .A1(n6230), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6217) );
  OAI22_X1 U7222 ( .A1(n6257), .A2(n6232), .B1(n6231), .B2(n6338), .ZN(n6215)
         );
  AOI21_X1 U7223 ( .B1(n6497), .B2(n6234), .A(n6215), .ZN(n6216) );
  OAI211_X1 U7224 ( .C1(n6237), .C2(n6500), .A(n6217), .B(n6216), .ZN(U3054)
         );
  NAND2_X1 U7225 ( .A1(n6230), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6220) );
  OAI22_X1 U7226 ( .A1(n6573), .A2(n6232), .B1(n6231), .B2(n6342), .ZN(n6218)
         );
  AOI21_X1 U7227 ( .B1(n6501), .B2(n6234), .A(n6218), .ZN(n6219) );
  OAI211_X1 U7228 ( .C1(n6237), .C2(n6574), .A(n6220), .B(n6219), .ZN(U3055)
         );
  NAND2_X1 U7229 ( .A1(n6230), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6223) );
  OAI22_X1 U7230 ( .A1(n6264), .A2(n6232), .B1(n6231), .B2(n6346), .ZN(n6221)
         );
  AOI21_X1 U7231 ( .B1(n6504), .B2(n6234), .A(n6221), .ZN(n6222) );
  OAI211_X1 U7232 ( .C1(n6237), .C2(n6507), .A(n6223), .B(n6222), .ZN(U3056)
         );
  NAND2_X1 U7233 ( .A1(n6230), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6226) );
  OAI22_X1 U7234 ( .A1(n6580), .A2(n6232), .B1(n6231), .B2(n6350), .ZN(n6224)
         );
  AOI21_X1 U7235 ( .B1(n6509), .B2(n6234), .A(n6224), .ZN(n6225) );
  OAI211_X1 U7236 ( .C1(n6237), .C2(n6581), .A(n6226), .B(n6225), .ZN(U3057)
         );
  NAND2_X1 U7237 ( .A1(n6230), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6229) );
  OAI22_X1 U7238 ( .A1(n6271), .A2(n6232), .B1(n6231), .B2(n6354), .ZN(n6227)
         );
  AOI21_X1 U7239 ( .B1(n6512), .B2(n6234), .A(n6227), .ZN(n6228) );
  OAI211_X1 U7240 ( .C1(n6237), .C2(n6515), .A(n6229), .B(n6228), .ZN(U3058)
         );
  NAND2_X1 U7241 ( .A1(n6230), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6236) );
  OAI22_X1 U7242 ( .A1(n6588), .A2(n6232), .B1(n6231), .B2(n6361), .ZN(n6233)
         );
  AOI21_X1 U7243 ( .B1(n6520), .B2(n6234), .A(n6233), .ZN(n6235) );
  OAI211_X1 U7244 ( .C1(n6237), .C2(n6589), .A(n6236), .B(n6235), .ZN(U3059)
         );
  NAND3_X1 U7245 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6610), .A3(n7013), .ZN(n6288) );
  NOR2_X1 U7246 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6288), .ZN(n6248)
         );
  INV_X1 U7247 ( .A(n6478), .ZN(n6241) );
  OAI211_X1 U7248 ( .C1(n6725), .C2(n6248), .A(n6241), .B(n6240), .ZN(n6247)
         );
  INV_X1 U7249 ( .A(n6551), .ZN(n6242) );
  NAND3_X1 U7250 ( .A1(n6314), .A2(n6484), .A3(n6242), .ZN(n6245) );
  INV_X1 U7251 ( .A(n6243), .ZN(n6282) );
  AND2_X1 U7252 ( .A1(n6282), .A2(n3087), .ZN(n6250) );
  AOI21_X1 U7253 ( .B1(n6245), .B2(n6244), .A(n6250), .ZN(n6246) );
  NAND2_X1 U7254 ( .A1(n6275), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6253) );
  INV_X1 U7255 ( .A(n6248), .ZN(n6277) );
  AOI22_X1 U7256 ( .A1(n6250), .A2(n6484), .B1(n6487), .B2(n6249), .ZN(n6276)
         );
  OAI22_X1 U7257 ( .A1(n6559), .A2(n6277), .B1(n6276), .B2(n6330), .ZN(n6251)
         );
  AOI21_X1 U7258 ( .B1(n6491), .B2(n6551), .A(n6251), .ZN(n6252) );
  OAI211_X1 U7259 ( .C1(n6560), .C2(n6314), .A(n6253), .B(n6252), .ZN(U3084)
         );
  NAND2_X1 U7260 ( .A1(n6275), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6256) );
  OAI22_X1 U7261 ( .A1(n6566), .A2(n6277), .B1(n6276), .B2(n6334), .ZN(n6254)
         );
  AOI21_X1 U7262 ( .B1(n6494), .B2(n6551), .A(n6254), .ZN(n6255) );
  OAI211_X1 U7263 ( .C1(n6567), .C2(n6314), .A(n6256), .B(n6255), .ZN(U3085)
         );
  NAND2_X1 U7264 ( .A1(n6275), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6260) );
  OAI22_X1 U7265 ( .A1(n6257), .A2(n6277), .B1(n6276), .B2(n6338), .ZN(n6258)
         );
  AOI21_X1 U7266 ( .B1(n6497), .B2(n6551), .A(n6258), .ZN(n6259) );
  OAI211_X1 U7267 ( .C1(n6500), .C2(n6314), .A(n6260), .B(n6259), .ZN(U3086)
         );
  NAND2_X1 U7268 ( .A1(n6275), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6263) );
  OAI22_X1 U7269 ( .A1(n6573), .A2(n6277), .B1(n6276), .B2(n6342), .ZN(n6261)
         );
  AOI21_X1 U7270 ( .B1(n6501), .B2(n6551), .A(n6261), .ZN(n6262) );
  OAI211_X1 U7271 ( .C1(n6574), .C2(n6314), .A(n6263), .B(n6262), .ZN(U3087)
         );
  NAND2_X1 U7272 ( .A1(n6275), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6267) );
  OAI22_X1 U7273 ( .A1(n6264), .A2(n6277), .B1(n6276), .B2(n6346), .ZN(n6265)
         );
  AOI21_X1 U7274 ( .B1(n6504), .B2(n6551), .A(n6265), .ZN(n6266) );
  OAI211_X1 U7275 ( .C1(n6507), .C2(n6314), .A(n6267), .B(n6266), .ZN(U3088)
         );
  NAND2_X1 U7276 ( .A1(n6275), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6270) );
  OAI22_X1 U7277 ( .A1(n6580), .A2(n6277), .B1(n6276), .B2(n6350), .ZN(n6268)
         );
  AOI21_X1 U7278 ( .B1(n6509), .B2(n6551), .A(n6268), .ZN(n6269) );
  OAI211_X1 U7279 ( .C1(n6581), .C2(n6314), .A(n6270), .B(n6269), .ZN(U3089)
         );
  NAND2_X1 U7280 ( .A1(n6275), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6274) );
  OAI22_X1 U7281 ( .A1(n6271), .A2(n6277), .B1(n6276), .B2(n6354), .ZN(n6272)
         );
  AOI21_X1 U7282 ( .B1(n6512), .B2(n6551), .A(n6272), .ZN(n6273) );
  OAI211_X1 U7283 ( .C1(n6515), .C2(n6314), .A(n6274), .B(n6273), .ZN(U3090)
         );
  NAND2_X1 U7284 ( .A1(n6275), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6280) );
  OAI22_X1 U7285 ( .A1(n6588), .A2(n6277), .B1(n6276), .B2(n6361), .ZN(n6278)
         );
  AOI21_X1 U7286 ( .B1(n6520), .B2(n6551), .A(n6278), .ZN(n6279) );
  OAI211_X1 U7287 ( .C1(n6589), .C2(n6314), .A(n6280), .B(n6279), .ZN(U3091)
         );
  AOI21_X1 U7288 ( .B1(n6292), .B2(STATEBS16_REG_SCAN_IN), .A(n6284), .ZN(
        n6287) );
  NOR2_X1 U7289 ( .A1(n6281), .A2(n6288), .ZN(n6310) );
  AOI21_X1 U7290 ( .B1(n6283), .B2(n6282), .A(n6310), .ZN(n6290) );
  AOI22_X1 U7291 ( .A1(n6287), .A2(n6290), .B1(n6284), .B2(n6288), .ZN(n6285)
         );
  NAND2_X1 U7292 ( .A1(n6286), .A2(n6285), .ZN(n6309) );
  INV_X1 U7293 ( .A(n6287), .ZN(n6289) );
  OAI22_X1 U7294 ( .A1(n6290), .A2(n6289), .B1(n6326), .B2(n6288), .ZN(n6308)
         );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6309), .B1(n6562), 
        .B2(n6308), .ZN(n6294) );
  AOI22_X1 U7296 ( .A1(n6359), .A2(n6525), .B1(n6524), .B2(n6310), .ZN(n6293)
         );
  OAI211_X1 U7297 ( .C1(n6314), .C2(n6565), .A(n6294), .B(n6293), .ZN(U3092)
         );
  AOI22_X1 U7298 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6309), .B1(n6569), 
        .B2(n6308), .ZN(n6296) );
  AOI22_X1 U7299 ( .A1(n6359), .A2(n6529), .B1(n6310), .B2(n6528), .ZN(n6295)
         );
  OAI211_X1 U7300 ( .C1(n6314), .C2(n6572), .A(n6296), .B(n6295), .ZN(U3093)
         );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6309), .B1(n6534), 
        .B2(n6308), .ZN(n6298) );
  AOI22_X1 U7302 ( .A1(n6359), .A2(n6533), .B1(n6310), .B2(n6532), .ZN(n6297)
         );
  OAI211_X1 U7303 ( .C1(n6314), .C2(n6537), .A(n6298), .B(n6297), .ZN(U3094)
         );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6309), .B1(n6576), 
        .B2(n6308), .ZN(n6300) );
  AOI22_X1 U7305 ( .A1(n6359), .A2(n6539), .B1(n6310), .B2(n6538), .ZN(n6299)
         );
  OAI211_X1 U7306 ( .C1(n6314), .C2(n6579), .A(n6300), .B(n6299), .ZN(U3095)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6309), .B1(n6544), 
        .B2(n6308), .ZN(n6302) );
  AOI22_X1 U7308 ( .A1(n6359), .A2(n6543), .B1(n6310), .B2(n6542), .ZN(n6301)
         );
  OAI211_X1 U7309 ( .C1(n6314), .C2(n6547), .A(n6302), .B(n6301), .ZN(U3096)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6309), .B1(n6583), 
        .B2(n6308), .ZN(n6305) );
  AOI22_X1 U7311 ( .A1(n6359), .A2(n6303), .B1(n6310), .B2(n6508), .ZN(n6304)
         );
  OAI211_X1 U7312 ( .C1(n6314), .C2(n6586), .A(n6305), .B(n6304), .ZN(U3097)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6309), .B1(n6553), 
        .B2(n6308), .ZN(n6307) );
  AOI22_X1 U7314 ( .A1(n6359), .A2(n6550), .B1(n6310), .B2(n6548), .ZN(n6306)
         );
  OAI211_X1 U7315 ( .C1(n6314), .C2(n6558), .A(n6307), .B(n6306), .ZN(U3098)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6309), .B1(n6593), 
        .B2(n6308), .ZN(n6313) );
  AOI22_X1 U7317 ( .A1(n6359), .A2(n6311), .B1(n6310), .B2(n6517), .ZN(n6312)
         );
  OAI211_X1 U7318 ( .C1(n6314), .C2(n6598), .A(n6313), .B(n6312), .ZN(U3099)
         );
  INV_X1 U7319 ( .A(n6597), .ZN(n6315) );
  OAI21_X1 U7320 ( .B1(n6359), .B2(n6315), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6316) );
  NOR2_X1 U7321 ( .A1(n6317), .A2(n6839), .ZN(n6318) );
  NOR2_X1 U7322 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6319), .ZN(n6356)
         );
  INV_X1 U7323 ( .A(n6320), .ZN(n6322) );
  INV_X1 U7324 ( .A(n6356), .ZN(n6321) );
  AOI22_X1 U7325 ( .A1(n6323), .A2(n6322), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6321), .ZN(n6324) );
  OAI211_X1 U7326 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6326), .A(n6325), .B(n6324), .ZN(n6355) );
  AOI22_X1 U7327 ( .A1(n6524), .A2(n6356), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n6355), .ZN(n6327) );
  OAI21_X1 U7328 ( .B1(n6597), .B2(n6560), .A(n6327), .ZN(n6328) );
  AOI21_X1 U7329 ( .B1(n6491), .B2(n6359), .A(n6328), .ZN(n6329) );
  OAI21_X1 U7330 ( .B1(n6362), .B2(n6330), .A(n6329), .ZN(U3100) );
  AOI22_X1 U7331 ( .A1(n6528), .A2(n6356), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n6355), .ZN(n6331) );
  OAI21_X1 U7332 ( .B1(n6597), .B2(n6567), .A(n6331), .ZN(n6332) );
  AOI21_X1 U7333 ( .B1(n6359), .B2(n6494), .A(n6332), .ZN(n6333) );
  OAI21_X1 U7334 ( .B1(n6362), .B2(n6334), .A(n6333), .ZN(U3101) );
  AOI22_X1 U7335 ( .A1(n6532), .A2(n6356), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n6355), .ZN(n6335) );
  OAI21_X1 U7336 ( .B1(n6597), .B2(n6500), .A(n6335), .ZN(n6336) );
  AOI21_X1 U7337 ( .B1(n6359), .B2(n6497), .A(n6336), .ZN(n6337) );
  OAI21_X1 U7338 ( .B1(n6362), .B2(n6338), .A(n6337), .ZN(U3102) );
  AOI22_X1 U7339 ( .A1(n6538), .A2(n6356), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n6355), .ZN(n6339) );
  OAI21_X1 U7340 ( .B1(n6597), .B2(n6574), .A(n6339), .ZN(n6340) );
  AOI21_X1 U7341 ( .B1(n6359), .B2(n6501), .A(n6340), .ZN(n6341) );
  OAI21_X1 U7342 ( .B1(n6362), .B2(n6342), .A(n6341), .ZN(U3103) );
  AOI22_X1 U7343 ( .A1(n6542), .A2(n6356), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n6355), .ZN(n6343) );
  OAI21_X1 U7344 ( .B1(n6597), .B2(n6507), .A(n6343), .ZN(n6344) );
  AOI21_X1 U7345 ( .B1(n6359), .B2(n6504), .A(n6344), .ZN(n6345) );
  OAI21_X1 U7346 ( .B1(n6362), .B2(n6346), .A(n6345), .ZN(U3104) );
  AOI22_X1 U7347 ( .A1(n6508), .A2(n6356), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n6355), .ZN(n6347) );
  OAI21_X1 U7348 ( .B1(n6597), .B2(n6581), .A(n6347), .ZN(n6348) );
  AOI21_X1 U7349 ( .B1(n6359), .B2(n6509), .A(n6348), .ZN(n6349) );
  OAI21_X1 U7350 ( .B1(n6362), .B2(n6350), .A(n6349), .ZN(U3105) );
  AOI22_X1 U7351 ( .A1(n6548), .A2(n6356), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n6355), .ZN(n6351) );
  OAI21_X1 U7352 ( .B1(n6597), .B2(n6515), .A(n6351), .ZN(n6352) );
  AOI21_X1 U7353 ( .B1(n6359), .B2(n6512), .A(n6352), .ZN(n6353) );
  OAI21_X1 U7354 ( .B1(n6362), .B2(n6354), .A(n6353), .ZN(U3106) );
  AOI22_X1 U7355 ( .A1(n6517), .A2(n6356), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n6355), .ZN(n6357) );
  OAI21_X1 U7356 ( .B1(n6597), .B2(n6589), .A(n6357), .ZN(n6358) );
  AOI21_X1 U7357 ( .B1(n6359), .B2(n6520), .A(n6358), .ZN(n6360) );
  OAI21_X1 U7358 ( .B1(n6362), .B2(n6361), .A(n6360), .ZN(U3107) );
  AND2_X1 U7359 ( .A1(n6746), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NAND3_X1 U7360 ( .A1(n6365), .A2(n6364), .A3(n6363), .ZN(n6366) );
  OAI22_X1 U7361 ( .A1(n6367), .A2(n6366), .B1(n6991), .B2(n6732), .ZN(U3455)
         );
  INV_X1 U7362 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6917) );
  OAI21_X1 U7363 ( .B1(n6719), .B2(n6917), .A(n6655), .ZN(U2789) );
  OAI21_X1 U7364 ( .B1(n6368), .B2(n6638), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6369) );
  OAI21_X1 U7365 ( .B1(n6370), .B2(n6642), .A(n6369), .ZN(U2790) );
  NOR2_X1 U7366 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6372) );
  OAI21_X1 U7367 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6372), .A(n6743), .ZN(n6371)
         );
  OAI21_X1 U7368 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6743), .A(n6371), .ZN(
        U2791) );
  OAI21_X1 U7369 ( .B1(BS16_N), .B2(n6372), .A(n6722), .ZN(n6721) );
  OAI21_X1 U7370 ( .B1(n6722), .B2(n6643), .A(n6721), .ZN(U2792) );
  NOR4_X1 U7371 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6376) );
  NOR4_X1 U7372 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6375) );
  NOR4_X1 U7373 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6374) );
  NOR4_X1 U7374 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6373) );
  NAND4_X1 U7375 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n6382)
         );
  NOR4_X1 U7376 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n6380) );
  AOI211_X1 U7377 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_29__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n6379) );
  NOR4_X1 U7378 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6378) );
  NOR4_X1 U7379 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6377) );
  NAND4_X1 U7380 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(n6381)
         );
  NOR2_X1 U7381 ( .A1(n6382), .A2(n6381), .ZN(n6738) );
  INV_X1 U7382 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6718) );
  NOR3_X1 U7383 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6384) );
  OAI21_X1 U7384 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6384), .A(n6738), .ZN(n6383)
         );
  OAI21_X1 U7385 ( .B1(n6738), .B2(n6718), .A(n6383), .ZN(U2794) );
  INV_X1 U7386 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6964) );
  AOI21_X1 U7387 ( .B1(n6944), .B2(n6964), .A(n6384), .ZN(n6386) );
  INV_X1 U7388 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6385) );
  INV_X1 U7389 ( .A(n6738), .ZN(n6741) );
  AOI22_X1 U7390 ( .A1(n6738), .A2(n6386), .B1(n6385), .B2(n6741), .ZN(U2795)
         );
  NOR3_X1 U7391 ( .A1(n6387), .A2(REIP_REG_10__SCAN_IN), .A3(n5488), .ZN(n6388) );
  AOI211_X1 U7392 ( .C1(n6390), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6389), 
        .B(n6388), .ZN(n6405) );
  INV_X1 U7393 ( .A(n6391), .ZN(n6392) );
  AOI22_X1 U7394 ( .A1(n6394), .A2(EBX_REG_10__SCAN_IN), .B1(n6393), .B2(n6392), .ZN(n6404) );
  AOI22_X1 U7395 ( .A1(n6398), .A2(n6397), .B1(n6396), .B2(n6395), .ZN(n6403)
         );
  INV_X1 U7396 ( .A(n6399), .ZN(n6400) );
  OAI21_X1 U7397 ( .B1(n6401), .B2(n6400), .A(REIP_REG_10__SCAN_IN), .ZN(n6402) );
  NAND4_X1 U7398 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(U2817)
         );
  INV_X1 U7399 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n7026) );
  AOI22_X1 U7400 ( .A1(n6409), .A2(EAX_REG_29__SCAN_IN), .B1(n6746), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6406) );
  OAI21_X1 U7401 ( .B1(n5208), .B2(n7026), .A(n6406), .ZN(U2894) );
  INV_X1 U7402 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U7403 ( .A1(n6409), .A2(EAX_REG_26__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U7404 ( .B1(n6408), .B2(n7009), .A(n6407), .ZN(U2897) );
  INV_X1 U7405 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6877) );
  AOI22_X1 U7406 ( .A1(n6409), .A2(EAX_REG_23__SCAN_IN), .B1(n6746), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n6410) );
  OAI21_X1 U7407 ( .B1(n5208), .B2(n6877), .A(n6410), .ZN(U2900) );
  INV_X1 U7408 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7409 ( .A1(n6746), .A2(DATAO_REG_14__SCAN_IN), .B1(n6745), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6411) );
  OAI21_X1 U7410 ( .B1(n5208), .B2(n6884), .A(n6411), .ZN(U2909) );
  INV_X1 U7411 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7412 ( .A1(n6746), .A2(DATAO_REG_13__SCAN_IN), .B1(n6745), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6412) );
  OAI21_X1 U7413 ( .B1(n5208), .B2(n6827), .A(n6412), .ZN(U2910) );
  AOI22_X1 U7414 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U7415 ( .A1(n6415), .A2(DATAI_10_), .ZN(n6417) );
  NAND2_X1 U7416 ( .A1(n6413), .A2(n6417), .ZN(U2934) );
  AOI22_X1 U7417 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U7418 ( .A1(n6415), .A2(DATAI_11_), .ZN(n6419) );
  NAND2_X1 U7419 ( .A1(n6414), .A2(n6419), .ZN(U2935) );
  AOI22_X1 U7420 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U7421 ( .A1(n6415), .A2(DATAI_14_), .ZN(n6422) );
  NAND2_X1 U7422 ( .A1(n6416), .A2(n6422), .ZN(U2938) );
  AOI22_X1 U7423 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U7424 ( .A1(n6418), .A2(n6417), .ZN(U2949) );
  AOI22_X1 U7425 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7426 ( .A1(n6420), .A2(n6419), .ZN(U2950) );
  AOI22_X1 U7427 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6421), .B1(n4692), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U7428 ( .A1(n6423), .A2(n6422), .ZN(U2953) );
  AOI22_X1 U7429 ( .A1(n5868), .A2(REIP_REG_2__SCAN_IN), .B1(n6424), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6434) );
  INV_X1 U7430 ( .A(n6425), .ZN(n6432) );
  INV_X1 U7431 ( .A(n6426), .ZN(n6428) );
  NAND2_X1 U7432 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  XNOR2_X1 U7433 ( .A(n6430), .B(n6429), .ZN(n6467) );
  AOI22_X1 U7434 ( .A1(n6432), .A2(n6431), .B1(n4424), .B2(n6467), .ZN(n6433)
         );
  OAI211_X1 U7435 ( .C1(n6436), .C2(n6435), .A(n6434), .B(n6433), .ZN(U2984)
         );
  AOI21_X1 U7436 ( .B1(n6463), .B2(n6438), .A(n6437), .ZN(n6442) );
  AOI22_X1 U7437 ( .A1(n6440), .A2(n4444), .B1(n6439), .B2(n6443), .ZN(n6441)
         );
  OAI211_X1 U7438 ( .C1(n6444), .C2(n6443), .A(n6442), .B(n6441), .ZN(U3007)
         );
  INV_X1 U7439 ( .A(n6445), .ZN(n6452) );
  AOI21_X1 U7440 ( .B1(n6463), .B2(n6447), .A(n6446), .ZN(n6451) );
  AOI22_X1 U7441 ( .A1(n6449), .A2(n4444), .B1(n6448), .B2(n6801), .ZN(n6450)
         );
  OAI211_X1 U7442 ( .C1(n6452), .C2(n6801), .A(n6451), .B(n6450), .ZN(U3009)
         );
  NAND2_X1 U7443 ( .A1(n6453), .A2(n4444), .ZN(n6457) );
  AOI21_X1 U7444 ( .B1(n6463), .B2(n6455), .A(n6454), .ZN(n6456) );
  OAI211_X1 U7445 ( .C1(n6458), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6457), 
        .B(n6456), .ZN(n6459) );
  INV_X1 U7446 ( .A(n6459), .ZN(n6460) );
  OAI21_X1 U7447 ( .B1(n6461), .B2(n3650), .A(n6460), .ZN(U3011) );
  AOI22_X1 U7448 ( .A1(n6463), .A2(n6462), .B1(n5868), .B2(REIP_REG_2__SCAN_IN), .ZN(n6474) );
  NAND3_X1 U7449 ( .A1(n6464), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U7450 ( .A1(n6466), .A2(n6465), .ZN(n6468) );
  AOI22_X1 U7451 ( .A1(n6468), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n4444), 
        .B2(n6467), .ZN(n6473) );
  OR3_X1 U7452 ( .A1(n6470), .A2(n6469), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6471) );
  NAND4_X1 U7453 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(U3016)
         );
  NOR2_X1 U7454 ( .A1(n6614), .A2(n6475), .ZN(U3019) );
  INV_X1 U7455 ( .A(n6476), .ZN(n6480) );
  NAND3_X1 U7456 ( .A1(n6478), .A2(n6477), .A3(n6839), .ZN(n6479) );
  OAI21_X1 U7457 ( .B1(n6480), .B2(n3087), .A(n6479), .ZN(n6518) );
  NOR2_X1 U7458 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6481), .ZN(n6516)
         );
  AOI22_X1 U7459 ( .A1(n6518), .A2(n6562), .B1(n6524), .B2(n6516), .ZN(n6493)
         );
  INV_X1 U7460 ( .A(n6557), .ZN(n6482) );
  OAI21_X1 U7461 ( .B1(n6519), .B2(n6482), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6483) );
  NAND3_X1 U7462 ( .A1(n6485), .A2(n6484), .A3(n6483), .ZN(n6490) );
  INV_X1 U7463 ( .A(n6516), .ZN(n6488) );
  AOI211_X1 U7464 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6488), .A(n6487), .B(
        n6486), .ZN(n6489) );
  NAND3_X1 U7465 ( .A1(n6839), .A2(n6490), .A3(n6489), .ZN(n6521) );
  AOI22_X1 U7466 ( .A1(n6521), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6491), 
        .B2(n6519), .ZN(n6492) );
  OAI211_X1 U7467 ( .C1(n6560), .C2(n6557), .A(n6493), .B(n6492), .ZN(U3068)
         );
  AOI22_X1 U7468 ( .A1(n6518), .A2(n6569), .B1(n6528), .B2(n6516), .ZN(n6496)
         );
  AOI22_X1 U7469 ( .A1(n6521), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6494), 
        .B2(n6519), .ZN(n6495) );
  OAI211_X1 U7470 ( .C1(n6567), .C2(n6557), .A(n6496), .B(n6495), .ZN(U3069)
         );
  AOI22_X1 U7471 ( .A1(n6518), .A2(n6534), .B1(n6532), .B2(n6516), .ZN(n6499)
         );
  AOI22_X1 U7472 ( .A1(n6521), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6497), 
        .B2(n6519), .ZN(n6498) );
  OAI211_X1 U7473 ( .C1(n6500), .C2(n6557), .A(n6499), .B(n6498), .ZN(U3070)
         );
  AOI22_X1 U7474 ( .A1(n6518), .A2(n6576), .B1(n6538), .B2(n6516), .ZN(n6503)
         );
  AOI22_X1 U7475 ( .A1(n6521), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6501), 
        .B2(n6519), .ZN(n6502) );
  OAI211_X1 U7476 ( .C1(n6574), .C2(n6557), .A(n6503), .B(n6502), .ZN(U3071)
         );
  AOI22_X1 U7477 ( .A1(n6518), .A2(n6544), .B1(n6542), .B2(n6516), .ZN(n6506)
         );
  AOI22_X1 U7478 ( .A1(n6521), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6504), 
        .B2(n6519), .ZN(n6505) );
  OAI211_X1 U7479 ( .C1(n6507), .C2(n6557), .A(n6506), .B(n6505), .ZN(U3072)
         );
  AOI22_X1 U7480 ( .A1(n6518), .A2(n6583), .B1(n6508), .B2(n6516), .ZN(n6511)
         );
  AOI22_X1 U7481 ( .A1(n6521), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6509), 
        .B2(n6519), .ZN(n6510) );
  OAI211_X1 U7482 ( .C1(n6581), .C2(n6557), .A(n6511), .B(n6510), .ZN(U3073)
         );
  AOI22_X1 U7483 ( .A1(n6518), .A2(n6553), .B1(n6548), .B2(n6516), .ZN(n6514)
         );
  AOI22_X1 U7484 ( .A1(n6521), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6512), 
        .B2(n6519), .ZN(n6513) );
  OAI211_X1 U7485 ( .C1(n6515), .C2(n6557), .A(n6514), .B(n6513), .ZN(U3074)
         );
  AOI22_X1 U7486 ( .A1(n6518), .A2(n6593), .B1(n6517), .B2(n6516), .ZN(n6523)
         );
  AOI22_X1 U7487 ( .A1(n6521), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6520), 
        .B2(n6519), .ZN(n6522) );
  OAI211_X1 U7488 ( .C1(n6589), .C2(n6557), .A(n6523), .B(n6522), .ZN(U3075)
         );
  AOI22_X1 U7489 ( .A1(n6551), .A2(n6525), .B1(n6549), .B2(n6524), .ZN(n6527)
         );
  AOI22_X1 U7490 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6554), .B1(n6562), 
        .B2(n6552), .ZN(n6526) );
  OAI211_X1 U7491 ( .C1(n6565), .C2(n6557), .A(n6527), .B(n6526), .ZN(U3076)
         );
  AOI22_X1 U7492 ( .A1(n6551), .A2(n6529), .B1(n6549), .B2(n6528), .ZN(n6531)
         );
  AOI22_X1 U7493 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6554), .B1(n6569), 
        .B2(n6552), .ZN(n6530) );
  OAI211_X1 U7494 ( .C1(n6572), .C2(n6557), .A(n6531), .B(n6530), .ZN(U3077)
         );
  AOI22_X1 U7495 ( .A1(n6551), .A2(n6533), .B1(n6549), .B2(n6532), .ZN(n6536)
         );
  AOI22_X1 U7496 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6554), .B1(n6534), 
        .B2(n6552), .ZN(n6535) );
  OAI211_X1 U7497 ( .C1(n6537), .C2(n6557), .A(n6536), .B(n6535), .ZN(U3078)
         );
  AOI22_X1 U7498 ( .A1(n6551), .A2(n6539), .B1(n6549), .B2(n6538), .ZN(n6541)
         );
  AOI22_X1 U7499 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6554), .B1(n6576), 
        .B2(n6552), .ZN(n6540) );
  OAI211_X1 U7500 ( .C1(n6579), .C2(n6557), .A(n6541), .B(n6540), .ZN(U3079)
         );
  AOI22_X1 U7501 ( .A1(n6551), .A2(n6543), .B1(n6549), .B2(n6542), .ZN(n6546)
         );
  AOI22_X1 U7502 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6554), .B1(n6544), 
        .B2(n6552), .ZN(n6545) );
  OAI211_X1 U7503 ( .C1(n6547), .C2(n6557), .A(n6546), .B(n6545), .ZN(U3080)
         );
  AOI22_X1 U7504 ( .A1(n6551), .A2(n6550), .B1(n6549), .B2(n6548), .ZN(n6556)
         );
  AOI22_X1 U7505 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6554), .B1(n6553), 
        .B2(n6552), .ZN(n6555) );
  OAI211_X1 U7506 ( .C1(n6558), .C2(n6557), .A(n6556), .B(n6555), .ZN(U3082)
         );
  OAI22_X1 U7507 ( .A1(n6590), .A2(n6560), .B1(n6559), .B2(n6587), .ZN(n6561)
         );
  INV_X1 U7508 ( .A(n6561), .ZN(n6564) );
  AOI22_X1 U7509 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6594), .B1(n6562), 
        .B2(n6592), .ZN(n6563) );
  OAI211_X1 U7510 ( .C1(n6565), .C2(n6597), .A(n6564), .B(n6563), .ZN(U3108)
         );
  OAI22_X1 U7511 ( .A1(n6590), .A2(n6567), .B1(n6566), .B2(n6587), .ZN(n6568)
         );
  INV_X1 U7512 ( .A(n6568), .ZN(n6571) );
  AOI22_X1 U7513 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6594), .B1(n6569), 
        .B2(n6592), .ZN(n6570) );
  OAI211_X1 U7514 ( .C1(n6572), .C2(n6597), .A(n6571), .B(n6570), .ZN(U3109)
         );
  OAI22_X1 U7515 ( .A1(n6590), .A2(n6574), .B1(n6573), .B2(n6587), .ZN(n6575)
         );
  INV_X1 U7516 ( .A(n6575), .ZN(n6578) );
  AOI22_X1 U7517 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6594), .B1(n6576), 
        .B2(n6592), .ZN(n6577) );
  OAI211_X1 U7518 ( .C1(n6579), .C2(n6597), .A(n6578), .B(n6577), .ZN(U3111)
         );
  OAI22_X1 U7519 ( .A1(n6590), .A2(n6581), .B1(n6580), .B2(n6587), .ZN(n6582)
         );
  INV_X1 U7520 ( .A(n6582), .ZN(n6585) );
  AOI22_X1 U7521 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6594), .B1(n6583), 
        .B2(n6592), .ZN(n6584) );
  OAI211_X1 U7522 ( .C1(n6586), .C2(n6597), .A(n6585), .B(n6584), .ZN(U3113)
         );
  OAI22_X1 U7523 ( .A1(n6590), .A2(n6589), .B1(n6588), .B2(n6587), .ZN(n6591)
         );
  INV_X1 U7524 ( .A(n6591), .ZN(n6596) );
  AOI22_X1 U7525 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6594), .B1(n6593), 
        .B2(n6592), .ZN(n6595) );
  OAI211_X1 U7526 ( .C1(n6598), .C2(n6597), .A(n6596), .B(n6595), .ZN(U3115)
         );
  AOI22_X1 U7527 ( .A1(n3895), .A2(n6600), .B1(n6599), .B2(n6727), .ZN(n6730)
         );
  NAND2_X1 U7528 ( .A1(n6601), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6735) );
  NAND3_X1 U7529 ( .A1(n6730), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6735), .ZN(n6605) );
  INV_X1 U7530 ( .A(n6602), .ZN(n6603) );
  OAI211_X1 U7531 ( .C1(n7013), .C2(n6605), .A(n6604), .B(n6603), .ZN(n6607)
         );
  NAND2_X1 U7532 ( .A1(n6605), .A2(n7013), .ZN(n6606) );
  NAND2_X1 U7533 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  AOI222_X1 U7534 ( .A1(n6610), .A2(n6609), .B1(n6610), .B2(n6608), .C1(n6609), 
        .C2(n6608), .ZN(n6613) );
  OR2_X1 U7535 ( .A1(n6613), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6612)
         );
  NAND2_X1 U7536 ( .A1(n6612), .A2(n6611), .ZN(n6616) );
  NAND2_X1 U7537 ( .A1(n6613), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6615) );
  NAND3_X1 U7538 ( .A1(n6616), .A2(n6615), .A3(n6614), .ZN(n6626) );
  NOR2_X1 U7539 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6620) );
  OAI211_X1 U7540 ( .C1(n6620), .C2(n6619), .A(n6618), .B(n6617), .ZN(n6621)
         );
  NOR2_X1 U7541 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  AND2_X1 U7542 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  NAND2_X1 U7543 ( .A1(n6639), .A2(n6640), .ZN(n6628) );
  NAND2_X1 U7544 ( .A1(READY_N), .A2(n6744), .ZN(n6627) );
  NAND2_X1 U7545 ( .A1(n6628), .A2(n6627), .ZN(n6632) );
  OR2_X1 U7546 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  OAI21_X1 U7547 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4465), .A(n6724), .ZN(
        n6645) );
  AOI221_X1 U7548 ( .B1(n6634), .B2(STATE2_REG_0__SCAN_IN), .C1(n6645), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6633), .ZN(n6637) );
  OAI211_X1 U7549 ( .C1(n6650), .C2(n6635), .A(n6724), .B(n6642), .ZN(n6636)
         );
  OAI211_X1 U7550 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n6636), .ZN(U3148)
         );
  NOR2_X1 U7551 ( .A1(n6642), .A2(n6734), .ZN(n6641) );
  AOI21_X1 U7552 ( .B1(n6641), .B2(n4465), .A(n6640), .ZN(n6647) );
  NAND2_X1 U7553 ( .A1(n6642), .A2(n6326), .ZN(n6644) );
  INV_X1 U7554 ( .A(n6644), .ZN(n6653) );
  OAI221_X1 U7555 ( .B1(n6653), .B2(n6645), .C1(n6644), .C2(n6643), .A(
        STATE2_REG_1__SCAN_IN), .ZN(n6646) );
  OAI21_X1 U7556 ( .B1(n6648), .B2(n6647), .A(n6646), .ZN(U3149) );
  INV_X1 U7557 ( .A(n6649), .ZN(n6723) );
  OAI211_X1 U7558 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4465), .A(n6723), .B(
        n6650), .ZN(n6652) );
  OAI21_X1 U7559 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(U3150) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6655), .ZN(U3151) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6655), .ZN(U3152) );
  INV_X1 U7562 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6984) );
  NOR2_X1 U7563 ( .A1(n6722), .A2(n6984), .ZN(U3153) );
  AND2_X1 U7564 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6655), .ZN(U3154) );
  AND2_X1 U7565 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6655), .ZN(U3155) );
  AND2_X1 U7566 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6655), .ZN(U3156) );
  AND2_X1 U7567 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6655), .ZN(U3157) );
  AND2_X1 U7568 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6655), .ZN(U3158) );
  AND2_X1 U7569 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6655), .ZN(U3159) );
  AND2_X1 U7570 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6655), .ZN(U3160) );
  AND2_X1 U7571 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6655), .ZN(U3161) );
  AND2_X1 U7572 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6655), .ZN(U3162) );
  AND2_X1 U7573 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6655), .ZN(U3163) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6655), .ZN(U3164) );
  AND2_X1 U7575 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6655), .ZN(U3165) );
  AND2_X1 U7576 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6655), .ZN(U3166) );
  AND2_X1 U7577 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6654), .ZN(U3167) );
  AND2_X1 U7578 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6654), .ZN(U3168) );
  AND2_X1 U7579 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6654), .ZN(U3169) );
  AND2_X1 U7580 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6654), .ZN(U3170) );
  AND2_X1 U7581 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6654), .ZN(U3171) );
  AND2_X1 U7582 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6654), .ZN(U3172) );
  INV_X1 U7583 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U7584 ( .A1(n6722), .A2(n6925), .ZN(U3173) );
  AND2_X1 U7585 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6654), .ZN(U3174) );
  AND2_X1 U7586 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6654), .ZN(U3175) );
  AND2_X1 U7587 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6654), .ZN(U3176) );
  AND2_X1 U7588 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6654), .ZN(U3177) );
  AND2_X1 U7589 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6654), .ZN(U3178) );
  AND2_X1 U7590 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6655), .ZN(U3179) );
  INV_X1 U7591 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U7592 ( .A1(n6722), .A2(n6873), .ZN(U3180) );
  NAND2_X1 U7593 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6659) );
  NAND2_X1 U7594 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6657) );
  INV_X1 U7595 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U7596 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6660) );
  OAI21_X1 U7597 ( .B1(n4465), .B2(n6668), .A(n6660), .ZN(n6656) );
  INV_X1 U7598 ( .A(NA_N), .ZN(n6870) );
  AOI221_X1 U7599 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6870), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6671) );
  AOI21_X1 U7600 ( .B1(n6657), .B2(n6656), .A(n6671), .ZN(n6658) );
  OAI221_X1 U7601 ( .B1(n6719), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6719), 
        .C2(n6659), .A(n6658), .ZN(U3181) );
  INV_X1 U7602 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6667) );
  NOR2_X1 U7603 ( .A1(n3752), .A2(n6667), .ZN(n6662) );
  INV_X1 U7604 ( .A(n6659), .ZN(n6661) );
  OAI21_X1 U7605 ( .B1(n6662), .B2(n6661), .A(n6660), .ZN(n6663) );
  OAI211_X1 U7606 ( .C1(n6668), .C2(n4465), .A(n6664), .B(n6663), .ZN(U3182)
         );
  NAND2_X1 U7607 ( .A1(READY_N), .A2(n6870), .ZN(n6666) );
  AOI21_X1 U7608 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6666), .A(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n6665) );
  AOI221_X1 U7609 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6665), .C2(HOLD), .A(n3752), .ZN(n6672) );
  OR4_X1 U7610 ( .A1(n3752), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6670) );
  NAND3_X1 U7611 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .A3(
        STATE_REG_2__SCAN_IN), .ZN(n6669) );
  OAI211_X1 U7612 ( .C1(n6672), .C2(n6671), .A(n6670), .B(n6669), .ZN(U3183)
         );
  NOR2_X1 U7613 ( .A1(n6673), .A2(n6743), .ZN(n6709) );
  NAND2_X1 U7614 ( .A1(n6673), .A2(n6719), .ZN(n6711) );
  INV_X1 U7615 ( .A(n6711), .ZN(n6714) );
  AOI22_X1 U7616 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6743), .ZN(n6674) );
  OAI21_X1 U7617 ( .B1(n6944), .B2(n6716), .A(n6674), .ZN(U3184) );
  AOI22_X1 U7618 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6743), .ZN(n6675) );
  OAI21_X1 U7619 ( .B1(n5566), .B2(n6705), .A(n6675), .ZN(U3185) );
  INV_X1 U7620 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6677) );
  AOI22_X1 U7621 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6743), .ZN(n6676) );
  OAI21_X1 U7622 ( .B1(n6677), .B2(n6705), .A(n6676), .ZN(U3186) );
  INV_X1 U7623 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6679) );
  AOI22_X1 U7624 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6743), .ZN(n6678) );
  OAI21_X1 U7625 ( .B1(n6679), .B2(n6705), .A(n6678), .ZN(U3187) );
  AOI22_X1 U7626 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6743), .ZN(n6680) );
  OAI21_X1 U7627 ( .B1(n5530), .B2(n6705), .A(n6680), .ZN(U3188) );
  AOI22_X1 U7628 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6743), .ZN(n6681) );
  OAI21_X1 U7629 ( .B1(n5502), .B2(n6705), .A(n6681), .ZN(U3189) );
  INV_X1 U7630 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6836) );
  OAI222_X1 U7631 ( .A1(n6705), .A2(n6682), .B1(n6836), .B2(n6719), .C1(n6683), 
        .C2(n6711), .ZN(U3190) );
  INV_X1 U7632 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6821) );
  OAI222_X1 U7633 ( .A1(n6711), .A2(n5488), .B1(n6821), .B2(n6719), .C1(n6683), 
        .C2(n6705), .ZN(U3191) );
  AOI22_X1 U7634 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6743), .ZN(n6684) );
  OAI21_X1 U7635 ( .B1(n5488), .B2(n6705), .A(n6684), .ZN(U3192) );
  INV_X1 U7636 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6869) );
  OAI222_X1 U7637 ( .A1(n6705), .A2(n6830), .B1(n6869), .B2(n6719), .C1(n6686), 
        .C2(n6711), .ZN(U3193) );
  AOI22_X1 U7638 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6743), .ZN(n6685) );
  OAI21_X1 U7639 ( .B1(n6686), .B2(n6705), .A(n6685), .ZN(U3194) );
  AOI22_X1 U7640 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6743), .ZN(n6687) );
  OAI21_X1 U7641 ( .B1(n6809), .B2(n6705), .A(n6687), .ZN(U3195) );
  INV_X1 U7642 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6921) );
  OAI222_X1 U7643 ( .A1(n6705), .A2(n6688), .B1(n6921), .B2(n6719), .C1(n6690), 
        .C2(n6711), .ZN(U3196) );
  AOI22_X1 U7644 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6743), .ZN(n6689) );
  OAI21_X1 U7645 ( .B1(n6690), .B2(n6705), .A(n6689), .ZN(U3197) );
  INV_X1 U7646 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6842) );
  OAI222_X1 U7647 ( .A1(n6705), .A2(n6691), .B1(n6842), .B2(n6719), .C1(n7004), 
        .C2(n6711), .ZN(U3198) );
  AOI22_X1 U7648 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6743), .ZN(n6692) );
  OAI21_X1 U7649 ( .B1(n7004), .B2(n6705), .A(n6692), .ZN(U3199) );
  INV_X1 U7650 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6794) );
  OAI222_X1 U7651 ( .A1(n6711), .A2(n6998), .B1(n6794), .B2(n6719), .C1(n5380), 
        .C2(n6705), .ZN(U3200) );
  INV_X1 U7652 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6795) );
  OAI222_X1 U7653 ( .A1(n6711), .A2(n6694), .B1(n6795), .B2(n6719), .C1(n6998), 
        .C2(n6705), .ZN(U3201) );
  AOI22_X1 U7654 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6743), .ZN(n6693) );
  OAI21_X1 U7655 ( .B1(n6694), .B2(n6716), .A(n6693), .ZN(U3202) );
  INV_X1 U7656 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6695) );
  INV_X1 U7657 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6800) );
  INV_X1 U7658 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6697) );
  OAI222_X1 U7659 ( .A1(n6716), .A2(n6695), .B1(n6800), .B2(n6719), .C1(n6697), 
        .C2(n6711), .ZN(U3203) );
  AOI22_X1 U7660 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6743), .ZN(n6696) );
  OAI21_X1 U7661 ( .B1(n6697), .B2(n6716), .A(n6696), .ZN(U3204) );
  INV_X1 U7662 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6699) );
  AOI22_X1 U7663 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6743), .ZN(n6698) );
  OAI21_X1 U7664 ( .B1(n6699), .B2(n6716), .A(n6698), .ZN(U3205) );
  AOI22_X1 U7665 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6709), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6743), .ZN(n6700) );
  OAI21_X1 U7666 ( .B1(n6701), .B2(n6711), .A(n6700), .ZN(U3206) );
  AOI22_X1 U7667 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6709), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6743), .ZN(n6702) );
  OAI21_X1 U7668 ( .B1(n6936), .B2(n6711), .A(n6702), .ZN(U3207) );
  INV_X1 U7669 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U7670 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6709), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6743), .ZN(n6703) );
  OAI21_X1 U7671 ( .B1(n6706), .B2(n6711), .A(n6703), .ZN(U3208) );
  AOI22_X1 U7672 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6743), .ZN(n6704) );
  OAI21_X1 U7673 ( .B1(n6706), .B2(n6705), .A(n6704), .ZN(U3209) );
  INV_X1 U7674 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6862) );
  OAI222_X1 U7675 ( .A1(n6716), .A2(n6708), .B1(n6862), .B2(n6719), .C1(n6707), 
        .C2(n6711), .ZN(U3210) );
  AOI22_X1 U7676 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6709), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6743), .ZN(n6710) );
  OAI21_X1 U7677 ( .B1(n6713), .B2(n6711), .A(n6710), .ZN(U3211) );
  AOI22_X1 U7678 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6743), .ZN(n6712) );
  OAI21_X1 U7679 ( .B1(n6713), .B2(n6716), .A(n6712), .ZN(U3212) );
  AOI22_X1 U7680 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6714), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6743), .ZN(n6715) );
  OAI21_X1 U7681 ( .B1(n6717), .B2(n6716), .A(n6715), .ZN(U3213) );
  MUX2_X1 U7682 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6743), .Z(U3445) );
  MUX2_X1 U7683 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6743), .Z(U3446) );
  INV_X1 U7684 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U7685 ( .A1(n6719), .A2(n6718), .B1(n6845), .B2(n6743), .ZN(U3447)
         );
  MUX2_X1 U7686 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6743), .Z(U3448) );
  OAI21_X1 U7687 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6722), .A(n6721), .ZN(
        n6720) );
  INV_X1 U7688 ( .A(n6720), .ZN(U3451) );
  OAI21_X1 U7689 ( .B1(n6722), .B2(n6964), .A(n6721), .ZN(U3452) );
  OAI221_X1 U7690 ( .B1(n6725), .B2(STATE2_REG_0__SCAN_IN), .C1(n6725), .C2(
        n6724), .A(n6723), .ZN(U3453) );
  AOI22_X1 U7691 ( .A1(n6728), .A2(n6727), .B1(STATE2_REG_1__SCAN_IN), .B2(
        n6726), .ZN(n6729) );
  OAI211_X1 U7692 ( .C1(n6730), .C2(n6734), .A(n6732), .B(n6729), .ZN(n6731)
         );
  OAI21_X1 U7693 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6732), .A(n6731), 
        .ZN(n6733) );
  OAI21_X1 U7694 ( .B1(n6735), .B2(n6734), .A(n6733), .ZN(U3461) );
  AOI21_X1 U7695 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7696 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6736), .B2(n6944), .ZN(n6737) );
  INV_X1 U7697 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7698 ( .A1(n6738), .A2(n6737), .B1(n6829), .B2(n6741), .ZN(U3468)
         );
  INV_X1 U7699 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6742) );
  NOR2_X1 U7700 ( .A1(n6741), .A2(REIP_REG_1__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U7701 ( .A1(n6742), .A2(n6741), .B1(n6740), .B2(n6739), .ZN(U3469)
         );
  MUX2_X1 U7702 ( .A(n6803), .B(W_R_N_REG_SCAN_IN), .S(n6743), .Z(U3470) );
  MUX2_X1 U7703 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6743), .Z(U3473) );
  AOI222_X1 U7704 ( .A1(n6746), .A2(DATAO_REG_10__SCAN_IN), .B1(n6745), .B2(
        EAX_REG_10__SCAN_IN), .C1(n6744), .C2(LWORD_REG_10__SCAN_IN), .ZN(
        n7045) );
  INV_X1 U7705 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6885) );
  NAND4_X1 U7706 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(
        INSTQUEUE_REG_11__2__SCAN_IN), .A3(INSTQUEUE_REG_10__2__SCAN_IN), .A4(
        n6885), .ZN(n6767) );
  INV_X1 U7707 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n7010) );
  INV_X1 U7708 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6810) );
  NAND4_X1 U7709 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(
        INSTQUEUE_REG_15__6__SCAN_IN), .A3(n7010), .A4(n6810), .ZN(n6766) );
  NAND4_X1 U7710 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(
        INSTQUEUE_REG_12__3__SCAN_IN), .A3(LWORD_REG_12__SCAN_IN), .A4(n3650), 
        .ZN(n6747) );
  NOR3_X1 U7711 ( .A1(DATAO_REG_19__SCAN_IN), .A2(n6998), .A3(n6747), .ZN(
        n6753) );
  NAND4_X1 U7712 ( .A1(DATAI_6_), .A2(n6975), .A3(n6974), .A4(n6979), .ZN(
        n6751) );
  INV_X1 U7713 ( .A(DATAI_30_), .ZN(n6995) );
  NAND4_X1 U7714 ( .A1(EAX_REG_3__SCAN_IN), .A2(DATAI_8_), .A3(
        DATAWIDTH_REG_29__SCAN_IN), .A4(n6995), .ZN(n6750) );
  NAND4_X1 U7715 ( .A1(EAX_REG_5__SCAN_IN), .A2(DATAI_17_), .A3(n7004), .A4(
        n5502), .ZN(n6749) );
  NAND4_X1 U7716 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(EBX_REG_20__SCAN_IN), .A3(UWORD_REG_13__SCAN_IN), .A4(n7028), .ZN(n6748) );
  NOR4_X1 U7717 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6752)
         );
  INV_X1 U7718 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n7022) );
  NAND4_X1 U7719 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6753), .A3(n6752), 
        .A4(n7022), .ZN(n6765) );
  NAND4_X1 U7720 ( .A1(DATAO_REG_5__SCAN_IN), .A2(DATAO_REG_22__SCAN_IN), .A3(
        n3942), .A4(n6809), .ZN(n6754) );
  NOR3_X1 U7721 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(READREQUEST_REG_SCAN_IN), 
        .A3(n6754), .ZN(n6763) );
  NAND4_X1 U7722 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        REIP_REG_25__SCAN_IN), .A3(ADS_N_REG_SCAN_IN), .A4(n6919), .ZN(n6761)
         );
  NAND4_X1 U7723 ( .A1(DATAO_REG_26__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), 
        .A3(n7012), .A4(n6932), .ZN(n6760) );
  NOR4_X1 U7724 ( .A1(DATAI_28_), .A2(DATAI_9_), .A3(DATAO_REG_25__SCAN_IN), 
        .A4(n6964), .ZN(n6758) );
  NOR4_X1 U7725 ( .A1(ADDRESS_REG_12__SCAN_IN), .A2(BS16_N), .A3(
        DATAO_REG_2__SCAN_IN), .A4(n6925), .ZN(n6757) );
  NOR4_X1 U7726 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(ADDRESS_REG_17__SCAN_IN), .A4(ADDRESS_REG_16__SCAN_IN), .ZN(n6756) );
  NOR4_X1 U7727 ( .A1(EBX_REG_30__SCAN_IN), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .A3(EAX_REG_21__SCAN_IN), .A4(DATAO_REG_7__SCAN_IN), .ZN(n6755) );
  NAND4_X1 U7728 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6759)
         );
  NOR3_X1 U7729 ( .A1(n6761), .A2(n6760), .A3(n6759), .ZN(n6762) );
  NAND4_X1 U7730 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6763), .A3(n6762), .A4(
        n6801), .ZN(n6764) );
  NOR4_X1 U7731 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6791)
         );
  NOR4_X1 U7732 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUE_REG_7__4__SCAN_IN), .A3(INSTQUEUE_REG_2__4__SCAN_IN), .A4(
        INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6768) );
  NAND4_X1 U7733 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6980), .A3(
        INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n6768), .ZN(n6789) );
  INV_X1 U7734 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6769) );
  NAND4_X1 U7735 ( .A1(n6769), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .A3(
        INSTQUEUE_REG_3__0__SCAN_IN), .A4(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n6770) );
  NOR3_X1 U7736 ( .A1(n6770), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .A3(
        INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6777) );
  INV_X1 U7737 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6934) );
  NAND4_X1 U7738 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(
        INSTQUEUE_REG_12__1__SCAN_IN), .A3(INSTQUEUE_REG_10__1__SCAN_IN), .A4(
        n6934), .ZN(n6775) );
  INV_X1 U7739 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6774) );
  INV_X1 U7740 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6890) );
  INV_X1 U7741 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6938) );
  AND4_X1 U7742 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(
        INSTQUEUE_REG_10__5__SCAN_IN), .A3(INSTQUEUE_REG_1__7__SCAN_IN), .A4(
        INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6771) );
  NAND4_X1 U7743 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n6890), .A3(n6938), 
        .A4(n6771), .ZN(n6773) );
  OR4_X1 U7744 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6888), .A3(
        INSTQUEUE_REG_0__1__SCAN_IN), .A4(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n6772) );
  NOR4_X1 U7745 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6776)
         );
  INV_X1 U7746 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6826) );
  NAND4_X1 U7747 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n6777), .A3(n6776), 
        .A4(n6826), .ZN(n6788) );
  NAND4_X1 U7748 ( .A1(UWORD_REG_6__SCAN_IN), .A2(ADDRESS_REG_9__SCAN_IN), 
        .A3(n6878), .A4(n6873), .ZN(n6781) );
  INV_X1 U7749 ( .A(DATAI_13_), .ZN(n6860) );
  NAND4_X1 U7750 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(NA_N), .A3(n6863), .A4(
        n6860), .ZN(n6780) );
  NAND4_X1 U7751 ( .A1(EBX_REG_29__SCAN_IN), .A2(EBX_REG_16__SCAN_IN), .A3(
        PHYADDRPOINTER_REG_6__SCAN_IN), .A4(LWORD_REG_6__SCAN_IN), .ZN(n6779)
         );
  NAND4_X1 U7752 ( .A1(EAX_REG_25__SCAN_IN), .A2(EBX_REG_26__SCAN_IN), .A3(
        LWORD_REG_14__SCAN_IN), .A4(n6877), .ZN(n6778) );
  OR4_X1 U7753 ( .A1(n6781), .A2(n6780), .A3(n6779), .A4(n6778), .ZN(n6787) );
  NOR4_X1 U7754 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6830), .A3(n6823), .A4(
        n6829), .ZN(n6785) );
  INV_X1 U7755 ( .A(DATAI_20_), .ZN(n6813) );
  NOR4_X1 U7756 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .A3(ADDRESS_REG_7__SCAN_IN), .A4(n6813), .ZN(n6784) );
  NOR4_X1 U7757 ( .A1(EBX_REG_27__SCAN_IN), .A2(EBX_REG_8__SCAN_IN), .A3(
        EAX_REG_18__SCAN_IN), .A4(BE_N_REG_1__SCAN_IN), .ZN(n6783) );
  NOR4_X1 U7758 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        REIP_REG_17__SCAN_IN), .A3(ADDRESS_REG_6__SCAN_IN), .A4(n6842), .ZN(
        n6782) );
  NAND4_X1 U7759 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6786)
         );
  NOR4_X1 U7760 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6790)
         );
  AOI21_X1 U7761 ( .B1(n6791), .B2(n6790), .A(keyinput29), .ZN(n7043) );
  INV_X1 U7762 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6793) );
  AOI22_X1 U7763 ( .A1(n6794), .A2(keyinput64), .B1(n6793), .B2(keyinput39), 
        .ZN(n6792) );
  OAI221_X1 U7764 ( .B1(n6794), .B2(keyinput64), .C1(n6793), .C2(keyinput39), 
        .A(n6792), .ZN(n6798) );
  XNOR2_X1 U7765 ( .A(n6795), .B(keyinput59), .ZN(n6797) );
  XOR2_X1 U7766 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .B(keyinput95), .Z(n6796)
         );
  OR3_X1 U7767 ( .A1(n6798), .A2(n6797), .A3(n6796), .ZN(n6806) );
  AOI22_X1 U7768 ( .A1(n6801), .A2(keyinput26), .B1(keyinput31), .B2(n6800), 
        .ZN(n6799) );
  OAI221_X1 U7769 ( .B1(n6801), .B2(keyinput26), .C1(n6800), .C2(keyinput31), 
        .A(n6799), .ZN(n6805) );
  AOI22_X1 U7770 ( .A1(n6803), .A2(keyinput90), .B1(keyinput100), .B2(n4542), 
        .ZN(n6802) );
  OAI221_X1 U7771 ( .B1(n6803), .B2(keyinput90), .C1(n4542), .C2(keyinput100), 
        .A(n6802), .ZN(n6804) );
  NOR3_X1 U7772 ( .A1(n6806), .A2(n6805), .A3(n6804), .ZN(n6853) );
  AOI22_X1 U7773 ( .A1(n4570), .A2(keyinput53), .B1(n3942), .B2(keyinput9), 
        .ZN(n6807) );
  OAI221_X1 U7774 ( .B1(n4570), .B2(keyinput53), .C1(n3942), .C2(keyinput9), 
        .A(n6807), .ZN(n6818) );
  AOI22_X1 U7775 ( .A1(n6810), .A2(keyinput92), .B1(keyinput67), .B2(n6809), 
        .ZN(n6808) );
  OAI221_X1 U7776 ( .B1(n6810), .B2(keyinput92), .C1(n6809), .C2(keyinput67), 
        .A(n6808), .ZN(n6817) );
  AOI22_X1 U7777 ( .A1(n4841), .A2(keyinput81), .B1(keyinput33), .B2(n6774), 
        .ZN(n6811) );
  OAI221_X1 U7778 ( .B1(n4841), .B2(keyinput81), .C1(n6774), .C2(keyinput33), 
        .A(n6811), .ZN(n6816) );
  AOI22_X1 U7779 ( .A1(n6814), .A2(keyinput51), .B1(keyinput10), .B2(n6813), 
        .ZN(n6812) );
  OAI221_X1 U7780 ( .B1(n6814), .B2(keyinput51), .C1(n6813), .C2(keyinput10), 
        .A(n6812), .ZN(n6815) );
  NOR4_X1 U7781 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n6852)
         );
  INV_X1 U7782 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U7783 ( .A1(n6821), .A2(keyinput87), .B1(n6820), .B2(keyinput57), 
        .ZN(n6819) );
  OAI221_X1 U7784 ( .B1(n6821), .B2(keyinput87), .C1(n6820), .C2(keyinput57), 
        .A(n6819), .ZN(n6834) );
  AOI22_X1 U7785 ( .A1(n6824), .A2(keyinput94), .B1(n6823), .B2(keyinput71), 
        .ZN(n6822) );
  OAI221_X1 U7786 ( .B1(n6824), .B2(keyinput94), .C1(n6823), .C2(keyinput71), 
        .A(n6822), .ZN(n6833) );
  AOI22_X1 U7787 ( .A1(n6827), .A2(keyinput15), .B1(n6826), .B2(keyinput85), 
        .ZN(n6825) );
  OAI221_X1 U7788 ( .B1(n6827), .B2(keyinput15), .C1(n6826), .C2(keyinput85), 
        .A(n6825), .ZN(n6832) );
  AOI22_X1 U7789 ( .A1(n6830), .A2(keyinput78), .B1(keyinput84), .B2(n6829), 
        .ZN(n6828) );
  OAI221_X1 U7790 ( .B1(n6830), .B2(keyinput78), .C1(n6829), .C2(keyinput84), 
        .A(n6828), .ZN(n6831) );
  NOR4_X1 U7791 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .ZN(n6851)
         );
  AOI22_X1 U7792 ( .A1(n6837), .A2(keyinput38), .B1(keyinput97), .B2(n6836), 
        .ZN(n6835) );
  OAI221_X1 U7793 ( .B1(n6837), .B2(keyinput38), .C1(n6836), .C2(keyinput97), 
        .A(n6835), .ZN(n6849) );
  INV_X1 U7794 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U7795 ( .A1(n6840), .A2(keyinput24), .B1(n6839), .B2(keyinput13), 
        .ZN(n6838) );
  OAI221_X1 U7796 ( .B1(n6840), .B2(keyinput24), .C1(n6839), .C2(keyinput13), 
        .A(n6838), .ZN(n6848) );
  AOI22_X1 U7797 ( .A1(n5380), .A2(keyinput120), .B1(keyinput60), .B2(n6842), 
        .ZN(n6841) );
  OAI221_X1 U7798 ( .B1(n5380), .B2(keyinput120), .C1(n6842), .C2(keyinput60), 
        .A(n6841), .ZN(n6847) );
  AOI22_X1 U7799 ( .A1(n6845), .A2(keyinput32), .B1(n6844), .B2(keyinput112), 
        .ZN(n6843) );
  OAI221_X1 U7800 ( .B1(n6845), .B2(keyinput32), .C1(n6844), .C2(keyinput112), 
        .A(n6843), .ZN(n6846) );
  NOR4_X1 U7801 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6850)
         );
  NAND4_X1 U7802 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n7041)
         );
  AOI22_X1 U7803 ( .A1(n5110), .A2(keyinput74), .B1(keyinput30), .B2(n6855), 
        .ZN(n6854) );
  OAI221_X1 U7804 ( .B1(n5110), .B2(keyinput74), .C1(n6855), .C2(keyinput30), 
        .A(n6854), .ZN(n6867) );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6858) );
  INV_X1 U7806 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n6857) );
  AOI22_X1 U7807 ( .A1(n6858), .A2(keyinput19), .B1(keyinput34), .B2(n6857), 
        .ZN(n6856) );
  OAI221_X1 U7808 ( .B1(n6858), .B2(keyinput19), .C1(n6857), .C2(keyinput34), 
        .A(n6856), .ZN(n6866) );
  AOI22_X1 U7809 ( .A1(n4131), .A2(keyinput63), .B1(keyinput127), .B2(n6860), 
        .ZN(n6859) );
  OAI221_X1 U7810 ( .B1(n4131), .B2(keyinput63), .C1(n6860), .C2(keyinput127), 
        .A(n6859), .ZN(n6865) );
  AOI22_X1 U7811 ( .A1(n6863), .A2(keyinput61), .B1(keyinput52), .B2(n6862), 
        .ZN(n6861) );
  OAI221_X1 U7812 ( .B1(n6863), .B2(keyinput61), .C1(n6862), .C2(keyinput52), 
        .A(n6861), .ZN(n6864) );
  NOR4_X1 U7813 ( .A1(n6867), .A2(n6866), .A3(n6865), .A4(n6864), .ZN(n6914)
         );
  AOI22_X1 U7814 ( .A1(n6870), .A2(keyinput126), .B1(keyinput5), .B2(n6869), 
        .ZN(n6868) );
  OAI221_X1 U7815 ( .B1(n6870), .B2(keyinput126), .C1(n6869), .C2(keyinput5), 
        .A(n6868), .ZN(n6882) );
  INV_X1 U7816 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6872) );
  AOI22_X1 U7817 ( .A1(n6873), .A2(keyinput82), .B1(n6872), .B2(keyinput56), 
        .ZN(n6871) );
  OAI221_X1 U7818 ( .B1(n6873), .B2(keyinput82), .C1(n6872), .C2(keyinput56), 
        .A(n6871), .ZN(n6881) );
  INV_X1 U7819 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6875) );
  AOI22_X1 U7820 ( .A1(n4573), .A2(keyinput119), .B1(n6875), .B2(keyinput11), 
        .ZN(n6874) );
  OAI221_X1 U7821 ( .B1(n4573), .B2(keyinput119), .C1(n6875), .C2(keyinput11), 
        .A(n6874), .ZN(n6880) );
  AOI22_X1 U7822 ( .A1(n6878), .A2(keyinput50), .B1(keyinput105), .B2(n6877), 
        .ZN(n6876) );
  OAI221_X1 U7823 ( .B1(n6878), .B2(keyinput50), .C1(n6877), .C2(keyinput105), 
        .A(n6876), .ZN(n6879) );
  NOR4_X1 U7824 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n6913)
         );
  AOI22_X1 U7825 ( .A1(n6885), .A2(keyinput109), .B1(keyinput22), .B2(n6884), 
        .ZN(n6883) );
  OAI221_X1 U7826 ( .B1(n6885), .B2(keyinput109), .C1(n6884), .C2(keyinput22), 
        .A(n6883), .ZN(n6897) );
  AOI22_X1 U7827 ( .A1(n6888), .A2(keyinput6), .B1(keyinput118), .B2(n6887), 
        .ZN(n6886) );
  OAI221_X1 U7828 ( .B1(n6888), .B2(keyinput6), .C1(n6887), .C2(keyinput118), 
        .A(n6886), .ZN(n6896) );
  AOI22_X1 U7829 ( .A1(n5106), .A2(keyinput8), .B1(keyinput66), .B2(n6890), 
        .ZN(n6889) );
  OAI221_X1 U7830 ( .B1(n5106), .B2(keyinput8), .C1(n6890), .C2(keyinput66), 
        .A(n6889), .ZN(n6895) );
  INV_X1 U7831 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6893) );
  AOI22_X1 U7832 ( .A1(n6893), .A2(keyinput93), .B1(n6892), .B2(keyinput49), 
        .ZN(n6891) );
  OAI221_X1 U7833 ( .B1(n6893), .B2(keyinput93), .C1(n6892), .C2(keyinput49), 
        .A(n6891), .ZN(n6894) );
  NOR4_X1 U7834 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6912)
         );
  AOI22_X1 U7835 ( .A1(n6899), .A2(keyinput98), .B1(keyinput16), .B2(n4551), 
        .ZN(n6898) );
  OAI221_X1 U7836 ( .B1(n6899), .B2(keyinput98), .C1(n4551), .C2(keyinput16), 
        .A(n6898), .ZN(n6910) );
  INV_X1 U7837 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6901) );
  AOI22_X1 U7838 ( .A1(n6902), .A2(keyinput103), .B1(n6901), .B2(keyinput101), 
        .ZN(n6900) );
  OAI221_X1 U7839 ( .B1(n6902), .B2(keyinput103), .C1(n6901), .C2(keyinput101), 
        .A(n6900), .ZN(n6909) );
  INV_X1 U7840 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6903) );
  XOR2_X1 U7841 ( .A(n6903), .B(keyinput68), .Z(n6907) );
  XNOR2_X1 U7842 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .B(keyinput99), .ZN(n6906)
         );
  XNOR2_X1 U7843 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .B(keyinput27), .ZN(n6905) );
  XNOR2_X1 U7844 ( .A(EBX_REG_29__SCAN_IN), .B(keyinput14), .ZN(n6904) );
  NAND4_X1 U7845 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6908)
         );
  NOR3_X1 U7846 ( .A1(n6910), .A2(n6909), .A3(n6908), .ZN(n6911) );
  NAND4_X1 U7847 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n7040)
         );
  INV_X1 U7848 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6916) );
  AOI22_X1 U7849 ( .A1(n6917), .A2(keyinput88), .B1(n6916), .B2(keyinput116), 
        .ZN(n6915) );
  OAI221_X1 U7850 ( .B1(n6917), .B2(keyinput88), .C1(n6916), .C2(keyinput116), 
        .A(n6915), .ZN(n6929) );
  AOI22_X1 U7851 ( .A1(n6919), .A2(keyinput3), .B1(n5159), .B2(keyinput114), 
        .ZN(n6918) );
  OAI221_X1 U7852 ( .B1(n6919), .B2(keyinput3), .C1(n5159), .C2(keyinput114), 
        .A(n6918), .ZN(n6928) );
  INV_X1 U7853 ( .A(BS16_N), .ZN(n6922) );
  AOI22_X1 U7854 ( .A1(n6922), .A2(keyinput40), .B1(keyinput17), .B2(n6921), 
        .ZN(n6920) );
  OAI221_X1 U7855 ( .B1(n6922), .B2(keyinput40), .C1(n6921), .C2(keyinput17), 
        .A(n6920), .ZN(n6927) );
  INV_X1 U7856 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6924) );
  AOI22_X1 U7857 ( .A1(n6925), .A2(keyinput89), .B1(n6924), .B2(keyinput76), 
        .ZN(n6923) );
  OAI221_X1 U7858 ( .B1(n6925), .B2(keyinput89), .C1(n6924), .C2(keyinput76), 
        .A(n6923), .ZN(n6926) );
  NOR4_X1 U7859 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6972)
         );
  INV_X1 U7860 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U7861 ( .A1(n6932), .A2(keyinput123), .B1(n6931), .B2(keyinput43), 
        .ZN(n6930) );
  OAI221_X1 U7862 ( .B1(n6932), .B2(keyinput123), .C1(n6931), .C2(keyinput43), 
        .A(n6930), .ZN(n6942) );
  AOI22_X1 U7863 ( .A1(n4546), .A2(keyinput124), .B1(n6934), .B2(keyinput28), 
        .ZN(n6933) );
  OAI221_X1 U7864 ( .B1(n4546), .B2(keyinput124), .C1(n6934), .C2(keyinput28), 
        .A(n6933), .ZN(n6941) );
  AOI22_X1 U7865 ( .A1(n6936), .A2(keyinput69), .B1(n6769), .B2(keyinput111), 
        .ZN(n6935) );
  OAI221_X1 U7866 ( .B1(n6936), .B2(keyinput69), .C1(n6769), .C2(keyinput111), 
        .A(n6935), .ZN(n6940) );
  AOI22_X1 U7867 ( .A1(n6938), .A2(keyinput7), .B1(keyinput55), .B2(n4437), 
        .ZN(n6937) );
  OAI221_X1 U7868 ( .B1(n6938), .B2(keyinput7), .C1(n4437), .C2(keyinput55), 
        .A(n6937), .ZN(n6939) );
  NOR4_X1 U7869 ( .A1(n6942), .A2(n6941), .A3(n6940), .A4(n6939), .ZN(n6971)
         );
  INV_X1 U7870 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7871 ( .A1(n6945), .A2(keyinput20), .B1(keyinput121), .B2(n6944), 
        .ZN(n6943) );
  OAI221_X1 U7872 ( .B1(n6945), .B2(keyinput20), .C1(n6944), .C2(keyinput121), 
        .A(n6943), .ZN(n6955) );
  INV_X1 U7873 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6948) );
  INV_X1 U7874 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6947) );
  AOI22_X1 U7875 ( .A1(n6948), .A2(keyinput72), .B1(keyinput2), .B2(n6947), 
        .ZN(n6946) );
  OAI221_X1 U7876 ( .B1(n6948), .B2(keyinput72), .C1(n6947), .C2(keyinput2), 
        .A(n6946), .ZN(n6954) );
  AOI22_X1 U7877 ( .A1(n5441), .A2(keyinput104), .B1(n5769), .B2(keyinput25), 
        .ZN(n6949) );
  OAI221_X1 U7878 ( .B1(n5441), .B2(keyinput104), .C1(n5769), .C2(keyinput25), 
        .A(n6949), .ZN(n6953) );
  XNOR2_X1 U7879 ( .A(EBX_REG_30__SCAN_IN), .B(keyinput110), .ZN(n6951) );
  XNOR2_X1 U7880 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput107), .ZN(n6950) );
  NAND2_X1 U7881 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  NOR4_X1 U7882 ( .A1(n6955), .A2(n6954), .A3(n6953), .A4(n6952), .ZN(n6970)
         );
  INV_X1 U7883 ( .A(DATAI_28_), .ZN(n6957) );
  AOI22_X1 U7884 ( .A1(n4548), .A2(keyinput102), .B1(n6957), .B2(keyinput70), 
        .ZN(n6956) );
  OAI221_X1 U7885 ( .B1(n4548), .B2(keyinput102), .C1(n6957), .C2(keyinput70), 
        .A(n6956), .ZN(n6968) );
  AOI22_X1 U7886 ( .A1(n4544), .A2(keyinput83), .B1(n6959), .B2(keyinput125), 
        .ZN(n6958) );
  OAI221_X1 U7887 ( .B1(n4544), .B2(keyinput83), .C1(n6959), .C2(keyinput125), 
        .A(n6958), .ZN(n6967) );
  INV_X1 U7888 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6961) );
  AOI22_X1 U7889 ( .A1(n4538), .A2(keyinput117), .B1(n6961), .B2(keyinput113), 
        .ZN(n6960) );
  OAI221_X1 U7890 ( .B1(n4538), .B2(keyinput117), .C1(n6961), .C2(keyinput113), 
        .A(n6960), .ZN(n6966) );
  INV_X1 U7891 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6963) );
  AOI22_X1 U7892 ( .A1(n6964), .A2(keyinput108), .B1(n6963), .B2(keyinput122), 
        .ZN(n6962) );
  OAI221_X1 U7893 ( .B1(n6964), .B2(keyinput108), .C1(n6963), .C2(keyinput122), 
        .A(n6962), .ZN(n6965) );
  NOR4_X1 U7894 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n6969)
         );
  NAND4_X1 U7895 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n7039)
         );
  AOI22_X1 U7896 ( .A1(n6975), .A2(keyinput23), .B1(keyinput96), .B2(n6974), 
        .ZN(n6973) );
  OAI221_X1 U7897 ( .B1(n6975), .B2(keyinput23), .C1(n6974), .C2(keyinput96), 
        .A(n6973), .ZN(n6988) );
  AOI22_X1 U7898 ( .A1(n6978), .A2(keyinput65), .B1(n6977), .B2(keyinput77), 
        .ZN(n6976) );
  OAI221_X1 U7899 ( .B1(n6978), .B2(keyinput65), .C1(n6977), .C2(keyinput77), 
        .A(n6976), .ZN(n6987) );
  XOR2_X1 U7900 ( .A(n6979), .B(keyinput45), .Z(n6983) );
  XNOR2_X1 U7901 ( .A(n6980), .B(keyinput86), .ZN(n6982) );
  XNOR2_X1 U7902 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput44), .ZN(n6981)
         );
  NAND3_X1 U7903 ( .A1(n6983), .A2(n6982), .A3(n6981), .ZN(n6986) );
  XNOR2_X1 U7904 ( .A(n6984), .B(keyinput41), .ZN(n6985) );
  NOR4_X1 U7905 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n7037)
         );
  INV_X1 U7906 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U7907 ( .A1(n6990), .A2(keyinput18), .ZN(n6989) );
  OAI221_X1 U7908 ( .B1(n6991), .B2(keyinput29), .C1(n6990), .C2(keyinput18), 
        .A(n6989), .ZN(n7002) );
  INV_X1 U7909 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6993) );
  AOI22_X1 U7910 ( .A1(n3650), .A2(keyinput37), .B1(n6993), .B2(keyinput42), 
        .ZN(n6992) );
  OAI221_X1 U7911 ( .B1(n3650), .B2(keyinput37), .C1(n6993), .C2(keyinput42), 
        .A(n6992), .ZN(n7001) );
  INV_X1 U7912 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U7913 ( .A1(n6996), .A2(keyinput79), .B1(keyinput54), .B2(n6995), 
        .ZN(n6994) );
  OAI221_X1 U7914 ( .B1(n6996), .B2(keyinput79), .C1(n6995), .C2(keyinput54), 
        .A(n6994), .ZN(n7000) );
  AOI22_X1 U7915 ( .A1(n6998), .A2(keyinput115), .B1(keyinput47), .B2(n4540), 
        .ZN(n6997) );
  OAI221_X1 U7916 ( .B1(n6998), .B2(keyinput115), .C1(n4540), .C2(keyinput47), 
        .A(n6997), .ZN(n6999) );
  NOR4_X1 U7917 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .ZN(n7036)
         );
  AOI22_X1 U7918 ( .A1(n5502), .A2(keyinput62), .B1(keyinput58), .B2(n7004), 
        .ZN(n7003) );
  OAI221_X1 U7919 ( .B1(n5502), .B2(keyinput62), .C1(n7004), .C2(keyinput58), 
        .A(n7003), .ZN(n7017) );
  INV_X1 U7920 ( .A(DATAI_17_), .ZN(n7007) );
  AOI22_X1 U7921 ( .A1(n7007), .A2(keyinput46), .B1(n7006), .B2(keyinput75), 
        .ZN(n7005) );
  OAI221_X1 U7922 ( .B1(n7007), .B2(keyinput46), .C1(n7006), .C2(keyinput75), 
        .A(n7005), .ZN(n7016) );
  AOI22_X1 U7923 ( .A1(n7010), .A2(keyinput12), .B1(keyinput91), .B2(n7009), 
        .ZN(n7008) );
  OAI221_X1 U7924 ( .B1(n7010), .B2(keyinput12), .C1(n7009), .C2(keyinput91), 
        .A(n7008), .ZN(n7015) );
  AOI22_X1 U7925 ( .A1(n7013), .A2(keyinput21), .B1(keyinput80), .B2(n7012), 
        .ZN(n7011) );
  OAI221_X1 U7926 ( .B1(n7013), .B2(keyinput21), .C1(n7012), .C2(keyinput80), 
        .A(n7011), .ZN(n7014) );
  NOR4_X1 U7927 ( .A1(n7017), .A2(n7016), .A3(n7015), .A4(n7014), .ZN(n7035)
         );
  INV_X1 U7928 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n7020) );
  AOI22_X1 U7929 ( .A1(n7020), .A2(keyinput0), .B1(keyinput48), .B2(n7019), 
        .ZN(n7018) );
  OAI221_X1 U7930 ( .B1(n7020), .B2(keyinput0), .C1(n7019), .C2(keyinput48), 
        .A(n7018), .ZN(n7033) );
  AOI22_X1 U7931 ( .A1(n7023), .A2(keyinput4), .B1(n7022), .B2(keyinput35), 
        .ZN(n7021) );
  OAI221_X1 U7932 ( .B1(n7023), .B2(keyinput4), .C1(n7022), .C2(keyinput35), 
        .A(n7021), .ZN(n7032) );
  INV_X1 U7933 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n7025) );
  AOI22_X1 U7934 ( .A1(n7026), .A2(keyinput106), .B1(n7025), .B2(keyinput36), 
        .ZN(n7024) );
  OAI221_X1 U7935 ( .B1(n7026), .B2(keyinput106), .C1(n7025), .C2(keyinput36), 
        .A(n7024), .ZN(n7031) );
  AOI22_X1 U7936 ( .A1(n7029), .A2(keyinput73), .B1(keyinput1), .B2(n7028), 
        .ZN(n7027) );
  OAI221_X1 U7937 ( .B1(n7029), .B2(keyinput73), .C1(n7028), .C2(keyinput1), 
        .A(n7027), .ZN(n7030) );
  NOR4_X1 U7938 ( .A1(n7033), .A2(n7032), .A3(n7031), .A4(n7030), .ZN(n7034)
         );
  NAND4_X1 U7939 ( .A1(n7037), .A2(n7036), .A3(n7035), .A4(n7034), .ZN(n7038)
         );
  NOR4_X1 U7940 ( .A1(n7041), .A2(n7040), .A3(n7039), .A4(n7038), .ZN(n7042)
         );
  OAI21_X1 U7941 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7043), .A(n7042), 
        .ZN(n7044) );
  XOR2_X1 U7942 ( .A(n7045), .B(n7044), .Z(U2913) );
  AND4_X1 U4377 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3318)
         );
  BUF_X1 U3611 ( .A(n3384), .Z(n3393) );
  CLKBUF_X1 U3532 ( .A(n4317), .Z(n4356) );
  CLKBUF_X2 U3538 ( .A(n3518), .Z(n3557) );
  INV_X1 U3544 ( .A(n3384), .ZN(n3896) );
  CLKBUF_X1 U3554 ( .A(n3894), .Z(n3895) );
  NAND2_X2 U3562 ( .A1(n4628), .A2(n3780), .ZN(n3787) );
  CLKBUF_X1 U4044 ( .A(n3671), .Z(n5832) );
  CLKBUF_X1 U4144 ( .A(n4701), .Z(n3087) );
  CLKBUF_X1 U4961 ( .A(n3787), .Z(n5214) );
endmodule

