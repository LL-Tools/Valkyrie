

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943;

  INV_X1 U2294 ( .A(n2260), .ZN(n2740) );
  CLKBUF_X2 U2297 ( .A(IR_REG_0__SCAN_IN), .Z(n2614) );
  INV_X1 U2298 ( .A(n3458), .ZN(n3440) );
  INV_X1 U2299 ( .A(n2259), .ZN(n2737) );
  NAND2_X1 U2300 ( .A1(n3484), .A2(n3387), .ZN(n3483) );
  OAI21_X2 U2301 ( .B1(n4019), .B2(n3856), .A(n3855), .ZN(n3955) );
  NOR2_X2 U2302 ( .A1(n2561), .A2(n2560), .ZN(n2566) );
  BUF_X4 U2303 ( .A(n2695), .Z(n2259) );
  NAND2_X1 U2304 ( .A1(n2599), .A2(n2597), .ZN(n2695) );
  AOI21_X2 U2305 ( .B1(n3483), .B2(n3402), .A(n3403), .ZN(n3533) );
  NAND2_X4 U2306 ( .A1(n2788), .A2(n2767), .ZN(n3401) );
  AND2_X1 U2307 ( .A1(n2600), .A2(n2599), .ZN(n3007) );
  OR2_X1 U2308 ( .A1(n3557), .A2(n3559), .ZN(n2499) );
  OAI21_X1 U2309 ( .B1(n3917), .B2(n3860), .A(n3859), .ZN(n3904) );
  NAND2_X1 U2310 ( .A1(n2456), .A2(n2457), .ZN(n3206) );
  NAND2_X1 U2311 ( .A1(n2321), .A2(n2325), .ZN(n2320) );
  NAND2_X1 U2312 ( .A1(n2933), .A2(n2686), .ZN(n4741) );
  INV_X4 U2313 ( .A(n3401), .ZN(n2263) );
  INV_X2 U2314 ( .A(n3401), .ZN(n3437) );
  INV_X2 U2315 ( .A(n2689), .ZN(n2788) );
  XNOR2_X1 U2316 ( .A(n2569), .B(n2568), .ZN(n2632) );
  NAND2_X1 U2317 ( .A1(n2643), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U2318 ( .A1(n2643), .A2(n2645), .ZN(n3808) );
  NAND2_X1 U2319 ( .A1(n2784), .A2(n2805), .ZN(n3615) );
  NAND2_X1 U2320 ( .A1(n2550), .A2(n2280), .ZN(n2561) );
  AOI21_X1 U2321 ( .B1(n2572), .B2(n2575), .A(n2954), .ZN(n2592) );
  AND3_X1 U2322 ( .A1(n2398), .A2(n2464), .A3(n2500), .ZN(n2572) );
  CLKBUF_X1 U2323 ( .A(n2903), .Z(n2905) );
  XNOR2_X1 U2324 ( .A(n2712), .B(IR_REG_2__SCAN_IN), .ZN(n4682) );
  NOR2_X2 U2325 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2607)
         );
  NOR2_X1 U2326 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2455)
         );
  AOI21_X2 U2327 ( .B1(n3522), .B2(n3524), .A(n3523), .ZN(n3552) );
  INV_X1 U2328 ( .A(n3401), .ZN(n2262) );
  NAND2_X1 U2329 ( .A1(n4668), .A2(n4663), .ZN(n2264) );
  AOI21_X1 U2330 ( .B1(n2474), .B2(n2470), .A(n3261), .ZN(n2469) );
  NOR2_X1 U2331 ( .A1(n2470), .A2(n3262), .ZN(n2472) );
  AND2_X1 U2332 ( .A1(n2449), .A2(n2301), .ZN(n2448) );
  OAI21_X1 U2333 ( .B1(n2414), .B2(n3743), .A(n2413), .ZN(n3745) );
  NAND2_X1 U2334 ( .A1(n2989), .A2(n2268), .ZN(n2414) );
  OAI21_X1 U2335 ( .B1(n3743), .B2(n2418), .A(n2417), .ZN(n2413) );
  INV_X1 U2336 ( .A(n3977), .ZN(n2369) );
  AOI21_X1 U2337 ( .B1(n2349), .B2(n4753), .A(n2296), .ZN(n2348) );
  INV_X1 U2338 ( .A(n4754), .ZN(n2349) );
  INV_X1 U2339 ( .A(IR_REG_25__SCAN_IN), .ZN(n2502) );
  AND2_X1 U2340 ( .A1(n3285), .A2(n3284), .ZN(n3511) );
  INV_X1 U2341 ( .A(n3993), .ZN(n3833) );
  INV_X1 U2342 ( .A(n2693), .ZN(n3464) );
  XNOR2_X1 U2343 ( .A(n2652), .B(n2420), .ZN(n2615) );
  XNOR2_X1 U2344 ( .A(n3754), .B(n2435), .ZN(n2971) );
  INV_X1 U2345 ( .A(n2436), .ZN(n3765) );
  OAI21_X1 U2346 ( .B1(n4594), .B2(n4593), .A(n2438), .ZN(n2436) );
  NAND2_X1 U2347 ( .A1(n4603), .A2(n3267), .ZN(n4602) );
  OAI21_X1 U2348 ( .B1(n4221), .B2(n3166), .A(n3165), .ZN(n4784) );
  NAND2_X1 U2349 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2577) );
  INV_X1 U2350 ( .A(n3170), .ZN(n2341) );
  INV_X1 U2351 ( .A(n2340), .ZN(n2339) );
  OAI21_X1 U2352 ( .B1(n3168), .B2(n2341), .A(n4134), .ZN(n2340) );
  INV_X1 U2353 ( .A(n3634), .ZN(n2326) );
  INV_X1 U2354 ( .A(n2646), .ZN(n2640) );
  INV_X1 U2355 ( .A(n2680), .ZN(n2682) );
  AND2_X1 U2356 ( .A1(n2375), .A2(n2288), .ZN(n2959) );
  OAI21_X1 U2357 ( .B1(n2411), .B2(n4582), .A(n2410), .ZN(n3748) );
  NAND2_X1 U2358 ( .A1(n3747), .A2(n2412), .ZN(n2411) );
  OAI21_X1 U2359 ( .B1(n3794), .B2(n2390), .A(n2386), .ZN(n2392) );
  AOI21_X1 U2360 ( .B1(n2389), .B2(n2388), .A(n2387), .ZN(n2386) );
  NOR2_X1 U2361 ( .A1(n2277), .A2(n2362), .ZN(n2361) );
  INV_X1 U2362 ( .A(n3839), .ZN(n2362) );
  AOI21_X1 U2363 ( .B1(n3830), .B2(n2369), .A(n2367), .ZN(n2366) );
  NOR2_X1 U2364 ( .A1(n3960), .A2(n3980), .ZN(n2367) );
  NAND2_X1 U2365 ( .A1(n4000), .A2(n3829), .ZN(n3830) );
  NOR2_X1 U2366 ( .A1(n2329), .A2(n3686), .ZN(n2328) );
  INV_X1 U2367 ( .A(n3852), .ZN(n2329) );
  AND2_X1 U2368 ( .A1(n2401), .A2(n4089), .ZN(n2400) );
  NAND2_X1 U2369 ( .A1(n2339), .A2(n2341), .ZN(n2337) );
  AND2_X1 U2370 ( .A1(n3877), .A2(n4852), .ZN(n2401) );
  AND2_X1 U2371 ( .A1(n3706), .A2(n3574), .ZN(n3643) );
  OR2_X1 U2372 ( .A1(n4850), .A2(n4123), .ZN(n3846) );
  OR2_X1 U2373 ( .A1(n3737), .A2(n3195), .ZN(n3648) );
  OR2_X1 U2374 ( .A1(n4225), .A2(n3175), .ZN(n3696) );
  AOI21_X1 U2375 ( .B1(n2325), .B2(n2324), .A(n2323), .ZN(n2322) );
  INV_X1 U2376 ( .A(n3631), .ZN(n2323) );
  INV_X1 U2377 ( .A(n3632), .ZN(n2324) );
  INV_X1 U2378 ( .A(n3626), .ZN(n2314) );
  INV_X1 U2379 ( .A(n3639), .ZN(n2312) );
  INV_X1 U2380 ( .A(IR_REG_26__SCAN_IN), .ZN(n2575) );
  AND2_X1 U2381 ( .A1(n2275), .A2(n2555), .ZN(n2500) );
  NOR2_X1 U2382 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2528)
         );
  NAND2_X1 U2383 ( .A1(n2535), .A2(IR_REG_31__SCAN_IN), .ZN(n2538) );
  INV_X1 U2384 ( .A(IR_REG_22__SCAN_IN), .ZN(n2555) );
  NOR2_X1 U2385 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2949)
         );
  NOR2_X1 U2386 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2518)
         );
  NOR2_X1 U2387 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2519)
         );
  INV_X1 U2388 ( .A(IR_REG_5__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U2389 ( .A1(n3238), .A2(n3237), .ZN(n2484) );
  AND2_X1 U2390 ( .A1(n3092), .A2(n3091), .ZN(n3089) );
  INV_X1 U2391 ( .A(n2497), .ZN(n2496) );
  INV_X1 U2392 ( .A(n2290), .ZN(n2493) );
  AOI21_X1 U2393 ( .B1(n2497), .B2(n3559), .A(n2495), .ZN(n2494) );
  INV_X1 U2394 ( .A(n3447), .ZN(n2495) );
  NOR2_X1 U2395 ( .A1(n2467), .A2(n2298), .ZN(n2465) );
  NOR2_X1 U2396 ( .A1(n4838), .A2(n3511), .ZN(n3286) );
  XNOR2_X1 U2397 ( .A(n2735), .B(n3458), .ZN(n2750) );
  OAI21_X1 U2398 ( .B1(n3495), .B2(n2461), .A(n2460), .ZN(n2459) );
  NAND2_X1 U2399 ( .A1(n3368), .A2(n3335), .ZN(n2461) );
  AOI21_X1 U2400 ( .B1(n2284), .B2(n3368), .A(n3367), .ZN(n2460) );
  NAND2_X1 U2401 ( .A1(n3116), .A2(n3118), .ZN(n3119) );
  NAND2_X1 U2402 ( .A1(n2567), .A2(n2524), .ZN(n2643) );
  INV_X1 U2403 ( .A(n2644), .ZN(n2567) );
  OR2_X1 U2404 ( .A1(n3451), .A2(n3912), .ZN(n3434) );
  OR2_X1 U2405 ( .A1(n2740), .A2(n2723), .ZN(n2724) );
  OR2_X1 U2406 ( .A1(n2693), .A2(n2617), .ZN(n2651) );
  NAND2_X1 U2407 ( .A1(n2614), .A2(n2282), .ZN(n2378) );
  OR2_X1 U2408 ( .A1(n4629), .A2(n4628), .ZN(n2375) );
  NOR2_X1 U2409 ( .A1(n2652), .A2(n2420), .ZN(n2419) );
  XNOR2_X1 U2410 ( .A(n2959), .B(n4694), .ZN(n4510) );
  NOR2_X1 U2411 ( .A1(n2722), .A2(n4510), .ZN(n4509) );
  NOR2_X1 U2412 ( .A1(n4513), .A2(n2978), .ZN(n2979) );
  INV_X1 U2413 ( .A(n4519), .ZN(n2450) );
  OR2_X1 U2414 ( .A1(n4652), .A2(n2452), .ZN(n2451) );
  OR2_X1 U2415 ( .A1(n4519), .A2(n2738), .ZN(n2452) );
  OAI21_X1 U2416 ( .B1(n4720), .B2(n4541), .A(n2964), .ZN(n2968) );
  NAND2_X1 U2417 ( .A1(n2509), .A2(n4720), .ZN(n2434) );
  NAND2_X1 U2418 ( .A1(n4564), .A2(n2970), .ZN(n3754) );
  NAND2_X1 U2419 ( .A1(n2971), .A2(REG2_REG_10__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U2420 ( .A1(n2393), .A2(n2394), .ZN(n3792) );
  AOI21_X1 U2421 ( .B1(n3765), .B2(n2395), .A(n2306), .ZN(n2394) );
  NAND2_X1 U2422 ( .A1(n4602), .A2(n3786), .ZN(n3800) );
  INV_X1 U2423 ( .A(n2428), .ZN(n2373) );
  NOR2_X1 U2424 ( .A1(n3903), .A2(n3862), .ZN(n3887) );
  AND4_X1 U2425 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3888)
         );
  NAND2_X1 U2426 ( .A1(n3938), .A2(n3838), .ZN(n3839) );
  INV_X1 U2427 ( .A(n3861), .ZN(n3905) );
  NAND2_X1 U2428 ( .A1(n3391), .A2(REG3_REG_24__SCAN_IN), .ZN(n3405) );
  AOI21_X1 U2429 ( .B1(n3834), .B2(n3832), .A(n2513), .ZN(n3941) );
  AOI21_X1 U2430 ( .B1(n4043), .B2(n3825), .A(n3824), .ZN(n4032) );
  NOR2_X1 U2431 ( .A1(n4074), .A2(n4057), .ZN(n4056) );
  INV_X1 U2432 ( .A(n2354), .ZN(n2353) );
  AOI21_X1 U2433 ( .B1(n2354), .B2(n2352), .A(n2294), .ZN(n2351) );
  AOI21_X1 U2434 ( .B1(n4118), .B2(n3820), .A(n2295), .ZN(n2354) );
  AOI21_X1 U2435 ( .B1(n2348), .B2(n2350), .A(n2267), .ZN(n2347) );
  INV_X1 U2436 ( .A(n4862), .ZN(n4737) );
  AND2_X1 U2437 ( .A1(n2793), .A2(n3721), .ZN(n4663) );
  NAND2_X1 U2438 ( .A1(n3874), .A2(n3873), .ZN(n4157) );
  AND2_X1 U2439 ( .A1(n3872), .A2(n3871), .ZN(n3873) );
  NAND2_X1 U2440 ( .A1(n3866), .A2(n4731), .ZN(n3874) );
  NAND2_X1 U2441 ( .A1(n4668), .A2(n4663), .ZN(n4887) );
  NAND4_X1 U2442 ( .A1(n2398), .A2(n2464), .A3(n2612), .A4(n2265), .ZN(n2579)
         );
  AND2_X1 U2443 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2560)
         );
  NAND2_X1 U2444 ( .A1(n2548), .A2(IR_REG_31__SCAN_IN), .ZN(n3214) );
  NOR2_X1 U2445 ( .A1(n3475), .A2(n2498), .ZN(n2497) );
  OAI211_X1 U2446 ( .C1(n2481), .C2(n2479), .A(n3064), .B(n2476), .ZN(n3068)
         );
  NAND2_X1 U2447 ( .A1(n2485), .A2(n2480), .ZN(n2479) );
  OR2_X1 U2448 ( .A1(n2259), .A2(n3418), .ZN(n3419) );
  NAND4_X1 U2449 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n4861)
         );
  NAND2_X1 U2450 ( .A1(n2631), .A2(n2504), .ZN(n3742) );
  AND2_X1 U2451 ( .A1(n2384), .A2(n2509), .ZN(n4541) );
  XNOR2_X1 U2452 ( .A(n2968), .B(n2984), .ZN(n4551) );
  NAND2_X1 U2453 ( .A1(n4551), .A2(REG2_REG_8__SCAN_IN), .ZN(n4550) );
  AND2_X1 U2454 ( .A1(n2416), .A2(n2990), .ZN(n3744) );
  AND2_X1 U2455 ( .A1(n2989), .A2(REG1_REG_10__SCAN_IN), .ZN(n2416) );
  OAI211_X1 U2456 ( .C1(n4594), .C2(n2444), .A(n2439), .B(n2437), .ZN(n3760)
         );
  NAND2_X1 U2457 ( .A1(n2445), .A2(n2447), .ZN(n2444) );
  AND2_X1 U2458 ( .A1(n2440), .A2(n2443), .ZN(n2439) );
  NOR2_X1 U2459 ( .A1(n4133), .A2(n3760), .ZN(n3766) );
  AND2_X1 U2460 ( .A1(n2426), .A2(n2372), .ZN(n2371) );
  NAND2_X1 U2461 ( .A1(n2427), .A2(REG1_REG_19__SCAN_IN), .ZN(n2426) );
  AOI21_X1 U2462 ( .B1(n2373), .B2(n3326), .A(n3803), .ZN(n2372) );
  INV_X1 U2463 ( .A(n2429), .ZN(n2427) );
  INV_X1 U2464 ( .A(n2425), .ZN(n2424) );
  OAI22_X1 U2465 ( .A1(n2428), .A2(n4609), .B1(n2429), .B2(n4609), .ZN(n2425)
         );
  INV_X1 U2466 ( .A(n2423), .ZN(n2422) );
  OAI22_X1 U2467 ( .A1(n2428), .A2(n3326), .B1(REG1_REG_19__SCAN_IN), .B2(
        n2429), .ZN(n2423) );
  INV_X1 U2469 ( .A(IR_REG_30__SCAN_IN), .ZN(n3200) );
  INV_X1 U2470 ( .A(n4590), .ZN(n2412) );
  AND2_X1 U2471 ( .A1(n2412), .A2(n3130), .ZN(n2409) );
  INV_X1 U2472 ( .A(n3806), .ZN(n2387) );
  INV_X1 U2473 ( .A(n3795), .ZN(n2388) );
  AND2_X1 U2474 ( .A1(n3954), .A2(n3680), .ZN(n3857) );
  AOI21_X1 U2475 ( .B1(n3905), .B2(n2333), .A(n3864), .ZN(n2332) );
  OR2_X1 U2476 ( .A1(n3494), .A2(n3334), .ZN(n2462) );
  NOR2_X1 U2477 ( .A1(n4918), .A2(n4917), .ZN(n3367) );
  INV_X1 U2478 ( .A(n3345), .ZN(n3460) );
  AND2_X1 U2479 ( .A1(n2945), .A2(n2677), .ZN(n2680) );
  INV_X1 U2480 ( .A(n2474), .ZN(n2471) );
  AND2_X1 U2481 ( .A1(n3688), .A2(n3933), .ZN(n3858) );
  NAND2_X1 U2482 ( .A1(n2442), .A2(n4466), .ZN(n2441) );
  INV_X1 U2483 ( .A(n2446), .ZN(n2442) );
  INV_X1 U2484 ( .A(n3770), .ZN(n2395) );
  NOR2_X1 U2485 ( .A1(n3780), .A2(n3782), .ZN(n3783) );
  INV_X1 U2486 ( .A(n2432), .ZN(n2391) );
  AND2_X1 U2487 ( .A1(n3934), .A2(n3858), .ZN(n3917) );
  OR2_X1 U2488 ( .A1(n4091), .A2(n4069), .ZN(n4048) );
  INV_X1 U2489 ( .A(n3820), .ZN(n2352) );
  OR2_X1 U2490 ( .A1(n4861), .A2(n3877), .ZN(n3687) );
  NAND2_X1 U2491 ( .A1(n3849), .A2(n3848), .ZN(n4854) );
  INV_X1 U2492 ( .A(n4857), .ZN(n3848) );
  INV_X1 U2493 ( .A(n4858), .ZN(n3849) );
  NOR2_X1 U2494 ( .A1(n2404), .A2(n3169), .ZN(n2403) );
  NAND2_X1 U2495 ( .A1(n3195), .A2(n3177), .ZN(n2404) );
  XNOR2_X1 U2496 ( .A(n2334), .B(n3865), .ZN(n3866) );
  OAI21_X1 U2497 ( .B1(n3904), .B2(n2331), .A(n2330), .ZN(n2334) );
  AOI21_X1 U2498 ( .B1(n2332), .B2(n3862), .A(n3863), .ZN(n2330) );
  INV_X1 U2499 ( .A(n2332), .ZN(n2331) );
  NOR2_X1 U2500 ( .A1(n2856), .A2(n3252), .ZN(n2855) );
  AND2_X1 U2501 ( .A1(n2276), .A2(n3172), .ZN(n2463) );
  NOR2_X1 U2502 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2526)
         );
  NOR2_X1 U2503 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2525)
         );
  INV_X1 U2504 ( .A(IR_REG_2__SCAN_IN), .ZN(n4431) );
  AND2_X1 U2505 ( .A1(n3319), .A2(n3318), .ZN(n3320) );
  AND3_X1 U2506 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2843) );
  XNOR2_X1 U2507 ( .A(n2749), .B(n3458), .ZN(n2825) );
  NAND2_X1 U2508 ( .A1(n3019), .A2(n2486), .ZN(n2485) );
  INV_X1 U2509 ( .A(n3020), .ZN(n2486) );
  INV_X1 U2510 ( .A(n3065), .ZN(n2480) );
  INV_X1 U2511 ( .A(n2484), .ZN(n2482) );
  NAND2_X1 U2512 ( .A1(n2637), .A2(n2636), .ZN(n3256) );
  NAND2_X1 U2513 ( .A1(n2642), .A2(n2641), .ZN(n3257) );
  NAND2_X1 U2514 ( .A1(n3742), .A2(n3437), .ZN(n2642) );
  AND2_X1 U2515 ( .A1(n3366), .A2(n3365), .ZN(n4901) );
  INV_X1 U2516 ( .A(n3320), .ZN(n3549) );
  AND2_X1 U2517 ( .A1(n3002), .A2(n3001), .ZN(n3237) );
  OAI21_X1 U2518 ( .B1(n2592), .B2(IR_REG_28__SCAN_IN), .A(n2591), .ZN(n2594)
         );
  NAND2_X1 U2519 ( .A1(n2592), .A2(IR_REG_27__SCAN_IN), .ZN(n2591) );
  NOR2_X1 U2520 ( .A1(n2682), .A2(n2678), .ZN(n2691) );
  OR2_X1 U2521 ( .A1(n3451), .A2(n3927), .ZN(n3420) );
  NAND2_X1 U2522 ( .A1(n2737), .A2(REG1_REG_0__SCAN_IN), .ZN(n2630) );
  NAND3_X1 U2523 ( .A1(n4463), .A2(n2675), .A3(n4464), .ZN(n2767) );
  NOR2_X1 U2524 ( .A1(n2615), .A2(n2616), .ZN(n2974) );
  OR2_X1 U2525 ( .A1(n4632), .A2(n4631), .ZN(n2421) );
  NAND2_X1 U2526 ( .A1(n2421), .A2(n2975), .ZN(n2976) );
  NOR2_X1 U2527 ( .A1(n2960), .A2(n4509), .ZN(n2961) );
  INV_X1 U2528 ( .A(n4932), .ZN(n4637) );
  OR2_X1 U2529 ( .A1(n4652), .A2(n2738), .ZN(n2454) );
  NAND2_X1 U2530 ( .A1(n2379), .A2(n2908), .ZN(n2383) );
  NAND2_X1 U2531 ( .A1(n2380), .A2(n2908), .ZN(n2381) );
  NAND4_X1 U2532 ( .A1(n2381), .A2(REG2_REG_6__SCAN_IN), .A3(n2383), .A4(n2382), .ZN(n2384) );
  INV_X1 U2533 ( .A(n4532), .ZN(n2406) );
  XNOR2_X1 U2534 ( .A(n2985), .B(n2984), .ZN(n4553) );
  OAI21_X1 U2535 ( .B1(n4532), .B2(n2407), .A(n2405), .ZN(n2985) );
  NAND2_X1 U2536 ( .A1(n2309), .A2(REG1_REG_6__SCAN_IN), .ZN(n2407) );
  OAI21_X1 U2537 ( .B1(n2983), .B2(n2408), .A(n2309), .ZN(n2405) );
  INV_X1 U2538 ( .A(n4544), .ZN(n2408) );
  XNOR2_X1 U2539 ( .A(n3746), .B(n4583), .ZN(n4582) );
  NAND2_X1 U2540 ( .A1(n4582), .A2(REG1_REG_12__SCAN_IN), .ZN(n4581) );
  INV_X1 U2541 ( .A(n2441), .ZN(n2438) );
  OR2_X1 U2542 ( .A1(n2441), .A2(n2447), .ZN(n2440) );
  NAND2_X1 U2543 ( .A1(n2446), .A2(n2445), .ZN(n2443) );
  NAND2_X1 U2544 ( .A1(n4584), .A2(n3758), .ZN(n4594) );
  INV_X1 U2545 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U2546 ( .A1(n4604), .A2(n3793), .ZN(n3794) );
  NAND2_X1 U2547 ( .A1(n2433), .A2(n4098), .ZN(n2432) );
  NAND2_X1 U2548 ( .A1(n3794), .A2(n3795), .ZN(n3804) );
  AND2_X1 U2549 ( .A1(n3800), .A2(n4893), .ZN(n3801) );
  NAND2_X1 U2550 ( .A1(n3811), .A2(n3808), .ZN(n2428) );
  OAI21_X1 U2551 ( .B1(n3810), .B2(n4650), .A(n2305), .ZN(n2429) );
  NAND2_X1 U2552 ( .A1(n3901), .A2(n2271), .ZN(n3893) );
  NAND2_X1 U2553 ( .A1(n2360), .A2(n2359), .ZN(n3885) );
  AOI21_X1 U2554 ( .B1(n2361), .B2(n2505), .A(n2293), .ZN(n2359) );
  AND4_X1 U2555 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3907)
         );
  OR2_X1 U2556 ( .A1(n3416), .A2(n3561), .ZN(n3430) );
  NOR2_X1 U2557 ( .A1(n3944), .A2(n3926), .ZN(n3901) );
  OR2_X1 U2558 ( .A1(n3943), .A2(n3936), .ZN(n3944) );
  INV_X1 U2559 ( .A(n3838), .ZN(n3926) );
  AND2_X1 U2560 ( .A1(n3678), .A2(n3859), .ZN(n3921) );
  AOI21_X1 U2561 ( .B1(n2366), .B2(n2368), .A(n2292), .ZN(n2364) );
  INV_X1 U2562 ( .A(n2366), .ZN(n2365) );
  NAND2_X1 U2563 ( .A1(n2369), .A2(n3974), .ZN(n2368) );
  OR2_X1 U2564 ( .A1(n3372), .A2(n3371), .ZN(n3392) );
  NOR2_X1 U2565 ( .A1(n4036), .A2(n2396), .ZN(n3979) );
  NAND2_X1 U2566 ( .A1(n3323), .A2(REG3_REG_20__SCAN_IN), .ZN(n3352) );
  OR2_X1 U2567 ( .A1(n3352), .A2(n4911), .ZN(n3372) );
  NAND2_X1 U2568 ( .A1(n2327), .A2(n3853), .ZN(n4019) );
  NAND2_X1 U2569 ( .A1(n4056), .A2(n4037), .ZN(n4036) );
  NAND2_X1 U2570 ( .A1(n4104), .A2(n2328), .ZN(n4027) );
  NAND2_X1 U2571 ( .A1(n3307), .A2(REG3_REG_18__SCAN_IN), .ZN(n3324) );
  AND2_X1 U2572 ( .A1(REG3_REG_17__SCAN_IN), .A2(n3296), .ZN(n3307) );
  NAND2_X1 U2573 ( .A1(n4846), .A2(n2270), .ZN(n4074) );
  NAND2_X1 U2574 ( .A1(n4846), .A2(n2400), .ZN(n4096) );
  NAND2_X1 U2575 ( .A1(n4104), .A2(n3851), .ZN(n4087) );
  AND2_X1 U2576 ( .A1(n3816), .A2(n2337), .ZN(n2336) );
  NAND2_X1 U2577 ( .A1(n4846), .A2(n2401), .ZN(n4110) );
  AND2_X1 U2578 ( .A1(n4846), .A2(n4852), .ZN(n4848) );
  NAND2_X1 U2579 ( .A1(n3217), .A2(REG3_REG_15__SCAN_IN), .ZN(n3264) );
  INV_X1 U2580 ( .A(n3815), .ZN(n4852) );
  INV_X1 U2581 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4398) );
  NOR2_X1 U2582 ( .A1(n3182), .A2(n4398), .ZN(n3217) );
  NOR2_X1 U2583 ( .A1(n4130), .A2(n4129), .ZN(n4846) );
  NAND2_X1 U2584 ( .A1(n3194), .A2(n2402), .ZN(n4130) );
  AND2_X1 U2585 ( .A1(n2403), .A2(n3576), .ZN(n2402) );
  NAND2_X1 U2586 ( .A1(n3151), .A2(REG3_REG_13__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U2587 ( .A1(n4218), .A2(n3168), .ZN(n2338) );
  NAND2_X1 U2588 ( .A1(n3194), .A2(n2403), .ZN(n4211) );
  INV_X1 U2589 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3094) );
  NOR2_X1 U2590 ( .A1(n3095), .A2(n3094), .ZN(n3131) );
  NOR2_X1 U2591 ( .A1(n4763), .A2(n2404), .ZN(n4796) );
  INV_X1 U2592 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4342) );
  NOR2_X1 U2593 ( .A1(n4763), .A2(n4224), .ZN(n4795) );
  NAND2_X1 U2594 ( .A1(n2320), .A2(n2318), .ZN(n3176) );
  AND2_X1 U2595 ( .A1(n2322), .A2(n2319), .ZN(n2318) );
  OR2_X1 U2596 ( .A1(n3031), .A2(n3030), .ZN(n3071) );
  NAND2_X1 U2597 ( .A1(n2320), .A2(n2322), .ZN(n4756) );
  INV_X1 U2598 ( .A(n3164), .ZN(n3054) );
  NAND2_X1 U2599 ( .A1(n4721), .A2(n3054), .ZN(n4764) );
  NOR2_X1 U2600 ( .A1(n2917), .A2(n2916), .ZN(n3009) );
  NOR2_X1 U2601 ( .A1(n4722), .A2(n4733), .ZN(n4721) );
  OR2_X1 U2602 ( .A1(n3739), .A2(n2909), .ZN(n2345) );
  NAND2_X1 U2603 ( .A1(n2890), .A2(n2343), .ZN(n2342) );
  NOR2_X1 U2604 ( .A1(n2910), .A2(n2344), .ZN(n2343) );
  INV_X1 U2605 ( .A(n2889), .ZN(n2344) );
  NAND2_X1 U2606 ( .A1(n2897), .A2(n2927), .ZN(n4722) );
  NAND2_X1 U2607 ( .A1(n2310), .A2(n2311), .ZN(n3048) );
  AOI21_X1 U2608 ( .B1(n2313), .B2(n2317), .A(n2312), .ZN(n2311) );
  NAND2_X1 U2609 ( .A1(n2315), .A2(n3626), .ZN(n2913) );
  NAND2_X1 U2610 ( .A1(n2316), .A2(n3623), .ZN(n2315) );
  INV_X1 U2611 ( .A(n2892), .ZN(n2316) );
  AND2_X1 U2612 ( .A1(n2855), .A2(n2874), .ZN(n2881) );
  NAND2_X1 U2613 ( .A1(n2854), .A2(n2787), .ZN(n2873) );
  OR2_X1 U2614 ( .A1(n2358), .A2(n2814), .ZN(n2357) );
  INV_X1 U2615 ( .A(n2786), .ZN(n2358) );
  NAND2_X1 U2616 ( .A1(n3616), .A2(n3618), .ZN(n2860) );
  NAND2_X1 U2617 ( .A1(n2853), .A2(n2860), .ZN(n2854) );
  INV_X1 U2618 ( .A(n2815), .ZN(n3692) );
  INV_X1 U2619 ( .A(n3705), .ZN(n3614) );
  INV_X1 U2620 ( .A(n4853), .ZN(n4787) );
  OR2_X1 U2621 ( .A1(n4664), .A2(n2805), .ZN(n2856) );
  INV_X1 U2622 ( .A(IR_REG_20__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U2623 ( .A1(n2790), .A2(n4664), .ZN(n3705) );
  AND2_X1 U2624 ( .A1(n2938), .A2(n2937), .ZN(n2946) );
  AND2_X1 U2625 ( .A1(n2587), .A2(n4463), .ZN(n2674) );
  AND2_X1 U2626 ( .A1(n2463), .A2(n2399), .ZN(n2398) );
  INV_X1 U2627 ( .A(IR_REG_21__SCAN_IN), .ZN(n2399) );
  AND2_X1 U2628 ( .A1(n2503), .A2(n2555), .ZN(n2501) );
  NAND2_X1 U2629 ( .A1(n2538), .A2(n2536), .ZN(n2540) );
  XNOR2_X1 U2630 ( .A(n2556), .B(n2555), .ZN(n2793) );
  INV_X1 U2631 ( .A(n3278), .ZN(n2550) );
  NAND2_X1 U2632 ( .A1(n2523), .A2(n2522), .ZN(n3273) );
  INV_X1 U2633 ( .A(IR_REG_15__SCAN_IN), .ZN(n2523) );
  INV_X1 U2634 ( .A(IR_REG_16__SCAN_IN), .ZN(n2522) );
  INV_X1 U2635 ( .A(IR_REG_13__SCAN_IN), .ZN(n3172) );
  AND4_X1 U2636 ( .A1(n2949), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n2520)
         );
  INV_X1 U2637 ( .A(IR_REG_9__SCAN_IN), .ZN(n2517) );
  AND2_X1 U2638 ( .A1(n3144), .A2(n3124), .ZN(n4570) );
  OR2_X1 U2639 ( .A1(n2951), .A2(IR_REG_9__SCAN_IN), .ZN(n3121) );
  INV_X1 U2640 ( .A(IR_REG_3__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U2641 ( .A1(n2483), .A2(n2484), .ZN(n3022) );
  NAND2_X1 U2642 ( .A1(n2499), .A2(n3558), .ZN(n3476) );
  NAND2_X1 U2643 ( .A1(n2473), .A2(n3227), .ZN(n3263) );
  OR2_X1 U2644 ( .A1(n3226), .A2(n3228), .ZN(n2473) );
  NAND2_X1 U2645 ( .A1(n3495), .A2(n3494), .ZN(n3493) );
  NOR2_X1 U2646 ( .A1(n2496), .A2(n2493), .ZN(n2488) );
  NAND2_X1 U2647 ( .A1(n2496), .A2(n2493), .ZN(n2491) );
  NAND2_X1 U2648 ( .A1(n2494), .A2(n2493), .ZN(n2492) );
  NAND2_X1 U2649 ( .A1(n2478), .A2(n2485), .ZN(n3066) );
  NAND2_X1 U2650 ( .A1(n2481), .A2(n2483), .ZN(n2478) );
  AOI21_X1 U2651 ( .B1(n2458), .B2(n3142), .A(n2302), .ZN(n2457) );
  INV_X1 U2652 ( .A(n3119), .ZN(n2458) );
  AND2_X1 U2653 ( .A1(n3293), .A2(n3514), .ZN(n3294) );
  CLKBUF_X1 U2654 ( .A(n3090), .Z(n3067) );
  CLKBUF_X1 U2655 ( .A(n3226), .Z(n3230) );
  CLKBUF_X1 U2656 ( .A(n3484), .Z(n3542) );
  NAND2_X1 U2657 ( .A1(n3120), .A2(n3119), .ZN(n3143) );
  NAND2_X1 U2658 ( .A1(n3000), .A2(n2999), .ZN(n3240) );
  INV_X1 U2659 ( .A(n4913), .ZN(n4899) );
  INV_X1 U2660 ( .A(n4830), .ZN(n4921) );
  INV_X1 U2661 ( .A(n4930), .ZN(n3565) );
  OR2_X1 U2662 ( .A1(n2692), .A2(n4932), .ZN(n4830) );
  INV_X1 U2663 ( .A(n3567), .ZN(n4925) );
  NAND4_X1 U2664 ( .A1(n3398), .A2(n3397), .A3(n3396), .A4(n3395), .ZN(n3993)
         );
  OR2_X1 U2665 ( .A1(n2259), .A2(n3394), .ZN(n3395) );
  OR2_X1 U2666 ( .A1(n2259), .A2(n3374), .ZN(n3375) );
  AND4_X1 U2667 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n4912)
         );
  NAND4_X1 U2668 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n4898)
         );
  NAND4_X1 U2669 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n4922)
         );
  NAND4_X1 U2670 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n4904)
         );
  NAND4_X1 U2671 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n4103)
         );
  NAND4_X1 U2672 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n4106)
         );
  NAND4_X1 U2673 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n4850)
         );
  NAND4_X1 U2674 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n4217)
         );
  NAND4_X1 U2675 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n4789)
         );
  NAND4_X1 U2676 ( .A1(n3101), .A2(n3100), .A3(n3099), .A4(n3098), .ZN(n3737)
         );
  NAND4_X1 U2677 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n4788)
         );
  NAND4_X1 U2678 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n4225)
         );
  NAND4_X1 U2679 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n4758)
         );
  OR2_X1 U2680 ( .A1(n2694), .A2(REG3_REG_3__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U2681 ( .A1(n2737), .A2(REG1_REG_3__SCAN_IN), .ZN(n2727) );
  NAND4_X1 U2682 ( .A1(n2699), .A2(n2698), .A3(n2697), .A4(n2696), .ZN(n3740)
         );
  OR2_X1 U2683 ( .A1(n2694), .A2(n2858), .ZN(n2697) );
  OR2_X1 U2684 ( .A1(n2693), .A2(n2957), .ZN(n2699) );
  OR2_X1 U2685 ( .A1(n2259), .A2(n4690), .ZN(n2696) );
  OR2_X1 U2686 ( .A1(n2694), .A2(n2817), .ZN(n2649) );
  NAND2_X1 U2687 ( .A1(n3007), .A2(REG0_REG_1__SCAN_IN), .ZN(n2650) );
  OR2_X1 U2688 ( .A1(n2259), .A2(n2420), .ZN(n2506) );
  AND2_X1 U2689 ( .A1(n2610), .A2(n2609), .ZN(n4505) );
  AND2_X1 U2690 ( .A1(n2289), .A2(n2378), .ZN(n2377) );
  NOR2_X1 U2691 ( .A1(n2956), .A2(n2376), .ZN(n4629) );
  AND2_X1 U2692 ( .A1(n4468), .A2(REG2_REG_1__SCAN_IN), .ZN(n2376) );
  INV_X1 U2693 ( .A(n2375), .ZN(n4627) );
  XNOR2_X1 U2694 ( .A(n2961), .B(n4703), .ZN(n4652) );
  INV_X1 U2695 ( .A(n2454), .ZN(n4651) );
  NOR2_X1 U2696 ( .A1(n4648), .A2(n2980), .ZN(n4523) );
  NAND2_X1 U2697 ( .A1(n4550), .A2(n2969), .ZN(n4565) );
  NAND2_X1 U2698 ( .A1(n3755), .A2(n3756), .ZN(n4576) );
  INV_X1 U2699 ( .A(n3744), .ZN(n2415) );
  NAND2_X1 U2700 ( .A1(n4581), .A2(n3747), .ZN(n4592) );
  NAND2_X1 U2701 ( .A1(n2273), .A2(n3749), .ZN(n3750) );
  INV_X1 U2702 ( .A(n2431), .ZN(n2430) );
  AND2_X1 U2703 ( .A1(n2431), .A2(n2273), .ZN(n3775) );
  NOR2_X1 U2704 ( .A1(n3766), .A2(n3765), .ZN(n3771) );
  XNOR2_X1 U2705 ( .A(n3792), .B(n4877), .ZN(n4605) );
  NAND2_X1 U2706 ( .A1(n4605), .A2(n4115), .ZN(n4604) );
  NAND2_X1 U2707 ( .A1(n3804), .A2(n2432), .ZN(n4613) );
  INV_X1 U2708 ( .A(n4607), .ZN(n4650) );
  AND2_X1 U2709 ( .A1(n4505), .A2(n4932), .ZN(n4656) );
  XNOR2_X1 U2710 ( .A(n4152), .B(n4146), .ZN(n4941) );
  OR2_X1 U2711 ( .A1(n4157), .A2(n3876), .ZN(n2512) );
  AOI211_X1 U2712 ( .C1(n3891), .C2(n4731), .A(n3890), .B(n3889), .ZN(n4162)
         );
  AND2_X1 U2713 ( .A1(n2363), .A2(n3839), .ZN(n3900) );
  OR2_X1 U2714 ( .A1(n3916), .A2(n2505), .ZN(n2363) );
  NAND2_X1 U2715 ( .A1(n4117), .A2(n3820), .ZN(n4086) );
  NAND2_X1 U2716 ( .A1(n2355), .A2(n3690), .ZN(n4117) );
  INV_X1 U2717 ( .A(n4119), .ZN(n2355) );
  NAND2_X1 U2718 ( .A1(n2890), .A2(n2889), .ZN(n2911) );
  NAND2_X1 U2719 ( .A1(n4674), .A2(n4727), .ZN(n4140) );
  NAND2_X1 U2720 ( .A1(n2815), .A2(n2814), .ZN(n2813) );
  INV_X1 U2721 ( .A(n4934), .ZN(n4940) );
  AND2_X1 U2722 ( .A1(n4674), .A2(n2804), .ZN(n4805) );
  NOR2_X1 U2723 ( .A1(n4157), .A2(n2511), .ZN(n4160) );
  AND2_X2 U2724 ( .A1(n2946), .A2(n2939), .ZN(n4897) );
  AND2_X1 U2725 ( .A1(n2766), .A2(STATE_REG_SCAN_IN), .ZN(n3729) );
  NAND2_X1 U2726 ( .A1(n3203), .A2(IR_REG_31__SCAN_IN), .ZN(n2581) );
  XNOR2_X1 U2727 ( .A(n2529), .B(IR_REG_26__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U2728 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2529) );
  INV_X1 U2729 ( .A(n2585), .ZN(n2675) );
  XNOR2_X1 U2730 ( .A(n2537), .B(IR_REG_24__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U2731 ( .A1(n2540), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  INV_X1 U2732 ( .A(n2793), .ZN(n3731) );
  OR2_X1 U2733 ( .A1(n2607), .A2(n2954), .ZN(n2712) );
  NAND2_X1 U2734 ( .A1(n2371), .A2(n2424), .ZN(n2370) );
  INV_X1 U2735 ( .A(n2736), .ZN(n3457) );
  AND2_X2 U2736 ( .A1(n3345), .A2(n2264), .ZN(n2736) );
  AND2_X1 U2737 ( .A1(n2275), .A2(n2501), .ZN(n2265) );
  AND2_X1 U2738 ( .A1(n2466), .A2(n2468), .ZN(n3510) );
  AND2_X1 U2739 ( .A1(n2415), .A2(n2990), .ZN(n2266) );
  INV_X1 U2740 ( .A(n3862), .ZN(n2333) );
  AND2_X1 U2741 ( .A1(n4225), .A2(n4765), .ZN(n2267) );
  AND2_X1 U2742 ( .A1(n2417), .A2(REG1_REG_10__SCAN_IN), .ZN(n2268) );
  NOR2_X1 U2743 ( .A1(n2303), .A2(n2983), .ZN(n2269) );
  INV_X1 U2744 ( .A(n4593), .ZN(n2447) );
  AND2_X1 U2745 ( .A1(n2400), .A2(n4069), .ZN(n2270) );
  AND2_X1 U2746 ( .A1(n3894), .A2(n3906), .ZN(n2271) );
  AND2_X1 U2747 ( .A1(n2271), .A2(n3879), .ZN(n2272) );
  NAND4_X1 U2748 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .ZN(n2778)
         );
  NAND4_X1 U2749 ( .A1(n2727), .A2(n2726), .A3(n2725), .A4(n2724), .ZN(n2757)
         );
  AOI21_X1 U2750 ( .B1(n4032), .B2(n3828), .A(n3827), .ZN(n3973) );
  OR2_X1 U2751 ( .A1(n3748), .A2(n2445), .ZN(n2273) );
  INV_X1 U2752 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2420) );
  AND2_X1 U2753 ( .A1(n2398), .A2(n2464), .ZN(n2545) );
  OAI21_X1 U2754 ( .B1(n3594), .B2(n2634), .A(n2633), .ZN(n4664) );
  NAND2_X1 U2755 ( .A1(n3493), .A2(n3335), .ZN(n4900) );
  OR2_X1 U2756 ( .A1(n2599), .A2(n2600), .ZN(n2694) );
  OR2_X1 U2757 ( .A1(n3238), .A2(n3237), .ZN(n2274) );
  AND2_X1 U2758 ( .A1(n2528), .A2(n2502), .ZN(n2275) );
  XNOR2_X1 U2759 ( .A(n2577), .B(n2576), .ZN(n2600) );
  AND4_X1 U2760 ( .A1(n2527), .A2(n2526), .A3(n2525), .A4(n2524), .ZN(n2276)
         );
  AND2_X1 U2761 ( .A1(n3840), .A2(n3906), .ZN(n2277) );
  NAND2_X1 U2762 ( .A1(n2464), .A2(n2463), .ZN(n2543) );
  NAND2_X1 U2763 ( .A1(n2534), .A2(n2528), .ZN(n2530) );
  OR2_X1 U2764 ( .A1(n3800), .A2(n4893), .ZN(n2278) );
  INV_X1 U2765 ( .A(IR_REG_31__SCAN_IN), .ZN(n2954) );
  NOR2_X1 U2766 ( .A1(n3771), .A2(n3770), .ZN(n2279) );
  NAND2_X1 U2767 ( .A1(n3273), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  INV_X1 U2768 ( .A(n3623), .ZN(n2317) );
  AND2_X1 U2769 ( .A1(n3804), .A2(n2389), .ZN(n2281) );
  AND2_X1 U2770 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2282)
         );
  AND2_X1 U2771 ( .A1(n2499), .A2(n2497), .ZN(n2283) );
  INV_X1 U2772 ( .A(n3262), .ZN(n2475) );
  NAND2_X1 U2773 ( .A1(n2462), .A2(n4915), .ZN(n2284) );
  OR2_X1 U2774 ( .A1(n2469), .A2(n2472), .ZN(n2285) );
  NOR2_X1 U2775 ( .A1(n2912), .A2(n2314), .ZN(n2313) );
  AND2_X1 U2776 ( .A1(n3089), .A2(n3142), .ZN(n2286) );
  AND2_X1 U2777 ( .A1(n2510), .A2(n2345), .ZN(n2287) );
  NAND2_X1 U2778 ( .A1(n4682), .A2(REG2_REG_2__SCAN_IN), .ZN(n2288) );
  OR2_X1 U2779 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2289)
         );
  NAND2_X1 U2780 ( .A1(n3240), .A2(n2274), .ZN(n2483) );
  XOR2_X1 U2781 ( .A(n3462), .B(n3461), .Z(n2290) );
  OR3_X1 U2782 ( .A1(n4036), .A2(n4923), .A3(n4008), .ZN(n2291) );
  NAND2_X1 U2783 ( .A1(n2338), .A2(n3170), .ZN(n3814) );
  NOR2_X1 U2784 ( .A1(n2988), .A2(n2435), .ZN(n3743) );
  OAI21_X1 U2785 ( .B1(n3973), .B2(n2365), .A(n2364), .ZN(n3953) );
  AND2_X1 U2786 ( .A1(n3960), .A2(n3980), .ZN(n2292) );
  INV_X1 U2787 ( .A(n3558), .ZN(n2498) );
  AND2_X1 U2788 ( .A1(n3922), .A2(n3902), .ZN(n2293) );
  NAND2_X1 U2789 ( .A1(n3090), .A2(n3089), .ZN(n3120) );
  AND2_X1 U2790 ( .A1(n4103), .A2(n4094), .ZN(n2294) );
  INV_X1 U2791 ( .A(n3169), .ZN(n4212) );
  INV_X1 U2792 ( .A(n3686), .ZN(n3851) );
  NAND2_X1 U2793 ( .A1(n2608), .A2(n2377), .ZN(n2652) );
  NOR2_X1 U2794 ( .A1(n4103), .A2(n4094), .ZN(n2295) );
  NOR2_X1 U2795 ( .A1(n4225), .A2(n4765), .ZN(n2296) );
  INV_X1 U2796 ( .A(n2397), .ZN(n4015) );
  NOR2_X1 U2797 ( .A1(n4036), .A2(n4923), .ZN(n2397) );
  AND2_X1 U2798 ( .A1(n2430), .A2(n2273), .ZN(n2297) );
  OR2_X1 U2799 ( .A1(n3287), .A2(n3286), .ZN(n2298) );
  INV_X1 U2800 ( .A(IR_REG_28__SCAN_IN), .ZN(n2612) );
  AND2_X1 U2801 ( .A1(n3321), .A2(n3549), .ZN(n2299) );
  AND2_X1 U2802 ( .A1(n3907), .A2(n3842), .ZN(n3863) );
  INV_X1 U2803 ( .A(n3633), .ZN(n2319) );
  AND2_X1 U2804 ( .A1(n2328), .A2(n3702), .ZN(n2300) );
  INV_X1 U2805 ( .A(n2468), .ZN(n2467) );
  AOI22_X1 U2806 ( .A1(n2469), .A2(n2471), .B1(n2472), .B2(n3228), .ZN(n2468)
         );
  NAND2_X1 U2807 ( .A1(n2981), .A2(REG2_REG_5__SCAN_IN), .ZN(n2301) );
  INV_X1 U2808 ( .A(IR_REG_29__SCAN_IN), .ZN(n2576) );
  INV_X1 U2809 ( .A(n4467), .ZN(n2435) );
  NAND2_X1 U2810 ( .A1(n2342), .A2(n2345), .ZN(n3042) );
  INV_X1 U2811 ( .A(n3227), .ZN(n2470) );
  OAI22_X1 U2812 ( .A1(n2873), .A2(n2872), .B1(n3620), .B2(n2874), .ZN(n2887)
         );
  NOR2_X1 U2813 ( .A1(n4764), .A2(n4765), .ZN(n3194) );
  INV_X1 U2814 ( .A(n4753), .ZN(n2350) );
  AND2_X1 U2815 ( .A1(n3127), .A2(n3126), .ZN(n2302) );
  AND2_X1 U2816 ( .A1(n2406), .A2(REG1_REG_6__SCAN_IN), .ZN(n2303) );
  INV_X1 U2817 ( .A(n2390), .ZN(n2389) );
  OR2_X1 U2818 ( .A1(n4614), .A2(n2391), .ZN(n2390) );
  INV_X1 U2819 ( .A(n4569), .ZN(n2418) );
  INV_X1 U2820 ( .A(n4020), .ZN(n4923) );
  NOR2_X1 U2821 ( .A1(n3759), .A2(REG1_REG_13__SCAN_IN), .ZN(n2304) );
  INV_X1 U2822 ( .A(n3805), .ZN(n2433) );
  NOR2_X1 U2823 ( .A1(n2896), .A2(n2909), .ZN(n2897) );
  NOR2_X1 U2824 ( .A1(n4656), .A2(n3808), .ZN(n2305) );
  AND2_X1 U2825 ( .A1(n4505), .A2(n4639), .ZN(n4609) );
  NAND2_X1 U2826 ( .A1(n2357), .A2(n2356), .ZN(n2853) );
  AND2_X1 U2827 ( .A1(n4465), .A2(REG2_REG_15__SCAN_IN), .ZN(n2306) );
  AND2_X1 U2828 ( .A1(n2454), .A2(n2453), .ZN(n2307) );
  AND2_X1 U2829 ( .A1(n2272), .A2(n3606), .ZN(n2308) );
  OR2_X1 U2830 ( .A1(n4538), .A2(REG1_REG_7__SCAN_IN), .ZN(n2309) );
  INV_X1 U2831 ( .A(IR_REG_4__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U2832 ( .A1(n2892), .A2(n2313), .ZN(n2310) );
  INV_X1 U2833 ( .A(n4730), .ZN(n2321) );
  OAI21_X1 U2834 ( .B1(n4730), .B2(n3050), .A(n3632), .ZN(n3174) );
  AOI21_X1 U2835 ( .B1(n3050), .B2(n3632), .A(n2326), .ZN(n2325) );
  NAND2_X1 U2836 ( .A1(n4104), .A2(n2300), .ZN(n2327) );
  NOR2_X2 U2837 ( .A1(n3904), .A2(n3905), .ZN(n3903) );
  NAND2_X1 U2838 ( .A1(n2335), .A2(n2336), .ZN(n3819) );
  NAND2_X1 U2839 ( .A1(n4218), .A2(n2339), .ZN(n2335) );
  NAND2_X1 U2840 ( .A1(n2342), .A2(n2287), .ZN(n3044) );
  NAND2_X1 U2841 ( .A1(n3163), .A2(n2348), .ZN(n2346) );
  NAND2_X1 U2842 ( .A1(n2346), .A2(n2347), .ZN(n4221) );
  OAI21_X1 U2843 ( .B1(n4119), .B2(n2353), .A(n2351), .ZN(n4081) );
  NAND3_X1 U2844 ( .A1(n3615), .A2(n2786), .A3(n3612), .ZN(n2356) );
  NAND2_X1 U2845 ( .A1(n3615), .A2(n3612), .ZN(n2815) );
  NAND2_X1 U2846 ( .A1(n3916), .A2(n2361), .ZN(n2360) );
  INV_X1 U2847 ( .A(n3953), .ZN(n3834) );
  NAND3_X1 U2848 ( .A1(n2398), .A2(n2464), .A3(n2265), .ZN(n2611) );
  NAND3_X1 U2849 ( .A1(n2374), .A2(n2370), .A3(n3813), .ZN(U3259) );
  NAND3_X1 U2850 ( .A1(n2422), .A2(n2424), .A3(n3803), .ZN(n2374) );
  NAND3_X1 U2851 ( .A1(n2451), .A2(n4718), .A3(n2448), .ZN(n2382) );
  INV_X1 U2852 ( .A(n2448), .ZN(n2379) );
  INV_X1 U2853 ( .A(n2451), .ZN(n2380) );
  NAND3_X1 U2854 ( .A1(n2382), .A2(n2383), .A3(n2381), .ZN(n4529) );
  NAND2_X1 U2855 ( .A1(n2451), .A2(n2448), .ZN(n2385) );
  INV_X1 U2856 ( .A(n2384), .ZN(n4528) );
  NAND2_X1 U2857 ( .A1(n2385), .A2(n2908), .ZN(n2509) );
  INV_X1 U2858 ( .A(n2392), .ZN(n3807) );
  NAND2_X1 U2859 ( .A1(n3766), .A2(n2395), .ZN(n2393) );
  NAND3_X1 U2860 ( .A1(n4020), .A2(n3831), .A3(n3991), .ZN(n2396) );
  NAND2_X1 U2861 ( .A1(n3901), .A2(n2272), .ZN(n4150) );
  NAND2_X1 U2862 ( .A1(n3901), .A2(n2308), .ZN(n4152) );
  AND2_X1 U2863 ( .A1(n3901), .A2(n3906), .ZN(n3892) );
  NAND2_X1 U2864 ( .A1(n4080), .A2(n3823), .ZN(n4043) );
  AOI22_X1 U2865 ( .A1(n3885), .A2(n3886), .B1(n3842), .B2(n3841), .ZN(n3843)
         );
  AOI21_X1 U2866 ( .B1(n3747), .B2(n2409), .A(n2304), .ZN(n2410) );
  NAND2_X1 U2867 ( .A1(n2990), .A2(n2989), .ZN(n2991) );
  NAND2_X1 U2868 ( .A1(n4783), .A2(n3097), .ZN(n2417) );
  NOR2_X1 U2869 ( .A1(n2974), .A2(n2419), .ZN(n4632) );
  INV_X1 U2870 ( .A(n2421), .ZN(n4630) );
  NAND2_X1 U2871 ( .A1(n3749), .A2(REG1_REG_14__SCAN_IN), .ZN(n2431) );
  OAI21_X1 U2872 ( .B1(n4528), .B2(n2434), .A(REG2_REG_7__SCAN_IN), .ZN(n2964)
         );
  NAND2_X1 U2873 ( .A1(n4594), .A2(n2438), .ZN(n2437) );
  INV_X1 U2874 ( .A(n4466), .ZN(n2445) );
  NOR2_X1 U2875 ( .A1(n3759), .A2(REG2_REG_13__SCAN_IN), .ZN(n2446) );
  INV_X1 U2876 ( .A(n2962), .ZN(n2453) );
  NAND2_X1 U2877 ( .A1(n2451), .A2(n2449), .ZN(n4518) );
  NAND2_X1 U2878 ( .A1(n2962), .A2(n2450), .ZN(n2449) );
  NAND3_X1 U2879 ( .A1(n2607), .A2(n2514), .A3(n2455), .ZN(n2830) );
  INV_X1 U2880 ( .A(n2830), .ZN(n2516) );
  NAND2_X1 U2881 ( .A1(n3090), .A2(n2286), .ZN(n2456) );
  INV_X1 U2882 ( .A(n2459), .ZN(n3541) );
  NAND2_X1 U2883 ( .A1(n2464), .A2(n3172), .ZN(n2548) );
  INV_X2 U2884 ( .A(n3171), .ZN(n2464) );
  NAND2_X1 U2885 ( .A1(n2466), .A2(n2465), .ZN(n3295) );
  NAND2_X1 U2886 ( .A1(n3226), .A2(n2285), .ZN(n2466) );
  AOI21_X1 U2887 ( .B1(n3228), .B2(n3227), .A(n2475), .ZN(n2474) );
  NAND3_X1 U2888 ( .A1(n2477), .A2(n2274), .A3(n3240), .ZN(n2476) );
  INV_X1 U2889 ( .A(n2479), .ZN(n2477) );
  NOR2_X1 U2890 ( .A1(n3021), .A2(n2482), .ZN(n2481) );
  OAI211_X1 U2891 ( .C1(n3557), .C2(n2492), .A(n2489), .B(n2487), .ZN(n3474)
         );
  NAND2_X1 U2892 ( .A1(n3557), .A2(n2488), .ZN(n2487) );
  OAI21_X1 U2893 ( .B1(n2494), .B2(n2290), .A(n2490), .ZN(n2489) );
  NAND2_X1 U2894 ( .A1(n2494), .A2(n2491), .ZN(n2490) );
  AND2_X1 U2895 ( .A1(n2545), .A2(n2555), .ZN(n2534) );
  OAI21_X1 U2896 ( .B1(n4682), .B2(REG1_REG_2__SCAN_IN), .A(n2975), .ZN(n4631)
         );
  NAND2_X1 U2897 ( .A1(n4682), .A2(REG1_REG_2__SCAN_IN), .ZN(n2975) );
  OR2_X1 U2898 ( .A1(n2652), .A2(n2617), .ZN(n2619) );
  NOR2_X1 U2899 ( .A1(n3784), .A2(n3783), .ZN(n3785) );
  OAI21_X1 U2900 ( .B1(n3093), .B2(n4783), .A(n4575), .ZN(n3757) );
  NAND2_X1 U2901 ( .A1(n3748), .A2(n2445), .ZN(n3749) );
  NAND4_X1 U2902 ( .A1(n2651), .A2(n2506), .A3(n2650), .A4(n2649), .ZN(n2657)
         );
  NOR2_X1 U2903 ( .A1(n2621), .A2(n4635), .ZN(n2956) );
  OAI21_X1 U2904 ( .B1(n3594), .B2(n2652), .A(n2653), .ZN(n2805) );
  NAND2_X1 U2905 ( .A1(n3594), .A2(DATAI_0_), .ZN(n2633) );
  XNOR2_X1 U2906 ( .A(n2707), .B(n2708), .ZN(n2705) );
  AOI22_X1 U2907 ( .A1(n2657), .A2(n2736), .B1(n2263), .B2(n2805), .ZN(n2708)
         );
  XNOR2_X1 U2908 ( .A(n2656), .B(n3458), .ZN(n2707) );
  NAND2_X1 U2909 ( .A1(n3810), .A2(n4607), .ZN(n3811) );
  AOI21_X2 U2910 ( .B1(n3552), .B2(n3322), .A(n2299), .ZN(n3495) );
  NAND2_X2 U2911 ( .A1(n2803), .A2(n4741), .ZN(n4674) );
  INV_X2 U2912 ( .A(n4674), .ZN(n4939) );
  AND2_X1 U2913 ( .A1(n2575), .A2(n2574), .ZN(n2503) );
  AND3_X1 U2914 ( .A1(n2630), .A2(n2629), .A3(n2628), .ZN(n2504) );
  INV_X1 U2915 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3782) );
  AND2_X1 U2916 ( .A1(n3909), .A2(n3926), .ZN(n2505) );
  OR2_X1 U2917 ( .A1(n3802), .A2(n4205), .ZN(n2507) );
  OR2_X1 U2918 ( .A1(n3835), .A2(n3936), .ZN(n2508) );
  NAND4_X1 U2919 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3922)
         );
  INV_X1 U2920 ( .A(n3922), .ZN(n3840) );
  AND2_X1 U2921 ( .A1(n3700), .A2(n3987), .ZN(n4002) );
  INV_X1 U2922 ( .A(n4668), .ZN(n2570) );
  AND2_X1 U2923 ( .A1(n3584), .A2(n4044), .ZN(n3852) );
  INV_X1 U2924 ( .A(n3821), .ZN(n4082) );
  INV_X1 U2925 ( .A(n2614), .ZN(n2634) );
  INV_X1 U2926 ( .A(n3515), .ZN(n3287) );
  INV_X1 U2927 ( .A(n3808), .ZN(n3809) );
  OR2_X1 U2928 ( .A1(n4734), .A2(n3244), .ZN(n2510) );
  NOR2_X1 U2929 ( .A1(n4156), .A2(n4887), .ZN(n2511) );
  AND2_X1 U2930 ( .A1(n3280), .A2(n3279), .ZN(n4465) );
  NAND4_X1 U2931 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3960)
         );
  AND2_X1 U2932 ( .A1(n3833), .A2(n3968), .ZN(n2513) );
  INV_X1 U2933 ( .A(n3945), .ZN(n3936) );
  INV_X1 U2934 ( .A(IR_REG_19__SCAN_IN), .ZN(n2524) );
  INV_X1 U2935 ( .A(IR_REG_27__SCAN_IN), .ZN(n2574) );
  INV_X1 U2936 ( .A(n3975), .ZN(n3829) );
  NAND2_X1 U2937 ( .A1(n3993), .A2(n3959), .ZN(n3832) );
  NOR2_X1 U2938 ( .A1(n2767), .A2(n2638), .ZN(n2639) );
  OR2_X1 U2939 ( .A1(n3287), .A2(n3288), .ZN(n3293) );
  INV_X1 U2940 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2617) );
  AND2_X1 U2941 ( .A1(n4861), .A2(n3877), .ZN(n3686) );
  INV_X1 U2942 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3030) );
  INV_X1 U2943 ( .A(n4113), .ZN(n3877) );
  INV_X1 U2944 ( .A(n3621), .ZN(n2874) );
  INV_X1 U2945 ( .A(n3141), .ZN(n3142) );
  NOR2_X1 U2946 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  OR2_X1 U2947 ( .A1(n3449), .A2(n4408), .ZN(n3875) );
  NOR2_X1 U2948 ( .A1(n3875), .A2(n4741), .ZN(n3876) );
  AND2_X1 U2949 ( .A1(n4922), .A2(n4905), .ZN(n3827) );
  NOR2_X1 U2950 ( .A1(n3264), .A2(n4413), .ZN(n3296) );
  AND2_X1 U2951 ( .A1(n3131), .A2(REG3_REG_12__SCAN_IN), .ZN(n3151) );
  OR2_X1 U2952 ( .A1(n4788), .A2(n3177), .ZN(n3710) );
  INV_X1 U2953 ( .A(n3831), .ZN(n4008) );
  INV_X1 U2954 ( .A(n4798), .ZN(n3195) );
  INV_X1 U2955 ( .A(n2888), .ZN(n2880) );
  INV_X1 U2956 ( .A(n3742), .ZN(n2790) );
  NAND2_X1 U2957 ( .A1(n3415), .A2(n3414), .ZN(n3557) );
  AND2_X1 U2958 ( .A1(n3485), .A2(n3486), .ZN(n3387) );
  XNOR2_X1 U2959 ( .A(n3412), .B(n3458), .ZN(n3502) );
  NAND2_X1 U2960 ( .A1(n2776), .A2(n2777), .ZN(n2754) );
  NOR2_X1 U2961 ( .A1(n3324), .A2(n4405), .ZN(n3323) );
  AND2_X1 U2962 ( .A1(n2687), .A2(n4741), .ZN(n4834) );
  OR2_X1 U2963 ( .A1(n3451), .A2(n3947), .ZN(n3409) );
  INV_X1 U2964 ( .A(n4749), .ZN(n2984) );
  INV_X1 U2965 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U2966 ( .A1(n3835), .A2(n3936), .ZN(n3836) );
  AND2_X1 U2967 ( .A1(n3851), .A2(n3687), .ZN(n4118) );
  AND2_X1 U2968 ( .A1(n3731), .A2(n3613), .ZN(n2795) );
  OR2_X1 U2969 ( .A1(n3071), .A2(n4342), .ZN(n3095) );
  INV_X1 U2970 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2916) );
  OR2_X1 U2971 ( .A1(n4075), .A2(n4887), .ZN(n4934) );
  INV_X1 U2972 ( .A(n4125), .ZN(n4138) );
  AND2_X1 U2973 ( .A1(n3725), .A2(n2794), .ZN(n4856) );
  INV_X1 U2974 ( .A(n2572), .ZN(n2532) );
  OR2_X1 U2975 ( .A1(n2686), .A2(n3733), .ZN(n2609) );
  INV_X1 U2976 ( .A(n4834), .ZN(n4924) );
  AND4_X1 U2977 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3962)
         );
  AND2_X1 U2978 ( .A1(n4505), .A2(n2620), .ZN(n4607) );
  OR2_X1 U2979 ( .A1(n3864), .A2(n3863), .ZN(n3886) );
  INV_X1 U2980 ( .A(n4213), .ZN(n4849) );
  AND2_X1 U2981 ( .A1(n4932), .A2(n2795), .ZN(n4862) );
  INV_X1 U2982 ( .A(n4856), .ZN(n4731) );
  NOR2_X1 U2983 ( .A1(n4696), .A2(n3613), .ZN(n2933) );
  AND2_X1 U2984 ( .A1(n2662), .A2(n2661), .ZN(n2945) );
  OR3_X1 U2985 ( .A1(n2570), .A2(n3731), .A3(n3808), .ZN(n4696) );
  INV_X1 U2986 ( .A(n4879), .ZN(n4888) );
  INV_X1 U2987 ( .A(n4887), .ZN(n4883) );
  INV_X1 U2988 ( .A(n2945), .ZN(n2939) );
  AND2_X1 U2989 ( .A1(n2767), .A2(n3729), .ZN(n2686) );
  INV_X1 U2990 ( .A(n3721), .ZN(n3613) );
  AND2_X1 U2991 ( .A1(n2596), .A2(n2609), .ZN(n4646) );
  OR2_X1 U2992 ( .A1(n2692), .A2(n4637), .ZN(n4913) );
  NAND2_X1 U2993 ( .A1(n2691), .A2(n2679), .ZN(n3567) );
  NAND4_X1 U2994 ( .A1(n3422), .A2(n3421), .A3(n3420), .A4(n3419), .ZN(n3909)
         );
  NAND4_X1 U2995 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n4091)
         );
  INV_X1 U2996 ( .A(n4609), .ZN(n4647) );
  INV_X1 U2997 ( .A(n4656), .ZN(n4612) );
  AND2_X1 U2998 ( .A1(n3193), .A2(n3192), .ZN(n4826) );
  INV_X1 U2999 ( .A(n4894), .ZN(n4892) );
  AND2_X2 U3000 ( .A1(n2946), .A2(n2945), .ZN(n4894) );
  AND2_X1 U3001 ( .A1(n4826), .A2(n4825), .ZN(n4828) );
  INV_X1 U3002 ( .A(n4897), .ZN(n4895) );
  XNOR2_X1 U3003 ( .A(n2613), .B(n2612), .ZN(n4932) );
  INV_X1 U3004 ( .A(n4570), .ZN(n4783) );
  INV_X1 U3005 ( .A(n4655), .ZN(n4703) );
  NAND2_X1 U3006 ( .A1(n2516), .A2(n2515), .ZN(n2903) );
  INV_X1 U3007 ( .A(n2903), .ZN(n2521) );
  NAND2_X1 U3008 ( .A1(n2521), .A2(n2520), .ZN(n3171) );
  INV_X1 U3009 ( .A(n3273), .ZN(n2527) );
  NAND2_X1 U3010 ( .A1(n2530), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  MUX2_X1 U3011 ( .A(IR_REG_31__SCAN_IN), .B(n2531), .S(IR_REG_25__SCAN_IN), 
        .Z(n2533) );
  NAND2_X1 U3012 ( .A1(n2533), .A2(n2532), .ZN(n2585) );
  INV_X1 U3013 ( .A(n2534), .ZN(n2535) );
  INV_X1 U3014 ( .A(IR_REG_23__SCAN_IN), .ZN(n2536) );
  INV_X1 U3015 ( .A(n2538), .ZN(n2539) );
  NAND2_X1 U3016 ( .A1(n2539), .A2(IR_REG_23__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U3017 ( .A1(n2541), .A2(n2540), .ZN(n2766) );
  INV_X1 U3018 ( .A(n3729), .ZN(n2542) );
  OR2_X2 U3019 ( .A1(n2767), .A2(n2542), .ZN(n3741) );
  INV_X1 U3020 ( .A(n3741), .ZN(U4043) );
  INV_X2 U3021 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3022 ( .A(DATAI_21_), .ZN(n4363) );
  NAND2_X1 U3023 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2544) );
  MUX2_X1 U3024 ( .A(IR_REG_31__SCAN_IN), .B(n2544), .S(IR_REG_21__SCAN_IN), 
        .Z(n2546) );
  INV_X1 U3025 ( .A(n2545), .ZN(n2554) );
  NAND2_X1 U3026 ( .A1(n2546), .A2(n2554), .ZN(n3721) );
  NAND2_X1 U3027 ( .A1(n3613), .A2(STATE_REG_SCAN_IN), .ZN(n2547) );
  OAI21_X1 U3028 ( .B1(STATE_REG_SCAN_IN), .B2(n4363), .A(n2547), .ZN(U3331)
         );
  INV_X1 U3029 ( .A(DATAI_17_), .ZN(n2553) );
  NAND2_X1 U3030 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U3031 ( .A1(n3214), .A2(n2549), .ZN(n3278) );
  INV_X1 U3032 ( .A(IR_REG_17__SCAN_IN), .ZN(n2551) );
  XNOR2_X1 U3033 ( .A(n2561), .B(n2551), .ZN(n3805) );
  NAND2_X1 U3034 ( .A1(n3805), .A2(STATE_REG_SCAN_IN), .ZN(n2552) );
  OAI21_X1 U3035 ( .B1(STATE_REG_SCAN_IN), .B2(n2553), .A(n2552), .ZN(U3335)
         );
  INV_X1 U3036 ( .A(DATAI_22_), .ZN(n4261) );
  NAND2_X1 U3037 ( .A1(n2554), .A2(IR_REG_31__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U3038 ( .A1(n3731), .A2(STATE_REG_SCAN_IN), .ZN(n2557) );
  OAI21_X1 U3039 ( .B1(STATE_REG_SCAN_IN), .B2(n4261), .A(n2557), .ZN(U3330)
         );
  INV_X1 U3040 ( .A(DATAI_25_), .ZN(n2559) );
  NAND2_X1 U3041 ( .A1(n2675), .A2(STATE_REG_SCAN_IN), .ZN(n2558) );
  OAI21_X1 U3042 ( .B1(STATE_REG_SCAN_IN), .B2(n2559), .A(n2558), .ZN(U3327)
         );
  INV_X1 U3043 ( .A(DATAI_18_), .ZN(n4265) );
  INV_X1 U3044 ( .A(n2566), .ZN(n2563) );
  INV_X1 U3045 ( .A(IR_REG_18__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U3046 ( .A(n2563), .B(n2562), .ZN(n4621) );
  NAND2_X1 U3047 ( .A1(n4621), .A2(STATE_REG_SCAN_IN), .ZN(n2564) );
  OAI21_X1 U3048 ( .B1(STATE_REG_SCAN_IN), .B2(n4265), .A(n2564), .ZN(U3334)
         );
  INV_X1 U3049 ( .A(DATAI_20_), .ZN(n4249) );
  NAND2_X1 U3050 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U3051 ( .A1(n2566), .A2(n2565), .ZN(n2644) );
  NAND2_X1 U3052 ( .A1(n2570), .A2(STATE_REG_SCAN_IN), .ZN(n2571) );
  OAI21_X1 U3053 ( .B1(STATE_REG_SCAN_IN), .B2(n4249), .A(n2571), .ZN(U3332)
         );
  INV_X1 U3054 ( .A(DATAI_27_), .ZN(n4357) );
  XNOR2_X1 U3055 ( .A(n2592), .B(IR_REG_27__SCAN_IN), .ZN(n4639) );
  INV_X1 U3056 ( .A(n4639), .ZN(n4503) );
  NAND2_X1 U3057 ( .A1(n4503), .A2(STATE_REG_SCAN_IN), .ZN(n2573) );
  OAI21_X1 U3058 ( .B1(STATE_REG_SCAN_IN), .B2(n4357), .A(n2573), .ZN(U3325)
         );
  INV_X1 U3059 ( .A(DATAI_29_), .ZN(n4350) );
  NAND2_X1 U3060 ( .A1(n2597), .A2(STATE_REG_SCAN_IN), .ZN(n2578) );
  OAI21_X1 U3061 ( .B1(STATE_REG_SCAN_IN), .B2(n4350), .A(n2578), .ZN(U3323)
         );
  INV_X1 U3062 ( .A(DATAI_30_), .ZN(n2584) );
  INV_X1 U3063 ( .A(n2579), .ZN(n2580) );
  NAND2_X1 U3064 ( .A1(n2580), .A2(n2576), .ZN(n3203) );
  XNOR2_X2 U3065 ( .A(n2581), .B(n3200), .ZN(n2599) );
  INV_X1 U3066 ( .A(n2599), .ZN(n2582) );
  NAND2_X1 U3067 ( .A1(n2582), .A2(STATE_REG_SCAN_IN), .ZN(n2583) );
  OAI21_X1 U3068 ( .B1(STATE_REG_SCAN_IN), .B2(n2584), .A(n2583), .ZN(U3322)
         );
  NAND2_X1 U3069 ( .A1(n2585), .A2(B_REG_SCAN_IN), .ZN(n2586) );
  MUX2_X1 U3070 ( .A(n2586), .B(B_REG_SCAN_IN), .S(n4464), .Z(n2587) );
  INV_X1 U3071 ( .A(n2674), .ZN(n2588) );
  AND2_X2 U3072 ( .A1(n2588), .A2(n2686), .ZN(n4501) );
  INV_X1 U3073 ( .A(n4463), .ZN(n2660) );
  INV_X1 U3074 ( .A(n4464), .ZN(n2659) );
  NAND3_X1 U3075 ( .A1(n2660), .A2(n3729), .A3(n2659), .ZN(n2589) );
  OAI21_X1 U3076 ( .B1(n4501), .B2(D_REG_0__SCAN_IN), .A(n2589), .ZN(n2590) );
  INV_X1 U3077 ( .A(n2590), .ZN(U3458) );
  NAND2_X1 U3078 ( .A1(n2612), .A2(IR_REG_27__SCAN_IN), .ZN(n2593) );
  NAND2_X4 U3079 ( .A1(n2594), .A2(n2593), .ZN(n3594) );
  NAND2_X1 U3080 ( .A1(n2795), .A2(n2766), .ZN(n2595) );
  AND2_X1 U3081 ( .A1(n3594), .A2(n2595), .ZN(n2610) );
  INV_X1 U3082 ( .A(n2610), .ZN(n2596) );
  OR2_X1 U3083 ( .A1(n2766), .A2(U3149), .ZN(n4469) );
  INV_X1 U3084 ( .A(n4469), .ZN(n3733) );
  NOR2_X1 U3085 ( .A1(n4646), .A2(U4043), .ZN(U3148) );
  INV_X1 U3086 ( .A(n2600), .ZN(n2597) );
  OR2_X2 U3087 ( .A1(n2599), .A2(n2597), .ZN(n2693) );
  NAND2_X1 U3088 ( .A1(n3464), .A2(REG2_REG_22__SCAN_IN), .ZN(n2605) );
  INV_X1 U3089 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2598) );
  OR2_X1 U3090 ( .A1(n2259), .A2(n2598), .ZN(n2604) );
  NAND2_X1 U3091 ( .A1(n2843), .A2(REG3_REG_6__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U3092 ( .A1(n3009), .A2(REG3_REG_8__SCAN_IN), .ZN(n3031) );
  INV_X1 U3093 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4911) );
  INV_X1 U3094 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3370) );
  XNOR2_X1 U3095 ( .A(n3372), .B(n3370), .ZN(n4009) );
  OR2_X1 U3096 ( .A1(n3451), .A2(n4009), .ZN(n2603) );
  INV_X1 U3097 ( .A(REG0_REG_22__SCAN_IN), .ZN(n2601) );
  OR2_X1 U3098 ( .A1(n2740), .A2(n2601), .ZN(n2602) );
  NAND2_X1 U3099 ( .A1(n3741), .A2(DATAO_REG_22__SCAN_IN), .ZN(n2606) );
  OAI21_X1 U3100 ( .B1(n4912), .B2(n3741), .A(n2606), .ZN(U3572) );
  INV_X1 U3101 ( .A(n2607), .ZN(n2608) );
  NAND2_X1 U3102 ( .A1(n2611), .A2(IR_REG_31__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3103 ( .A1(n2614), .A2(REG1_REG_0__SCAN_IN), .ZN(n2616) );
  AOI211_X1 U3104 ( .C1(n2616), .C2(n2615), .A(n2974), .B(n4647), .ZN(n2623)
         );
  NAND2_X1 U3105 ( .A1(n2614), .A2(REG2_REG_0__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U3106 ( .A1(n2652), .A2(n2617), .ZN(n2618) );
  NAND2_X1 U3107 ( .A1(n2619), .A2(n2618), .ZN(n2621) );
  NOR2_X1 U3108 ( .A1(n4639), .A2(n4932), .ZN(n2620) );
  AOI211_X1 U3109 ( .C1(n4635), .C2(n2621), .A(n2956), .B(n4650), .ZN(n2622)
         );
  NOR2_X1 U3110 ( .A1(n2623), .A2(n2622), .ZN(n2625) );
  AOI22_X1 U3111 ( .A1(n4646), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n2624) );
  OAI211_X1 U3112 ( .C1(n2652), .C2(n4612), .A(n2625), .B(n2624), .ZN(U3241)
         );
  INV_X1 U3113 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2626) );
  OR2_X1 U3114 ( .A1(n2694), .A2(n2626), .ZN(n2631) );
  INV_X1 U3115 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2627) );
  OR2_X1 U3116 ( .A1(n2693), .A2(n2627), .ZN(n2629) );
  NAND2_X1 U3117 ( .A1(n2261), .A2(REG0_REG_0__SCAN_IN), .ZN(n2628) );
  NAND2_X2 U3118 ( .A1(n2632), .A2(n3613), .ZN(n2689) );
  AND2_X4 U3119 ( .A1(n2689), .A2(n2767), .ZN(n3345) );
  NAND2_X1 U3120 ( .A1(n3742), .A2(n2736), .ZN(n2637) );
  NOR2_X1 U3121 ( .A1(n2767), .A2(n2634), .ZN(n2635) );
  AOI21_X1 U3122 ( .B1(n4664), .B2(n3437), .A(n2635), .ZN(n2636) );
  NAND2_X1 U3123 ( .A1(n4664), .A2(n3345), .ZN(n2646) );
  INV_X1 U3124 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3125 ( .A1(n3256), .A2(n3257), .ZN(n2648) );
  NAND2_X1 U3126 ( .A1(n2644), .A2(IR_REG_19__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3127 ( .A1(n3808), .A2(n3731), .ZN(n2688) );
  NAND2_X4 U3128 ( .A1(n2689), .A2(n2688), .ZN(n3458) );
  NAND2_X1 U3129 ( .A1(n2646), .A2(n3440), .ZN(n2647) );
  NAND2_X1 U3130 ( .A1(n2648), .A2(n2647), .ZN(n2706) );
  INV_X1 U3131 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2817) );
  NAND2_X1 U3132 ( .A1(n2657), .A2(n2262), .ZN(n2655) );
  INV_X1 U3133 ( .A(n2652), .ZN(n4468) );
  NAND2_X1 U3134 ( .A1(n3594), .A2(DATAI_1_), .ZN(n2653) );
  NAND2_X1 U3135 ( .A1(n2805), .A2(n3345), .ZN(n2654) );
  NAND2_X1 U3136 ( .A1(n2655), .A2(n2654), .ZN(n2656) );
  XNOR2_X1 U3137 ( .A(n2706), .B(n2705), .ZN(n2704) );
  INV_X1 U3138 ( .A(D_REG_0__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3139 ( .A1(n2674), .A2(n2658), .ZN(n2662) );
  NAND2_X1 U3140 ( .A1(n2660), .A2(n2659), .ZN(n2661) );
  NOR4_X1 U3141 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2671) );
  NOR4_X1 U3142 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2670) );
  INV_X1 U3143 ( .A(D_REG_31__SCAN_IN), .ZN(n4500) );
  INV_X1 U3144 ( .A(D_REG_30__SCAN_IN), .ZN(n4499) );
  INV_X1 U3145 ( .A(D_REG_29__SCAN_IN), .ZN(n4498) );
  INV_X1 U3146 ( .A(D_REG_28__SCAN_IN), .ZN(n4497) );
  NAND4_X1 U3147 ( .A1(n4500), .A2(n4499), .A3(n4498), .A4(n4497), .ZN(n2668)
         );
  NOR4_X1 U31480 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2666) );
  NOR4_X1 U31490 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2665) );
  NOR4_X1 U3150 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2664) );
  NOR4_X1 U3151 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2663) );
  NAND4_X1 U3152 ( .A1(n2666), .A2(n2665), .A3(n2664), .A4(n2663), .ZN(n2667)
         );
  NOR4_X1 U3153 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(n2668), 
        .A4(n2667), .ZN(n2669) );
  NAND3_X1 U3154 ( .A1(n2671), .A2(n2670), .A3(n2669), .ZN(n2672) );
  AND2_X1 U3155 ( .A1(n2674), .A2(n2672), .ZN(n2936) );
  INV_X1 U3156 ( .A(D_REG_1__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3157 ( .A1(n2674), .A2(n2673), .ZN(n2676) );
  OR2_X1 U3158 ( .A1(n2675), .A2(n4463), .ZN(n4462) );
  NAND2_X1 U3159 ( .A1(n2676), .A2(n4462), .ZN(n2937) );
  NOR2_X1 U3160 ( .A1(n2936), .A2(n2937), .ZN(n2677) );
  INV_X1 U3161 ( .A(n2686), .ZN(n2678) );
  NAND2_X1 U3162 ( .A1(n4668), .A2(n3808), .ZN(n2681) );
  AOI21_X1 U3163 ( .B1(n2681), .B2(n4663), .A(n2795), .ZN(n2679) );
  NAND2_X1 U3164 ( .A1(n2570), .A2(n4663), .ZN(n4853) );
  NOR3_X1 U3165 ( .A1(n2680), .A2(U3149), .A3(n4853), .ZN(n2769) );
  INV_X1 U3166 ( .A(n2769), .ZN(n2685) );
  NAND2_X1 U3167 ( .A1(n2681), .A2(n2795), .ZN(n2765) );
  NAND2_X1 U3168 ( .A1(n2686), .A2(n2765), .ZN(n2934) );
  INV_X1 U3169 ( .A(n2934), .ZN(n2684) );
  INV_X1 U3170 ( .A(n4663), .ZN(n2683) );
  OAI21_X1 U3171 ( .B1(n3808), .B2(n2683), .A(n2682), .ZN(n2768) );
  NAND3_X1 U3172 ( .A1(n2685), .A2(n2684), .A3(n2768), .ZN(n3258) );
  NAND2_X1 U3173 ( .A1(n2691), .A2(n4787), .ZN(n2687) );
  INV_X1 U3174 ( .A(n2805), .ZN(n2785) );
  NOR2_X1 U3175 ( .A1(n4834), .A2(n2785), .ZN(n2702) );
  NOR2_X1 U3176 ( .A1(n2689), .A2(n2688), .ZN(n2690) );
  NAND2_X1 U3177 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U3178 ( .A1(n2261), .A2(REG0_REG_2__SCAN_IN), .ZN(n2698) );
  INV_X1 U3179 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2858) );
  INV_X1 U3180 ( .A(n3740), .ZN(n2700) );
  OAI22_X1 U3181 ( .A1(n2790), .A2(n4830), .B1(n4913), .B2(n2700), .ZN(n2701)
         );
  AOI211_X1 U3182 ( .C1(REG3_REG_1__SCAN_IN), .C2(n3258), .A(n2702), .B(n2701), 
        .ZN(n2703) );
  OAI21_X1 U3183 ( .B1(n2704), .B2(n3567), .A(n2703), .ZN(U3219) );
  NAND2_X1 U3184 ( .A1(n2706), .A2(n2705), .ZN(n2711) );
  INV_X1 U3185 ( .A(n2707), .ZN(n2709) );
  OR2_X1 U3186 ( .A1(n2709), .A2(n2708), .ZN(n2710) );
  NAND2_X1 U3187 ( .A1(n2711), .A2(n2710), .ZN(n3248) );
  INV_X1 U3188 ( .A(n3248), .ZN(n2720) );
  NAND2_X1 U3189 ( .A1(n3740), .A2(n2263), .ZN(n2714) );
  MUX2_X1 U3190 ( .A(n4682), .B(DATAI_2_), .S(n3594), .Z(n3252) );
  NAND2_X1 U3191 ( .A1(n3252), .A2(n3345), .ZN(n2713) );
  NAND2_X1 U3192 ( .A1(n2714), .A2(n2713), .ZN(n2715) );
  XNOR2_X1 U3193 ( .A(n2715), .B(n3440), .ZN(n2717) );
  AOI22_X1 U3194 ( .A1(n3740), .A2(n2736), .B1(n3437), .B2(n3252), .ZN(n2716)
         );
  NAND2_X1 U3195 ( .A1(n2717), .A2(n2716), .ZN(n2721) );
  OR2_X1 U3196 ( .A1(n2717), .A2(n2716), .ZN(n2718) );
  NAND2_X1 U3197 ( .A1(n2721), .A2(n2718), .ZN(n3251) );
  INV_X1 U3198 ( .A(n3251), .ZN(n2719) );
  NAND2_X1 U3199 ( .A1(n2720), .A2(n2719), .ZN(n3249) );
  NAND2_X1 U3200 ( .A1(n3249), .A2(n2721), .ZN(n2776) );
  INV_X1 U3201 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2722) );
  OR2_X1 U3202 ( .A1(n2693), .A2(n2722), .ZN(n2726) );
  INV_X1 U3203 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3204 ( .A1(n2757), .A2(n3437), .ZN(n2734) );
  NAND2_X1 U3205 ( .A1(n2607), .A2(n4431), .ZN(n2728) );
  NAND2_X1 U3206 ( .A1(n2728), .A2(IR_REG_31__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3207 ( .A1(n2730), .A2(n2729), .ZN(n2745) );
  OR2_X1 U3208 ( .A1(n2730), .A2(n2729), .ZN(n2731) );
  NAND2_X1 U3209 ( .A1(n2745), .A2(n2731), .ZN(n4694) );
  INV_X1 U32100 ( .A(n4694), .ZN(n2732) );
  MUX2_X1 U32110 ( .A(n2732), .B(DATAI_3_), .S(n3594), .Z(n3621) );
  NAND2_X1 U32120 ( .A1(n3621), .A2(n3345), .ZN(n2733) );
  NAND2_X1 U32130 ( .A1(n2734), .A2(n2733), .ZN(n2735) );
  AOI22_X1 U32140 ( .A1(n2757), .A2(n2736), .B1(n2263), .B2(n3621), .ZN(n2751)
         );
  XNOR2_X1 U32150 ( .A(n2750), .B(n2751), .ZN(n2777) );
  NAND2_X1 U32160 ( .A1(n2737), .A2(REG1_REG_4__SCAN_IN), .ZN(n2744) );
  INV_X1 U32170 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2738) );
  OR2_X1 U32180 ( .A1(n2693), .A2(n2738), .ZN(n2743) );
  XNOR2_X1 U32190 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(
        n2882) );
  OR2_X1 U32200 ( .A1(n2694), .A2(n2882), .ZN(n2742) );
  INV_X1 U32210 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2739) );
  OR2_X1 U32220 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  NAND2_X1 U32230 ( .A1(n2778), .A2(n3437), .ZN(n2748) );
  NAND2_X1 U32240 ( .A1(n2745), .A2(IR_REG_31__SCAN_IN), .ZN(n2746) );
  XNOR2_X1 U32250 ( .A(n2746), .B(IR_REG_4__SCAN_IN), .ZN(n4655) );
  MUX2_X1 U32260 ( .A(n4655), .B(DATAI_4_), .S(n3594), .Z(n2888) );
  NAND2_X1 U32270 ( .A1(n2888), .A2(n3345), .ZN(n2747) );
  NAND2_X1 U32280 ( .A1(n2748), .A2(n2747), .ZN(n2749) );
  AOI22_X1 U32290 ( .A1(n2778), .A2(n2736), .B1(n3437), .B2(n2888), .ZN(n2826)
         );
  XNOR2_X1 U32300 ( .A(n2825), .B(n2826), .ZN(n2755) );
  INV_X1 U32310 ( .A(n2750), .ZN(n2752) );
  NAND2_X1 U32320 ( .A1(n2752), .A2(n2751), .ZN(n2756) );
  AND2_X1 U32330 ( .A1(n2755), .A2(n2756), .ZN(n2753) );
  NAND2_X1 U32340 ( .A1(n2754), .A2(n2753), .ZN(n2829) );
  NAND2_X1 U32350 ( .A1(n2829), .A2(n4925), .ZN(n2775) );
  AOI21_X1 U32360 ( .B1(n2754), .B2(n2756), .A(n2755), .ZN(n2774) );
  INV_X1 U32370 ( .A(n2694), .ZN(n2915) );
  AOI21_X1 U32380 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2758) );
  NOR2_X1 U32390 ( .A1(n2758), .A2(n2843), .ZN(n2898) );
  NAND2_X1 U32400 ( .A1(n2915), .A2(n2898), .ZN(n2764) );
  INV_X1 U32410 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2759) );
  OR2_X1 U32420 ( .A1(n2740), .A2(n2759), .ZN(n2763) );
  OR2_X1 U32430 ( .A1(n2693), .A2(n2963), .ZN(n2762) );
  INV_X1 U32440 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2760) );
  OR2_X1 U32450 ( .A1(n2259), .A2(n2760), .ZN(n2761) );
  NAND4_X1 U32460 ( .A1(n2764), .A2(n2763), .A3(n2762), .A4(n2761), .ZN(n3739)
         );
  AOI22_X1 U32470 ( .A1(n4921), .A2(n2757), .B1(n4899), .B2(n3739), .ZN(n2773)
         );
  INV_X1 U32480 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4423) );
  NOR2_X1 U32490 ( .A1(STATE_REG_SCAN_IN), .A2(n4423), .ZN(n4645) );
  NAND4_X1 U32500 ( .A1(n2768), .A2(n2767), .A3(n2766), .A4(n2765), .ZN(n2770)
         );
  AOI21_X2 U32510 ( .B1(STATE_REG_SCAN_IN), .B2(n2770), .A(n2769), .ZN(n4930)
         );
  NOR2_X1 U32520 ( .A1(n4930), .A2(n2882), .ZN(n2771) );
  AOI211_X1 U32530 ( .C1(n2888), .C2(n4924), .A(n4645), .B(n2771), .ZN(n2772)
         );
  OAI211_X1 U32540 ( .C1(n2775), .C2(n2774), .A(n2773), .B(n2772), .ZN(U3227)
         );
  OAI21_X1 U32550 ( .B1(n2777), .B2(n2776), .A(n2754), .ZN(n2782) );
  AOI22_X1 U32560 ( .A1(n4921), .A2(n3740), .B1(n4899), .B2(n2778), .ZN(n2780)
         );
  INV_X1 U32570 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4401) );
  NOR2_X1 U32580 ( .A1(STATE_REG_SCAN_IN), .A2(n4401), .ZN(n4511) );
  AOI21_X1 U32590 ( .B1(n4924), .B2(n3621), .A(n4511), .ZN(n2779) );
  OAI211_X1 U32600 ( .C1(n4930), .C2(REG3_REG_3__SCAN_IN), .A(n2780), .B(n2779), .ZN(n2781) );
  AOI21_X1 U32610 ( .B1(n2782), .B2(n4925), .A(n2781), .ZN(n2783) );
  INV_X1 U32620 ( .A(n2783), .ZN(U3215) );
  INV_X1 U32630 ( .A(n2657), .ZN(n2784) );
  NAND2_X1 U32640 ( .A1(n2657), .A2(n2785), .ZN(n3612) );
  AND2_X1 U32650 ( .A1(n3742), .A2(n4664), .ZN(n2814) );
  NAND2_X1 U32660 ( .A1(n2657), .A2(n2805), .ZN(n2786) );
  INV_X1 U32670 ( .A(n3252), .ZN(n2864) );
  OR2_X1 U32680 ( .A1(n3740), .A2(n2864), .ZN(n3616) );
  NAND2_X1 U32690 ( .A1(n3740), .A2(n2864), .ZN(n3618) );
  OR2_X1 U32700 ( .A1(n3740), .A2(n3252), .ZN(n2787) );
  XNOR2_X1 U32710 ( .A(n2757), .B(n3621), .ZN(n3691) );
  XNOR2_X1 U32720 ( .A(n2873), .B(n3691), .ZN(n4697) );
  XNOR2_X1 U32730 ( .A(n2788), .B(n2793), .ZN(n2789) );
  NAND2_X1 U32740 ( .A1(n2789), .A2(n3808), .ZN(n4660) );
  INV_X1 U32750 ( .A(n4664), .ZN(n3611) );
  NAND2_X1 U32760 ( .A1(n3692), .A2(n3614), .ZN(n2818) );
  NAND2_X1 U32770 ( .A1(n2818), .A2(n3615), .ZN(n2791) );
  INV_X1 U32780 ( .A(n2860), .ZN(n3693) );
  NAND2_X1 U32790 ( .A1(n2791), .A2(n3693), .ZN(n2859) );
  NAND2_X1 U32800 ( .A1(n2859), .A2(n3616), .ZN(n2792) );
  NAND2_X1 U32810 ( .A1(n2792), .A2(n3691), .ZN(n2875) );
  OAI21_X1 U32820 ( .B1(n3691), .B2(n2792), .A(n2875), .ZN(n2799) );
  NAND2_X1 U32830 ( .A1(n2570), .A2(n3613), .ZN(n3725) );
  OR2_X1 U32840 ( .A1(n3808), .A2(n2793), .ZN(n2794) );
  INV_X1 U32850 ( .A(n2778), .ZN(n2797) );
  NAND2_X1 U32860 ( .A1(n4637), .A2(n2795), .ZN(n4213) );
  AOI22_X1 U32870 ( .A1(n3740), .A2(n4849), .B1(n4787), .B2(n3621), .ZN(n2796)
         );
  OAI21_X1 U32880 ( .B1(n2797), .B2(n4737), .A(n2796), .ZN(n2798) );
  AOI21_X1 U32890 ( .B1(n2799), .B2(n4731), .A(n2798), .ZN(n2800) );
  OAI21_X1 U32900 ( .B1(n4697), .B2(n4660), .A(n2800), .ZN(n4699) );
  INV_X1 U32910 ( .A(n4699), .ZN(n2811) );
  INV_X1 U32920 ( .A(n2937), .ZN(n2802) );
  NOR2_X1 U32930 ( .A1(n2936), .A2(n2934), .ZN(n2801) );
  NAND3_X1 U32940 ( .A1(n2939), .A2(n2802), .A3(n2801), .ZN(n2803) );
  INV_X1 U32950 ( .A(n4697), .ZN(n2809) );
  NAND2_X1 U32960 ( .A1(n2788), .A2(n3809), .ZN(n2816) );
  INV_X1 U32970 ( .A(n2816), .ZN(n2804) );
  NOR2_X1 U32980 ( .A1(n2855), .A2(n2874), .ZN(n2806) );
  OR2_X1 U32990 ( .A1(n2881), .A2(n2806), .ZN(n4695) );
  NAND2_X1 U33000 ( .A1(n4674), .A2(n3808), .ZN(n4075) );
  INV_X1 U33010 ( .A(n4741), .ZN(n4867) );
  AOI22_X1 U33020 ( .A1(n4939), .A2(REG2_REG_3__SCAN_IN), .B1(n4867), .B2(
        n4401), .ZN(n2807) );
  OAI21_X1 U33030 ( .B1(n4695), .B2(n4934), .A(n2807), .ZN(n2808) );
  AOI21_X1 U33040 ( .B1(n2809), .B2(n4805), .A(n2808), .ZN(n2810) );
  OAI21_X1 U33050 ( .B1(n2811), .B2(n4939), .A(n2810), .ZN(U3287) );
  NAND2_X1 U33060 ( .A1(n4664), .A2(n2805), .ZN(n2812) );
  AND2_X1 U33070 ( .A1(n2856), .A2(n2812), .ZN(n4679) );
  OAI21_X1 U33080 ( .B1(n2815), .B2(n2814), .A(n2813), .ZN(n4676) );
  NAND2_X1 U33090 ( .A1(n4660), .A2(n2816), .ZN(n4727) );
  OAI22_X1 U33100 ( .A1(n4676), .A2(n4140), .B1(n2817), .B2(n4741), .ZN(n2823)
         );
  OAI21_X1 U33110 ( .B1(n3692), .B2(n3614), .A(n2818), .ZN(n2819) );
  NAND2_X1 U33120 ( .A1(n2819), .A2(n4731), .ZN(n2821) );
  AOI22_X1 U33130 ( .A1(n3740), .A2(n4862), .B1(n4787), .B2(n2805), .ZN(n2820)
         );
  OAI211_X1 U33140 ( .C1(n2790), .C2(n4213), .A(n2821), .B(n2820), .ZN(n4677)
         );
  MUX2_X1 U33150 ( .A(n4677), .B(REG2_REG_1__SCAN_IN), .S(n4939), .Z(n2822) );
  AOI211_X1 U33160 ( .C1(n4940), .C2(n4679), .A(n2823), .B(n2822), .ZN(n2824)
         );
  INV_X1 U33170 ( .A(n2824), .ZN(U3289) );
  INV_X1 U33180 ( .A(n2825), .ZN(n2827) );
  OR2_X1 U33190 ( .A1(n2827), .A2(n2826), .ZN(n2828) );
  NAND2_X1 U33200 ( .A1(n2829), .A2(n2828), .ZN(n2995) );
  NAND2_X1 U33210 ( .A1(n3739), .A2(n3437), .ZN(n2833) );
  NAND2_X1 U33220 ( .A1(n2830), .A2(IR_REG_31__SCAN_IN), .ZN(n2831) );
  XNOR2_X1 U33230 ( .A(n2831), .B(IR_REG_5__SCAN_IN), .ZN(n2981) );
  MUX2_X1 U33240 ( .A(n2981), .B(DATAI_5_), .S(n3594), .Z(n2909) );
  NAND2_X1 U33250 ( .A1(n2909), .A2(n3345), .ZN(n2832) );
  NAND2_X1 U33260 ( .A1(n2833), .A2(n2832), .ZN(n2834) );
  XNOR2_X1 U33270 ( .A(n2834), .B(n3458), .ZN(n2840) );
  INV_X1 U33280 ( .A(n2840), .ZN(n2838) );
  NAND2_X1 U33290 ( .A1(n3739), .A2(n2736), .ZN(n2836) );
  NAND2_X1 U33300 ( .A1(n2909), .A2(n3437), .ZN(n2835) );
  NAND2_X1 U33310 ( .A1(n2836), .A2(n2835), .ZN(n2839) );
  INV_X1 U33320 ( .A(n2839), .ZN(n2837) );
  NAND2_X1 U33330 ( .A1(n2838), .A2(n2837), .ZN(n2999) );
  INV_X1 U33340 ( .A(n2999), .ZN(n2841) );
  AND2_X1 U33350 ( .A1(n2840), .A2(n2839), .ZN(n2996) );
  NOR2_X1 U33360 ( .A1(n2841), .A2(n2996), .ZN(n2842) );
  XNOR2_X1 U33370 ( .A(n2995), .B(n2842), .ZN(n2852) );
  NAND2_X1 U33380 ( .A1(n2737), .A2(REG1_REG_6__SCAN_IN), .ZN(n2848) );
  INV_X1 U33390 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2928) );
  OR2_X1 U33400 ( .A1(n2693), .A2(n2928), .ZN(n2847) );
  OAI21_X1 U33410 ( .B1(n2843), .B2(REG3_REG_6__SCAN_IN), .A(n2917), .ZN(n3242) );
  OR2_X1 U33420 ( .A1(n3451), .A2(n3242), .ZN(n2846) );
  INV_X1 U33430 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2844) );
  OR2_X1 U33440 ( .A1(n2740), .A2(n2844), .ZN(n2845) );
  NAND4_X1 U33450 ( .A1(n2848), .A2(n2847), .A3(n2846), .A4(n2845), .ZN(n4734)
         );
  AOI22_X1 U33460 ( .A1(n4899), .A2(n4734), .B1(n4921), .B2(n2778), .ZN(n2851)
         );
  INV_X1 U33470 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4338) );
  NOR2_X1 U33480 ( .A1(STATE_REG_SCAN_IN), .A2(n4338), .ZN(n4520) );
  INV_X1 U33490 ( .A(n2909), .ZN(n2891) );
  NOR2_X1 U33500 ( .A1(n4834), .A2(n2891), .ZN(n2849) );
  AOI211_X1 U33510 ( .C1(n3565), .C2(n2898), .A(n4520), .B(n2849), .ZN(n2850)
         );
  OAI211_X1 U33520 ( .C1(n2852), .C2(n3567), .A(n2851), .B(n2850), .ZN(U3224)
         );
  OAI21_X1 U3353 ( .B1(n2853), .B2(n2860), .A(n2854), .ZN(n4689) );
  INV_X1 U33540 ( .A(n2855), .ZN(n4686) );
  NAND2_X1 U3355 ( .A1(n2856), .A2(n3252), .ZN(n4685) );
  NAND3_X1 U3356 ( .A1(n4940), .A2(n4686), .A3(n4685), .ZN(n2857) );
  OAI21_X1 U3357 ( .B1(n4741), .B2(n2858), .A(n2857), .ZN(n2870) );
  NAND3_X1 U3358 ( .A1(n2818), .A2(n2860), .A3(n3615), .ZN(n2861) );
  NAND2_X1 U3359 ( .A1(n2859), .A2(n2861), .ZN(n2866) );
  NAND2_X1 U3360 ( .A1(n2757), .A2(n4862), .ZN(n2863) );
  NAND2_X1 U3361 ( .A1(n2657), .A2(n4849), .ZN(n2862) );
  OAI211_X1 U3362 ( .C1(n4853), .C2(n2864), .A(n2863), .B(n2862), .ZN(n2865)
         );
  AOI21_X1 U3363 ( .B1(n2866), .B2(n4731), .A(n2865), .ZN(n2868) );
  INV_X1 U3364 ( .A(n4660), .ZN(n4794) );
  NAND2_X1 U3365 ( .A1(n4689), .A2(n4794), .ZN(n2867) );
  NAND2_X1 U3366 ( .A1(n2868), .A2(n2867), .ZN(n4687) );
  MUX2_X1 U3367 ( .A(REG2_REG_2__SCAN_IN), .B(n4687), .S(n4674), .Z(n2869) );
  AOI211_X1 U3368 ( .C1(n4805), .C2(n4689), .A(n2870), .B(n2869), .ZN(n2871)
         );
  INV_X1 U3369 ( .A(n2871), .ZN(U3288) );
  NOR2_X1 U3370 ( .A1(n2757), .A2(n3621), .ZN(n2872) );
  INV_X1 U3371 ( .A(n2757), .ZN(n3620) );
  OR2_X1 U3372 ( .A1(n2778), .A2(n2880), .ZN(n3623) );
  NAND2_X1 U3373 ( .A1(n2778), .A2(n2880), .ZN(n3626) );
  NAND2_X1 U3374 ( .A1(n3623), .A2(n3626), .ZN(n3699) );
  XNOR2_X1 U3375 ( .A(n2887), .B(n3699), .ZN(n2884) );
  OAI22_X1 U3376 ( .A1(n3620), .A2(n4213), .B1(n2880), .B2(n4853), .ZN(n2878)
         );
  OR2_X1 U3377 ( .A1(n2757), .A2(n2874), .ZN(n3622) );
  NAND2_X1 U3378 ( .A1(n2875), .A2(n3622), .ZN(n2892) );
  XNOR2_X1 U3379 ( .A(n2892), .B(n3699), .ZN(n2876) );
  NOR2_X1 U3380 ( .A1(n2876), .A2(n4856), .ZN(n2877) );
  AOI211_X1 U3381 ( .C1(n4862), .C2(n3739), .A(n2878), .B(n2877), .ZN(n2879)
         );
  OAI21_X1 U3382 ( .B1(n4660), .B2(n2884), .A(n2879), .ZN(n4705) );
  NAND2_X1 U3383 ( .A1(n2881), .A2(n2880), .ZN(n2896) );
  OAI211_X1 U3384 ( .C1(n2881), .C2(n2880), .A(n4883), .B(n2896), .ZN(n4704)
         );
  OAI22_X1 U3385 ( .A1(n4704), .A2(n3809), .B1(n4741), .B2(n2882), .ZN(n2883)
         );
  OAI21_X1 U3386 ( .B1(n4705), .B2(n2883), .A(n4674), .ZN(n2886) );
  INV_X1 U3387 ( .A(n2884), .ZN(n4707) );
  AOI22_X1 U3388 ( .A1(n4707), .A2(n4805), .B1(REG2_REG_4__SCAN_IN), .B2(n4939), .ZN(n2885) );
  NAND2_X1 U3389 ( .A1(n2886), .A2(n2885), .ZN(U3286) );
  NAND2_X1 U3390 ( .A1(n2887), .A2(n3699), .ZN(n2890) );
  NAND2_X1 U3391 ( .A1(n2778), .A2(n2888), .ZN(n2889) );
  AND2_X1 U3392 ( .A1(n3739), .A2(n2891), .ZN(n2912) );
  INV_X1 U3393 ( .A(n2912), .ZN(n3625) );
  OR2_X1 U3394 ( .A1(n3739), .A2(n2891), .ZN(n3639) );
  NAND2_X1 U3395 ( .A1(n3625), .A2(n3639), .ZN(n3695) );
  XNOR2_X1 U3396 ( .A(n2911), .B(n3695), .ZN(n4712) );
  XOR2_X1 U3397 ( .A(n3695), .B(n2913), .Z(n2895) );
  AOI22_X1 U3398 ( .A1(n2778), .A2(n4849), .B1(n2909), .B2(n4787), .ZN(n2894)
         );
  NAND2_X1 U3399 ( .A1(n4734), .A2(n4862), .ZN(n2893) );
  OAI211_X1 U3400 ( .C1(n2895), .C2(n4856), .A(n2894), .B(n2893), .ZN(n4713)
         );
  NAND2_X1 U3401 ( .A1(n4713), .A2(n4674), .ZN(n2902) );
  AOI21_X1 U3402 ( .B1(n2909), .B2(n2896), .A(n2897), .ZN(n4715) );
  INV_X1 U3403 ( .A(n2898), .ZN(n2899) );
  OAI22_X1 U3404 ( .A1(n4674), .A2(n2963), .B1(n2899), .B2(n4741), .ZN(n2900)
         );
  AOI21_X1 U3405 ( .B1(n4715), .B2(n4940), .A(n2900), .ZN(n2901) );
  OAI211_X1 U3406 ( .C1(n4712), .C2(n4140), .A(n2902), .B(n2901), .ZN(U3285)
         );
  NAND2_X1 U3407 ( .A1(n2905), .A2(IR_REG_31__SCAN_IN), .ZN(n2904) );
  MUX2_X1 U3408 ( .A(IR_REG_31__SCAN_IN), .B(n2904), .S(IR_REG_6__SCAN_IN), 
        .Z(n2907) );
  NOR2_X1 U3409 ( .A1(n2905), .A2(IR_REG_6__SCAN_IN), .ZN(n2955) );
  INV_X1 U3410 ( .A(n2955), .ZN(n2906) );
  NAND2_X1 U3411 ( .A1(n2907), .A2(n2906), .ZN(n4718) );
  INV_X1 U3412 ( .A(n4718), .ZN(n2908) );
  MUX2_X1 U3413 ( .A(n2908), .B(DATAI_6_), .S(n3594), .Z(n3244) );
  INV_X1 U3414 ( .A(n3244), .ZN(n2927) );
  OR2_X1 U3415 ( .A1(n4734), .A2(n2927), .ZN(n3628) );
  NAND2_X1 U3416 ( .A1(n4734), .A2(n2927), .ZN(n3638) );
  NAND2_X1 U3417 ( .A1(n3628), .A2(n3638), .ZN(n3698) );
  AND2_X1 U3418 ( .A1(n3739), .A2(n2909), .ZN(n2910) );
  XOR2_X1 U3419 ( .A(n3698), .B(n3042), .Z(n2941) );
  XNOR2_X1 U3420 ( .A(n3048), .B(n3698), .ZN(n2926) );
  AOI22_X1 U3421 ( .A1(n3739), .A2(n4849), .B1(n4787), .B2(n3244), .ZN(n2925)
         );
  NAND2_X1 U3422 ( .A1(n3464), .A2(REG2_REG_7__SCAN_IN), .ZN(n2923) );
  INV_X1 U3423 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2914) );
  OR2_X1 U3424 ( .A1(n2259), .A2(n2914), .ZN(n2922) );
  INV_X1 U3425 ( .A(n2915), .ZN(n3451) );
  AND2_X1 U3426 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  OR2_X1 U3427 ( .A1(n2918), .A2(n3009), .ZN(n4742) );
  OR2_X1 U3428 ( .A1(n3451), .A2(n4742), .ZN(n2921) );
  INV_X1 U3429 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2919) );
  OR2_X1 U3430 ( .A1(n2740), .A2(n2919), .ZN(n2920) );
  NAND4_X1 U3431 ( .A1(n2923), .A2(n2922), .A3(n2921), .A4(n2920), .ZN(n3738)
         );
  NAND2_X1 U3432 ( .A1(n3738), .A2(n4862), .ZN(n2924) );
  OAI211_X1 U3433 ( .C1(n2926), .C2(n4856), .A(n2925), .B(n2924), .ZN(n2942)
         );
  NAND2_X1 U3434 ( .A1(n2942), .A2(n4674), .ZN(n2932) );
  OAI21_X1 U3435 ( .B1(n2897), .B2(n2927), .A(n4722), .ZN(n2940) );
  INV_X1 U3436 ( .A(n2940), .ZN(n2930) );
  OAI22_X1 U3437 ( .A1(n4674), .A2(n2928), .B1(n3242), .B2(n4741), .ZN(n2929)
         );
  AOI21_X1 U3438 ( .B1(n2930), .B2(n4940), .A(n2929), .ZN(n2931) );
  OAI211_X1 U3439 ( .C1(n2941), .C2(n4140), .A(n2932), .B(n2931), .ZN(U3284)
         );
  OR2_X1 U3440 ( .A1(n2934), .A2(n2933), .ZN(n2935) );
  NOR2_X1 U3441 ( .A1(n2936), .A2(n2935), .ZN(n2938) );
  NAND2_X1 U3442 ( .A1(n4660), .A2(n4696), .ZN(n4879) );
  OAI22_X1 U3443 ( .A1(n2941), .A2(n4888), .B1(n4887), .B2(n2940), .ZN(n2943)
         );
  OR2_X1 U3444 ( .A1(n2943), .A2(n2942), .ZN(n2947) );
  NAND2_X1 U3445 ( .A1(n2947), .A2(n4897), .ZN(n2944) );
  OAI21_X1 U3446 ( .B1(n4897), .B2(n2844), .A(n2944), .ZN(U3479) );
  INV_X1 U3447 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U3448 ( .A1(n2947), .A2(n4894), .ZN(n2948) );
  OAI21_X1 U3449 ( .B1(n4894), .B2(n4533), .A(n2948), .ZN(U3524) );
  NAND2_X1 U3450 ( .A1(n2955), .A2(n2949), .ZN(n2951) );
  NAND2_X1 U3451 ( .A1(n3121), .A2(IR_REG_31__SCAN_IN), .ZN(n2950) );
  XNOR2_X1 U3452 ( .A(n2950), .B(IR_REG_10__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U3453 ( .A1(n2951), .A2(IR_REG_31__SCAN_IN), .ZN(n2952) );
  XNOR2_X1 U3454 ( .A(n2952), .B(IR_REG_9__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U3455 ( .A1(n4558), .A2(REG2_REG_9__SCAN_IN), .ZN(n2970) );
  INV_X1 U3456 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2953) );
  INV_X1 U3457 ( .A(n4558), .ZN(n4752) );
  AOI22_X1 U34580 ( .A1(n4558), .A2(REG2_REG_9__SCAN_IN), .B1(n2953), .B2(
        n4752), .ZN(n4566) );
  OR2_X1 U34590 ( .A1(n2955), .A2(n2954), .ZN(n2965) );
  XNOR2_X1 U3460 ( .A(n2965), .B(IR_REG_7__SCAN_IN), .ZN(n4538) );
  INV_X1 U3461 ( .A(n4538), .ZN(n4720) );
  INV_X1 U3462 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2957) );
  MUX2_X1 U3463 ( .A(REG2_REG_2__SCAN_IN), .B(n2957), .S(n4682), .Z(n2958) );
  INV_X1 U3464 ( .A(n2958), .ZN(n4628) );
  NOR2_X1 U3465 ( .A1(n2959), .A2(n4694), .ZN(n2960) );
  NOR2_X1 U3466 ( .A1(n2961), .A2(n4703), .ZN(n2962) );
  INV_X1 U34670 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2963) );
  INV_X1 U3468 ( .A(n2981), .ZN(n4711) );
  AOI22_X1 U34690 ( .A1(n2981), .A2(n2963), .B1(REG2_REG_5__SCAN_IN), .B2(
        n4711), .ZN(n4519) );
  INV_X1 U3470 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4537) );
  INV_X1 U34710 ( .A(IR_REG_7__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U3472 ( .A1(n2965), .A2(n4439), .ZN(n2966) );
  NAND2_X1 U34730 ( .A1(n2966), .A2(IR_REG_31__SCAN_IN), .ZN(n2967) );
  XNOR2_X1 U3474 ( .A(n2967), .B(IR_REG_8__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U34750 ( .A1(n4749), .A2(n2968), .ZN(n2969) );
  NAND2_X1 U3476 ( .A1(n4566), .A2(n4565), .ZN(n4564) );
  OAI211_X1 U34770 ( .C1(n2971), .C2(REG2_REG_10__SCAN_IN), .A(n4607), .B(
        n3755), .ZN(n2973) );
  NOR2_X1 U3478 ( .A1(STATE_REG_SCAN_IN), .A2(n4342), .ZN(n3102) );
  AOI21_X1 U34790 ( .B1(n4646), .B2(ADDR_REG_10__SCAN_IN), .A(n3102), .ZN(
        n2972) );
  OAI211_X1 U3480 ( .C1(n4612), .C2(n2435), .A(n2973), .B(n2972), .ZN(n2994)
         );
  INV_X1 U34810 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2992) );
  INV_X1 U3482 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4708) );
  XNOR2_X1 U34830 ( .A(n2976), .B(n2732), .ZN(n4514) );
  INV_X1 U3484 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4700) );
  NOR2_X1 U34850 ( .A1(n4514), .A2(n4700), .ZN(n4513) );
  INV_X1 U3486 ( .A(n2976), .ZN(n2977) );
  NOR2_X1 U34870 ( .A1(n2977), .A2(n4694), .ZN(n2978) );
  XNOR2_X1 U3488 ( .A(n2979), .B(n4703), .ZN(n4649) );
  NOR2_X1 U34890 ( .A1(n4708), .A2(n4649), .ZN(n4648) );
  NOR2_X1 U3490 ( .A1(n2979), .A2(n4703), .ZN(n2980) );
  AOI22_X1 U34910 ( .A1(n2981), .A2(n2760), .B1(REG1_REG_5__SCAN_IN), .B2(
        n4711), .ZN(n4524) );
  NOR2_X1 U3492 ( .A1(n4523), .A2(n4524), .ZN(n4522) );
  AOI21_X1 U34930 ( .B1(REG1_REG_5__SCAN_IN), .B2(n2981), .A(n4522), .ZN(n2982) );
  NOR2_X1 U3494 ( .A1(n2982), .A2(n4718), .ZN(n2983) );
  XNOR2_X1 U34950 ( .A(n4718), .B(n2982), .ZN(n4532) );
  NAND2_X1 U3496 ( .A1(n4538), .A2(REG1_REG_7__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U34970 ( .A1(n4749), .A2(n2985), .ZN(n2986) );
  NAND2_X1 U3498 ( .A1(n4553), .A2(REG1_REG_8__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U34990 ( .A1(n2986), .A2(n4552), .ZN(n4560) );
  AND2_X1 U3500 ( .A1(n4560), .A2(REG1_REG_9__SCAN_IN), .ZN(n2987) );
  OAI22_X1 U35010 ( .A1(n2987), .A2(n4558), .B1(REG1_REG_9__SCAN_IN), .B2(
        n4560), .ZN(n2988) );
  INV_X1 U3502 ( .A(n3743), .ZN(n2990) );
  NAND2_X1 U35030 ( .A1(n2988), .A2(n2435), .ZN(n2989) );
  AOI211_X1 U3504 ( .C1(n2992), .C2(n2991), .A(n3744), .B(n4647), .ZN(n2993)
         );
  OR2_X1 U35050 ( .A1(n2994), .A2(n2993), .ZN(U3250) );
  INV_X1 U35060 ( .A(n2995), .ZN(n2998) );
  INV_X1 U35070 ( .A(n2996), .ZN(n2997) );
  NAND2_X1 U35080 ( .A1(n2998), .A2(n2997), .ZN(n3000) );
  NAND2_X1 U35090 ( .A1(n4734), .A2(n2736), .ZN(n3002) );
  NAND2_X1 U35100 ( .A1(n3244), .A2(n2263), .ZN(n3001) );
  AOI22_X1 U35110 ( .A1(n4734), .A2(n3437), .B1(n3345), .B2(n3244), .ZN(n3003)
         );
  XNOR2_X1 U35120 ( .A(n3003), .B(n3458), .ZN(n3238) );
  MUX2_X1 U35130 ( .A(n4538), .B(DATAI_7_), .S(n3594), .Z(n4733) );
  AOI22_X1 U35140 ( .A1(n3738), .A2(n2736), .B1(n3437), .B2(n4733), .ZN(n3020)
         );
  NAND2_X1 U35150 ( .A1(n3738), .A2(n2263), .ZN(n3005) );
  NAND2_X1 U35160 ( .A1(n4733), .A2(n3345), .ZN(n3004) );
  NAND2_X1 U35170 ( .A1(n3005), .A2(n3004), .ZN(n3006) );
  XNOR2_X1 U35180 ( .A(n3006), .B(n3458), .ZN(n3019) );
  XOR2_X1 U35190 ( .A(n3020), .B(n3019), .Z(n3021) );
  XNOR2_X1 U35200 ( .A(n3022), .B(n3021), .ZN(n3018) );
  NAND2_X1 U35210 ( .A1(n2261), .A2(REG0_REG_8__SCAN_IN), .ZN(n3014) );
  INV_X1 U35220 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3056) );
  OR2_X1 U35230 ( .A1(n2693), .A2(n3056), .ZN(n3013) );
  INV_X1 U35240 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3008) );
  OR2_X1 U35250 ( .A1(n2259), .A2(n3008), .ZN(n3012) );
  OR2_X1 U35260 ( .A1(n3009), .A2(REG3_REG_8__SCAN_IN), .ZN(n3010) );
  NAND2_X1 U35270 ( .A1(n3031), .A2(n3010), .ZN(n3055) );
  OR2_X1 U35280 ( .A1(n3451), .A2(n3055), .ZN(n3011) );
  AOI22_X1 U35290 ( .A1(n4921), .A2(n4734), .B1(n4899), .B2(n4758), .ZN(n3017)
         );
  NOR2_X1 U35300 ( .A1(STATE_REG_SCAN_IN), .A2(n2916), .ZN(n4542) );
  NOR2_X1 U35310 ( .A1(n4930), .A2(n4742), .ZN(n3015) );
  AOI211_X1 U35320 ( .C1(n4733), .C2(n4924), .A(n4542), .B(n3015), .ZN(n3016)
         );
  OAI211_X1 U35330 ( .C1(n3018), .C2(n3567), .A(n3017), .B(n3016), .ZN(U3210)
         );
  NAND2_X1 U35340 ( .A1(n4758), .A2(n2263), .ZN(n3024) );
  MUX2_X1 U35350 ( .A(n4749), .B(DATAI_8_), .S(n3594), .Z(n3164) );
  NAND2_X1 U35360 ( .A1(n3164), .A2(n3345), .ZN(n3023) );
  NAND2_X1 U35370 ( .A1(n3024), .A2(n3023), .ZN(n3025) );
  XNOR2_X1 U35380 ( .A(n3025), .B(n3440), .ZN(n3027) );
  AOI22_X1 U35390 ( .A1(n4758), .A2(n2736), .B1(n2263), .B2(n3164), .ZN(n3026)
         );
  NOR2_X1 U35400 ( .A1(n3027), .A2(n3026), .ZN(n3065) );
  NAND2_X1 U35410 ( .A1(n3027), .A2(n3026), .ZN(n3064) );
  INV_X1 U35420 ( .A(n3064), .ZN(n3028) );
  NOR2_X1 U35430 ( .A1(n3065), .A2(n3028), .ZN(n3029) );
  XNOR2_X1 U35440 ( .A(n3066), .B(n3029), .ZN(n3041) );
  NAND2_X1 U35450 ( .A1(n2737), .A2(REG1_REG_9__SCAN_IN), .ZN(n3037) );
  OR2_X1 U35460 ( .A1(n2693), .A2(n2953), .ZN(n3036) );
  NAND2_X1 U35470 ( .A1(n3031), .A2(n3030), .ZN(n3032) );
  NAND2_X1 U35480 ( .A1(n3071), .A2(n3032), .ZN(n4769) );
  OR2_X1 U35490 ( .A1(n3451), .A2(n4769), .ZN(n3035) );
  INV_X1 U35500 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3033) );
  OR2_X1 U35510 ( .A1(n2740), .A2(n3033), .ZN(n3034) );
  AOI22_X1 U35520 ( .A1(n4899), .A2(n4225), .B1(n4921), .B2(n3738), .ZN(n3040)
         );
  INV_X1 U35530 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4304) );
  NOR2_X1 U35540 ( .A1(STATE_REG_SCAN_IN), .A2(n4304), .ZN(n4549) );
  NOR2_X1 U35550 ( .A1(n4930), .A2(n3055), .ZN(n3038) );
  AOI211_X1 U35560 ( .C1(n3164), .C2(n4924), .A(n4549), .B(n3038), .ZN(n3039)
         );
  OAI211_X1 U35570 ( .C1(n3041), .C2(n3567), .A(n3040), .B(n3039), .ZN(U3218)
         );
  NAND2_X1 U35580 ( .A1(n4734), .A2(n3244), .ZN(n3043) );
  NAND2_X1 U35590 ( .A1(n3044), .A2(n3043), .ZN(n4725) );
  INV_X1 U35600 ( .A(n4733), .ZN(n3045) );
  OR2_X1 U35610 ( .A1(n3738), .A2(n3045), .ZN(n3629) );
  NAND2_X1 U35620 ( .A1(n3738), .A2(n3045), .ZN(n3632) );
  NAND2_X1 U35630 ( .A1(n3629), .A2(n3632), .ZN(n4726) );
  NAND2_X1 U35640 ( .A1(n4725), .A2(n4726), .ZN(n3047) );
  NAND2_X1 U35650 ( .A1(n3738), .A2(n4733), .ZN(n3046) );
  NAND2_X1 U35660 ( .A1(n3047), .A2(n3046), .ZN(n3163) );
  OR2_X1 U35670 ( .A1(n4758), .A2(n3054), .ZN(n3634) );
  NAND2_X1 U35680 ( .A1(n4758), .A2(n3054), .ZN(n3631) );
  NAND2_X1 U35690 ( .A1(n3634), .A2(n3631), .ZN(n3711) );
  XNOR2_X1 U35700 ( .A(n3163), .B(n3711), .ZN(n3109) );
  NAND2_X1 U35710 ( .A1(n3048), .A2(n3638), .ZN(n3049) );
  NAND2_X1 U35720 ( .A1(n3049), .A2(n3628), .ZN(n4730) );
  INV_X1 U35730 ( .A(n3629), .ZN(n3050) );
  XOR2_X1 U35740 ( .A(n3174), .B(n3711), .Z(n3053) );
  AOI22_X1 U35750 ( .A1(n3738), .A2(n4849), .B1(n3164), .B2(n4787), .ZN(n3052)
         );
  NAND2_X1 U35760 ( .A1(n4225), .A2(n4862), .ZN(n3051) );
  OAI211_X1 U35770 ( .C1(n3053), .C2(n4856), .A(n3052), .B(n3051), .ZN(n3111)
         );
  NAND2_X1 U35780 ( .A1(n3111), .A2(n4674), .ZN(n3060) );
  OAI21_X1 U35790 ( .B1(n4721), .B2(n3054), .A(n4764), .ZN(n3108) );
  INV_X1 U35800 ( .A(n3108), .ZN(n3058) );
  OAI22_X1 U35810 ( .A1(n4674), .A2(n3056), .B1(n3055), .B2(n4741), .ZN(n3057)
         );
  AOI21_X1 U3582 ( .B1(n3058), .B2(n4940), .A(n3057), .ZN(n3059) );
  OAI211_X1 U3583 ( .C1(n3109), .C2(n4140), .A(n3060), .B(n3059), .ZN(U3282)
         );
  NAND2_X1 U3584 ( .A1(n4225), .A2(n3437), .ZN(n3062) );
  MUX2_X1 U3585 ( .A(n4558), .B(DATAI_9_), .S(n3594), .Z(n4765) );
  NAND2_X1 U3586 ( .A1(n4765), .A2(n3345), .ZN(n3061) );
  NAND2_X1 U3587 ( .A1(n3062), .A2(n3061), .ZN(n3063) );
  XNOR2_X1 U3588 ( .A(n3063), .B(n3458), .ZN(n3083) );
  AOI22_X1 U3589 ( .A1(n4225), .A2(n2736), .B1(n3437), .B2(n4765), .ZN(n3084)
         );
  XNOR2_X1 U3590 ( .A(n3083), .B(n3084), .ZN(n3069) );
  NAND2_X1 U3591 ( .A1(n3068), .A2(n3069), .ZN(n3090) );
  OAI21_X1 U3592 ( .B1(n3069), .B2(n3068), .A(n3067), .ZN(n3081) );
  NAND2_X1 U3593 ( .A1(n2260), .A2(REG0_REG_10__SCAN_IN), .ZN(n3077) );
  INV_X1 U3594 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3070) );
  OR2_X1 U3595 ( .A1(n2693), .A2(n3070), .ZN(n3076) );
  NAND2_X1 U3596 ( .A1(n3071), .A2(n4342), .ZN(n3072) );
  AND2_X1 U3597 ( .A1(n3095), .A2(n3072), .ZN(n4776) );
  INV_X1 U3598 ( .A(n4776), .ZN(n3073) );
  OR2_X1 U3599 ( .A1(n3451), .A2(n3073), .ZN(n3075) );
  OR2_X1 U3600 ( .A1(n2259), .A2(n2992), .ZN(n3074) );
  AOI22_X1 U3601 ( .A1(n4921), .A2(n4758), .B1(n4899), .B2(n4788), .ZN(n3079)
         );
  AND2_X1 U3602 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4562) );
  AOI21_X1 U3603 ( .B1(n4924), .B2(n4765), .A(n4562), .ZN(n3078) );
  OAI211_X1 U3604 ( .C1(n4930), .C2(n4769), .A(n3079), .B(n3078), .ZN(n3080)
         );
  AOI21_X1 U3605 ( .B1(n3081), .B2(n4925), .A(n3080), .ZN(n3082) );
  INV_X1 U3606 ( .A(n3082), .ZN(U3228) );
  INV_X1 U3607 ( .A(n3083), .ZN(n3085) );
  NAND2_X1 U3608 ( .A1(n3085), .A2(n3084), .ZN(n3092) );
  NAND2_X1 U3609 ( .A1(n4788), .A2(n2263), .ZN(n3087) );
  MUX2_X1 U3610 ( .A(n4467), .B(DATAI_10_), .S(n3594), .Z(n4224) );
  NAND2_X1 U3611 ( .A1(n4224), .A2(n3345), .ZN(n3086) );
  NAND2_X1 U3612 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  XNOR2_X1 U3613 ( .A(n3088), .B(n3458), .ZN(n3116) );
  AOI22_X1 U3614 ( .A1(n4788), .A2(n2736), .B1(n3437), .B2(n4224), .ZN(n3117)
         );
  XNOR2_X1 U3615 ( .A(n3116), .B(n3117), .ZN(n3091) );
  NAND2_X1 U3616 ( .A1(n3120), .A2(n4925), .ZN(n3107) );
  AOI21_X1 U3617 ( .B1(n3067), .B2(n3092), .A(n3091), .ZN(n3106) );
  NAND2_X1 U3618 ( .A1(n2260), .A2(REG0_REG_11__SCAN_IN), .ZN(n3101) );
  INV_X1 U3619 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3093) );
  OR2_X1 U3620 ( .A1(n2693), .A2(n3093), .ZN(n3100) );
  AND2_X1 U3621 ( .A1(n3095), .A2(n3094), .ZN(n3096) );
  OR2_X1 U3622 ( .A1(n3096), .A2(n3131), .ZN(n4802) );
  OR2_X1 U3623 ( .A1(n3451), .A2(n4802), .ZN(n3099) );
  INV_X1 U3624 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3097) );
  OR2_X1 U3625 ( .A1(n2259), .A2(n3097), .ZN(n3098) );
  AOI22_X1 U3626 ( .A1(n4921), .A2(n4225), .B1(n4899), .B2(n3737), .ZN(n3105)
         );
  INV_X1 U3627 ( .A(n4224), .ZN(n3177) );
  NOR2_X1 U3628 ( .A1(n4834), .A2(n3177), .ZN(n3103) );
  AOI211_X1 U3629 ( .C1(n3565), .C2(n4776), .A(n3103), .B(n3102), .ZN(n3104)
         );
  OAI211_X1 U3630 ( .C1(n3107), .C2(n3106), .A(n3105), .B(n3104), .ZN(U3214)
         );
  INV_X1 U3631 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3113) );
  OAI22_X1 U3632 ( .A1(n3109), .A2(n4888), .B1(n4887), .B2(n3108), .ZN(n3110)
         );
  OR2_X1 U3633 ( .A1(n3111), .A2(n3110), .ZN(n3114) );
  NAND2_X1 U3634 ( .A1(n3114), .A2(n4897), .ZN(n3112) );
  OAI21_X1 U3635 ( .B1(n4897), .B2(n3113), .A(n3112), .ZN(U3483) );
  NAND2_X1 U3636 ( .A1(n3114), .A2(n4894), .ZN(n3115) );
  OAI21_X1 U3637 ( .B1(n4894), .B2(n3008), .A(n3115), .ZN(U3526) );
  INV_X1 U3638 ( .A(n3117), .ZN(n3118) );
  OAI21_X1 U3639 ( .B1(n3121), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3123) );
  INV_X1 U3640 ( .A(IR_REG_11__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U3641 ( .A1(n3123), .A2(n3122), .ZN(n3144) );
  OR2_X1 U3642 ( .A1(n3123), .A2(n3122), .ZN(n3124) );
  MUX2_X1 U3643 ( .A(n4570), .B(DATAI_11_), .S(n3594), .Z(n4798) );
  AOI22_X1 U3644 ( .A1(n3737), .A2(n3437), .B1(n3345), .B2(n4798), .ZN(n3125)
         );
  XOR2_X1 U3645 ( .A(n3458), .B(n3125), .Z(n3127) );
  INV_X1 U3646 ( .A(n3737), .ZN(n4227) );
  OAI22_X1 U3647 ( .A1(n4227), .A2(n3457), .B1(n3401), .B2(n3195), .ZN(n3126)
         );
  NOR2_X1 U3648 ( .A1(n3127), .A2(n3126), .ZN(n3141) );
  NOR2_X1 U3649 ( .A1(n3141), .A2(n2302), .ZN(n3128) );
  XNOR2_X1 U3650 ( .A(n3143), .B(n3128), .ZN(n3140) );
  NAND2_X1 U3651 ( .A1(n2260), .A2(REG0_REG_12__SCAN_IN), .ZN(n3136) );
  INV_X1 U3652 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3129) );
  OR2_X1 U3653 ( .A1(n2693), .A2(n3129), .ZN(n3135) );
  INV_X1 U3654 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3130) );
  OR2_X1 U3655 ( .A1(n2259), .A2(n3130), .ZN(n3134) );
  NOR2_X1 U3656 ( .A1(n3131), .A2(REG3_REG_12__SCAN_IN), .ZN(n3132) );
  OR2_X1 U3657 ( .A1(n3151), .A2(n3132), .ZN(n3158) );
  OR2_X1 U3658 ( .A1(n3451), .A2(n3158), .ZN(n3133) );
  AOI22_X1 U3659 ( .A1(n4921), .A2(n4788), .B1(n4899), .B2(n4789), .ZN(n3139)
         );
  AND2_X1 U3660 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4573) );
  NOR2_X1 U3661 ( .A1(n4930), .A2(n4802), .ZN(n3137) );
  AOI211_X1 U3662 ( .C1(n4798), .C2(n4924), .A(n4573), .B(n3137), .ZN(n3138)
         );
  OAI211_X1 U3663 ( .C1(n3140), .C2(n3567), .A(n3139), .B(n3138), .ZN(U3233)
         );
  NAND2_X1 U3664 ( .A1(n3144), .A2(IR_REG_31__SCAN_IN), .ZN(n3145) );
  XNOR2_X1 U3665 ( .A(n3145), .B(IR_REG_12__SCAN_IN), .ZN(n4583) );
  MUX2_X1 U3666 ( .A(n4583), .B(DATAI_12_), .S(n3594), .Z(n3169) );
  AOI22_X1 U3667 ( .A1(n4789), .A2(n3437), .B1(n3345), .B2(n3169), .ZN(n3146)
         );
  XOR2_X1 U3668 ( .A(n3458), .B(n3146), .Z(n3204) );
  INV_X1 U3669 ( .A(n4789), .ZN(n3147) );
  OAI22_X1 U3670 ( .A1(n3147), .A2(n3457), .B1(n3401), .B2(n4212), .ZN(n3205)
         );
  INV_X1 U3671 ( .A(n3205), .ZN(n3148) );
  XNOR2_X1 U3672 ( .A(n3204), .B(n3148), .ZN(n3149) );
  XNOR2_X1 U3673 ( .A(n3206), .B(n3149), .ZN(n3162) );
  NAND2_X1 U3674 ( .A1(n2261), .A2(REG0_REG_13__SCAN_IN), .ZN(n3157) );
  INV_X1 U3675 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3150) );
  OR2_X1 U3676 ( .A1(n2693), .A2(n3150), .ZN(n3156) );
  OR2_X1 U3677 ( .A1(n3151), .A2(REG3_REG_13__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U3678 ( .A1(n3152), .A2(n3182), .ZN(n3231) );
  OR2_X1 U3679 ( .A1(n3451), .A2(n3231), .ZN(n3155) );
  INV_X1 U3680 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3153) );
  OR2_X1 U3681 ( .A1(n2259), .A2(n3153), .ZN(n3154) );
  AOI22_X1 U3682 ( .A1(n4921), .A2(n3737), .B1(n4899), .B2(n4217), .ZN(n3161)
         );
  INV_X1 U3683 ( .A(n3158), .ZN(n4812) );
  INV_X1 U3684 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4410) );
  NOR2_X1 U3685 ( .A1(STATE_REG_SCAN_IN), .A2(n4410), .ZN(n4580) );
  NOR2_X1 U3686 ( .A1(n4834), .A2(n4212), .ZN(n3159) );
  AOI211_X1 U3687 ( .C1(n3565), .C2(n4812), .A(n4580), .B(n3159), .ZN(n3160)
         );
  OAI211_X1 U3688 ( .C1(n3162), .C2(n3567), .A(n3161), .B(n3160), .ZN(U3221)
         );
  OR2_X1 U3689 ( .A1(n4758), .A2(n3164), .ZN(n4754) );
  NAND2_X1 U3690 ( .A1(n4758), .A2(n3164), .ZN(n4753) );
  AND2_X1 U3691 ( .A1(n4788), .A2(n4224), .ZN(n3166) );
  OR2_X1 U3692 ( .A1(n4788), .A2(n4224), .ZN(n3165) );
  NAND2_X1 U3693 ( .A1(n3737), .A2(n3195), .ZN(n3642) );
  NAND2_X1 U3694 ( .A1(n3648), .A2(n3642), .ZN(n4785) );
  NOR2_X1 U3695 ( .A1(n3737), .A2(n4798), .ZN(n3167) );
  AOI21_X1 U3696 ( .B1(n4784), .B2(n4785), .A(n3167), .ZN(n4218) );
  OR2_X1 U3697 ( .A1(n4789), .A2(n3169), .ZN(n3168) );
  NAND2_X1 U3698 ( .A1(n4789), .A2(n3169), .ZN(n3170) );
  NAND2_X1 U3699 ( .A1(n3171), .A2(IR_REG_31__SCAN_IN), .ZN(n3173) );
  XNOR2_X1 U3700 ( .A(n3173), .B(n3172), .ZN(n4820) );
  INV_X1 U3701 ( .A(n4820), .ZN(n3759) );
  MUX2_X1 U3702 ( .A(n3759), .B(DATAI_13_), .S(n3594), .Z(n3233) );
  OR2_X1 U3703 ( .A1(n4217), .A2(n3233), .ZN(n4134) );
  NAND2_X1 U3704 ( .A1(n4217), .A2(n3233), .ZN(n4136) );
  NAND2_X1 U3705 ( .A1(n4134), .A2(n4136), .ZN(n3180) );
  XNOR2_X1 U3706 ( .A(n3814), .B(n3180), .ZN(n4824) );
  NAND2_X1 U3707 ( .A1(n4824), .A2(n4794), .ZN(n3193) );
  INV_X1 U3708 ( .A(n4765), .ZN(n3175) );
  AND2_X1 U3709 ( .A1(n4225), .A2(n3175), .ZN(n3633) );
  NAND2_X1 U3710 ( .A1(n3176), .A2(n3696), .ZN(n4222) );
  NAND2_X1 U3711 ( .A1(n4788), .A2(n3177), .ZN(n3709) );
  NAND2_X1 U3712 ( .A1(n4222), .A2(n3709), .ZN(n3178) );
  NAND2_X1 U3713 ( .A1(n3178), .A2(n3710), .ZN(n4786) );
  NAND2_X1 U3714 ( .A1(n4786), .A2(n3642), .ZN(n3179) );
  NAND2_X1 U3715 ( .A1(n3179), .A2(n3648), .ZN(n3575) );
  NOR2_X1 U3716 ( .A1(n4789), .A2(n4212), .ZN(n3708) );
  NAND2_X1 U3717 ( .A1(n4789), .A2(n4212), .ZN(n3706) );
  OAI21_X1 U3718 ( .B1(n3575), .B2(n3708), .A(n3706), .ZN(n3181) );
  INV_X1 U3719 ( .A(n3180), .ZN(n3689) );
  XNOR2_X1 U3720 ( .A(n3181), .B(n3689), .ZN(n3191) );
  INV_X1 U3721 ( .A(n3233), .ZN(n3576) );
  NAND2_X1 U3722 ( .A1(n2261), .A2(REG0_REG_14__SCAN_IN), .ZN(n3187) );
  INV_X1 U3723 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4133) );
  OR2_X1 U3724 ( .A1(n2693), .A2(n4133), .ZN(n3186) );
  INV_X1 U3725 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3751) );
  OR2_X1 U3726 ( .A1(n2259), .A2(n3751), .ZN(n3185) );
  AOI21_X1 U3727 ( .B1(n3182), .B2(n4398), .A(n3217), .ZN(n3183) );
  INV_X1 U3728 ( .A(n3183), .ZN(n4132) );
  OR2_X1 U3729 ( .A1(n3451), .A2(n4132), .ZN(n3184) );
  NAND2_X1 U3730 ( .A1(n4850), .A2(n4862), .ZN(n3189) );
  NAND2_X1 U3731 ( .A1(n4789), .A2(n4849), .ZN(n3188) );
  OAI211_X1 U3732 ( .C1(n4853), .C2(n3576), .A(n3189), .B(n3188), .ZN(n3190)
         );
  AOI21_X1 U3733 ( .B1(n3191), .B2(n4731), .A(n3190), .ZN(n3192) );
  INV_X1 U3734 ( .A(n3194), .ZN(n4763) );
  NAND2_X1 U3735 ( .A1(n4211), .A2(n3233), .ZN(n3196) );
  NAND2_X1 U3736 ( .A1(n4130), .A2(n3196), .ZN(n4821) );
  NOR2_X1 U3737 ( .A1(n4821), .A2(n4934), .ZN(n3198) );
  OAI22_X1 U3738 ( .A1(n4674), .A2(n3150), .B1(n3231), .B2(n4741), .ZN(n3197)
         );
  AOI211_X1 U3739 ( .C1(n4824), .C2(n4805), .A(n3198), .B(n3197), .ZN(n3199)
         );
  OAI21_X1 U3740 ( .B1(n4826), .B2(n4939), .A(n3199), .ZN(U3277) );
  NAND3_X1 U3741 ( .A1(n3200), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3202) );
  INV_X1 U3742 ( .A(DATAI_31_), .ZN(n3201) );
  OAI22_X1 U3743 ( .A1(n3203), .A2(n3202), .B1(STATE_REG_SCAN_IN), .B2(n3201), 
        .ZN(U3321) );
  NAND2_X1 U3744 ( .A1(n3206), .A2(n3205), .ZN(n3208) );
  OAI21_X1 U3745 ( .B1(n3206), .B2(n3205), .A(n3204), .ZN(n3207) );
  NAND2_X1 U3746 ( .A1(n3208), .A2(n3207), .ZN(n3226) );
  NAND2_X1 U3747 ( .A1(n4217), .A2(n2263), .ZN(n3210) );
  NAND2_X1 U3748 ( .A1(n3233), .A2(n3345), .ZN(n3209) );
  NAND2_X1 U3749 ( .A1(n3210), .A2(n3209), .ZN(n3211) );
  XNOR2_X1 U3750 ( .A(n3211), .B(n3440), .ZN(n3213) );
  AOI22_X1 U3751 ( .A1(n4217), .A2(n2736), .B1(n2263), .B2(n3233), .ZN(n3212)
         );
  NOR2_X1 U3752 ( .A1(n3213), .A2(n3212), .ZN(n3228) );
  NAND2_X1 U3753 ( .A1(n3213), .A2(n3212), .ZN(n3227) );
  XNOR2_X1 U3754 ( .A(n3214), .B(IR_REG_14__SCAN_IN), .ZN(n4466) );
  MUX2_X1 U3755 ( .A(n4466), .B(DATAI_14_), .S(n3594), .Z(n4129) );
  AOI22_X1 U3756 ( .A1(n4850), .A2(n2263), .B1(n3345), .B2(n4129), .ZN(n3215)
         );
  XNOR2_X1 U3757 ( .A(n3215), .B(n3458), .ZN(n3261) );
  AOI22_X1 U3758 ( .A1(n4850), .A2(n2736), .B1(n2263), .B2(n4129), .ZN(n3262)
         );
  XNOR2_X1 U3759 ( .A(n3261), .B(n3262), .ZN(n3216) );
  XNOR2_X1 U3760 ( .A(n3263), .B(n3216), .ZN(n3225) );
  NAND2_X1 U3761 ( .A1(n2260), .A2(REG0_REG_15__SCAN_IN), .ZN(n3221) );
  INV_X1 U3762 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3767) );
  OR2_X1 U3763 ( .A1(n2693), .A2(n3767), .ZN(n3220) );
  OAI21_X1 U3764 ( .B1(n3217), .B2(REG3_REG_15__SCAN_IN), .A(n3264), .ZN(n4866) );
  OR2_X1 U3765 ( .A1(n3451), .A2(n4866), .ZN(n3219) );
  OR2_X1 U3766 ( .A1(n2259), .A2(n3782), .ZN(n3218) );
  AOI22_X1 U3767 ( .A1(n4899), .A2(n4106), .B1(n4921), .B2(n4217), .ZN(n3224)
         );
  NOR2_X1 U3768 ( .A1(STATE_REG_SCAN_IN), .A2(n4398), .ZN(n3752) );
  NOR2_X1 U3769 ( .A1(n4930), .A2(n4132), .ZN(n3222) );
  AOI211_X1 U3770 ( .C1(n4129), .C2(n4924), .A(n3752), .B(n3222), .ZN(n3223)
         );
  OAI211_X1 U3771 ( .C1(n3225), .C2(n3567), .A(n3224), .B(n3223), .ZN(U3212)
         );
  NOR2_X1 U3772 ( .A1(n3228), .A2(n2470), .ZN(n3229) );
  XNOR2_X1 U3773 ( .A(n3230), .B(n3229), .ZN(n3236) );
  AOI22_X1 U3774 ( .A1(n4899), .A2(n4850), .B1(n4921), .B2(n4789), .ZN(n3235)
         );
  INV_X1 U3775 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4317) );
  NOR2_X1 U3776 ( .A1(STATE_REG_SCAN_IN), .A2(n4317), .ZN(n4598) );
  NOR2_X1 U3777 ( .A1(n4930), .A2(n3231), .ZN(n3232) );
  AOI211_X1 U3778 ( .C1(n3233), .C2(n4924), .A(n4598), .B(n3232), .ZN(n3234)
         );
  OAI211_X1 U3779 ( .C1(n3236), .C2(n3567), .A(n3235), .B(n3234), .ZN(U3231)
         );
  XNOR2_X1 U3780 ( .A(n3238), .B(n3237), .ZN(n3239) );
  XNOR2_X1 U3781 ( .A(n3240), .B(n3239), .ZN(n3247) );
  AOI22_X1 U3782 ( .A1(n4899), .A2(n3738), .B1(n4921), .B2(n3739), .ZN(n3246)
         );
  INV_X1 U3783 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3241) );
  NOR2_X1 U3784 ( .A1(STATE_REG_SCAN_IN), .A2(n3241), .ZN(n4530) );
  NOR2_X1 U3785 ( .A1(n4930), .A2(n3242), .ZN(n3243) );
  AOI211_X1 U3786 ( .C1(n3244), .C2(n4924), .A(n4530), .B(n3243), .ZN(n3245)
         );
  OAI211_X1 U3787 ( .C1(n3247), .C2(n3567), .A(n3246), .B(n3245), .ZN(U3236)
         );
  INV_X1 U3788 ( .A(n3249), .ZN(n3250) );
  AOI21_X1 U3789 ( .B1(n3248), .B2(n3251), .A(n3250), .ZN(n3255) );
  AOI22_X1 U3790 ( .A1(n3258), .A2(REG3_REG_2__SCAN_IN), .B1(n4924), .B2(n3252), .ZN(n3254) );
  AOI22_X1 U3791 ( .A1(n4899), .A2(n2757), .B1(n4921), .B2(n2657), .ZN(n3253)
         );
  OAI211_X1 U3792 ( .C1(n3255), .C2(n3567), .A(n3254), .B(n3253), .ZN(U3234)
         );
  XOR2_X1 U3793 ( .A(n3257), .B(n3256), .Z(n4636) );
  NAND2_X1 U3794 ( .A1(n4636), .A2(n4925), .ZN(n3260) );
  AOI22_X1 U3795 ( .A1(n3258), .A2(REG3_REG_0__SCAN_IN), .B1(n4924), .B2(n4664), .ZN(n3259) );
  OAI211_X1 U3796 ( .C1(n2784), .C2(n4913), .A(n3260), .B(n3259), .ZN(U3229)
         );
  NAND2_X1 U3797 ( .A1(n2261), .A2(REG0_REG_16__SCAN_IN), .ZN(n3271) );
  INV_X1 U3798 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4115) );
  OR2_X1 U3799 ( .A1(n2693), .A2(n4115), .ZN(n3270) );
  NAND2_X1 U3800 ( .A1(n3264), .A2(n4413), .ZN(n3266) );
  INV_X1 U3801 ( .A(n3296), .ZN(n3265) );
  NAND2_X1 U3802 ( .A1(n3266), .A2(n3265), .ZN(n4114) );
  OR2_X1 U3803 ( .A1(n3451), .A2(n4114), .ZN(n3269) );
  INV_X1 U3804 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3267) );
  OR2_X1 U3805 ( .A1(n2259), .A2(n3267), .ZN(n3268) );
  OR2_X1 U3806 ( .A1(n3278), .A2(IR_REG_15__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U3807 ( .A1(n3280), .A2(IR_REG_31__SCAN_IN), .ZN(n3272) );
  MUX2_X1 U3808 ( .A(IR_REG_31__SCAN_IN), .B(n3272), .S(IR_REG_16__SCAN_IN), 
        .Z(n3275) );
  OR2_X1 U3809 ( .A1(n3278), .A2(n3273), .ZN(n3274) );
  NAND2_X1 U3810 ( .A1(n3275), .A2(n3274), .ZN(n4877) );
  INV_X1 U3811 ( .A(n4877), .ZN(n3276) );
  MUX2_X1 U3812 ( .A(n3276), .B(DATAI_16_), .S(n3594), .Z(n4113) );
  AOI22_X1 U3813 ( .A1(n4861), .A2(n2262), .B1(n3345), .B2(n4113), .ZN(n3277)
         );
  XOR2_X1 U3814 ( .A(n3458), .B(n3277), .Z(n3289) );
  INV_X1 U3815 ( .A(n4861), .ZN(n4831) );
  OAI22_X1 U3816 ( .A1(n4831), .A2(n3457), .B1(n3401), .B2(n3877), .ZN(n3290)
         );
  NAND2_X1 U3817 ( .A1(n3289), .A2(n3290), .ZN(n3515) );
  NAND2_X1 U3818 ( .A1(n4106), .A2(n2263), .ZN(n3282) );
  NAND2_X1 U3819 ( .A1(n3278), .A2(IR_REG_15__SCAN_IN), .ZN(n3279) );
  MUX2_X1 U3820 ( .A(n4465), .B(DATAI_15_), .S(n3594), .Z(n3815) );
  NAND2_X1 U3821 ( .A1(n3815), .A2(n3345), .ZN(n3281) );
  NAND2_X1 U3822 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  XNOR2_X1 U3823 ( .A(n3283), .B(n3440), .ZN(n4838) );
  NAND2_X1 U3824 ( .A1(n4106), .A2(n2736), .ZN(n3285) );
  NAND2_X1 U3825 ( .A1(n3815), .A2(n2263), .ZN(n3284) );
  NAND2_X1 U3826 ( .A1(n4838), .A2(n3511), .ZN(n3288) );
  INV_X1 U3827 ( .A(n3289), .ZN(n3292) );
  INV_X1 U3828 ( .A(n3290), .ZN(n3291) );
  NAND2_X1 U3829 ( .A1(n3292), .A2(n3291), .ZN(n3514) );
  NAND2_X1 U3830 ( .A1(n3295), .A2(n3294), .ZN(n3522) );
  NAND2_X1 U3831 ( .A1(n2737), .A2(REG1_REG_17__SCAN_IN), .ZN(n3301) );
  INV_X1 U3832 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4098) );
  OR2_X1 U3833 ( .A1(n2693), .A2(n4098), .ZN(n3300) );
  XNOR2_X1 U3834 ( .A(REG3_REG_17__SCAN_IN), .B(n3296), .ZN(n4097) );
  OR2_X1 U3835 ( .A1(n3451), .A2(n4097), .ZN(n3299) );
  INV_X1 U3836 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3297) );
  OR2_X1 U3837 ( .A1(n2740), .A2(n3297), .ZN(n3298) );
  NAND2_X1 U3838 ( .A1(n4103), .A2(n3437), .ZN(n3303) );
  MUX2_X1 U3839 ( .A(n3805), .B(DATAI_17_), .S(n3594), .Z(n4094) );
  NAND2_X1 U3840 ( .A1(n4094), .A2(n3345), .ZN(n3302) );
  NAND2_X1 U3841 ( .A1(n3303), .A2(n3302), .ZN(n3304) );
  XNOR2_X1 U3842 ( .A(n3304), .B(n3440), .ZN(n3306) );
  AOI22_X1 U3843 ( .A1(n4103), .A2(n2736), .B1(n3437), .B2(n4094), .ZN(n3305)
         );
  OR2_X1 U3844 ( .A1(n3306), .A2(n3305), .ZN(n3524) );
  AND2_X1 U3845 ( .A1(n3306), .A2(n3305), .ZN(n3523) );
  NAND2_X1 U3846 ( .A1(n3464), .A2(REG2_REG_18__SCAN_IN), .ZN(n3314) );
  INV_X1 U3847 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4205) );
  OR2_X1 U3848 ( .A1(n2259), .A2(n4205), .ZN(n3313) );
  INV_X1 U3849 ( .A(n3307), .ZN(n3309) );
  INV_X1 U3850 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U3851 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  NAND2_X1 U3852 ( .A1(n3324), .A2(n3310), .ZN(n4076) );
  OR2_X1 U3853 ( .A1(n3451), .A2(n4076), .ZN(n3312) );
  INV_X1 U3854 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4457) );
  OR2_X1 U3855 ( .A1(n2740), .A2(n4457), .ZN(n3311) );
  NAND2_X1 U3856 ( .A1(n4091), .A2(n2263), .ZN(n3316) );
  MUX2_X1 U3857 ( .A(n4621), .B(DATAI_18_), .S(n3594), .Z(n4072) );
  NAND2_X1 U3858 ( .A1(n4072), .A2(n3345), .ZN(n3315) );
  NAND2_X1 U3859 ( .A1(n3316), .A2(n3315), .ZN(n3317) );
  XNOR2_X1 U3860 ( .A(n3317), .B(n3440), .ZN(n3550) );
  NAND2_X1 U3861 ( .A1(n4091), .A2(n2736), .ZN(n3319) );
  NAND2_X1 U3862 ( .A1(n4072), .A2(n2263), .ZN(n3318) );
  NAND2_X1 U3863 ( .A1(n3550), .A2(n3320), .ZN(n3322) );
  INV_X1 U3864 ( .A(n3550), .ZN(n3321) );
  NAND2_X1 U3865 ( .A1(n2261), .A2(REG0_REG_19__SCAN_IN), .ZN(n3330) );
  INV_X1 U3866 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4061) );
  OR2_X1 U3867 ( .A1(n2693), .A2(n4061), .ZN(n3329) );
  INV_X1 U3868 ( .A(n3323), .ZN(n3338) );
  NAND2_X1 U3869 ( .A1(n3324), .A2(n4405), .ZN(n3325) );
  NAND2_X1 U3870 ( .A1(n3338), .A2(n3325), .ZN(n4060) );
  OR2_X1 U3871 ( .A1(n3451), .A2(n4060), .ZN(n3328) );
  INV_X1 U3872 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3326) );
  OR2_X1 U3873 ( .A1(n2259), .A2(n3326), .ZN(n3327) );
  MUX2_X1 U3874 ( .A(n3809), .B(DATAI_19_), .S(n3594), .Z(n4057) );
  AOI22_X1 U3875 ( .A1(n4904), .A2(n3437), .B1(n3345), .B2(n4057), .ZN(n3331)
         );
  XOR2_X1 U3876 ( .A(n3458), .B(n3331), .Z(n3333) );
  INV_X1 U3877 ( .A(n4904), .ZN(n4030) );
  INV_X1 U3878 ( .A(n4057), .ZN(n3682) );
  OAI22_X1 U3879 ( .A1(n4030), .A2(n3457), .B1(n3401), .B2(n3682), .ZN(n3332)
         );
  NOR2_X1 U3880 ( .A1(n3333), .A2(n3332), .ZN(n3334) );
  AOI21_X1 U3881 ( .B1(n3333), .B2(n3332), .A(n3334), .ZN(n3494) );
  INV_X1 U3882 ( .A(n3334), .ZN(n3335) );
  NAND2_X1 U3883 ( .A1(n3464), .A2(REG2_REG_20__SCAN_IN), .ZN(n3344) );
  INV_X1 U3884 ( .A(REG1_REG_20__SCAN_IN), .ZN(n3336) );
  OR2_X1 U3885 ( .A1(n2259), .A2(n3336), .ZN(n3343) );
  INV_X1 U3886 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U3887 ( .A1(n3338), .A2(n3337), .ZN(n3339) );
  NAND2_X1 U3888 ( .A1(n3352), .A2(n3339), .ZN(n4910) );
  OR2_X1 U3889 ( .A1(n3451), .A2(n4910), .ZN(n3342) );
  INV_X1 U3890 ( .A(REG0_REG_20__SCAN_IN), .ZN(n3340) );
  OR2_X1 U3891 ( .A1(n2740), .A2(n3340), .ZN(n3341) );
  NAND2_X1 U3892 ( .A1(n4922), .A2(n2263), .ZN(n3347) );
  NAND2_X1 U3893 ( .A1(n3594), .A2(DATAI_20_), .ZN(n4037) );
  OR2_X1 U3894 ( .A1(n4037), .A2(n3460), .ZN(n3346) );
  NAND2_X1 U3895 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  XNOR2_X1 U3896 ( .A(n3348), .B(n3458), .ZN(n3363) );
  NAND2_X1 U3897 ( .A1(n4922), .A2(n2736), .ZN(n3350) );
  OR2_X1 U3898 ( .A1(n4037), .A2(n3401), .ZN(n3349) );
  NAND2_X1 U3899 ( .A1(n3350), .A2(n3349), .ZN(n3364) );
  NAND2_X1 U3900 ( .A1(n3363), .A2(n3364), .ZN(n4915) );
  NAND2_X1 U3901 ( .A1(n3464), .A2(REG2_REG_21__SCAN_IN), .ZN(n3358) );
  INV_X1 U3902 ( .A(REG1_REG_21__SCAN_IN), .ZN(n3351) );
  OR2_X1 U3903 ( .A1(n2259), .A2(n3351), .ZN(n3357) );
  NAND2_X1 U3904 ( .A1(n3352), .A2(n4911), .ZN(n3353) );
  NAND2_X1 U3905 ( .A1(n3372), .A2(n3353), .ZN(n4929) );
  OR2_X1 U3906 ( .A1(n3451), .A2(n4929), .ZN(n3356) );
  INV_X1 U3907 ( .A(REG0_REG_21__SCAN_IN), .ZN(n3354) );
  OR2_X1 U3908 ( .A1(n2740), .A2(n3354), .ZN(n3355) );
  NAND2_X1 U3909 ( .A1(n3594), .A2(DATAI_21_), .ZN(n4020) );
  NOR2_X1 U3910 ( .A1(n4020), .A2(n3401), .ZN(n3359) );
  AOI21_X1 U3911 ( .B1(n4898), .B2(n2736), .A(n3359), .ZN(n4917) );
  NAND2_X1 U3912 ( .A1(n4898), .A2(n2263), .ZN(n3361) );
  OR2_X1 U3913 ( .A1(n4020), .A2(n3460), .ZN(n3360) );
  NAND2_X1 U3914 ( .A1(n3361), .A2(n3360), .ZN(n3362) );
  XNOR2_X1 U3915 ( .A(n3362), .B(n3440), .ZN(n4918) );
  INV_X1 U3916 ( .A(n3363), .ZN(n3366) );
  INV_X1 U3917 ( .A(n3364), .ZN(n3365) );
  AOI21_X1 U3918 ( .B1(n4917), .B2(n4918), .A(n4901), .ZN(n3368) );
  NAND2_X1 U3919 ( .A1(n3594), .A2(DATAI_22_), .ZN(n3831) );
  OAI22_X1 U3920 ( .A1(n4912), .A2(n3457), .B1(n3401), .B2(n3831), .ZN(n3384)
         );
  OAI22_X1 U3921 ( .A1(n4912), .A2(n3401), .B1(n3460), .B2(n3831), .ZN(n3369)
         );
  XNOR2_X1 U3922 ( .A(n3369), .B(n3458), .ZN(n3383) );
  XOR2_X1 U3923 ( .A(n3384), .B(n3383), .Z(n3543) );
  NAND2_X1 U3924 ( .A1(n3541), .A2(n3543), .ZN(n3484) );
  NAND2_X1 U3925 ( .A1(n2260), .A2(REG0_REG_23__SCAN_IN), .ZN(n3378) );
  INV_X1 U3926 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3982) );
  OR2_X1 U3927 ( .A1(n2693), .A2(n3982), .ZN(n3377) );
  INV_X1 U3928 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4343) );
  OAI21_X1 U3929 ( .B1(n3372), .B2(n3370), .A(n4343), .ZN(n3373) );
  NAND2_X1 U3930 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n3371) );
  NAND2_X1 U3931 ( .A1(n3373), .A2(n3392), .ZN(n3981) );
  OR2_X1 U3932 ( .A1(n3451), .A2(n3981), .ZN(n3376) );
  INV_X1 U3933 ( .A(REG1_REG_23__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U3934 ( .A1(n3960), .A2(n2263), .ZN(n3380) );
  NAND2_X1 U3935 ( .A1(n3594), .A2(DATAI_23_), .ZN(n3991) );
  OR2_X1 U3936 ( .A1(n3991), .A2(n3460), .ZN(n3379) );
  NAND2_X1 U3937 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  XNOR2_X1 U3938 ( .A(n3381), .B(n3458), .ZN(n3388) );
  NOR2_X1 U3939 ( .A1(n3991), .A2(n3401), .ZN(n3382) );
  AOI21_X1 U3940 ( .B1(n3960), .B2(n2736), .A(n3382), .ZN(n3389) );
  XNOR2_X1 U3941 ( .A(n3388), .B(n3389), .ZN(n3485) );
  INV_X1 U3942 ( .A(n3383), .ZN(n3386) );
  INV_X1 U3943 ( .A(n3384), .ZN(n3385) );
  NAND2_X1 U3944 ( .A1(n3386), .A2(n3385), .ZN(n3486) );
  INV_X1 U3945 ( .A(n3388), .ZN(n3390) );
  OR2_X1 U3946 ( .A1(n3390), .A2(n3389), .ZN(n3402) );
  NAND2_X1 U3947 ( .A1(n2261), .A2(REG0_REG_24__SCAN_IN), .ZN(n3398) );
  INV_X1 U3948 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3966) );
  OR2_X1 U3949 ( .A1(n2693), .A2(n3966), .ZN(n3397) );
  INV_X1 U3950 ( .A(n3392), .ZN(n3391) );
  INV_X1 U3951 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U3952 ( .A1(n3392), .A2(n4421), .ZN(n3393) );
  NAND2_X1 U3953 ( .A1(n3405), .A2(n3393), .ZN(n3965) );
  OR2_X1 U3954 ( .A1(n3451), .A2(n3965), .ZN(n3396) );
  INV_X1 U3955 ( .A(REG1_REG_24__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U3956 ( .A1(n3594), .A2(DATAI_24_), .ZN(n3968) );
  NOR2_X1 U3957 ( .A1(n3968), .A2(n3460), .ZN(n3399) );
  AOI21_X1 U3958 ( .B1(n3993), .B2(n3437), .A(n3399), .ZN(n3400) );
  XNOR2_X1 U3959 ( .A(n3400), .B(n3458), .ZN(n3403) );
  OAI22_X1 U3960 ( .A1(n3833), .A2(n3457), .B1(n3401), .B2(n3968), .ZN(n3534)
         );
  NAND3_X1 U3961 ( .A1(n3483), .A2(n3403), .A3(n3402), .ZN(n3531) );
  OAI21_X1 U3962 ( .B1(n3533), .B2(n3534), .A(n3531), .ZN(n3504) );
  INV_X1 U3963 ( .A(n3504), .ZN(n3413) );
  NAND2_X1 U3964 ( .A1(n3464), .A2(REG2_REG_25__SCAN_IN), .ZN(n3411) );
  INV_X1 U3965 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4240) );
  OR2_X1 U3966 ( .A1(n2740), .A2(n4240), .ZN(n3410) );
  INV_X1 U3967 ( .A(n3405), .ZN(n3404) );
  NAND2_X1 U3968 ( .A1(n3404), .A2(REG3_REG_25__SCAN_IN), .ZN(n3416) );
  INV_X1 U3969 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U3970 ( .A1(n3405), .A2(n4412), .ZN(n3406) );
  NAND2_X1 U3971 ( .A1(n3416), .A2(n3406), .ZN(n3947) );
  INV_X1 U3972 ( .A(REG1_REG_25__SCAN_IN), .ZN(n3407) );
  OR2_X1 U3973 ( .A1(n2259), .A2(n3407), .ZN(n3408) );
  NAND2_X1 U3974 ( .A1(n3594), .A2(DATAI_25_), .ZN(n3945) );
  OAI22_X1 U3975 ( .A1(n3962), .A2(n3401), .B1(n3460), .B2(n3945), .ZN(n3412)
         );
  OAI22_X1 U3976 ( .A1(n3962), .A2(n3457), .B1(n3401), .B2(n3945), .ZN(n3501)
         );
  OAI21_X1 U3977 ( .B1(n3413), .B2(n3502), .A(n3501), .ZN(n3415) );
  NAND2_X1 U3978 ( .A1(n3413), .A2(n3502), .ZN(n3414) );
  NAND2_X1 U3979 ( .A1(n2260), .A2(REG0_REG_26__SCAN_IN), .ZN(n3422) );
  INV_X1 U3980 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3928) );
  OR2_X1 U3981 ( .A1(n2693), .A2(n3928), .ZN(n3421) );
  INV_X1 U3982 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U3983 ( .A1(n3416), .A2(n3561), .ZN(n3417) );
  NAND2_X1 U3984 ( .A1(n3430), .A2(n3417), .ZN(n3927) );
  INV_X1 U3985 ( .A(REG1_REG_26__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U3986 ( .A1(n3594), .A2(DATAI_26_), .ZN(n3838) );
  NOR2_X1 U3987 ( .A1(n3838), .A2(n3460), .ZN(n3423) );
  AOI21_X1 U3988 ( .B1(n3909), .B2(n3437), .A(n3423), .ZN(n3424) );
  XNOR2_X1 U3989 ( .A(n3424), .B(n3458), .ZN(n3427) );
  NOR2_X1 U3990 ( .A1(n3838), .A2(n3401), .ZN(n3425) );
  AOI21_X1 U3991 ( .B1(n3909), .B2(n2736), .A(n3425), .ZN(n3426) );
  NOR2_X1 U3992 ( .A1(n3427), .A2(n3426), .ZN(n3559) );
  NAND2_X1 U3993 ( .A1(n3427), .A2(n3426), .ZN(n3558) );
  NAND2_X1 U3994 ( .A1(n3464), .A2(REG2_REG_27__SCAN_IN), .ZN(n3436) );
  INV_X1 U3995 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3428) );
  OR2_X1 U3996 ( .A1(n2259), .A2(n3428), .ZN(n3435) );
  INV_X1 U3997 ( .A(n3430), .ZN(n3429) );
  NAND2_X1 U3998 ( .A1(n3429), .A2(REG3_REG_27__SCAN_IN), .ZN(n3449) );
  INV_X1 U3999 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4245) );
  NAND2_X1 U4000 ( .A1(n3430), .A2(n4245), .ZN(n3431) );
  NAND2_X1 U4001 ( .A1(n3449), .A2(n3431), .ZN(n3912) );
  INV_X1 U4002 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3432) );
  OR2_X1 U4003 ( .A1(n2740), .A2(n3432), .ZN(n3433) );
  NAND2_X1 U4004 ( .A1(n3922), .A2(n2263), .ZN(n3439) );
  NAND2_X1 U4005 ( .A1(n3594), .A2(DATAI_27_), .ZN(n3906) );
  OR2_X1 U4006 ( .A1(n3906), .A2(n3460), .ZN(n3438) );
  NAND2_X1 U4007 ( .A1(n3439), .A2(n3438), .ZN(n3441) );
  XNOR2_X1 U4008 ( .A(n3441), .B(n3440), .ZN(n3444) );
  INV_X1 U4009 ( .A(n3444), .ZN(n3446) );
  NOR2_X1 U4010 ( .A1(n3906), .A2(n3401), .ZN(n3442) );
  AOI21_X1 U4011 ( .B1(n3922), .B2(n2736), .A(n3442), .ZN(n3443) );
  INV_X1 U4012 ( .A(n3443), .ZN(n3445) );
  OR2_X1 U4013 ( .A1(n3444), .A2(n3443), .ZN(n3447) );
  OAI21_X1 U4014 ( .B1(n3446), .B2(n3445), .A(n3447), .ZN(n3475) );
  NAND2_X1 U4015 ( .A1(n3464), .A2(REG2_REG_28__SCAN_IN), .ZN(n3456) );
  INV_X1 U4016 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3448) );
  OR2_X1 U4017 ( .A1(n2740), .A2(n3448), .ZN(n3455) );
  INV_X1 U4018 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U4019 ( .A1(n3449), .A2(n4408), .ZN(n3450) );
  NAND2_X1 U4020 ( .A1(n3875), .A2(n3450), .ZN(n3463) );
  OR2_X1 U4021 ( .A1(n3451), .A2(n3463), .ZN(n3454) );
  INV_X1 U4022 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3452) );
  OR2_X1 U4023 ( .A1(n2259), .A2(n3452), .ZN(n3453) );
  NAND2_X1 U4024 ( .A1(n3594), .A2(DATAI_28_), .ZN(n3894) );
  OAI22_X1 U4025 ( .A1(n3907), .A2(n3457), .B1(n3401), .B2(n3894), .ZN(n3459)
         );
  XNOR2_X1 U4026 ( .A(n3459), .B(n3458), .ZN(n3462) );
  OAI22_X1 U4027 ( .A1(n3907), .A2(n3401), .B1(n3460), .B2(n3894), .ZN(n3461)
         );
  INV_X1 U4028 ( .A(n3463), .ZN(n3895) );
  OAI22_X1 U4029 ( .A1(n4834), .A2(n3894), .B1(STATE_REG_SCAN_IN), .B2(n4408), 
        .ZN(n3472) );
  NAND2_X1 U4030 ( .A1(n3464), .A2(REG2_REG_29__SCAN_IN), .ZN(n3470) );
  INV_X1 U4031 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3465) );
  OR2_X1 U4032 ( .A1(n2740), .A2(n3465), .ZN(n3469) );
  OR2_X1 U4033 ( .A1(n3451), .A2(n3875), .ZN(n3468) );
  INV_X1 U4034 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3466) );
  OR2_X1 U4035 ( .A1(n2259), .A2(n3466), .ZN(n3467) );
  OAI22_X1 U4036 ( .A1(n3888), .A2(n4913), .B1(n4830), .B2(n3840), .ZN(n3471)
         );
  AOI211_X1 U4037 ( .C1(n3565), .C2(n3895), .A(n3472), .B(n3471), .ZN(n3473)
         );
  OAI21_X1 U4038 ( .B1(n3474), .B2(n3567), .A(n3473), .ZN(U3217) );
  AOI21_X1 U4039 ( .B1(n3476), .B2(n3475), .A(n3567), .ZN(n3477) );
  INV_X1 U4040 ( .A(n3477), .ZN(n3482) );
  INV_X1 U4041 ( .A(n3912), .ZN(n3480) );
  OAI22_X1 U4042 ( .A1(n4834), .A2(n3906), .B1(STATE_REG_SCAN_IN), .B2(n4245), 
        .ZN(n3479) );
  INV_X1 U40430 ( .A(n3909), .ZN(n3938) );
  OAI22_X1 U4044 ( .A1(n3907), .A2(n4913), .B1(n4830), .B2(n3938), .ZN(n3478)
         );
  AOI211_X1 U4045 ( .C1(n3565), .C2(n3480), .A(n3479), .B(n3478), .ZN(n3481)
         );
  OAI21_X1 U4046 ( .B1(n3482), .B2(n2283), .A(n3481), .ZN(U3211) );
  NAND2_X1 U4047 ( .A1(n3483), .A2(n4925), .ZN(n3492) );
  AOI21_X1 U4048 ( .B1(n3542), .B2(n3486), .A(n3485), .ZN(n3491) );
  INV_X1 U4049 ( .A(n3981), .ZN(n3489) );
  OAI22_X1 U4050 ( .A1(n4834), .A2(n3991), .B1(STATE_REG_SCAN_IN), .B2(n4343), 
        .ZN(n3488) );
  OAI22_X1 U4051 ( .A1(n3833), .A2(n4913), .B1(n4830), .B2(n4912), .ZN(n3487)
         );
  AOI211_X1 U4052 ( .C1(n3565), .C2(n3489), .A(n3488), .B(n3487), .ZN(n3490)
         );
  OAI21_X1 U4053 ( .B1(n3492), .B2(n3491), .A(n3490), .ZN(U3213) );
  OAI21_X1 U4054 ( .B1(n3495), .B2(n3494), .A(n3493), .ZN(n3499) );
  AOI22_X1 U4055 ( .A1(n4899), .A2(n4922), .B1(n4921), .B2(n4091), .ZN(n3497)
         );
  NOR2_X1 U4056 ( .A1(STATE_REG_SCAN_IN), .A2(n4405), .ZN(n3812) );
  AOI21_X1 U4057 ( .B1(n4924), .B2(n4057), .A(n3812), .ZN(n3496) );
  OAI211_X1 U4058 ( .C1(n4930), .C2(n4060), .A(n3497), .B(n3496), .ZN(n3498)
         );
  AOI21_X1 U4059 ( .B1(n3499), .B2(n4925), .A(n3498), .ZN(n3500) );
  INV_X1 U4060 ( .A(n3500), .ZN(U3216) );
  XNOR2_X1 U4061 ( .A(n3502), .B(n3501), .ZN(n3503) );
  XNOR2_X1 U4062 ( .A(n3504), .B(n3503), .ZN(n3509) );
  INV_X1 U4063 ( .A(n3947), .ZN(n3507) );
  OAI22_X1 U4064 ( .A1(n4834), .A2(n3945), .B1(STATE_REG_SCAN_IN), .B2(n4412), 
        .ZN(n3506) );
  OAI22_X1 U4065 ( .A1(n3833), .A2(n4830), .B1(n4913), .B2(n3938), .ZN(n3505)
         );
  AOI211_X1 U4066 ( .C1(n3565), .C2(n3507), .A(n3506), .B(n3505), .ZN(n3508)
         );
  OAI21_X1 U4067 ( .B1(n3509), .B2(n3567), .A(n3508), .ZN(U3222) );
  INV_X1 U4068 ( .A(n3510), .ZN(n3513) );
  INV_X1 U4069 ( .A(n3511), .ZN(n4837) );
  AOI21_X1 U4070 ( .B1(n3510), .B2(n3511), .A(n4838), .ZN(n3512) );
  AOI21_X1 U4071 ( .B1(n3513), .B2(n4837), .A(n3512), .ZN(n3517) );
  NAND2_X1 U4072 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  XNOR2_X1 U4073 ( .A(n3517), .B(n3516), .ZN(n3521) );
  AOI22_X1 U4074 ( .A1(n4921), .A2(n4106), .B1(n4899), .B2(n4103), .ZN(n3520)
         );
  NOR2_X1 U4075 ( .A1(STATE_REG_SCAN_IN), .A2(n4413), .ZN(n4601) );
  NOR2_X1 U4076 ( .A1(n4930), .A2(n4114), .ZN(n3518) );
  AOI211_X1 U4077 ( .C1(n4113), .C2(n4924), .A(n4601), .B(n3518), .ZN(n3519)
         );
  OAI211_X1 U4078 ( .C1(n3521), .C2(n3567), .A(n3520), .B(n3519), .ZN(U3223)
         );
  INV_X1 U4079 ( .A(n3523), .ZN(n3525) );
  NAND2_X1 U4080 ( .A1(n3525), .A2(n3524), .ZN(n3526) );
  XNOR2_X1 U4081 ( .A(n3522), .B(n3526), .ZN(n3530) );
  AOI22_X1 U4082 ( .A1(n4921), .A2(n4861), .B1(n4899), .B2(n4091), .ZN(n3529)
         );
  INV_X1 U4083 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4339) );
  NOR2_X1 U4084 ( .A1(STATE_REG_SCAN_IN), .A2(n4339), .ZN(n3790) );
  NOR2_X1 U4085 ( .A1(n4930), .A2(n4097), .ZN(n3527) );
  AOI211_X1 U4086 ( .C1(n4094), .C2(n4924), .A(n3790), .B(n3527), .ZN(n3528)
         );
  OAI211_X1 U4087 ( .C1(n3530), .C2(n3567), .A(n3529), .B(n3528), .ZN(U3225)
         );
  INV_X1 U4088 ( .A(n3531), .ZN(n3532) );
  NOR2_X1 U4089 ( .A1(n3533), .A2(n3532), .ZN(n3535) );
  XNOR2_X1 U4090 ( .A(n3535), .B(n3534), .ZN(n3540) );
  INV_X1 U4091 ( .A(n3965), .ZN(n3538) );
  OAI22_X1 U4092 ( .A1(n4834), .A2(n3968), .B1(STATE_REG_SCAN_IN), .B2(n4421), 
        .ZN(n3537) );
  INV_X1 U4093 ( .A(n3960), .ZN(n4005) );
  OAI22_X1 U4094 ( .A1(n4005), .A2(n4830), .B1(n4913), .B2(n3962), .ZN(n3536)
         );
  AOI211_X1 U4095 ( .C1(n3565), .C2(n3538), .A(n3537), .B(n3536), .ZN(n3539)
         );
  OAI21_X1 U4096 ( .B1(n3540), .B2(n3567), .A(n3539), .ZN(U3226) );
  OAI21_X1 U4097 ( .B1(n3543), .B2(n3541), .A(n3542), .ZN(n3547) );
  AOI22_X1 U4098 ( .A1(n4899), .A2(n3960), .B1(n4921), .B2(n4898), .ZN(n3545)
         );
  AOI22_X1 U4099 ( .A1(n4924), .A2(n4008), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3544) );
  OAI211_X1 U4100 ( .C1(n4930), .C2(n4009), .A(n3545), .B(n3544), .ZN(n3546)
         );
  AOI21_X1 U4101 ( .B1(n3547), .B2(n4925), .A(n3546), .ZN(n3548) );
  INV_X1 U4102 ( .A(n3548), .ZN(U3232) );
  XNOR2_X1 U4103 ( .A(n3550), .B(n3549), .ZN(n3551) );
  XNOR2_X1 U4104 ( .A(n3552), .B(n3551), .ZN(n3556) );
  AOI22_X1 U4105 ( .A1(n4921), .A2(n4103), .B1(n4899), .B2(n4904), .ZN(n3555)
         );
  AND2_X1 U4106 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4616) );
  NOR2_X1 U4107 ( .A1(n4930), .A2(n4076), .ZN(n3553) );
  AOI211_X1 U4108 ( .C1(n4072), .C2(n4924), .A(n4616), .B(n3553), .ZN(n3554)
         );
  OAI211_X1 U4109 ( .C1(n3556), .C2(n3567), .A(n3555), .B(n3554), .ZN(U3235)
         );
  NOR2_X1 U4110 ( .A1(n3559), .A2(n2498), .ZN(n3560) );
  XNOR2_X1 U4111 ( .A(n3557), .B(n3560), .ZN(n3568) );
  INV_X1 U4112 ( .A(n3927), .ZN(n3564) );
  OAI22_X1 U4113 ( .A1(n4834), .A2(n3838), .B1(STATE_REG_SCAN_IN), .B2(n3561), 
        .ZN(n3563) );
  OAI22_X1 U4114 ( .A1(n3962), .A2(n4830), .B1(n4913), .B2(n3840), .ZN(n3562)
         );
  AOI211_X1 U4115 ( .C1(n3565), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3566)
         );
  OAI21_X1 U4116 ( .B1(n3568), .B2(n3567), .A(n3566), .ZN(U3237) );
  INV_X1 U4117 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3572) );
  NAND2_X1 U4118 ( .A1(n2260), .A2(REG0_REG_31__SCAN_IN), .ZN(n3571) );
  INV_X1 U4119 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3569) );
  OR2_X1 U4120 ( .A1(n2259), .A2(n3569), .ZN(n3570) );
  OAI211_X1 U4121 ( .C1(n2693), .C2(n3572), .A(n3571), .B(n3570), .ZN(n4145)
         );
  INV_X1 U4122 ( .A(n4145), .ZN(n3605) );
  NAND2_X1 U4123 ( .A1(n3594), .A2(DATAI_30_), .ZN(n3606) );
  INV_X1 U4124 ( .A(n3606), .ZN(n4155) );
  OR2_X1 U4125 ( .A1(n3962), .A2(n3936), .ZN(n3688) );
  NAND2_X1 U4126 ( .A1(n3993), .A2(n3968), .ZN(n3933) );
  INV_X1 U4127 ( .A(n4072), .ZN(n4069) );
  NAND2_X1 U4128 ( .A1(n4091), .A2(n4069), .ZN(n4049) );
  NAND2_X1 U4129 ( .A1(n4904), .A2(n3682), .ZN(n3573) );
  AND2_X1 U4130 ( .A1(n4049), .A2(n3573), .ZN(n3584) );
  INV_X1 U4131 ( .A(n4094), .ZN(n4089) );
  NAND2_X1 U4132 ( .A1(n4103), .A2(n4089), .ZN(n4044) );
  NAND2_X1 U4133 ( .A1(n4217), .A2(n3576), .ZN(n3574) );
  NAND2_X1 U4134 ( .A1(n3575), .A2(n3643), .ZN(n3578) );
  NOR2_X1 U4135 ( .A1(n4217), .A2(n3576), .ZN(n3577) );
  AOI21_X1 U4136 ( .B1(n3643), .B2(n3708), .A(n3577), .ZN(n3646) );
  NAND2_X1 U4137 ( .A1(n3578), .A2(n3646), .ZN(n3845) );
  INV_X1 U4138 ( .A(n4129), .ZN(n4123) );
  OR2_X1 U4139 ( .A1(n4106), .A2(n4852), .ZN(n3701) );
  NAND2_X1 U4140 ( .A1(n3846), .A2(n3701), .ZN(n3652) );
  NAND2_X1 U4141 ( .A1(n4850), .A2(n4123), .ZN(n3697) );
  INV_X1 U4142 ( .A(n3697), .ZN(n3580) );
  NAND2_X1 U4143 ( .A1(n4106), .A2(n4852), .ZN(n3850) );
  INV_X1 U4144 ( .A(n3850), .ZN(n3579) );
  AOI21_X1 U4145 ( .B1(n3580), .B2(n3701), .A(n3579), .ZN(n3650) );
  OAI21_X1 U4146 ( .B1(n3845), .B2(n3652), .A(n3650), .ZN(n3581) );
  NAND2_X1 U4147 ( .A1(n4922), .A2(n4037), .ZN(n3702) );
  INV_X1 U4148 ( .A(n3702), .ZN(n3854) );
  AOI211_X1 U4149 ( .C1(n3581), .C2(n3687), .A(n3686), .B(n3854), .ZN(n3587)
         );
  OR2_X1 U4150 ( .A1(n4103), .A2(n4089), .ZN(n4046) );
  NAND2_X1 U4151 ( .A1(n4048), .A2(n4046), .ZN(n3583) );
  NOR2_X1 U4152 ( .A1(n4904), .A2(n3682), .ZN(n3582) );
  AOI21_X1 U4153 ( .B1(n3584), .B2(n3583), .A(n3582), .ZN(n4026) );
  OR2_X1 U4154 ( .A1(n4922), .A2(n4037), .ZN(n3703) );
  NAND2_X1 U4155 ( .A1(n4026), .A2(n3703), .ZN(n3585) );
  NAND2_X1 U4156 ( .A1(n3585), .A2(n3702), .ZN(n3853) );
  INV_X1 U4157 ( .A(n3853), .ZN(n3586) );
  NAND2_X1 U4158 ( .A1(n4912), .A2(n4008), .ZN(n3987) );
  OR2_X1 U4159 ( .A1(n4898), .A2(n4020), .ZN(n3984) );
  NAND2_X1 U4160 ( .A1(n3987), .A2(n3984), .ZN(n3856) );
  AOI211_X1 U4161 ( .C1(n3852), .C2(n3587), .A(n3586), .B(n3856), .ZN(n3590)
         );
  AND2_X1 U4162 ( .A1(n4898), .A2(n4020), .ZN(n3985) );
  AND2_X1 U4163 ( .A1(n3987), .A2(n3985), .ZN(n3588) );
  OR2_X1 U4164 ( .A1(n4912), .A2(n4008), .ZN(n3700) );
  NAND2_X1 U4165 ( .A1(n3960), .A2(n3991), .ZN(n3679) );
  NAND2_X1 U4166 ( .A1(n3700), .A2(n3679), .ZN(n3661) );
  NOR2_X1 U4167 ( .A1(n3588), .A2(n3661), .ZN(n3855) );
  INV_X1 U4168 ( .A(n3855), .ZN(n3589) );
  OR2_X1 U4169 ( .A1(n3960), .A2(n3991), .ZN(n3954) );
  OR2_X1 U4170 ( .A1(n3993), .A2(n3968), .ZN(n3680) );
  OAI21_X1 U4171 ( .B1(n3590), .B2(n3589), .A(n3857), .ZN(n3597) );
  INV_X1 U4172 ( .A(n3888), .ZN(n3736) );
  NAND2_X1 U4173 ( .A1(n3594), .A2(DATAI_29_), .ZN(n3879) );
  INV_X1 U4174 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U4175 ( .A1(n2261), .A2(REG0_REG_30__SCAN_IN), .ZN(n3593) );
  INV_X1 U4176 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3591) );
  OR2_X1 U4177 ( .A1(n2259), .A2(n3591), .ZN(n3592) );
  OAI211_X1 U4178 ( .C1(n2693), .C2(n4933), .A(n3593), .B(n3592), .ZN(n3868)
         );
  INV_X1 U4179 ( .A(n3868), .ZN(n3596) );
  NAND2_X1 U4180 ( .A1(n3594), .A2(DATAI_31_), .ZN(n4146) );
  NAND2_X1 U4181 ( .A1(n4145), .A2(n4146), .ZN(n3672) );
  INV_X1 U4182 ( .A(n3672), .ZN(n3595) );
  AOI21_X1 U4183 ( .B1(n4155), .B2(n3596), .A(n3595), .ZN(n3684) );
  OAI21_X1 U4184 ( .B1(n3736), .B2(n3879), .A(n3684), .ZN(n3599) );
  INV_X1 U4185 ( .A(n3894), .ZN(n3842) );
  NOR2_X1 U4186 ( .A1(n3922), .A2(n3906), .ZN(n3862) );
  OR2_X1 U4187 ( .A1(n3863), .A2(n3862), .ZN(n3600) );
  AOI211_X1 U4188 ( .C1(n3858), .C2(n3597), .A(n3599), .B(n3600), .ZN(n3603)
         );
  NAND2_X1 U4189 ( .A1(n3962), .A2(n3936), .ZN(n3918) );
  OR2_X1 U4190 ( .A1(n3909), .A2(n3838), .ZN(n3678) );
  NAND2_X1 U4191 ( .A1(n3918), .A2(n3678), .ZN(n3860) );
  INV_X1 U4192 ( .A(n3860), .ZN(n3664) );
  NOR2_X1 U4193 ( .A1(n3907), .A2(n3842), .ZN(n3864) );
  INV_X1 U4194 ( .A(n3879), .ZN(n3878) );
  NOR2_X1 U4195 ( .A1(n3888), .A2(n3878), .ZN(n3598) );
  OR2_X1 U4196 ( .A1(n3864), .A2(n3598), .ZN(n3666) );
  INV_X1 U4197 ( .A(n3666), .ZN(n3601) );
  AOI21_X1 U4198 ( .B1(n3600), .B2(n3601), .A(n3599), .ZN(n3671) );
  INV_X1 U4199 ( .A(n3906), .ZN(n3902) );
  XNOR2_X1 U4200 ( .A(n3922), .B(n3902), .ZN(n3861) );
  NAND2_X1 U4201 ( .A1(n3909), .A2(n3838), .ZN(n3859) );
  NAND3_X1 U4202 ( .A1(n3861), .A2(n3601), .A3(n3859), .ZN(n3602) );
  AOI22_X1 U4203 ( .A1(n3603), .A2(n3664), .B1(n3671), .B2(n3602), .ZN(n3604)
         );
  AOI21_X1 U4204 ( .B1(n3605), .B2(n4155), .A(n3604), .ZN(n3610) );
  OR2_X1 U4205 ( .A1(n4145), .A2(n4146), .ZN(n3608) );
  NAND2_X1 U4206 ( .A1(n3868), .A2(n3606), .ZN(n3607) );
  NAND2_X1 U4207 ( .A1(n3608), .A2(n3607), .ZN(n3673) );
  INV_X1 U4208 ( .A(n3673), .ZN(n3685) );
  NOR2_X1 U4209 ( .A1(n3685), .A2(n4146), .ZN(n3609) );
  NOR2_X1 U4210 ( .A1(n3610), .A2(n3609), .ZN(n3726) );
  INV_X1 U4211 ( .A(n3687), .ZN(n3658) );
  NAND2_X1 U4212 ( .A1(n3742), .A2(n3611), .ZN(n3704) );
  OAI211_X1 U4213 ( .C1(n3614), .C2(n3613), .A(n3704), .B(n3612), .ZN(n3617)
         );
  NAND3_X1 U4214 ( .A1(n3617), .A2(n3616), .A3(n3615), .ZN(n3619) );
  OAI211_X1 U4215 ( .C1(n3621), .C2(n3620), .A(n3619), .B(n3618), .ZN(n3624)
         );
  NAND3_X1 U4216 ( .A1(n3624), .A2(n3623), .A3(n3622), .ZN(n3627) );
  NAND4_X1 U4217 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3638), .ZN(n3630)
         );
  NAND3_X1 U4218 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n3636) );
  AND3_X1 U4219 ( .A1(n2319), .A2(n3632), .A3(n3631), .ZN(n3637) );
  AOI21_X1 U4220 ( .B1(n3696), .B2(n3634), .A(n3633), .ZN(n3635) );
  AOI21_X1 U4221 ( .B1(n3636), .B2(n3637), .A(n3635), .ZN(n3656) );
  INV_X1 U4222 ( .A(n3643), .ZN(n3649) );
  INV_X1 U4223 ( .A(n3637), .ZN(n3641) );
  INV_X1 U4224 ( .A(n3638), .ZN(n3640) );
  NOR3_X1 U4225 ( .A1(n3641), .A2(n3640), .A3(n3639), .ZN(n3645) );
  INV_X1 U4226 ( .A(n3710), .ZN(n3644) );
  AND3_X1 U4227 ( .A1(n3643), .A2(n3642), .A3(n3709), .ZN(n3653) );
  OAI21_X1 U4228 ( .B1(n3645), .B2(n3644), .A(n3653), .ZN(n3647) );
  OAI211_X1 U4229 ( .C1(n3649), .C2(n3648), .A(n3647), .B(n3646), .ZN(n3651)
         );
  OAI21_X1 U4230 ( .B1(n3652), .B2(n3651), .A(n3650), .ZN(n3655) );
  NAND3_X1 U4231 ( .A1(n3653), .A2(n3697), .A3(n3850), .ZN(n3654) );
  AOI221_X1 U4232 ( .B1(n3656), .B2(n3655), .C1(n3654), .C2(n3655), .A(n3686), 
        .ZN(n3657) );
  OAI211_X1 U4233 ( .C1(n3658), .C2(n3657), .A(n3852), .B(n3702), .ZN(n3659)
         );
  AOI21_X1 U4234 ( .B1(n3659), .B2(n3853), .A(n3985), .ZN(n3660) );
  NOR2_X1 U4235 ( .A1(n3660), .A2(n3856), .ZN(n3662) );
  OAI21_X1 U4236 ( .B1(n3662), .B2(n3661), .A(n3857), .ZN(n3663) );
  NAND2_X1 U4237 ( .A1(n3663), .A2(n3858), .ZN(n3665) );
  NAND2_X1 U4238 ( .A1(n3665), .A2(n3664), .ZN(n3670) );
  NOR2_X1 U4239 ( .A1(n3902), .A2(n3840), .ZN(n3668) );
  INV_X1 U4240 ( .A(n3859), .ZN(n3667) );
  NOR4_X1 U4241 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3673), .ZN(n3669)
         );
  NAND2_X1 U4242 ( .A1(n3670), .A2(n3669), .ZN(n3677) );
  INV_X1 U4243 ( .A(n3671), .ZN(n3675) );
  NAND2_X1 U4244 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  NAND2_X1 U4245 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  AOI21_X1 U4246 ( .B1(n3677), .B2(n3676), .A(n2570), .ZN(n3724) );
  NAND2_X1 U4247 ( .A1(n3954), .A2(n3679), .ZN(n3990) );
  NAND2_X1 U4248 ( .A1(n3680), .A2(n3933), .ZN(n3956) );
  INV_X1 U4249 ( .A(n3985), .ZN(n3681) );
  NAND2_X1 U4250 ( .A1(n3681), .A2(n3984), .ZN(n4018) );
  XNOR2_X1 U4251 ( .A(n4904), .B(n3682), .ZN(n4052) );
  NOR4_X1 U4252 ( .A1(n3990), .A2(n3956), .A3(n4018), .A4(n4052), .ZN(n3683)
         );
  NAND4_X1 U4253 ( .A1(n3921), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3718)
         );
  INV_X1 U4254 ( .A(n4118), .ZN(n3690) );
  NAND2_X1 U4255 ( .A1(n3688), .A2(n3918), .ZN(n3942) );
  NOR3_X1 U4256 ( .A1(n3690), .A2(n3689), .A3(n3942), .ZN(n3694) );
  NAND4_X1 U4257 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3717)
         );
  NAND2_X1 U4258 ( .A1(n4048), .A2(n4049), .ZN(n3821) );
  NOR4_X1 U4259 ( .A1(n3695), .A2(n3821), .A3(n4785), .A4(n4726), .ZN(n3715)
         );
  NAND2_X1 U4260 ( .A1(n2319), .A2(n3696), .ZN(n4757) );
  NAND2_X1 U4261 ( .A1(n3846), .A2(n3697), .ZN(n4125) );
  NOR4_X1 U4262 ( .A1(n4757), .A2(n3699), .A3(n4125), .A4(n3698), .ZN(n3714)
         );
  INV_X1 U4263 ( .A(n4002), .ZN(n4000) );
  NAND2_X1 U4264 ( .A1(n3701), .A2(n3850), .ZN(n4857) );
  NAND2_X1 U4265 ( .A1(n3703), .A2(n3702), .ZN(n4031) );
  NAND2_X1 U4266 ( .A1(n3705), .A2(n3704), .ZN(n4672) );
  NOR4_X1 U4267 ( .A1(n4000), .A2(n4857), .A3(n4031), .A4(n4672), .ZN(n3713)
         );
  NAND2_X1 U4268 ( .A1(n4046), .A2(n4044), .ZN(n4088) );
  INV_X1 U4269 ( .A(n3706), .ZN(n3707) );
  OR2_X1 U4270 ( .A1(n3708), .A2(n3707), .ZN(n4219) );
  NAND2_X1 U4271 ( .A1(n3710), .A2(n3709), .ZN(n4223) );
  NOR4_X1 U4272 ( .A1(n4088), .A2(n4219), .A3(n4223), .A4(n3711), .ZN(n3712)
         );
  NAND4_X1 U4273 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3716)
         );
  NOR3_X1 U4274 ( .A1(n3718), .A2(n3717), .A3(n3716), .ZN(n3720) );
  XNOR2_X1 U4275 ( .A(n3888), .B(n3879), .ZN(n3865) );
  INV_X1 U4276 ( .A(n3886), .ZN(n3719) );
  NAND4_X1 U4277 ( .A1(n3720), .A2(n3865), .A3(n3719), .A4(n3861), .ZN(n3722)
         );
  AOI21_X1 U4278 ( .B1(n3722), .B2(n3721), .A(n4668), .ZN(n3723) );
  OAI22_X1 U4279 ( .A1(n3726), .A2(n3725), .B1(n3724), .B2(n3723), .ZN(n3727)
         );
  INV_X1 U4280 ( .A(n3727), .ZN(n3728) );
  MUX2_X1 U4281 ( .A(n3728), .B(n3727), .S(n3808), .Z(n3735) );
  NAND2_X1 U4282 ( .A1(n3729), .A2(n3808), .ZN(n3730) );
  NOR4_X1 U4283 ( .A1(n3401), .A2(n4639), .A3(n4932), .A4(n3730), .ZN(n3732)
         );
  MUX2_X1 U4284 ( .A(n3733), .B(n3732), .S(n3731), .Z(n3734) );
  INV_X1 U4285 ( .A(B_REG_SCAN_IN), .ZN(n3869) );
  OAI22_X1 U4286 ( .A1(n3735), .A2(n4469), .B1(n3734), .B2(n3869), .ZN(U3239)
         );
  MUX2_X1 U4287 ( .A(n4145), .B(DATAO_REG_31__SCAN_IN), .S(n3741), .Z(U3581)
         );
  MUX2_X1 U4288 ( .A(n3868), .B(DATAO_REG_30__SCAN_IN), .S(n3741), .Z(U3580)
         );
  MUX2_X1 U4289 ( .A(DATAO_REG_29__SCAN_IN), .B(n3736), .S(U4043), .Z(U3579)
         );
  INV_X1 U4290 ( .A(n3907), .ZN(n3841) );
  MUX2_X1 U4291 ( .A(DATAO_REG_28__SCAN_IN), .B(n3841), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4292 ( .A(n3922), .B(DATAO_REG_27__SCAN_IN), .S(n3741), .Z(U3577)
         );
  MUX2_X1 U4293 ( .A(n3909), .B(DATAO_REG_26__SCAN_IN), .S(n3741), .Z(U3576)
         );
  INV_X1 U4294 ( .A(n3962), .ZN(n3835) );
  MUX2_X1 U4295 ( .A(DATAO_REG_25__SCAN_IN), .B(n3835), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4296 ( .A(n3993), .B(DATAO_REG_24__SCAN_IN), .S(n3741), .Z(U3574)
         );
  MUX2_X1 U4297 ( .A(n3960), .B(DATAO_REG_23__SCAN_IN), .S(n3741), .Z(U3573)
         );
  MUX2_X1 U4298 ( .A(n4898), .B(DATAO_REG_21__SCAN_IN), .S(n3741), .Z(U3571)
         );
  MUX2_X1 U4299 ( .A(n4922), .B(DATAO_REG_20__SCAN_IN), .S(n3741), .Z(U3570)
         );
  MUX2_X1 U4300 ( .A(n4904), .B(DATAO_REG_19__SCAN_IN), .S(n3741), .Z(U3569)
         );
  MUX2_X1 U4301 ( .A(n4091), .B(DATAO_REG_18__SCAN_IN), .S(n3741), .Z(U3568)
         );
  MUX2_X1 U4302 ( .A(n4103), .B(DATAO_REG_17__SCAN_IN), .S(n3741), .Z(U3567)
         );
  MUX2_X1 U4303 ( .A(n4861), .B(DATAO_REG_16__SCAN_IN), .S(n3741), .Z(U3566)
         );
  MUX2_X1 U4304 ( .A(n4106), .B(DATAO_REG_15__SCAN_IN), .S(n3741), .Z(U3565)
         );
  MUX2_X1 U4305 ( .A(n4850), .B(DATAO_REG_14__SCAN_IN), .S(n3741), .Z(U3564)
         );
  MUX2_X1 U4306 ( .A(n4217), .B(DATAO_REG_13__SCAN_IN), .S(n3741), .Z(U3563)
         );
  MUX2_X1 U4307 ( .A(n4789), .B(DATAO_REG_12__SCAN_IN), .S(n3741), .Z(U3562)
         );
  MUX2_X1 U4308 ( .A(n3737), .B(DATAO_REG_11__SCAN_IN), .S(n3741), .Z(U3561)
         );
  MUX2_X1 U4309 ( .A(n4788), .B(DATAO_REG_10__SCAN_IN), .S(n3741), .Z(U3560)
         );
  MUX2_X1 U4310 ( .A(n4225), .B(DATAO_REG_9__SCAN_IN), .S(n3741), .Z(U3559) );
  MUX2_X1 U4311 ( .A(n4758), .B(DATAO_REG_8__SCAN_IN), .S(n3741), .Z(U3558) );
  MUX2_X1 U4312 ( .A(n3738), .B(DATAO_REG_7__SCAN_IN), .S(n3741), .Z(U3557) );
  MUX2_X1 U4313 ( .A(n4734), .B(DATAO_REG_6__SCAN_IN), .S(n3741), .Z(U3556) );
  MUX2_X1 U4314 ( .A(n3739), .B(DATAO_REG_5__SCAN_IN), .S(n3741), .Z(U3555) );
  MUX2_X1 U4315 ( .A(n2778), .B(DATAO_REG_4__SCAN_IN), .S(n3741), .Z(U3554) );
  MUX2_X1 U4316 ( .A(n2757), .B(DATAO_REG_3__SCAN_IN), .S(n3741), .Z(U3553) );
  MUX2_X1 U4317 ( .A(n3740), .B(DATAO_REG_2__SCAN_IN), .S(n3741), .Z(U3552) );
  MUX2_X1 U4318 ( .A(n2657), .B(DATAO_REG_1__SCAN_IN), .S(n3741), .Z(U3551) );
  MUX2_X1 U4319 ( .A(n3742), .B(DATAO_REG_0__SCAN_IN), .S(n3741), .Z(U3550) );
  NAND2_X1 U4320 ( .A1(n4570), .A2(REG1_REG_11__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U4321 ( .A1(n4583), .A2(n3745), .ZN(n3747) );
  INV_X1 U4322 ( .A(n3745), .ZN(n3746) );
  INV_X1 U4323 ( .A(n4583), .ZN(n4811) );
  NOR2_X1 U4324 ( .A1(n4820), .A2(n3153), .ZN(n4590) );
  AOI21_X1 U4325 ( .B1(n3751), .B2(n3750), .A(n2297), .ZN(n3763) );
  AOI21_X1 U4326 ( .B1(n4646), .B2(ADDR_REG_14__SCAN_IN), .A(n3752), .ZN(n3753) );
  OAI21_X1 U4327 ( .B1(n4612), .B2(n2445), .A(n3753), .ZN(n3762) );
  AOI22_X1 U4328 ( .A1(n4570), .A2(REG2_REG_11__SCAN_IN), .B1(n3093), .B2(
        n4783), .ZN(n4577) );
  NAND2_X1 U4329 ( .A1(n3754), .A2(n4467), .ZN(n3756) );
  NAND2_X1 U4330 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  XNOR2_X1 U4331 ( .A(n4811), .B(n3757), .ZN(n4585) );
  NAND2_X1 U4332 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U4333 ( .A1(n4583), .A2(n3757), .ZN(n3758) );
  NOR2_X1 U4334 ( .A1(n4820), .A2(n3150), .ZN(n4593) );
  AOI211_X1 U4335 ( .C1(n4133), .C2(n3760), .A(n3766), .B(n4650), .ZN(n3761)
         );
  AOI211_X1 U4336 ( .C1(n4609), .C2(n3763), .A(n3762), .B(n3761), .ZN(n3764)
         );
  INV_X1 U4337 ( .A(n3764), .ZN(U3254) );
  INV_X1 U4338 ( .A(n4465), .ZN(n3780) );
  AND2_X1 U4339 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4832) );
  OR2_X1 U4340 ( .A1(n4465), .A2(n3767), .ZN(n3769) );
  NAND2_X1 U4341 ( .A1(n4465), .A2(n3767), .ZN(n3768) );
  AND2_X1 U4342 ( .A1(n3769), .A2(n3768), .ZN(n3770) );
  AOI211_X1 U4343 ( .C1(n3771), .C2(n3770), .A(n2279), .B(n4650), .ZN(n3772)
         );
  AOI211_X1 U4344 ( .C1(n4646), .C2(ADDR_REG_15__SCAN_IN), .A(n4832), .B(n3772), .ZN(n3779) );
  OR2_X1 U4345 ( .A1(n4465), .A2(n3782), .ZN(n3774) );
  NAND2_X1 U4346 ( .A1(n4465), .A2(n3782), .ZN(n3773) );
  AND2_X1 U4347 ( .A1(n3774), .A2(n3773), .ZN(n3776) );
  NOR2_X1 U4348 ( .A1(n3775), .A2(n3776), .ZN(n3784) );
  AOI21_X1 U4349 ( .B1(n3776), .B2(n3775), .A(n3784), .ZN(n3777) );
  NAND2_X1 U4350 ( .A1(n4609), .A2(n3777), .ZN(n3778) );
  OAI211_X1 U4351 ( .C1(n4612), .C2(n3780), .A(n3779), .B(n3778), .ZN(U3255)
         );
  INV_X1 U4352 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4893) );
  NOR2_X1 U4353 ( .A1(n2433), .A2(n4893), .ZN(n3781) );
  AOI21_X1 U4354 ( .B1(n4893), .B2(n2433), .A(n3781), .ZN(n3788) );
  XNOR2_X1 U4355 ( .A(n3785), .B(n3276), .ZN(n4603) );
  NAND2_X1 U4356 ( .A1(n3785), .A2(n4877), .ZN(n3786) );
  NAND2_X1 U4357 ( .A1(n3800), .A2(n3788), .ZN(n3787) );
  OAI21_X1 U4358 ( .B1(n3788), .B2(n3800), .A(n3787), .ZN(n3789) );
  AOI22_X1 U4359 ( .A1(n3789), .A2(n4609), .B1(n4656), .B2(n3805), .ZN(n3799)
         );
  AOI21_X1 U4360 ( .B1(n4646), .B2(ADDR_REG_17__SCAN_IN), .A(n3790), .ZN(n3798) );
  XNOR2_X1 U4361 ( .A(n3805), .B(n4098), .ZN(n3795) );
  INV_X1 U4362 ( .A(n3792), .ZN(n3791) );
  NAND2_X1 U4363 ( .A1(n3791), .A2(n4877), .ZN(n3793) );
  OAI21_X1 U4364 ( .B1(n3795), .B2(n3794), .A(n3804), .ZN(n3796) );
  NAND2_X1 U4365 ( .A1(n4607), .A2(n3796), .ZN(n3797) );
  NAND3_X1 U4366 ( .A1(n3799), .A2(n3798), .A3(n3797), .ZN(U3257) );
  AOI21_X1 U4367 ( .B1(n2278), .B2(n2433), .A(n3801), .ZN(n4617) );
  XOR2_X1 U4368 ( .A(REG1_REG_18__SCAN_IN), .B(n4621), .Z(n4618) );
  NAND2_X1 U4369 ( .A1(n4617), .A2(n4618), .ZN(n4623) );
  INV_X1 U4370 ( .A(n4621), .ZN(n3802) );
  NAND2_X1 U4371 ( .A1(n4623), .A2(n2507), .ZN(n3803) );
  NAND2_X1 U4372 ( .A1(n4621), .A2(REG2_REG_18__SCAN_IN), .ZN(n3806) );
  OAI21_X1 U4373 ( .B1(n4621), .B2(REG2_REG_18__SCAN_IN), .A(n3806), .ZN(n4614) );
  XNOR2_X1 U4374 ( .A(n3807), .B(REG2_REG_19__SCAN_IN), .ZN(n3810) );
  AOI21_X1 U4375 ( .B1(n4646), .B2(ADDR_REG_19__SCAN_IN), .A(n3812), .ZN(n3813) );
  NAND2_X1 U4376 ( .A1(n4106), .A2(n3815), .ZN(n3817) );
  AND3_X1 U4377 ( .A1(n4125), .A2(n3817), .A3(n4136), .ZN(n3816) );
  NOR2_X1 U4378 ( .A1(n4850), .A2(n4129), .ZN(n4843) );
  INV_X1 U4379 ( .A(n4106), .ZN(n4124) );
  AOI22_X1 U4380 ( .A1(n4843), .A2(n3817), .B1(n4124), .B2(n4852), .ZN(n3818)
         );
  NAND2_X1 U4381 ( .A1(n3819), .A2(n3818), .ZN(n4119) );
  NAND2_X1 U4382 ( .A1(n4861), .A2(n4113), .ZN(n3820) );
  INV_X1 U4383 ( .A(n4081), .ZN(n3822) );
  NAND2_X1 U4384 ( .A1(n3822), .A2(n3821), .ZN(n4080) );
  OR2_X1 U4385 ( .A1(n4091), .A2(n4072), .ZN(n3823) );
  NAND2_X1 U4386 ( .A1(n4904), .A2(n4057), .ZN(n3825) );
  NOR2_X1 U4387 ( .A1(n4904), .A2(n4057), .ZN(n3824) );
  INV_X1 U4388 ( .A(n4922), .ZN(n3826) );
  NAND2_X1 U4389 ( .A1(n3826), .A2(n4037), .ZN(n3828) );
  INV_X1 U4390 ( .A(n4037), .ZN(n4905) );
  NAND2_X1 U4391 ( .A1(n4898), .A2(n4923), .ZN(n3974) );
  NOR2_X1 U4392 ( .A1(n4898), .A2(n4923), .ZN(n3975) );
  NOR2_X1 U4393 ( .A1(n4912), .A2(n3831), .ZN(n3977) );
  INV_X1 U4394 ( .A(n3991), .ZN(n3980) );
  INV_X1 U4395 ( .A(n3968), .ZN(n3959) );
  NAND2_X1 U4396 ( .A1(n3941), .A2(n2508), .ZN(n3837) );
  NAND2_X1 U4397 ( .A1(n3837), .A2(n3836), .ZN(n3916) );
  INV_X1 U4398 ( .A(n3843), .ZN(n3844) );
  XNOR2_X1 U4399 ( .A(n3844), .B(n3865), .ZN(n4158) );
  INV_X1 U4400 ( .A(n4158), .ZN(n3884) );
  NAND2_X1 U4401 ( .A1(n3845), .A2(n4138), .ZN(n3847) );
  NAND2_X1 U4402 ( .A1(n3847), .A2(n3846), .ZN(n4858) );
  NAND2_X1 U4403 ( .A1(n4854), .A2(n3850), .ZN(n4105) );
  NAND2_X1 U4404 ( .A1(n4105), .A2(n4118), .ZN(n4104) );
  NAND2_X1 U4405 ( .A1(n3955), .A2(n3857), .ZN(n3934) );
  OAI22_X1 U4406 ( .A1(n3907), .A2(n4213), .B1(n3879), .B2(n4853), .ZN(n3867)
         );
  INV_X1 U4407 ( .A(n3867), .ZN(n3872) );
  OR2_X1 U4408 ( .A1(n4639), .A2(n3869), .ZN(n3870) );
  AND2_X1 U4409 ( .A1(n3870), .A2(n4862), .ZN(n4144) );
  NAND2_X1 U4410 ( .A1(n3868), .A2(n4144), .ZN(n3871) );
  NAND2_X1 U4411 ( .A1(n3979), .A2(n3968), .ZN(n3943) );
  INV_X1 U4412 ( .A(n3893), .ZN(n3880) );
  OAI21_X1 U4413 ( .B1(n3880), .B2(n3879), .A(n4150), .ZN(n4156) );
  INV_X1 U4414 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3881) );
  OAI22_X1 U4415 ( .A1(n4156), .A2(n4934), .B1(n3881), .B2(n4674), .ZN(n3882)
         );
  AOI21_X1 U4416 ( .B1(n2512), .B2(n4674), .A(n3882), .ZN(n3883) );
  OAI21_X1 U4417 ( .B1(n3884), .B2(n4140), .A(n3883), .ZN(U3354) );
  XNOR2_X1 U4418 ( .A(n3885), .B(n3886), .ZN(n4163) );
  XNOR2_X1 U4419 ( .A(n3887), .B(n3886), .ZN(n3891) );
  NOR2_X1 U4420 ( .A1(n3888), .A2(n4737), .ZN(n3890) );
  OAI22_X1 U4421 ( .A1(n3840), .A2(n4213), .B1(n4853), .B2(n3894), .ZN(n3889)
         );
  INV_X1 U4422 ( .A(n4162), .ZN(n3898) );
  OAI211_X1 U4423 ( .C1(n3892), .C2(n3894), .A(n4883), .B(n3893), .ZN(n4161)
         );
  AOI22_X1 U4424 ( .A1(n4939), .A2(REG2_REG_28__SCAN_IN), .B1(n3895), .B2(
        n4867), .ZN(n3896) );
  OAI21_X1 U4425 ( .B1(n4161), .B2(n4075), .A(n3896), .ZN(n3897) );
  AOI21_X1 U4426 ( .B1(n3898), .B2(n4674), .A(n3897), .ZN(n3899) );
  OAI21_X1 U4427 ( .B1(n4163), .B2(n4140), .A(n3899), .ZN(U3262) );
  XNOR2_X1 U4428 ( .A(n3900), .B(n3905), .ZN(n4167) );
  INV_X1 U4429 ( .A(n3901), .ZN(n4169) );
  AOI21_X1 U4430 ( .B1(n3902), .B2(n4169), .A(n3892), .ZN(n4165) );
  AOI22_X1 U4431 ( .A1(n4165), .A2(n4940), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4939), .ZN(n3915) );
  AOI21_X1 U4432 ( .B1(n3905), .B2(n3904), .A(n3903), .ZN(n3911) );
  OAI22_X1 U4433 ( .A1(n3907), .A2(n4737), .B1(n3906), .B2(n4853), .ZN(n3908)
         );
  AOI21_X1 U4434 ( .B1(n4849), .B2(n3909), .A(n3908), .ZN(n3910) );
  OAI21_X1 U4435 ( .B1(n3911), .B2(n4856), .A(n3910), .ZN(n4164) );
  NOR2_X1 U4436 ( .A1(n4741), .A2(n3912), .ZN(n3913) );
  OAI21_X1 U4437 ( .B1(n4164), .B2(n3913), .A(n4674), .ZN(n3914) );
  OAI211_X1 U4438 ( .C1(n4167), .C2(n4140), .A(n3915), .B(n3914), .ZN(U3263)
         );
  XOR2_X1 U4439 ( .A(n3921), .B(n3916), .Z(n4172) );
  INV_X1 U4440 ( .A(n3918), .ZN(n3919) );
  NOR2_X1 U4441 ( .A1(n3917), .A2(n3919), .ZN(n3920) );
  XOR2_X1 U4442 ( .A(n3921), .B(n3920), .Z(n3925) );
  AOI22_X1 U4443 ( .A1(n3922), .A2(n4862), .B1(n4787), .B2(n3926), .ZN(n3923)
         );
  OAI21_X1 U4444 ( .B1(n3962), .B2(n4213), .A(n3923), .ZN(n3924) );
  AOI21_X1 U4445 ( .B1(n3925), .B2(n4731), .A(n3924), .ZN(n4171) );
  INV_X1 U4446 ( .A(n4171), .ZN(n3931) );
  NAND2_X1 U4447 ( .A1(n3944), .A2(n3926), .ZN(n4168) );
  AND3_X1 U4448 ( .A1(n4169), .A2(n4940), .A3(n4168), .ZN(n3930) );
  OAI22_X1 U4449 ( .A1(n4674), .A2(n3928), .B1(n3927), .B2(n4741), .ZN(n3929)
         );
  AOI211_X1 U4450 ( .C1(n3931), .C2(n4674), .A(n3930), .B(n3929), .ZN(n3932)
         );
  OAI21_X1 U4451 ( .B1(n4172), .B2(n4140), .A(n3932), .ZN(U3264) );
  NAND2_X1 U4452 ( .A1(n3934), .A2(n3933), .ZN(n3935) );
  XNOR2_X1 U4453 ( .A(n3935), .B(n3942), .ZN(n3940) );
  AOI22_X1 U4454 ( .A1(n3993), .A2(n4849), .B1(n3936), .B2(n4787), .ZN(n3937)
         );
  OAI21_X1 U4455 ( .B1(n3938), .B2(n4737), .A(n3937), .ZN(n3939) );
  AOI21_X1 U4456 ( .B1(n3940), .B2(n4731), .A(n3939), .ZN(n4173) );
  XOR2_X1 U4457 ( .A(n3942), .B(n3941), .Z(n4176) );
  INV_X1 U4458 ( .A(n4140), .ZN(n4871) );
  NAND2_X1 U4459 ( .A1(n4176), .A2(n4871), .ZN(n3952) );
  INV_X1 U4460 ( .A(n3943), .ZN(n3946) );
  OAI21_X1 U4461 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n4174) );
  INV_X1 U4462 ( .A(n4174), .ZN(n3950) );
  INV_X1 U4463 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3948) );
  OAI22_X1 U4464 ( .A1(n4674), .A2(n3948), .B1(n3947), .B2(n4741), .ZN(n3949)
         );
  AOI21_X1 U4465 ( .B1(n3950), .B2(n4940), .A(n3949), .ZN(n3951) );
  OAI211_X1 U4466 ( .C1(n4939), .C2(n4173), .A(n3952), .B(n3951), .ZN(U3265)
         );
  XNOR2_X1 U4467 ( .A(n3953), .B(n3956), .ZN(n4181) );
  NAND2_X1 U4468 ( .A1(n3955), .A2(n3954), .ZN(n3958) );
  INV_X1 U4469 ( .A(n3956), .ZN(n3957) );
  XNOR2_X1 U4470 ( .A(n3958), .B(n3957), .ZN(n3964) );
  AOI22_X1 U4471 ( .A1(n3960), .A2(n4849), .B1(n4787), .B2(n3959), .ZN(n3961)
         );
  OAI21_X1 U4472 ( .B1(n3962), .B2(n4737), .A(n3961), .ZN(n3963) );
  AOI21_X1 U4473 ( .B1(n3964), .B2(n4731), .A(n3963), .ZN(n4180) );
  OAI22_X1 U4474 ( .A1(n4674), .A2(n3966), .B1(n3965), .B2(n4741), .ZN(n3967)
         );
  INV_X1 U4475 ( .A(n3967), .ZN(n3970) );
  OR2_X1 U4476 ( .A1(n3979), .A2(n3968), .ZN(n4178) );
  NAND3_X1 U4477 ( .A1(n4178), .A2(n3943), .A3(n4940), .ZN(n3969) );
  OAI211_X1 U4478 ( .C1(n4180), .C2(n4939), .A(n3970), .B(n3969), .ZN(n3971)
         );
  INV_X1 U4479 ( .A(n3971), .ZN(n3972) );
  OAI21_X1 U4480 ( .B1(n4181), .B2(n4140), .A(n3972), .ZN(U3266) );
  OAI21_X1 U4481 ( .B1(n3973), .B2(n3975), .A(n3974), .ZN(n4001) );
  INV_X1 U4482 ( .A(n4001), .ZN(n3976) );
  NOR2_X1 U4483 ( .A1(n3976), .A2(n4002), .ZN(n3998) );
  NOR2_X1 U4484 ( .A1(n3998), .A2(n3977), .ZN(n3978) );
  XOR2_X1 U4485 ( .A(n3990), .B(n3978), .Z(n4185) );
  AOI21_X1 U4486 ( .B1(n3980), .B2(n2291), .A(n3979), .ZN(n4183) );
  OAI22_X1 U4487 ( .A1(n4674), .A2(n3982), .B1(n3981), .B2(n4741), .ZN(n3983)
         );
  AOI21_X1 U4488 ( .B1(n4183), .B2(n4940), .A(n3983), .ZN(n3997) );
  INV_X1 U4489 ( .A(n4019), .ZN(n3986) );
  OAI21_X1 U4490 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n4003) );
  INV_X1 U4491 ( .A(n3987), .ZN(n3988) );
  AOI21_X1 U4492 ( .B1(n4003), .B2(n4002), .A(n3988), .ZN(n3989) );
  XOR2_X1 U4493 ( .A(n3990), .B(n3989), .Z(n3995) );
  OAI22_X1 U4494 ( .A1(n4912), .A2(n4213), .B1(n4853), .B2(n3991), .ZN(n3992)
         );
  AOI21_X1 U4495 ( .B1(n4862), .B2(n3993), .A(n3992), .ZN(n3994) );
  OAI21_X1 U4496 ( .B1(n3995), .B2(n4856), .A(n3994), .ZN(n4182) );
  NAND2_X1 U4497 ( .A1(n4182), .A2(n4674), .ZN(n3996) );
  OAI211_X1 U4498 ( .C1(n4185), .C2(n4140), .A(n3997), .B(n3996), .ZN(U3267)
         );
  INV_X1 U4499 ( .A(n3998), .ZN(n3999) );
  OAI21_X1 U4500 ( .B1(n4001), .B2(n4000), .A(n3999), .ZN(n4189) );
  XNOR2_X1 U4501 ( .A(n4003), .B(n4002), .ZN(n4007) );
  AOI22_X1 U4502 ( .A1(n4898), .A2(n4849), .B1(n4008), .B2(n4787), .ZN(n4004)
         );
  OAI21_X1 U4503 ( .B1(n4005), .B2(n4737), .A(n4004), .ZN(n4006) );
  AOI21_X1 U4504 ( .B1(n4007), .B2(n4731), .A(n4006), .ZN(n4188) );
  INV_X1 U4505 ( .A(n4188), .ZN(n4013) );
  NAND2_X1 U4506 ( .A1(n4015), .A2(n4008), .ZN(n4186) );
  AND3_X1 U4507 ( .A1(n2291), .A2(n4940), .A3(n4186), .ZN(n4012) );
  INV_X1 U4508 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4010) );
  OAI22_X1 U4509 ( .A1(n4674), .A2(n4010), .B1(n4009), .B2(n4741), .ZN(n4011)
         );
  AOI211_X1 U4510 ( .C1(n4013), .C2(n4674), .A(n4012), .B(n4011), .ZN(n4014)
         );
  OAI21_X1 U4511 ( .B1(n4189), .B2(n4140), .A(n4014), .ZN(U3268) );
  XOR2_X1 U4512 ( .A(n4018), .B(n3973), .Z(n4193) );
  AOI21_X1 U4513 ( .B1(n4923), .B2(n4036), .A(n2397), .ZN(n4191) );
  INV_X1 U4514 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4016) );
  OAI22_X1 U4515 ( .A1(n4674), .A2(n4016), .B1(n4929), .B2(n4741), .ZN(n4017)
         );
  AOI21_X1 U4516 ( .B1(n4191), .B2(n4940), .A(n4017), .ZN(n4025) );
  XNOR2_X1 U4517 ( .A(n4019), .B(n4018), .ZN(n4023) );
  OAI22_X1 U4518 ( .A1(n4912), .A2(n4737), .B1(n4853), .B2(n4020), .ZN(n4021)
         );
  AOI21_X1 U4519 ( .B1(n4849), .B2(n4922), .A(n4021), .ZN(n4022) );
  OAI21_X1 U4520 ( .B1(n4023), .B2(n4856), .A(n4022), .ZN(n4190) );
  NAND2_X1 U4521 ( .A1(n4190), .A2(n4674), .ZN(n4024) );
  OAI211_X1 U4522 ( .C1(n4193), .C2(n4140), .A(n4025), .B(n4024), .ZN(U3269)
         );
  NAND2_X1 U4523 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  XOR2_X1 U4524 ( .A(n4031), .B(n4028), .Z(n4035) );
  AOI22_X1 U4525 ( .A1(n4898), .A2(n4862), .B1(n4905), .B2(n4787), .ZN(n4029)
         );
  OAI21_X1 U4526 ( .B1(n4030), .B2(n4213), .A(n4029), .ZN(n4034) );
  XNOR2_X1 U4527 ( .A(n4032), .B(n4031), .ZN(n4196) );
  NOR2_X1 U4528 ( .A1(n4196), .A2(n4660), .ZN(n4033) );
  AOI211_X1 U4529 ( .C1(n4035), .C2(n4731), .A(n4034), .B(n4033), .ZN(n4195)
         );
  INV_X1 U4530 ( .A(n4196), .ZN(n4041) );
  OAI211_X1 U4531 ( .C1(n4056), .C2(n4037), .A(n4883), .B(n4036), .ZN(n4194)
         );
  INV_X1 U4532 ( .A(n4910), .ZN(n4038) );
  AOI22_X1 U4533 ( .A1(n4939), .A2(REG2_REG_20__SCAN_IN), .B1(n4038), .B2(
        n4867), .ZN(n4039) );
  OAI21_X1 U4534 ( .B1(n4194), .B2(n4075), .A(n4039), .ZN(n4040) );
  AOI21_X1 U4535 ( .B1(n4041), .B2(n4805), .A(n4040), .ZN(n4042) );
  OAI21_X1 U4536 ( .B1(n4195), .B2(n4939), .A(n4042), .ZN(U3270) );
  XOR2_X1 U4537 ( .A(n4052), .B(n4043), .Z(n4198) );
  INV_X1 U4538 ( .A(n4044), .ZN(n4045) );
  OR2_X1 U4539 ( .A1(n4087), .A2(n4045), .ZN(n4047) );
  NAND2_X1 U4540 ( .A1(n4047), .A2(n4046), .ZN(n4066) );
  INV_X1 U4541 ( .A(n4048), .ZN(n4050) );
  OAI21_X1 U4542 ( .B1(n4066), .B2(n4050), .A(n4049), .ZN(n4051) );
  XOR2_X1 U4543 ( .A(n4052), .B(n4051), .Z(n4055) );
  AOI22_X1 U4544 ( .A1(n4922), .A2(n4862), .B1(n4057), .B2(n4787), .ZN(n4054)
         );
  NAND2_X1 U4545 ( .A1(n4091), .A2(n4849), .ZN(n4053) );
  OAI211_X1 U4546 ( .C1(n4055), .C2(n4856), .A(n4054), .B(n4053), .ZN(n4200)
         );
  NAND2_X1 U4547 ( .A1(n4200), .A2(n4674), .ZN(n4065) );
  INV_X1 U4548 ( .A(n4056), .ZN(n4059) );
  NAND2_X1 U4549 ( .A1(n4074), .A2(n4057), .ZN(n4058) );
  NAND2_X1 U4550 ( .A1(n4059), .A2(n4058), .ZN(n4197) );
  INV_X1 U4551 ( .A(n4197), .ZN(n4063) );
  OAI22_X1 U4552 ( .A1(n4674), .A2(n4061), .B1(n4060), .B2(n4741), .ZN(n4062)
         );
  AOI21_X1 U4553 ( .B1(n4063), .B2(n4940), .A(n4062), .ZN(n4064) );
  OAI211_X1 U4554 ( .C1(n4198), .C2(n4140), .A(n4065), .B(n4064), .ZN(U3271)
         );
  XNOR2_X1 U4555 ( .A(n4066), .B(n4082), .ZN(n4071) );
  NAND2_X1 U4556 ( .A1(n4103), .A2(n4849), .ZN(n4068) );
  NAND2_X1 U4557 ( .A1(n4904), .A2(n4862), .ZN(n4067) );
  OAI211_X1 U4558 ( .C1(n4853), .C2(n4069), .A(n4068), .B(n4067), .ZN(n4070)
         );
  AOI21_X1 U4559 ( .B1(n4071), .B2(n4731), .A(n4070), .ZN(n4204) );
  AOI21_X1 U4560 ( .B1(n4096), .B2(n4072), .A(n4887), .ZN(n4073) );
  AND2_X1 U4561 ( .A1(n4074), .A2(n4073), .ZN(n4201) );
  INV_X1 U4562 ( .A(n4075), .ZN(n4079) );
  INV_X1 U4563 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4077) );
  OAI22_X1 U4564 ( .A1(n4674), .A2(n4077), .B1(n4076), .B2(n4741), .ZN(n4078)
         );
  AOI21_X1 U4565 ( .B1(n4201), .B2(n4079), .A(n4078), .ZN(n4085) );
  NAND2_X1 U4566 ( .A1(n4081), .A2(n4082), .ZN(n4083) );
  NAND2_X1 U4567 ( .A1(n4080), .A2(n4083), .ZN(n4202) );
  NAND2_X1 U4568 ( .A1(n4202), .A2(n4871), .ZN(n4084) );
  OAI211_X1 U4569 ( .C1(n4204), .C2(n4939), .A(n4085), .B(n4084), .ZN(U3272)
         );
  XNOR2_X1 U4570 ( .A(n4086), .B(n4088), .ZN(n4889) );
  XOR2_X1 U4571 ( .A(n4088), .B(n4087), .Z(n4093) );
  OAI22_X1 U4572 ( .A1(n4831), .A2(n4213), .B1(n4089), .B2(n4853), .ZN(n4090)
         );
  AOI21_X1 U4573 ( .B1(n4862), .B2(n4091), .A(n4090), .ZN(n4092) );
  OAI21_X1 U4574 ( .B1(n4093), .B2(n4856), .A(n4092), .ZN(n4891) );
  NAND2_X1 U4575 ( .A1(n4891), .A2(n4674), .ZN(n4102) );
  NAND2_X1 U4576 ( .A1(n4110), .A2(n4094), .ZN(n4095) );
  NAND2_X1 U4577 ( .A1(n4096), .A2(n4095), .ZN(n4886) );
  INV_X1 U4578 ( .A(n4886), .ZN(n4100) );
  OAI22_X1 U4579 ( .A1(n4674), .A2(n4098), .B1(n4097), .B2(n4741), .ZN(n4099)
         );
  AOI21_X1 U4580 ( .B1(n4100), .B2(n4940), .A(n4099), .ZN(n4101) );
  OAI211_X1 U4581 ( .C1(n4140), .C2(n4889), .A(n4102), .B(n4101), .ZN(U3273)
         );
  INV_X1 U4582 ( .A(n4103), .ZN(n4109) );
  OAI211_X1 U4583 ( .C1(n4105), .C2(n4118), .A(n4104), .B(n4731), .ZN(n4108)
         );
  AOI22_X1 U4584 ( .A1(n4106), .A2(n4849), .B1(n4113), .B2(n4787), .ZN(n4107)
         );
  OAI211_X1 U4585 ( .C1(n4109), .C2(n4737), .A(n4108), .B(n4107), .ZN(n4880)
         );
  INV_X1 U4586 ( .A(n4880), .ZN(n4122) );
  INV_X1 U4587 ( .A(n4848), .ZN(n4112) );
  INV_X1 U4588 ( .A(n4110), .ZN(n4111) );
  AOI21_X1 U4589 ( .B1(n4113), .B2(n4112), .A(n4111), .ZN(n4882) );
  OAI22_X1 U4590 ( .A1(n4674), .A2(n4115), .B1(n4114), .B2(n4741), .ZN(n4116)
         );
  AOI21_X1 U4591 ( .B1(n4882), .B2(n4940), .A(n4116), .ZN(n4121) );
  NAND2_X1 U4592 ( .A1(n4119), .A2(n4118), .ZN(n4878) );
  NAND3_X1 U4593 ( .A1(n4117), .A2(n4878), .A3(n4871), .ZN(n4120) );
  OAI211_X1 U4594 ( .C1(n4122), .C2(n4939), .A(n4121), .B(n4120), .ZN(U3274)
         );
  OAI22_X1 U4595 ( .A1(n4124), .A2(n4737), .B1(n4123), .B2(n4853), .ZN(n4128)
         );
  XNOR2_X1 U4596 ( .A(n3845), .B(n4125), .ZN(n4126) );
  NOR2_X1 U4597 ( .A1(n4126), .A2(n4856), .ZN(n4127) );
  AOI211_X1 U4598 ( .C1(n4849), .C2(n4217), .A(n4128), .B(n4127), .ZN(n4209)
         );
  AND2_X1 U4599 ( .A1(n4130), .A2(n4129), .ZN(n4131) );
  NOR2_X1 U4600 ( .A1(n4846), .A2(n4131), .ZN(n4207) );
  OAI22_X1 U4601 ( .A1(n4674), .A2(n4133), .B1(n4741), .B2(n4132), .ZN(n4142)
         );
  INV_X1 U4602 ( .A(n3814), .ZN(n4137) );
  INV_X1 U4603 ( .A(n4134), .ZN(n4135) );
  AOI21_X1 U4604 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4139) );
  NOR2_X1 U4605 ( .A1(n4139), .A2(n4138), .ZN(n4844) );
  AOI21_X1 U4606 ( .B1(n4139), .B2(n4138), .A(n4844), .ZN(n4210) );
  NOR2_X1 U4607 ( .A1(n4210), .A2(n4140), .ZN(n4141) );
  AOI211_X1 U4608 ( .C1(n4207), .C2(n4940), .A(n4142), .B(n4141), .ZN(n4143)
         );
  OAI21_X1 U4609 ( .B1(n4939), .B2(n4209), .A(n4143), .ZN(U3276) );
  NAND2_X1 U4610 ( .A1(n4145), .A2(n4144), .ZN(n4153) );
  OR2_X1 U4611 ( .A1(n4146), .A2(n4853), .ZN(n4147) );
  AND2_X1 U4612 ( .A1(n4153), .A2(n4147), .ZN(n4943) );
  INV_X1 U4613 ( .A(n4943), .ZN(n4148) );
  AOI21_X1 U4614 ( .B1(n4941), .B2(n4883), .A(n4148), .ZN(n4231) );
  MUX2_X1 U4615 ( .A(n3569), .B(n4231), .S(n4894), .Z(n4149) );
  INV_X1 U4616 ( .A(n4149), .ZN(U3549) );
  NAND2_X1 U4617 ( .A1(n4150), .A2(n4155), .ZN(n4151) );
  NAND2_X1 U4618 ( .A1(n4152), .A2(n4151), .ZN(n4935) );
  INV_X1 U4619 ( .A(n4153), .ZN(n4154) );
  AOI21_X1 U4620 ( .B1(n4155), .B2(n4787), .A(n4154), .ZN(n4938) );
  OAI21_X1 U4621 ( .B1(n4935), .B2(n4887), .A(n4938), .ZN(n4234) );
  MUX2_X1 U4622 ( .A(n4234), .B(REG1_REG_30__SCAN_IN), .S(n4892), .Z(U3548) );
  NAND2_X1 U4623 ( .A1(n4158), .A2(n4879), .ZN(n4159) );
  NAND2_X1 U4624 ( .A1(n4160), .A2(n4159), .ZN(n4235) );
  MUX2_X1 U4625 ( .A(REG1_REG_29__SCAN_IN), .B(n4235), .S(n4894), .Z(U3547) );
  OAI211_X1 U4626 ( .C1(n4163), .C2(n4888), .A(n4162), .B(n4161), .ZN(n4236)
         );
  MUX2_X1 U4627 ( .A(REG1_REG_28__SCAN_IN), .B(n4236), .S(n4894), .Z(U3546) );
  AOI21_X1 U4628 ( .B1(n4883), .B2(n4165), .A(n4164), .ZN(n4166) );
  OAI21_X1 U4629 ( .B1(n4167), .B2(n4888), .A(n4166), .ZN(n4237) );
  MUX2_X1 U4630 ( .A(REG1_REG_27__SCAN_IN), .B(n4237), .S(n4894), .Z(U3545) );
  NAND3_X1 U4631 ( .A1(n4169), .A2(n4883), .A3(n4168), .ZN(n4170) );
  OAI211_X1 U4632 ( .C1(n4172), .C2(n4888), .A(n4171), .B(n4170), .ZN(n4238)
         );
  MUX2_X1 U4633 ( .A(REG1_REG_26__SCAN_IN), .B(n4238), .S(n4894), .Z(U3544) );
  OAI21_X1 U4634 ( .B1(n4887), .B2(n4174), .A(n4173), .ZN(n4175) );
  AOI21_X1 U4635 ( .B1(n4176), .B2(n4879), .A(n4175), .ZN(n4239) );
  NAND2_X1 U4636 ( .A1(n4892), .A2(REG1_REG_25__SCAN_IN), .ZN(n4177) );
  OAI21_X1 U4637 ( .B1(n4239), .B2(n4892), .A(n4177), .ZN(U3543) );
  NAND3_X1 U4638 ( .A1(n4178), .A2(n4883), .A3(n3943), .ZN(n4179) );
  OAI211_X1 U4639 ( .C1(n4181), .C2(n4888), .A(n4180), .B(n4179), .ZN(n4450)
         );
  MUX2_X1 U4640 ( .A(REG1_REG_24__SCAN_IN), .B(n4450), .S(n4894), .Z(U3542) );
  AOI21_X1 U4641 ( .B1(n4883), .B2(n4183), .A(n4182), .ZN(n4184) );
  OAI21_X1 U4642 ( .B1(n4185), .B2(n4888), .A(n4184), .ZN(n4451) );
  MUX2_X1 U4643 ( .A(REG1_REG_23__SCAN_IN), .B(n4451), .S(n4894), .Z(U3541) );
  NAND3_X1 U4644 ( .A1(n2291), .A2(n4883), .A3(n4186), .ZN(n4187) );
  OAI211_X1 U4645 ( .C1(n4189), .C2(n4888), .A(n4188), .B(n4187), .ZN(n4452)
         );
  MUX2_X1 U4646 ( .A(REG1_REG_22__SCAN_IN), .B(n4452), .S(n4894), .Z(U3540) );
  AOI21_X1 U4647 ( .B1(n4883), .B2(n4191), .A(n4190), .ZN(n4192) );
  OAI21_X1 U4648 ( .B1(n4193), .B2(n4888), .A(n4192), .ZN(n4453) );
  MUX2_X1 U4649 ( .A(REG1_REG_21__SCAN_IN), .B(n4453), .S(n4894), .Z(U3539) );
  OAI211_X1 U4650 ( .C1(n4196), .C2(n4696), .A(n4195), .B(n4194), .ZN(n4454)
         );
  MUX2_X1 U4651 ( .A(REG1_REG_20__SCAN_IN), .B(n4454), .S(n4894), .Z(U3538) );
  OAI22_X1 U4652 ( .A1(n4198), .A2(n4888), .B1(n4887), .B2(n4197), .ZN(n4199)
         );
  OR2_X1 U4653 ( .A1(n4200), .A2(n4199), .ZN(n4455) );
  MUX2_X1 U4654 ( .A(REG1_REG_19__SCAN_IN), .B(n4455), .S(n4894), .Z(U3537) );
  AOI21_X1 U4655 ( .B1(n4202), .B2(n4879), .A(n4201), .ZN(n4203) );
  AND2_X1 U4656 ( .A1(n4204), .A2(n4203), .ZN(n4456) );
  MUX2_X1 U4657 ( .A(n4205), .B(n4456), .S(n4894), .Z(n4206) );
  INV_X1 U4658 ( .A(n4206), .ZN(U3536) );
  NAND2_X1 U4659 ( .A1(n4207), .A2(n4883), .ZN(n4208) );
  OAI211_X1 U4660 ( .C1(n4210), .C2(n4888), .A(n4209), .B(n4208), .ZN(n4459)
         );
  MUX2_X1 U4661 ( .A(REG1_REG_14__SCAN_IN), .B(n4459), .S(n4894), .Z(U3532) );
  OAI21_X1 U4662 ( .B1(n4796), .B2(n4212), .A(n4211), .ZN(n4813) );
  OAI22_X1 U4663 ( .A1(n4227), .A2(n4213), .B1(n4212), .B2(n4853), .ZN(n4216)
         );
  XNOR2_X1 U4664 ( .A(n3575), .B(n4219), .ZN(n4214) );
  NOR2_X1 U4665 ( .A1(n4214), .A2(n4856), .ZN(n4215) );
  AOI211_X1 U4666 ( .C1(n4862), .C2(n4217), .A(n4216), .B(n4215), .ZN(n4818)
         );
  XOR2_X1 U4667 ( .A(n4219), .B(n4218), .Z(n4815) );
  NAND2_X1 U4668 ( .A1(n4815), .A2(n4879), .ZN(n4220) );
  OAI211_X1 U4669 ( .C1(n4887), .C2(n4813), .A(n4818), .B(n4220), .ZN(n4460)
         );
  MUX2_X1 U4670 ( .A(REG1_REG_12__SCAN_IN), .B(n4460), .S(n4894), .Z(U3530) );
  XOR2_X1 U4671 ( .A(n4223), .B(n4221), .Z(n4778) );
  AOI21_X1 U4672 ( .B1(n4224), .B2(n4763), .A(n4795), .ZN(n4777) );
  AOI22_X1 U4673 ( .A1(n4778), .A2(n4879), .B1(n4883), .B2(n4777), .ZN(n4230)
         );
  XOR2_X1 U4674 ( .A(n4223), .B(n4222), .Z(n4229) );
  AOI22_X1 U4675 ( .A1(n4225), .A2(n4849), .B1(n4224), .B2(n4787), .ZN(n4226)
         );
  OAI21_X1 U4676 ( .B1(n4227), .B2(n4737), .A(n4226), .ZN(n4228) );
  AOI21_X1 U4677 ( .B1(n4229), .B2(n4731), .A(n4228), .ZN(n4781) );
  NAND2_X1 U4678 ( .A1(n4230), .A2(n4781), .ZN(n4461) );
  MUX2_X1 U4679 ( .A(REG1_REG_10__SCAN_IN), .B(n4461), .S(n4894), .Z(U3528) );
  INV_X1 U4680 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4232) );
  MUX2_X1 U4681 ( .A(n4232), .B(n4231), .S(n4897), .Z(n4233) );
  INV_X1 U4682 ( .A(n4233), .ZN(U3517) );
  MUX2_X1 U4683 ( .A(n4234), .B(REG0_REG_30__SCAN_IN), .S(n4895), .Z(U3516) );
  MUX2_X1 U4684 ( .A(REG0_REG_29__SCAN_IN), .B(n4235), .S(n4897), .Z(U3515) );
  MUX2_X1 U4685 ( .A(REG0_REG_28__SCAN_IN), .B(n4236), .S(n4897), .Z(U3514) );
  MUX2_X1 U4686 ( .A(REG0_REG_27__SCAN_IN), .B(n4237), .S(n4897), .Z(U3513) );
  MUX2_X1 U4687 ( .A(REG0_REG_26__SCAN_IN), .B(n4238), .S(n4897), .Z(U3512) );
  MUX2_X1 U4688 ( .A(n4240), .B(n4239), .S(n4897), .Z(n4449) );
  INV_X1 U4689 ( .A(keyinput_123), .ZN(n4328) );
  AOI22_X1 U4690 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_116), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput_117), .ZN(n4241) );
  OAI221_X1 U4691 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_116), .C1(
        REG3_REG_20__SCAN_IN), .C2(keyinput_117), .A(n4241), .ZN(n4319) );
  OAI22_X1 U4692 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_114), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput_115), .ZN(n4242) );
  AOI221_X1 U4693 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_114), .C1(
        keyinput_115), .C2(REG3_REG_9__SCAN_IN), .A(n4242), .ZN(n4315) );
  OAI22_X1 U4694 ( .A1(n4339), .A2(keyinput_112), .B1(keyinput_111), .B2(
        REG3_REG_5__SCAN_IN), .ZN(n4243) );
  AOI221_X1 U4695 ( .B1(n4339), .B2(keyinput_112), .C1(REG3_REG_5__SCAN_IN), 
        .C2(keyinput_111), .A(n4243), .ZN(n4312) );
  INV_X1 U4696 ( .A(keyinput_104), .ZN(n4302) );
  INV_X1 U4697 ( .A(keyinput_103), .ZN(n4300) );
  INV_X1 U4698 ( .A(keyinput_102), .ZN(n4298) );
  OAI22_X1 U4699 ( .A1(n2916), .A2(keyinput_97), .B1(n4245), .B2(keyinput_98), 
        .ZN(n4244) );
  AOI221_X1 U4700 ( .B1(n2916), .B2(keyinput_97), .C1(keyinput_98), .C2(n4245), 
        .A(n4244), .ZN(n4296) );
  INV_X1 U4701 ( .A(keyinput_96), .ZN(n4291) );
  INV_X1 U4702 ( .A(keyinput_95), .ZN(n4289) );
  INV_X1 U4703 ( .A(DATAI_0_), .ZN(n4626) );
  AOI22_X1 U4704 ( .A1(DATAI_2_), .A2(keyinput_93), .B1(DATAI_3_), .B2(
        keyinput_92), .ZN(n4246) );
  OAI221_X1 U4705 ( .B1(DATAI_2_), .B2(keyinput_93), .C1(DATAI_3_), .C2(
        keyinput_92), .A(n4246), .ZN(n4287) );
  INV_X1 U4706 ( .A(keyinput_80), .ZN(n4271) );
  INV_X1 U4707 ( .A(DATAI_15_), .ZN(n4372) );
  INV_X1 U4708 ( .A(DATAI_19_), .ZN(n4248) );
  OAI22_X1 U4709 ( .A1(n4249), .A2(keyinput_75), .B1(n4248), .B2(keyinput_76), 
        .ZN(n4247) );
  AOI221_X1 U4710 ( .B1(n4249), .B2(keyinput_75), .C1(keyinput_76), .C2(n4248), 
        .A(n4247), .ZN(n4269) );
  INV_X1 U4711 ( .A(keyinput_74), .ZN(n4263) );
  INV_X1 U4712 ( .A(DATAI_23_), .ZN(n4470) );
  OAI22_X1 U4713 ( .A1(n4470), .A2(keyinput_72), .B1(DATAI_24_), .B2(
        keyinput_71), .ZN(n4250) );
  AOI221_X1 U4714 ( .B1(n4470), .B2(keyinput_72), .C1(keyinput_71), .C2(
        DATAI_24_), .A(n4250), .ZN(n4259) );
  AOI22_X1 U4715 ( .A1(DATAI_31_), .A2(keyinput_64), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n4251) );
  OAI221_X1 U4716 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(DATAI_30_), .C2(
        keyinput_65), .A(n4251), .ZN(n4254) );
  AOI22_X1 U4717 ( .A1(DATAI_28_), .A2(keyinput_67), .B1(DATAI_29_), .B2(
        keyinput_66), .ZN(n4252) );
  OAI221_X1 U4718 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(DATAI_29_), .C2(
        keyinput_66), .A(n4252), .ZN(n4253) );
  OAI22_X1 U4719 ( .A1(DATAI_27_), .A2(keyinput_68), .B1(n4254), .B2(n4253), 
        .ZN(n4257) );
  OAI22_X1 U4720 ( .A1(DATAI_26_), .A2(keyinput_69), .B1(DATAI_25_), .B2(
        keyinput_70), .ZN(n4255) );
  AOI221_X1 U4721 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(keyinput_70), .C2(
        DATAI_25_), .A(n4255), .ZN(n4256) );
  OAI221_X1 U4722 ( .B1(n4257), .B2(keyinput_68), .C1(n4257), .C2(DATAI_27_), 
        .A(n4256), .ZN(n4258) );
  AOI22_X1 U4723 ( .A1(keyinput_73), .A2(n4261), .B1(n4259), .B2(n4258), .ZN(
        n4260) );
  OAI21_X1 U4724 ( .B1(n4261), .B2(keyinput_73), .A(n4260), .ZN(n4262) );
  OAI221_X1 U4725 ( .B1(DATAI_21_), .B2(n4263), .C1(n4363), .C2(keyinput_74), 
        .A(n4262), .ZN(n4268) );
  XOR2_X1 U4726 ( .A(DATAI_17_), .B(keyinput_78), .Z(n4267) );
  AOI22_X1 U4727 ( .A1(DATAI_16_), .A2(keyinput_79), .B1(n4265), .B2(
        keyinput_77), .ZN(n4264) );
  OAI221_X1 U4728 ( .B1(DATAI_16_), .B2(keyinput_79), .C1(n4265), .C2(
        keyinput_77), .A(n4264), .ZN(n4266) );
  AOI211_X1 U4729 ( .C1(n4269), .C2(n4268), .A(n4267), .B(n4266), .ZN(n4270)
         );
  AOI221_X1 U4730 ( .B1(DATAI_15_), .B2(n4271), .C1(n4372), .C2(keyinput_80), 
        .A(n4270), .ZN(n4277) );
  XNOR2_X1 U4731 ( .A(DATAI_11_), .B(keyinput_84), .ZN(n4276) );
  INV_X1 U4732 ( .A(DATAI_14_), .ZN(n4375) );
  AOI22_X1 U4733 ( .A1(DATAI_13_), .A2(keyinput_82), .B1(n4375), .B2(
        keyinput_81), .ZN(n4272) );
  OAI221_X1 U4734 ( .B1(DATAI_13_), .B2(keyinput_82), .C1(n4375), .C2(
        keyinput_81), .A(n4272), .ZN(n4275) );
  INV_X1 U4735 ( .A(DATAI_12_), .ZN(n4810) );
  AOI22_X1 U4736 ( .A1(DATAI_10_), .A2(keyinput_85), .B1(n4810), .B2(
        keyinput_83), .ZN(n4273) );
  OAI221_X1 U4737 ( .B1(DATAI_10_), .B2(keyinput_85), .C1(n4810), .C2(
        keyinput_83), .A(n4273), .ZN(n4274) );
  NOR4_X1 U4738 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4284)
         );
  AOI22_X1 U4739 ( .A1(DATAI_7_), .A2(keyinput_88), .B1(DATAI_9_), .B2(
        keyinput_86), .ZN(n4278) );
  OAI221_X1 U4740 ( .B1(DATAI_7_), .B2(keyinput_88), .C1(DATAI_9_), .C2(
        keyinput_86), .A(n4278), .ZN(n4283) );
  INV_X1 U4741 ( .A(DATAI_4_), .ZN(n4702) );
  AOI22_X1 U4742 ( .A1(DATAI_6_), .A2(keyinput_89), .B1(n4702), .B2(
        keyinput_91), .ZN(n4279) );
  OAI221_X1 U4743 ( .B1(DATAI_6_), .B2(keyinput_89), .C1(n4702), .C2(
        keyinput_91), .A(n4279), .ZN(n4282) );
  INV_X1 U4744 ( .A(DATAI_5_), .ZN(n4710) );
  INV_X1 U4745 ( .A(DATAI_8_), .ZN(n4750) );
  AOI22_X1 U4746 ( .A1(n4710), .A2(keyinput_90), .B1(n4750), .B2(keyinput_87), 
        .ZN(n4280) );
  OAI221_X1 U4747 ( .B1(n4710), .B2(keyinput_90), .C1(n4750), .C2(keyinput_87), 
        .A(n4280), .ZN(n4281) );
  NOR4_X1 U4748 ( .A1(n4284), .A2(n4283), .A3(n4282), .A4(n4281), .ZN(n4286)
         );
  INV_X1 U4749 ( .A(DATAI_1_), .ZN(n4388) );
  NAND2_X1 U4750 ( .A1(n4388), .A2(keyinput_94), .ZN(n4285) );
  OAI221_X1 U4751 ( .B1(n4287), .B2(n4286), .C1(n4388), .C2(keyinput_94), .A(
        n4285), .ZN(n4288) );
  OAI221_X1 U4752 ( .B1(DATAI_0_), .B2(n4289), .C1(n4626), .C2(keyinput_95), 
        .A(n4288), .ZN(n4290) );
  OAI221_X1 U4753 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_96), .C1(U3149), .C2(
        n4291), .A(n4290), .ZN(n4295) );
  XOR2_X1 U4754 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_101), .Z(n4294) );
  AOI22_X1 U4755 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_100), .B1(
        REG3_REG_14__SCAN_IN), .B2(keyinput_99), .ZN(n4292) );
  OAI221_X1 U4756 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_100), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_99), .A(n4292), .ZN(n4293) );
  AOI211_X1 U4757 ( .C1(n4296), .C2(n4295), .A(n4294), .B(n4293), .ZN(n4297)
         );
  AOI221_X1 U4758 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_102), .C1(n4401), 
        .C2(n4298), .A(n4297), .ZN(n4299) );
  AOI221_X1 U4759 ( .B1(REG3_REG_19__SCAN_IN), .B2(n4300), .C1(n4405), .C2(
        keyinput_103), .A(n4299), .ZN(n4301) );
  AOI221_X1 U4760 ( .B1(REG3_REG_28__SCAN_IN), .B2(n4302), .C1(n4408), .C2(
        keyinput_104), .A(n4301), .ZN(n4310) );
  AOI22_X1 U4761 ( .A1(n4304), .A2(keyinput_105), .B1(keyinput_106), .B2(n2817), .ZN(n4303) );
  OAI221_X1 U4762 ( .B1(n4304), .B2(keyinput_105), .C1(n2817), .C2(
        keyinput_106), .A(n4303), .ZN(n4309) );
  OAI22_X1 U4763 ( .A1(n4410), .A2(keyinput_108), .B1(n4911), .B2(keyinput_107), .ZN(n4305) );
  AOI221_X1 U4764 ( .B1(n4410), .B2(keyinput_108), .C1(keyinput_107), .C2(
        n4911), .A(n4305), .ZN(n4308) );
  OAI22_X1 U4765 ( .A1(n4413), .A2(keyinput_110), .B1(n4412), .B2(keyinput_109), .ZN(n4306) );
  AOI221_X1 U4766 ( .B1(n4413), .B2(keyinput_110), .C1(keyinput_109), .C2(
        n4412), .A(n4306), .ZN(n4307) );
  OAI211_X1 U4767 ( .C1(n4310), .C2(n4309), .A(n4308), .B(n4307), .ZN(n4311)
         );
  AOI22_X1 U4768 ( .A1(n4312), .A2(n4311), .B1(keyinput_113), .B2(
        REG3_REG_24__SCAN_IN), .ZN(n4313) );
  OAI21_X1 U4769 ( .B1(keyinput_113), .B2(REG3_REG_24__SCAN_IN), .A(n4313), 
        .ZN(n4314) );
  AOI22_X1 U4770 ( .A1(n4315), .A2(n4314), .B1(keyinput_118), .B2(n4317), .ZN(
        n4316) );
  OAI21_X1 U4771 ( .B1(keyinput_118), .B2(n4317), .A(n4316), .ZN(n4318) );
  OAI22_X1 U4772 ( .A1(n4319), .A2(n4318), .B1(keyinput_119), .B2(n2614), .ZN(
        n4320) );
  AOI21_X1 U4773 ( .B1(keyinput_119), .B2(n2614), .A(n4320), .ZN(n4325) );
  INV_X1 U4774 ( .A(IR_REG_1__SCAN_IN), .ZN(n4321) );
  XOR2_X1 U4775 ( .A(n4321), .B(keyinput_120), .Z(n4323) );
  XNOR2_X1 U4776 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4322) );
  NAND2_X1 U4777 ( .A1(n4323), .A2(n4322), .ZN(n4324) );
  OAI22_X1 U4778 ( .A1(n4325), .A2(n4324), .B1(IR_REG_3__SCAN_IN), .B2(
        keyinput_122), .ZN(n4326) );
  AOI21_X1 U4779 ( .B1(keyinput_122), .B2(IR_REG_3__SCAN_IN), .A(n4326), .ZN(
        n4327) );
  AOI221_X1 U4780 ( .B1(IR_REG_4__SCAN_IN), .B2(n4328), .C1(n2514), .C2(
        keyinput_123), .A(n4327), .ZN(n4335) );
  INV_X1 U4781 ( .A(keyinput_124), .ZN(n4329) );
  MUX2_X1 U4782 ( .A(keyinput_124), .B(n4329), .S(IR_REG_5__SCAN_IN), .Z(n4334) );
  INV_X1 U4783 ( .A(IR_REG_6__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4784 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_126), .B1(n4331), .B2(
        keyinput_125), .ZN(n4330) );
  OAI221_X1 U4785 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_126), .C1(n4331), 
        .C2(keyinput_125), .A(n4330), .ZN(n4332) );
  INV_X1 U4786 ( .A(n4332), .ZN(n4333) );
  OAI21_X1 U4787 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n4447) );
  INV_X1 U4788 ( .A(IR_REG_8__SCAN_IN), .ZN(n4336) );
  MUX2_X1 U4789 ( .A(n4336), .B(keyinput_63), .S(keyinput_127), .Z(n4446) );
  INV_X1 U4790 ( .A(keyinput_59), .ZN(n4438) );
  INV_X1 U4791 ( .A(keyinput_55), .ZN(n4430) );
  AOI22_X1 U4792 ( .A1(n4339), .A2(keyinput_48), .B1(n4338), .B2(keyinput_47), 
        .ZN(n4337) );
  OAI221_X1 U4793 ( .B1(n4339), .B2(keyinput_48), .C1(n4338), .C2(keyinput_47), 
        .A(n4337), .ZN(n4419) );
  OAI22_X1 U4794 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_41), .B1(keyinput_42), .B2(REG3_REG_1__SCAN_IN), .ZN(n4340) );
  AOI221_X1 U4795 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_41), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput_42), .A(n4340), .ZN(n4417) );
  INV_X1 U4796 ( .A(keyinput_40), .ZN(n4407) );
  INV_X1 U4797 ( .A(keyinput_39), .ZN(n4404) );
  INV_X1 U4798 ( .A(keyinput_38), .ZN(n4402) );
  AOI22_X1 U4799 ( .A1(n4343), .A2(keyinput_36), .B1(n4342), .B2(keyinput_37), 
        .ZN(n4341) );
  OAI221_X1 U4800 ( .B1(n4343), .B2(keyinput_36), .C1(n4342), .C2(keyinput_37), 
        .A(n4341), .ZN(n4400) );
  OAI22_X1 U4801 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_33), .B1(keyinput_34), .B2(REG3_REG_27__SCAN_IN), .ZN(n4344) );
  AOI221_X1 U4802 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_33), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_34), .A(n4344), .ZN(n4396) );
  INV_X1 U4803 ( .A(keyinput_32), .ZN(n4394) );
  INV_X1 U4804 ( .A(keyinput_31), .ZN(n4392) );
  AOI22_X1 U4805 ( .A1(DATAI_2_), .A2(keyinput_29), .B1(DATAI_3_), .B2(
        keyinput_28), .ZN(n4345) );
  OAI221_X1 U4806 ( .B1(DATAI_2_), .B2(keyinput_29), .C1(DATAI_3_), .C2(
        keyinput_28), .A(n4345), .ZN(n4390) );
  INV_X1 U4807 ( .A(DATAI_10_), .ZN(n4346) );
  XNOR2_X1 U4808 ( .A(keyinput_21), .B(n4346), .ZN(n4379) );
  INV_X1 U4809 ( .A(keyinput_16), .ZN(n4371) );
  OAI22_X1 U4810 ( .A1(DATAI_20_), .A2(keyinput_11), .B1(keyinput_12), .B2(
        DATAI_19_), .ZN(n4347) );
  AOI221_X1 U4811 ( .B1(DATAI_20_), .B2(keyinput_11), .C1(DATAI_19_), .C2(
        keyinput_12), .A(n4347), .ZN(n4369) );
  INV_X1 U4812 ( .A(keyinput_10), .ZN(n4364) );
  OAI22_X1 U4813 ( .A1(n4470), .A2(keyinput_8), .B1(keyinput_7), .B2(DATAI_24_), .ZN(n4348) );
  AOI221_X1 U4814 ( .B1(n4470), .B2(keyinput_8), .C1(DATAI_24_), .C2(
        keyinput_7), .A(n4348), .ZN(n4360) );
  INV_X1 U4815 ( .A(DATAI_28_), .ZN(n4931) );
  AOI22_X1 U4816 ( .A1(n4350), .A2(keyinput_2), .B1(keyinput_3), .B2(n4931), 
        .ZN(n4349) );
  OAI221_X1 U4817 ( .B1(n4350), .B2(keyinput_2), .C1(n4931), .C2(keyinput_3), 
        .A(n4349), .ZN(n4353) );
  AOI22_X1 U4818 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n4351) );
  OAI221_X1 U4819 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n4351), .ZN(n4352) );
  OAI22_X1 U4820 ( .A1(keyinput_4), .A2(n4357), .B1(n4353), .B2(n4352), .ZN(
        n4358) );
  INV_X1 U4821 ( .A(DATAI_26_), .ZN(n4355) );
  OAI22_X1 U4822 ( .A1(n4355), .A2(keyinput_5), .B1(keyinput_6), .B2(DATAI_25_), .ZN(n4354) );
  AOI221_X1 U4823 ( .B1(n4355), .B2(keyinput_5), .C1(DATAI_25_), .C2(
        keyinput_6), .A(n4354), .ZN(n4356) );
  OAI221_X1 U4824 ( .B1(n4358), .B2(keyinput_4), .C1(n4358), .C2(n4357), .A(
        n4356), .ZN(n4359) );
  AOI22_X1 U4825 ( .A1(n4360), .A2(n4359), .B1(keyinput_9), .B2(DATAI_22_), 
        .ZN(n4361) );
  OAI21_X1 U4826 ( .B1(keyinput_9), .B2(DATAI_22_), .A(n4361), .ZN(n4362) );
  OAI221_X1 U4827 ( .B1(DATAI_21_), .B2(n4364), .C1(n4363), .C2(keyinput_10), 
        .A(n4362), .ZN(n4368) );
  XOR2_X1 U4828 ( .A(DATAI_18_), .B(keyinput_13), .Z(n4367) );
  INV_X1 U4829 ( .A(DATAI_16_), .ZN(n4876) );
  AOI22_X1 U4830 ( .A1(DATAI_17_), .A2(keyinput_14), .B1(n4876), .B2(
        keyinput_15), .ZN(n4365) );
  OAI221_X1 U4831 ( .B1(DATAI_17_), .B2(keyinput_14), .C1(n4876), .C2(
        keyinput_15), .A(n4365), .ZN(n4366) );
  AOI211_X1 U4832 ( .C1(n4369), .C2(n4368), .A(n4367), .B(n4366), .ZN(n4370)
         );
  AOI221_X1 U4833 ( .B1(DATAI_15_), .B2(keyinput_16), .C1(n4372), .C2(n4371), 
        .A(n4370), .ZN(n4378) );
  INV_X1 U4834 ( .A(DATAI_11_), .ZN(n4782) );
  AOI22_X1 U4835 ( .A1(n4782), .A2(keyinput_20), .B1(n4810), .B2(keyinput_19), 
        .ZN(n4373) );
  OAI221_X1 U4836 ( .B1(n4782), .B2(keyinput_20), .C1(n4810), .C2(keyinput_19), 
        .A(n4373), .ZN(n4377) );
  INV_X1 U4837 ( .A(DATAI_13_), .ZN(n4819) );
  AOI22_X1 U4838 ( .A1(n4819), .A2(keyinput_18), .B1(n4375), .B2(keyinput_17), 
        .ZN(n4374) );
  OAI221_X1 U4839 ( .B1(n4819), .B2(keyinput_18), .C1(n4375), .C2(keyinput_17), 
        .A(n4374), .ZN(n4376) );
  NOR4_X1 U4840 ( .A1(n4379), .A2(n4378), .A3(n4377), .A4(n4376), .ZN(n4386)
         );
  INV_X1 U4841 ( .A(DATAI_7_), .ZN(n4719) );
  AOI22_X1 U4842 ( .A1(DATAI_5_), .A2(keyinput_26), .B1(n4719), .B2(
        keyinput_24), .ZN(n4380) );
  OAI221_X1 U4843 ( .B1(DATAI_5_), .B2(keyinput_26), .C1(n4719), .C2(
        keyinput_24), .A(n4380), .ZN(n4385) );
  INV_X1 U4844 ( .A(DATAI_6_), .ZN(n4717) );
  AOI22_X1 U4845 ( .A1(DATAI_9_), .A2(keyinput_22), .B1(n4717), .B2(
        keyinput_25), .ZN(n4381) );
  OAI221_X1 U4846 ( .B1(DATAI_9_), .B2(keyinput_22), .C1(n4717), .C2(
        keyinput_25), .A(n4381), .ZN(n4384) );
  AOI22_X1 U4847 ( .A1(n4750), .A2(keyinput_23), .B1(keyinput_27), .B2(n4702), 
        .ZN(n4382) );
  OAI221_X1 U4848 ( .B1(n4750), .B2(keyinput_23), .C1(n4702), .C2(keyinput_27), 
        .A(n4382), .ZN(n4383) );
  NOR4_X1 U4849 ( .A1(n4386), .A2(n4385), .A3(n4384), .A4(n4383), .ZN(n4389)
         );
  NAND2_X1 U4850 ( .A1(n4388), .A2(keyinput_30), .ZN(n4387) );
  OAI221_X1 U4851 ( .B1(n4390), .B2(n4389), .C1(n4388), .C2(keyinput_30), .A(
        n4387), .ZN(n4391) );
  OAI221_X1 U4852 ( .B1(DATAI_0_), .B2(keyinput_31), .C1(n4626), .C2(n4392), 
        .A(n4391), .ZN(n4393) );
  OAI221_X1 U4853 ( .B1(STATE_REG_SCAN_IN), .B2(n4394), .C1(U3149), .C2(
        keyinput_32), .A(n4393), .ZN(n4395) );
  AOI22_X1 U4854 ( .A1(n4396), .A2(n4395), .B1(keyinput_35), .B2(n4398), .ZN(
        n4397) );
  OAI21_X1 U4855 ( .B1(keyinput_35), .B2(n4398), .A(n4397), .ZN(n4399) );
  OAI222_X1 U4856 ( .A1(REG3_REG_3__SCAN_IN), .A2(n4402), .B1(n4401), .B2(
        keyinput_38), .C1(n4400), .C2(n4399), .ZN(n4403) );
  OAI221_X1 U4857 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_39), .C1(n4405), 
        .C2(n4404), .A(n4403), .ZN(n4406) );
  OAI221_X1 U4858 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_40), .C1(n4408), 
        .C2(n4407), .A(n4406), .ZN(n4416) );
  AOI22_X1 U4859 ( .A1(n4410), .A2(keyinput_44), .B1(keyinput_43), .B2(n4911), 
        .ZN(n4409) );
  OAI221_X1 U4860 ( .B1(n4410), .B2(keyinput_44), .C1(n4911), .C2(keyinput_43), 
        .A(n4409), .ZN(n4415) );
  AOI22_X1 U4861 ( .A1(n4413), .A2(keyinput_46), .B1(keyinput_45), .B2(n4412), 
        .ZN(n4411) );
  OAI221_X1 U4862 ( .B1(n4413), .B2(keyinput_46), .C1(n4412), .C2(keyinput_45), 
        .A(n4411), .ZN(n4414) );
  AOI211_X1 U4863 ( .C1(n4417), .C2(n4416), .A(n4415), .B(n4414), .ZN(n4418)
         );
  OAI22_X1 U4864 ( .A1(keyinput_49), .A2(n4421), .B1(n4419), .B2(n4418), .ZN(
        n4420) );
  AOI21_X1 U4865 ( .B1(keyinput_49), .B2(n4421), .A(n4420), .ZN(n4428) );
  AOI22_X1 U4866 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_51), .B1(n4423), 
        .B2(keyinput_50), .ZN(n4422) );
  OAI221_X1 U4867 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_51), .C1(n4423), 
        .C2(keyinput_50), .A(n4422), .ZN(n4427) );
  OAI22_X1 U4868 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_54), .B1(
        keyinput_52), .B2(REG3_REG_0__SCAN_IN), .ZN(n4424) );
  AOI221_X1 U4869 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_54), .C1(
        REG3_REG_0__SCAN_IN), .C2(keyinput_52), .A(n4424), .ZN(n4426) );
  XNOR2_X1 U4870 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .ZN(n4425) );
  OAI211_X1 U4871 ( .C1(n4428), .C2(n4427), .A(n4426), .B(n4425), .ZN(n4429)
         );
  OAI221_X1 U4872 ( .B1(n2614), .B2(keyinput_55), .C1(n2634), .C2(n4430), .A(
        n4429), .ZN(n4435) );
  XNOR2_X1 U4873 ( .A(n4431), .B(keyinput_57), .ZN(n4433) );
  XNOR2_X1 U4874 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .ZN(n4432) );
  NOR2_X1 U4875 ( .A1(n4433), .A2(n4432), .ZN(n4434) );
  AOI22_X1 U4876 ( .A1(n4435), .A2(n4434), .B1(IR_REG_3__SCAN_IN), .B2(
        keyinput_58), .ZN(n4436) );
  OAI21_X1 U4877 ( .B1(keyinput_58), .B2(IR_REG_3__SCAN_IN), .A(n4436), .ZN(
        n4437) );
  OAI221_X1 U4878 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_59), .C1(n2514), .C2(
        n4438), .A(n4437), .ZN(n4443) );
  XNOR2_X1 U4879 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4442) );
  XNOR2_X1 U4880 ( .A(n4439), .B(keyinput_62), .ZN(n4441) );
  XNOR2_X1 U4881 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n4440) );
  AOI211_X1 U4882 ( .C1(n4443), .C2(n4442), .A(n4441), .B(n4440), .ZN(n4445)
         );
  XOR2_X1 U4883 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .Z(n4444) );
  AOI211_X1 U4884 ( .C1(n4447), .C2(n4446), .A(n4445), .B(n4444), .ZN(n4448)
         );
  XNOR2_X1 U4885 ( .A(n4449), .B(n4448), .ZN(U3511) );
  MUX2_X1 U4886 ( .A(REG0_REG_24__SCAN_IN), .B(n4450), .S(n4897), .Z(U3510) );
  MUX2_X1 U4887 ( .A(REG0_REG_23__SCAN_IN), .B(n4451), .S(n4897), .Z(U3509) );
  MUX2_X1 U4888 ( .A(REG0_REG_22__SCAN_IN), .B(n4452), .S(n4897), .Z(U3508) );
  MUX2_X1 U4889 ( .A(REG0_REG_21__SCAN_IN), .B(n4453), .S(n4897), .Z(U3507) );
  MUX2_X1 U4890 ( .A(REG0_REG_20__SCAN_IN), .B(n4454), .S(n4897), .Z(U3506) );
  MUX2_X1 U4891 ( .A(REG0_REG_19__SCAN_IN), .B(n4455), .S(n4897), .Z(U3505) );
  MUX2_X1 U4892 ( .A(n4457), .B(n4456), .S(n4897), .Z(n4458) );
  INV_X1 U4893 ( .A(n4458), .ZN(U3503) );
  MUX2_X1 U4894 ( .A(REG0_REG_14__SCAN_IN), .B(n4459), .S(n4897), .Z(U3495) );
  MUX2_X1 U4895 ( .A(REG0_REG_12__SCAN_IN), .B(n4460), .S(n4897), .Z(U3491) );
  MUX2_X1 U4896 ( .A(REG0_REG_10__SCAN_IN), .B(n4461), .S(n4897), .Z(U3487) );
  MUX2_X1 U4897 ( .A(D_REG_1__SCAN_IN), .B(n4462), .S(n4501), .Z(U3459) );
  MUX2_X1 U4898 ( .A(n4463), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4899 ( .A(n4464), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4900 ( .A(DATAI_19_), .B(n3809), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4901 ( .A(n4465), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U4902 ( .A(n4466), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U4903 ( .A(n4467), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U4904 ( .A(n4468), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI21_X1 U4905 ( .B1(STATE_REG_SCAN_IN), .B2(n4470), .A(n4469), .ZN(U3329)
         );
  INV_X1 U4906 ( .A(D_REG_2__SCAN_IN), .ZN(n4471) );
  NOR2_X1 U4907 ( .A1(n4501), .A2(n4471), .ZN(U3320) );
  INV_X1 U4908 ( .A(D_REG_3__SCAN_IN), .ZN(n4472) );
  NOR2_X1 U4909 ( .A1(n4501), .A2(n4472), .ZN(U3319) );
  INV_X1 U4910 ( .A(D_REG_4__SCAN_IN), .ZN(n4473) );
  NOR2_X1 U4911 ( .A1(n4501), .A2(n4473), .ZN(U3318) );
  INV_X1 U4912 ( .A(D_REG_5__SCAN_IN), .ZN(n4474) );
  NOR2_X1 U4913 ( .A1(n4501), .A2(n4474), .ZN(U3317) );
  INV_X1 U4914 ( .A(D_REG_6__SCAN_IN), .ZN(n4475) );
  NOR2_X1 U4915 ( .A1(n4501), .A2(n4475), .ZN(U3316) );
  INV_X1 U4916 ( .A(D_REG_7__SCAN_IN), .ZN(n4476) );
  NOR2_X1 U4917 ( .A1(n4501), .A2(n4476), .ZN(U3315) );
  INV_X1 U4918 ( .A(D_REG_8__SCAN_IN), .ZN(n4477) );
  NOR2_X1 U4919 ( .A1(n4501), .A2(n4477), .ZN(U3314) );
  INV_X1 U4920 ( .A(D_REG_9__SCAN_IN), .ZN(n4478) );
  NOR2_X1 U4921 ( .A1(n4501), .A2(n4478), .ZN(U3313) );
  INV_X1 U4922 ( .A(D_REG_10__SCAN_IN), .ZN(n4479) );
  NOR2_X1 U4923 ( .A1(n4501), .A2(n4479), .ZN(U3312) );
  INV_X1 U4924 ( .A(D_REG_11__SCAN_IN), .ZN(n4480) );
  NOR2_X1 U4925 ( .A1(n4501), .A2(n4480), .ZN(U3311) );
  INV_X1 U4926 ( .A(D_REG_12__SCAN_IN), .ZN(n4481) );
  NOR2_X1 U4927 ( .A1(n4501), .A2(n4481), .ZN(U3310) );
  INV_X1 U4928 ( .A(D_REG_13__SCAN_IN), .ZN(n4482) );
  NOR2_X1 U4929 ( .A1(n4501), .A2(n4482), .ZN(U3309) );
  INV_X1 U4930 ( .A(D_REG_14__SCAN_IN), .ZN(n4483) );
  NOR2_X1 U4931 ( .A1(n4501), .A2(n4483), .ZN(U3308) );
  INV_X1 U4932 ( .A(D_REG_15__SCAN_IN), .ZN(n4484) );
  NOR2_X1 U4933 ( .A1(n4501), .A2(n4484), .ZN(U3307) );
  INV_X1 U4934 ( .A(D_REG_16__SCAN_IN), .ZN(n4485) );
  NOR2_X1 U4935 ( .A1(n4501), .A2(n4485), .ZN(U3306) );
  INV_X1 U4936 ( .A(D_REG_17__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U4937 ( .A1(n4501), .A2(n4486), .ZN(U3305) );
  INV_X1 U4938 ( .A(D_REG_18__SCAN_IN), .ZN(n4487) );
  NOR2_X1 U4939 ( .A1(n4501), .A2(n4487), .ZN(U3304) );
  INV_X1 U4940 ( .A(D_REG_19__SCAN_IN), .ZN(n4488) );
  NOR2_X1 U4941 ( .A1(n4501), .A2(n4488), .ZN(U3303) );
  INV_X1 U4942 ( .A(D_REG_20__SCAN_IN), .ZN(n4489) );
  NOR2_X1 U4943 ( .A1(n4501), .A2(n4489), .ZN(U3302) );
  INV_X1 U4944 ( .A(D_REG_21__SCAN_IN), .ZN(n4490) );
  NOR2_X1 U4945 ( .A1(n4501), .A2(n4490), .ZN(U3301) );
  INV_X1 U4946 ( .A(D_REG_22__SCAN_IN), .ZN(n4491) );
  NOR2_X1 U4947 ( .A1(n4501), .A2(n4491), .ZN(U3300) );
  INV_X1 U4948 ( .A(D_REG_23__SCAN_IN), .ZN(n4492) );
  NOR2_X1 U4949 ( .A1(n4501), .A2(n4492), .ZN(U3299) );
  INV_X1 U4950 ( .A(D_REG_24__SCAN_IN), .ZN(n4493) );
  NOR2_X1 U4951 ( .A1(n4501), .A2(n4493), .ZN(U3298) );
  INV_X1 U4952 ( .A(D_REG_25__SCAN_IN), .ZN(n4494) );
  NOR2_X1 U4953 ( .A1(n4501), .A2(n4494), .ZN(U3297) );
  INV_X1 U4954 ( .A(D_REG_26__SCAN_IN), .ZN(n4495) );
  NOR2_X1 U4955 ( .A1(n4501), .A2(n4495), .ZN(U3296) );
  INV_X1 U4956 ( .A(D_REG_27__SCAN_IN), .ZN(n4496) );
  NOR2_X1 U4957 ( .A1(n4501), .A2(n4496), .ZN(U3295) );
  NOR2_X1 U4958 ( .A1(n4501), .A2(n4497), .ZN(U3294) );
  NOR2_X1 U4959 ( .A1(n4501), .A2(n4498), .ZN(U3293) );
  NOR2_X1 U4960 ( .A1(n4501), .A2(n4499), .ZN(U3292) );
  NOR2_X1 U4961 ( .A1(n4501), .A2(n4500), .ZN(U3291) );
  OR2_X1 U4962 ( .A1(n4639), .A2(REG2_REG_0__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U4963 ( .A1(n4502), .A2(n4637), .ZN(n4504) );
  INV_X1 U4964 ( .A(n4504), .ZN(n4642) );
  OAI211_X1 U4965 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4503), .A(n4505), .B(n4642), 
        .ZN(n4508) );
  AOI22_X1 U4966 ( .A1(n4505), .A2(n4504), .B1(n4609), .B2(n2638), .ZN(n4507)
         );
  AOI22_X1 U4967 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4646), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4506) );
  OAI221_X1 U4968 ( .B1(n2614), .B2(n4508), .C1(n2634), .C2(n4507), .A(n4506), 
        .ZN(U3240) );
  AOI211_X1 U4969 ( .C1(n2722), .C2(n4510), .A(n4509), .B(n4650), .ZN(n4512)
         );
  AOI211_X1 U4970 ( .C1(n4646), .C2(ADDR_REG_3__SCAN_IN), .A(n4512), .B(n4511), 
        .ZN(n4517) );
  AOI21_X1 U4971 ( .B1(n4700), .B2(n4514), .A(n4513), .ZN(n4515) );
  NAND2_X1 U4972 ( .A1(n4609), .A2(n4515), .ZN(n4516) );
  OAI211_X1 U4973 ( .C1(n4612), .C2(n4694), .A(n4517), .B(n4516), .ZN(U3243)
         );
  AOI211_X1 U4974 ( .C1(n2307), .C2(n4519), .A(n4518), .B(n4650), .ZN(n4521)
         );
  AOI211_X1 U4975 ( .C1(n4646), .C2(ADDR_REG_5__SCAN_IN), .A(n4521), .B(n4520), 
        .ZN(n4527) );
  AOI21_X1 U4976 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n4525) );
  NAND2_X1 U4977 ( .A1(n4609), .A2(n4525), .ZN(n4526) );
  OAI211_X1 U4978 ( .C1(n4612), .C2(n4711), .A(n4527), .B(n4526), .ZN(U3245)
         );
  AOI211_X1 U4979 ( .C1(n2928), .C2(n4529), .A(n4528), .B(n4650), .ZN(n4531)
         );
  AOI211_X1 U4980 ( .C1(n4646), .C2(ADDR_REG_6__SCAN_IN), .A(n4531), .B(n4530), 
        .ZN(n4536) );
  AOI21_X1 U4981 ( .B1(n4533), .B2(n4532), .A(n2303), .ZN(n4534) );
  NAND2_X1 U4982 ( .A1(n4609), .A2(n4534), .ZN(n4535) );
  OAI211_X1 U4983 ( .C1(n4612), .C2(n4718), .A(n4536), .B(n4535), .ZN(U3246)
         );
  AOI22_X1 U4984 ( .A1(n4538), .A2(n4537), .B1(REG2_REG_7__SCAN_IN), .B2(n4720), .ZN(n4540) );
  OAI21_X1 U4985 ( .B1(n4541), .B2(n4540), .A(n4607), .ZN(n4539) );
  AOI21_X1 U4986 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4543) );
  AOI211_X1 U4987 ( .C1(n4646), .C2(ADDR_REG_7__SCAN_IN), .A(n4543), .B(n4542), 
        .ZN(n4548) );
  NAND2_X1 U4988 ( .A1(n2309), .A2(n4544), .ZN(n4546) );
  AOI21_X1 U4989 ( .B1(n2269), .B2(n4546), .A(n4647), .ZN(n4545) );
  OAI21_X1 U4990 ( .B1(n2269), .B2(n4546), .A(n4545), .ZN(n4547) );
  OAI211_X1 U4991 ( .C1(n4612), .C2(n4720), .A(n4548), .B(n4547), .ZN(U3247)
         );
  AOI21_X1 U4992 ( .B1(n4646), .B2(ADDR_REG_8__SCAN_IN), .A(n4549), .ZN(n4557)
         );
  OAI211_X1 U4993 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4551), .A(n4607), .B(n4550), 
        .ZN(n4556) );
  NAND2_X1 U4994 ( .A1(n4749), .A2(n4656), .ZN(n4555) );
  OAI211_X1 U4995 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4553), .A(n4609), .B(n4552), 
        .ZN(n4554) );
  NAND4_X1 U4996 ( .A1(n4557), .A2(n4556), .A3(n4555), .A4(n4554), .ZN(U3248)
         );
  INV_X1 U4997 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U4998 ( .A1(n4558), .A2(REG1_REG_9__SCAN_IN), .B1(n4767), .B2(n4752), .ZN(n4561) );
  OAI21_X1 U4999 ( .B1(n4561), .B2(n4560), .A(n4609), .ZN(n4559) );
  AOI21_X1 U5000 ( .B1(n4561), .B2(n4560), .A(n4559), .ZN(n4563) );
  AOI211_X1 U5001 ( .C1(n4646), .C2(ADDR_REG_9__SCAN_IN), .A(n4563), .B(n4562), 
        .ZN(n4568) );
  OAI211_X1 U5002 ( .C1(n4566), .C2(n4565), .A(n4607), .B(n4564), .ZN(n4567)
         );
  OAI211_X1 U5003 ( .C1(n4612), .C2(n4752), .A(n4568), .B(n4567), .ZN(U3249)
         );
  OAI21_X1 U5004 ( .B1(n4570), .B2(REG1_REG_11__SCAN_IN), .A(n4569), .ZN(n4572) );
  OAI21_X1 U5005 ( .B1(n2266), .B2(n4572), .A(n4609), .ZN(n4571) );
  AOI21_X1 U5006 ( .B1(n2266), .B2(n4572), .A(n4571), .ZN(n4574) );
  AOI211_X1 U5007 ( .C1(n4646), .C2(ADDR_REG_11__SCAN_IN), .A(n4574), .B(n4573), .ZN(n4579) );
  OAI211_X1 U5008 ( .C1(n4577), .C2(n4576), .A(n4607), .B(n4575), .ZN(n4578)
         );
  OAI211_X1 U5009 ( .C1(n4612), .C2(n4783), .A(n4579), .B(n4578), .ZN(U3251)
         );
  AOI21_X1 U5010 ( .B1(n4646), .B2(ADDR_REG_12__SCAN_IN), .A(n4580), .ZN(n4589) );
  OAI211_X1 U5011 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4582), .A(n4609), .B(n4581), .ZN(n4588) );
  NAND2_X1 U5012 ( .A1(n4583), .A2(n4656), .ZN(n4587) );
  OAI211_X1 U5013 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4585), .A(n4607), .B(n4584), .ZN(n4586) );
  NAND4_X1 U5014 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(U3252)
         );
  AOI21_X1 U5015 ( .B1(n4820), .B2(n3153), .A(n4590), .ZN(n4591) );
  XNOR2_X1 U5016 ( .A(n4592), .B(n4591), .ZN(n4600) );
  AOI21_X1 U5017 ( .B1(n4820), .B2(n3150), .A(n4593), .ZN(n4595) );
  XNOR2_X1 U5018 ( .A(n4595), .B(n4594), .ZN(n4596) );
  OAI22_X1 U5019 ( .A1(n4820), .A2(n4612), .B1(n4650), .B2(n4596), .ZN(n4597)
         );
  AOI211_X1 U5020 ( .C1(n4646), .C2(ADDR_REG_13__SCAN_IN), .A(n4598), .B(n4597), .ZN(n4599) );
  OAI21_X1 U5021 ( .B1(n4600), .B2(n4647), .A(n4599), .ZN(U3253) );
  AOI21_X1 U5022 ( .B1(n4646), .B2(ADDR_REG_16__SCAN_IN), .A(n4601), .ZN(n4611) );
  OAI21_X1 U5023 ( .B1(n4603), .B2(n3267), .A(n4602), .ZN(n4608) );
  OAI21_X1 U5024 ( .B1(n4605), .B2(n4115), .A(n4604), .ZN(n4606) );
  AOI22_X1 U5025 ( .A1(n4609), .A2(n4608), .B1(n4607), .B2(n4606), .ZN(n4610)
         );
  OAI211_X1 U5026 ( .C1(n4877), .C2(n4612), .A(n4611), .B(n4610), .ZN(U3256)
         );
  AOI211_X1 U5027 ( .C1(n4614), .C2(n4613), .A(n2281), .B(n4650), .ZN(n4615)
         );
  AOI211_X1 U5028 ( .C1(n4646), .C2(ADDR_REG_18__SCAN_IN), .A(n4616), .B(n4615), .ZN(n4625) );
  INV_X1 U5029 ( .A(n4617), .ZN(n4620) );
  INV_X1 U5030 ( .A(n4618), .ZN(n4619) );
  AOI21_X1 U5031 ( .B1(n4620), .B2(n4619), .A(n4647), .ZN(n4622) );
  AOI22_X1 U5032 ( .A1(n4623), .A2(n4622), .B1(n4656), .B2(n4621), .ZN(n4624)
         );
  NAND2_X1 U5033 ( .A1(n4625), .A2(n4624), .ZN(U3258) );
  AOI22_X1 U5034 ( .A1(STATE_REG_SCAN_IN), .A2(n2634), .B1(n4626), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5035 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4646), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4644) );
  AOI211_X1 U5036 ( .C1(n4629), .C2(n4628), .A(n4627), .B(n4650), .ZN(n4634)
         );
  AOI211_X1 U5037 ( .C1(n4632), .C2(n4631), .A(n4630), .B(n4647), .ZN(n4633)
         );
  AOI211_X1 U5038 ( .C1(n4656), .C2(n4682), .A(n4634), .B(n4633), .ZN(n4643)
         );
  INV_X1 U5039 ( .A(n4635), .ZN(n4640) );
  NAND2_X1 U5040 ( .A1(n4636), .A2(n4639), .ZN(n4638) );
  OAI211_X1 U5041 ( .C1(n4640), .C2(n4639), .A(n4638), .B(n4637), .ZN(n4641)
         );
  OAI211_X1 U5042 ( .C1(n2614), .C2(n4642), .A(n4641), .B(U4043), .ZN(n4657)
         );
  NAND3_X1 U5043 ( .A1(n4644), .A2(n4643), .A3(n4657), .ZN(U3242) );
  AOI21_X1 U5044 ( .B1(n4646), .B2(ADDR_REG_4__SCAN_IN), .A(n4645), .ZN(n4659)
         );
  AOI211_X1 U5045 ( .C1(n4708), .C2(n4649), .A(n4648), .B(n4647), .ZN(n4654)
         );
  AOI211_X1 U5046 ( .C1(n2738), .C2(n4652), .A(n4651), .B(n4650), .ZN(n4653)
         );
  AOI211_X1 U5047 ( .C1(n4656), .C2(n4655), .A(n4654), .B(n4653), .ZN(n4658)
         );
  NAND3_X1 U5048 ( .A1(n4659), .A2(n4658), .A3(n4657), .ZN(U3244) );
  INV_X1 U5049 ( .A(n4696), .ZN(n4823) );
  NAND2_X1 U5050 ( .A1(n4660), .A2(n4856), .ZN(n4662) );
  AND2_X1 U5051 ( .A1(n2657), .A2(n4862), .ZN(n4661) );
  AOI21_X1 U5052 ( .B1(n4672), .B2(n4662), .A(n4661), .ZN(n4669) );
  NAND2_X1 U5053 ( .A1(n4664), .A2(n4663), .ZN(n4665) );
  NAND2_X1 U5054 ( .A1(n4669), .A2(n4665), .ZN(n4671) );
  AOI21_X1 U5055 ( .B1(n4823), .B2(n4672), .A(n4671), .ZN(n4667) );
  AOI22_X1 U5056 ( .A1(n4894), .A2(n4667), .B1(n2638), .B2(n4892), .ZN(U3518)
         );
  INV_X1 U5057 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5058 ( .A1(n4897), .A2(n4667), .B1(n4666), .B2(n4895), .ZN(U3467)
         );
  NAND3_X1 U5059 ( .A1(n4669), .A2(n3809), .A3(n4668), .ZN(n4670) );
  NAND2_X1 U5060 ( .A1(n4671), .A2(n4670), .ZN(n4675) );
  AOI22_X1 U5061 ( .A1(n4672), .A2(n4805), .B1(REG3_REG_0__SCAN_IN), .B2(n4867), .ZN(n4673) );
  OAI221_X1 U5062 ( .B1(n4939), .B2(n4675), .C1(n4674), .C2(n2627), .A(n4673), 
        .ZN(U3290) );
  NOR2_X1 U5063 ( .A1(n4676), .A2(n4888), .ZN(n4678) );
  AOI211_X1 U5064 ( .C1(n4883), .C2(n4679), .A(n4678), .B(n4677), .ZN(n4681)
         );
  AOI22_X1 U5065 ( .A1(n4894), .A2(n4681), .B1(n2420), .B2(n4892), .ZN(U3519)
         );
  INV_X1 U5066 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5067 ( .A1(n4897), .A2(n4681), .B1(n4680), .B2(n4895), .ZN(U3469)
         );
  INV_X1 U5068 ( .A(n4682), .ZN(n4684) );
  INV_X1 U5069 ( .A(DATAI_2_), .ZN(n4683) );
  AOI22_X1 U5070 ( .A1(STATE_REG_SCAN_IN), .A2(n4684), .B1(n4683), .B2(U3149), 
        .ZN(U3350) );
  AND3_X1 U5071 ( .A1(n4686), .A2(n4883), .A3(n4685), .ZN(n4688) );
  AOI211_X1 U5072 ( .C1(n4823), .C2(n4689), .A(n4688), .B(n4687), .ZN(n4692)
         );
  INV_X1 U5073 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5074 ( .A1(n4894), .A2(n4692), .B1(n4690), .B2(n4892), .ZN(U3520)
         );
  INV_X1 U5075 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5076 ( .A1(n4897), .A2(n4692), .B1(n4691), .B2(n4895), .ZN(U3471)
         );
  INV_X1 U5077 ( .A(DATAI_3_), .ZN(n4693) );
  AOI22_X1 U5078 ( .A1(STATE_REG_SCAN_IN), .A2(n4694), .B1(n4693), .B2(U3149), 
        .ZN(U3349) );
  OAI22_X1 U5079 ( .A1(n4697), .A2(n4696), .B1(n4887), .B2(n4695), .ZN(n4698)
         );
  NOR2_X1 U5080 ( .A1(n4699), .A2(n4698), .ZN(n4701) );
  AOI22_X1 U5081 ( .A1(n4894), .A2(n4701), .B1(n4700), .B2(n4892), .ZN(U3521)
         );
  AOI22_X1 U5082 ( .A1(n4897), .A2(n4701), .B1(n2723), .B2(n4895), .ZN(U3473)
         );
  AOI22_X1 U5083 ( .A1(STATE_REG_SCAN_IN), .A2(n4703), .B1(n4702), .B2(U3149), 
        .ZN(U3348) );
  INV_X1 U5084 ( .A(n4704), .ZN(n4706) );
  AOI211_X1 U5085 ( .C1(n4707), .C2(n4823), .A(n4706), .B(n4705), .ZN(n4709)
         );
  AOI22_X1 U5086 ( .A1(n4894), .A2(n4709), .B1(n4708), .B2(n4892), .ZN(U3522)
         );
  AOI22_X1 U5087 ( .A1(n4897), .A2(n4709), .B1(n2739), .B2(n4895), .ZN(U3475)
         );
  AOI22_X1 U5088 ( .A1(STATE_REG_SCAN_IN), .A2(n4711), .B1(n4710), .B2(U3149), 
        .ZN(U3347) );
  NOR2_X1 U5089 ( .A1(n4712), .A2(n4888), .ZN(n4714) );
  AOI211_X1 U5090 ( .C1(n4883), .C2(n4715), .A(n4714), .B(n4713), .ZN(n4716)
         );
  AOI22_X1 U5091 ( .A1(n4894), .A2(n4716), .B1(n2760), .B2(n4892), .ZN(U3523)
         );
  AOI22_X1 U5092 ( .A1(n4897), .A2(n4716), .B1(n2759), .B2(n4895), .ZN(U3477)
         );
  AOI22_X1 U5093 ( .A1(STATE_REG_SCAN_IN), .A2(n4718), .B1(n4717), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5094 ( .A1(STATE_REG_SCAN_IN), .A2(n4720), .B1(n4719), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5095 ( .A(n4721), .ZN(n4724) );
  AOI21_X1 U5096 ( .B1(n4722), .B2(n4733), .A(n4887), .ZN(n4723) );
  NAND2_X1 U5097 ( .A1(n4724), .A2(n4723), .ZN(n4743) );
  INV_X1 U5098 ( .A(n4726), .ZN(n4729) );
  XNOR2_X1 U5099 ( .A(n4725), .B(n4729), .ZN(n4744) );
  NAND2_X1 U5100 ( .A1(n4744), .A2(n4727), .ZN(n4728) );
  OAI211_X1 U5101 ( .C1(n3809), .C2(n4743), .A(n4728), .B(n4674), .ZN(n4739)
         );
  INV_X1 U5102 ( .A(n4758), .ZN(n4738) );
  XNOR2_X1 U5103 ( .A(n4730), .B(n4729), .ZN(n4732) );
  NAND2_X1 U5104 ( .A1(n4732), .A2(n4731), .ZN(n4736) );
  AOI22_X1 U5105 ( .A1(n4734), .A2(n4849), .B1(n4787), .B2(n4733), .ZN(n4735)
         );
  OAI211_X1 U5106 ( .C1(n4738), .C2(n4737), .A(n4736), .B(n4735), .ZN(n4747)
         );
  OAI22_X1 U5107 ( .A1(n4739), .A2(n4747), .B1(REG2_REG_7__SCAN_IN), .B2(n4674), .ZN(n4740) );
  OAI21_X1 U5108 ( .B1(n4742), .B2(n4741), .A(n4740), .ZN(U3283) );
  INV_X1 U5109 ( .A(n4743), .ZN(n4746) );
  AND2_X1 U5110 ( .A1(n4744), .A2(n4879), .ZN(n4745) );
  NOR3_X1 U5111 ( .A1(n4747), .A2(n4746), .A3(n4745), .ZN(n4748) );
  AOI22_X1 U5112 ( .A1(n4894), .A2(n4748), .B1(n2914), .B2(n4892), .ZN(U3525)
         );
  AOI22_X1 U5113 ( .A1(n4897), .A2(n4748), .B1(n2919), .B2(n4895), .ZN(U3481)
         );
  AOI22_X1 U5114 ( .A1(STATE_REG_SCAN_IN), .A2(n2984), .B1(n4750), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5115 ( .A(DATAI_9_), .ZN(n4751) );
  AOI22_X1 U5116 ( .A1(STATE_REG_SCAN_IN), .A2(n4752), .B1(n4751), .B2(U3149), 
        .ZN(U3343) );
  OAI21_X1 U5117 ( .B1(n3163), .B2(n2350), .A(n4754), .ZN(n4755) );
  XNOR2_X1 U5118 ( .A(n4755), .B(n4757), .ZN(n4772) );
  XOR2_X1 U5119 ( .A(n4757), .B(n4756), .Z(n4761) );
  AOI22_X1 U5120 ( .A1(n4758), .A2(n4849), .B1(n4787), .B2(n4765), .ZN(n4760)
         );
  NAND2_X1 U5121 ( .A1(n4788), .A2(n4862), .ZN(n4759) );
  OAI211_X1 U5122 ( .C1(n4761), .C2(n4856), .A(n4760), .B(n4759), .ZN(n4762)
         );
  AOI21_X1 U5123 ( .B1(n4794), .B2(n4772), .A(n4762), .ZN(n4775) );
  AOI21_X1 U5124 ( .B1(n4765), .B2(n4764), .A(n3194), .ZN(n4771) );
  AOI22_X1 U5125 ( .A1(n4772), .A2(n4823), .B1(n4883), .B2(n4771), .ZN(n4766)
         );
  AND2_X1 U5126 ( .A1(n4775), .A2(n4766), .ZN(n4768) );
  AOI22_X1 U5127 ( .A1(n4894), .A2(n4768), .B1(n4767), .B2(n4892), .ZN(U3527)
         );
  AOI22_X1 U5128 ( .A1(n4897), .A2(n4768), .B1(n3033), .B2(n4895), .ZN(U3485)
         );
  INV_X1 U5129 ( .A(n4769), .ZN(n4770) );
  AOI22_X1 U5130 ( .A1(n4770), .A2(n4867), .B1(REG2_REG_9__SCAN_IN), .B2(n4939), .ZN(n4774) );
  AOI22_X1 U5131 ( .A1(n4772), .A2(n4805), .B1(n4940), .B2(n4771), .ZN(n4773)
         );
  OAI211_X1 U5132 ( .C1(n4939), .C2(n4775), .A(n4774), .B(n4773), .ZN(U3281)
         );
  AOI22_X1 U5133 ( .A1(n4776), .A2(n4867), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4939), .ZN(n4780) );
  AOI22_X1 U5134 ( .A1(n4778), .A2(n4871), .B1(n4940), .B2(n4777), .ZN(n4779)
         );
  OAI211_X1 U5135 ( .C1(n4939), .C2(n4781), .A(n4780), .B(n4779), .ZN(U3280)
         );
  AOI22_X1 U5136 ( .A1(STATE_REG_SCAN_IN), .A2(n4783), .B1(n4782), .B2(U3149), 
        .ZN(U3341) );
  XNOR2_X1 U5137 ( .A(n4784), .B(n4785), .ZN(n4806) );
  XNOR2_X1 U5138 ( .A(n4786), .B(n4785), .ZN(n4792) );
  AOI22_X1 U5139 ( .A1(n4788), .A2(n4849), .B1(n4798), .B2(n4787), .ZN(n4791)
         );
  NAND2_X1 U5140 ( .A1(n4789), .A2(n4862), .ZN(n4790) );
  OAI211_X1 U5141 ( .C1(n4792), .C2(n4856), .A(n4791), .B(n4790), .ZN(n4793)
         );
  AOI21_X1 U5142 ( .B1(n4794), .B2(n4806), .A(n4793), .ZN(n4809) );
  INV_X1 U5143 ( .A(n4795), .ZN(n4797) );
  AOI21_X1 U5144 ( .B1(n4798), .B2(n4797), .A(n4796), .ZN(n4804) );
  AOI22_X1 U5145 ( .A1(n4806), .A2(n4823), .B1(n4883), .B2(n4804), .ZN(n4799)
         );
  AND2_X1 U5146 ( .A1(n4809), .A2(n4799), .ZN(n4801) );
  AOI22_X1 U5147 ( .A1(n4894), .A2(n4801), .B1(n3097), .B2(n4892), .ZN(U3529)
         );
  INV_X1 U5148 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4800) );
  AOI22_X1 U5149 ( .A1(n4897), .A2(n4801), .B1(n4800), .B2(n4895), .ZN(U3489)
         );
  INV_X1 U5150 ( .A(n4802), .ZN(n4803) );
  AOI22_X1 U5151 ( .A1(n4803), .A2(n4867), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4939), .ZN(n4808) );
  AOI22_X1 U5152 ( .A1(n4806), .A2(n4805), .B1(n4940), .B2(n4804), .ZN(n4807)
         );
  OAI211_X1 U5153 ( .C1(n4939), .C2(n4809), .A(n4808), .B(n4807), .ZN(U3279)
         );
  AOI22_X1 U5154 ( .A1(STATE_REG_SCAN_IN), .A2(n4811), .B1(n4810), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5155 ( .A1(n4812), .A2(n4867), .B1(REG2_REG_12__SCAN_IN), .B2(
        n4939), .ZN(n4817) );
  INV_X1 U5156 ( .A(n4813), .ZN(n4814) );
  AOI22_X1 U5157 ( .A1(n4815), .A2(n4871), .B1(n4940), .B2(n4814), .ZN(n4816)
         );
  OAI211_X1 U5158 ( .C1(n4939), .C2(n4818), .A(n4817), .B(n4816), .ZN(U3278)
         );
  AOI22_X1 U5159 ( .A1(STATE_REG_SCAN_IN), .A2(n4820), .B1(n4819), .B2(U3149), 
        .ZN(U3339) );
  NOR2_X1 U5160 ( .A1(n4821), .A2(n4887), .ZN(n4822) );
  AOI21_X1 U5161 ( .B1(n4824), .B2(n4823), .A(n4822), .ZN(n4825) );
  AOI22_X1 U5162 ( .A1(n4894), .A2(n4828), .B1(n3153), .B2(n4892), .ZN(U3531)
         );
  INV_X1 U5163 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U5164 ( .A1(n4897), .A2(n4828), .B1(n4827), .B2(n4895), .ZN(U3493)
         );
  INV_X1 U5165 ( .A(n4850), .ZN(n4829) );
  OAI22_X1 U5166 ( .A1(n4831), .A2(n4913), .B1(n4830), .B2(n4829), .ZN(n4836)
         );
  INV_X1 U5167 ( .A(n4832), .ZN(n4833) );
  OAI21_X1 U5168 ( .B1(n4834), .B2(n4852), .A(n4833), .ZN(n4835) );
  NOR2_X1 U5169 ( .A1(n4836), .A2(n4835), .ZN(n4842) );
  XNOR2_X1 U5170 ( .A(n4838), .B(n4837), .ZN(n4839) );
  XNOR2_X1 U5171 ( .A(n3510), .B(n4839), .ZN(n4840) );
  NAND2_X1 U5172 ( .A1(n4840), .A2(n4925), .ZN(n4841) );
  OAI211_X1 U5173 ( .C1(n4930), .C2(n4866), .A(n4842), .B(n4841), .ZN(U3238)
         );
  NOR2_X1 U5174 ( .A1(n4844), .A2(n4843), .ZN(n4845) );
  XOR2_X1 U5175 ( .A(n4857), .B(n4845), .Z(n4872) );
  NOR2_X1 U5176 ( .A1(n4846), .A2(n4852), .ZN(n4847) );
  OR2_X1 U5177 ( .A1(n4848), .A2(n4847), .ZN(n4869) );
  NAND2_X1 U5178 ( .A1(n4850), .A2(n4849), .ZN(n4851) );
  OAI21_X1 U5179 ( .B1(n4853), .B2(n4852), .A(n4851), .ZN(n4860) );
  INV_X1 U5180 ( .A(n4854), .ZN(n4855) );
  AOI211_X1 U5181 ( .C1(n4858), .C2(n4857), .A(n4856), .B(n4855), .ZN(n4859)
         );
  AOI211_X1 U5182 ( .C1(n4862), .C2(n4861), .A(n4860), .B(n4859), .ZN(n4875)
         );
  OAI21_X1 U5183 ( .B1(n4887), .B2(n4869), .A(n4875), .ZN(n4863) );
  AOI21_X1 U5184 ( .B1(n4879), .B2(n4872), .A(n4863), .ZN(n4865) );
  AOI22_X1 U5185 ( .A1(n4894), .A2(n4865), .B1(n3782), .B2(n4892), .ZN(U3533)
         );
  INV_X1 U5186 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U5187 ( .A1(n4897), .A2(n4865), .B1(n4864), .B2(n4895), .ZN(U3497)
         );
  INV_X1 U5188 ( .A(n4866), .ZN(n4868) );
  AOI22_X1 U5189 ( .A1(n4868), .A2(n4867), .B1(REG2_REG_15__SCAN_IN), .B2(
        n4939), .ZN(n4874) );
  INV_X1 U5190 ( .A(n4869), .ZN(n4870) );
  AOI22_X1 U5191 ( .A1(n4872), .A2(n4871), .B1(n4940), .B2(n4870), .ZN(n4873)
         );
  OAI211_X1 U5192 ( .C1(n4939), .C2(n4875), .A(n4874), .B(n4873), .ZN(U3275)
         );
  AOI22_X1 U5193 ( .A1(STATE_REG_SCAN_IN), .A2(n4877), .B1(n4876), .B2(U3149), 
        .ZN(U3336) );
  AND3_X1 U5194 ( .A1(n4117), .A2(n4879), .A3(n4878), .ZN(n4881) );
  AOI211_X1 U5195 ( .C1(n4883), .C2(n4882), .A(n4881), .B(n4880), .ZN(n4885)
         );
  AOI22_X1 U5196 ( .A1(n4894), .A2(n4885), .B1(n3267), .B2(n4892), .ZN(U3534)
         );
  INV_X1 U5197 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U5198 ( .A1(n4897), .A2(n4885), .B1(n4884), .B2(n4895), .ZN(U3499)
         );
  OAI22_X1 U5199 ( .A1(n4889), .A2(n4888), .B1(n4887), .B2(n4886), .ZN(n4890)
         );
  NOR2_X1 U5200 ( .A1(n4891), .A2(n4890), .ZN(n4896) );
  AOI22_X1 U5201 ( .A1(n4894), .A2(n4896), .B1(n4893), .B2(n4892), .ZN(U3535)
         );
  AOI22_X1 U5202 ( .A1(n4897), .A2(n4896), .B1(n3297), .B2(n4895), .ZN(U3501)
         );
  AOI22_X1 U5203 ( .A1(n4899), .A2(n4898), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4909) );
  OR2_X1 U5204 ( .A1(n4900), .A2(n4901), .ZN(n4916) );
  INV_X1 U5205 ( .A(n4915), .ZN(n4903) );
  OAI21_X1 U5206 ( .B1(n4903), .B2(n4901), .A(n4900), .ZN(n4902) );
  OAI211_X1 U5207 ( .C1(n4916), .C2(n4903), .A(n4925), .B(n4902), .ZN(n4907)
         );
  AOI22_X1 U5208 ( .A1(n4905), .A2(n4924), .B1(n4921), .B2(n4904), .ZN(n4906)
         );
  AND2_X1 U5209 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  OAI211_X1 U5210 ( .C1(n4930), .C2(n4910), .A(n4909), .B(n4908), .ZN(U3230)
         );
  OAI22_X1 U5211 ( .A1(n4913), .A2(n4912), .B1(STATE_REG_SCAN_IN), .B2(n4911), 
        .ZN(n4914) );
  INV_X1 U5212 ( .A(n4914), .ZN(n4928) );
  NAND2_X1 U5213 ( .A1(n4916), .A2(n4915), .ZN(n4920) );
  XNOR2_X1 U5214 ( .A(n4918), .B(n4917), .ZN(n4919) );
  XNOR2_X1 U5215 ( .A(n4920), .B(n4919), .ZN(n4926) );
  AOI222_X1 U5216 ( .A1(n4926), .A2(n4925), .B1(n4924), .B2(n4923), .C1(n4922), 
        .C2(n4921), .ZN(n4927) );
  OAI211_X1 U5217 ( .C1(n4930), .C2(n4929), .A(n4928), .B(n4927), .ZN(U3220)
         );
  AOI22_X1 U5218 ( .A1(STATE_REG_SCAN_IN), .A2(n4932), .B1(n4931), .B2(U3149), 
        .ZN(U3324) );
  OAI22_X1 U5219 ( .A1(n4935), .A2(n4934), .B1(n4933), .B2(n4674), .ZN(n4936)
         );
  INV_X1 U5220 ( .A(n4936), .ZN(n4937) );
  OAI21_X1 U5221 ( .B1(n4939), .B2(n4938), .A(n4937), .ZN(U3261) );
  AOI22_X1 U5222 ( .A1(n4941), .A2(n4940), .B1(n4939), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4942) );
  OAI21_X1 U5223 ( .B1(n4939), .B2(n4943), .A(n4942), .ZN(U3260) );
  CLKBUF_X1 U2295 ( .A(n3007), .Z(n2260) );
  CLKBUF_X1 U2296 ( .A(n3007), .Z(n2261) );
  CLKBUF_X1 U2468 ( .A(n2632), .Z(n4668) );
endmodule

