

module b22_C_gen_AntiSAT_k_128_1 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15400, n15401;

  NAND2_X2 U7213 ( .A1(n9592), .A2(P3_U3151), .ZN(n13125) );
  AOI211_X1 U7214 ( .C1(n13222), .C2(n13226), .A(n14926), .B(n13225), .ZN(
        n13227) );
  AOI21_X1 U7215 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(n13407) );
  OR2_X1 U7216 ( .A1(n13890), .A2(n13889), .ZN(n13891) );
  NAND2_X1 U7217 ( .A1(n7614), .A2(n7613), .ZN(n14205) );
  NAND2_X1 U7218 ( .A1(n9099), .A2(n9098), .ZN(n13702) );
  OR2_X1 U7219 ( .A1(n7558), .A2(n11336), .ZN(n7561) );
  CLKBUF_X2 U7220 ( .A(n10879), .Z(n12518) );
  INV_X2 U7222 ( .A(n6502), .ZN(n9471) );
  INV_X4 U7223 ( .A(n12548), .ZN(n6483) );
  NAND2_X1 U7224 ( .A1(n11560), .A2(n8102), .ZN(n11050) );
  OR2_X1 U7225 ( .A1(n9218), .A2(n11210), .ZN(n10662) );
  CLKBUF_X2 U7226 ( .A(n8357), .Z(n8083) );
  NAND2_X1 U7227 ( .A1(n7713), .A2(n7712), .ZN(n11600) );
  CLKBUF_X2 U7228 ( .A(n7852), .Z(n8358) );
  AND3_X1 U7229 ( .A1(n7702), .A2(n7701), .A3(n7700), .ZN(n14850) );
  XNOR2_X1 U7230 ( .A(n8849), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8820) );
  CLKBUF_X2 U7231 ( .A(n7851), .Z(n8356) );
  CLKBUF_X2 U7232 ( .A(n7853), .Z(n8357) );
  NAND2_X1 U7233 ( .A1(n10201), .A2(n10200), .ZN(n12028) );
  NAND4_X1 U7234 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n14086)
         );
  CLKBUF_X1 U7235 ( .A(n7675), .Z(n6504) );
  NOR2_X2 U7236 ( .A1(n11704), .A2(n8100), .ZN(n8202) );
  CLKBUF_X2 U7237 ( .A(n7675), .Z(n6503) );
  INV_X1 U7238 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9589) );
  AND2_X1 U7239 ( .A1(n10512), .A2(n9592), .ZN(n7685) );
  NOR2_X1 U7240 ( .A1(n8163), .A2(n7596), .ZN(n7597) );
  AND3_X1 U7241 ( .A1(n7587), .A2(n7586), .A3(n7585), .ZN(n7590) );
  AND2_X1 U7242 ( .A1(n7032), .A2(n7031), .ZN(n7591) );
  NOR2_X1 U7243 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7032) );
  NOR2_X1 U7244 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7031) );
  NAND2_X1 U7245 ( .A1(n13153), .A2(n6468), .ZN(n6465) );
  AND2_X2 U7246 ( .A1(n6465), .A2(n6466), .ZN(n13163) );
  OR2_X1 U7247 ( .A1(n6467), .A2(n13203), .ZN(n6466) );
  INV_X1 U7248 ( .A(n6601), .ZN(n6467) );
  AND2_X1 U7249 ( .A1(n13204), .A2(n6601), .ZN(n6468) );
  INV_X1 U7250 ( .A(n6663), .ZN(n6469) );
  NOR2_X1 U7251 ( .A1(n10702), .A2(n10701), .ZN(n10820) );
  NAND2_X1 U7252 ( .A1(n8113), .A2(n6473), .ZN(n6470) );
  AND2_X1 U7253 ( .A1(n6470), .A2(n6471), .ZN(n11885) );
  OR2_X1 U7254 ( .A1(n6472), .A2(n11870), .ZN(n6471) );
  INV_X1 U7255 ( .A(n8114), .ZN(n6472) );
  AND2_X1 U7256 ( .A1(n8112), .A2(n8114), .ZN(n6473) );
  CLKBUF_X1 U7257 ( .A(n11049), .Z(n6474) );
  NAND2_X1 U7258 ( .A1(n14323), .A2(n8129), .ZN(n6475) );
  NOR2_X1 U7259 ( .A1(n7092), .A2(n7686), .ZN(n6476) );
  NOR2_X1 U7260 ( .A1(n7092), .A2(n7686), .ZN(n7090) );
  INV_X4 U7261 ( .A(n15334), .ZN(n13001) );
  XOR2_X1 U7262 ( .A(n15284), .B(n11524), .Z(n15283) );
  AND3_X1 U7264 ( .A1(n9708), .A2(n9707), .A3(n9706), .ZN(n10837) );
  OR2_X1 U7265 ( .A1(n8882), .A2(n8881), .ZN(n11231) );
  CLKBUF_X3 U7266 ( .A(n10058), .Z(n10033) );
  CLKBUF_X2 U7267 ( .A(n9695), .Z(n10099) );
  OAI211_X1 U7268 ( .C1(n10033), .C2(SI_5_), .A(n9730), .B(n9729), .ZN(n11449)
         );
  INV_X1 U7269 ( .A(n10812), .ZN(n11089) );
  XNOR2_X1 U7270 ( .A(n10664), .B(n10665), .ZN(n10720) );
  INV_X2 U7271 ( .A(n8904), .ZN(n9206) );
  NAND2_X1 U7273 ( .A1(n8902), .A2(n8901), .ZN(n11306) );
  NAND2_X1 U7274 ( .A1(n7821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7826) );
  OAI211_X1 U7275 ( .C1(n10058), .C2(n7504), .A(n9688), .B(n9687), .ZN(n15326)
         );
  NAND2_X1 U7276 ( .A1(n10106), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10108) );
  AND2_X1 U7277 ( .A1(n11433), .A2(n11432), .ZN(n11437) );
  NAND2_X2 U7279 ( .A1(n9032), .A2(n9031), .ZN(n14656) );
  NAND2_X1 U7280 ( .A1(n8808), .A2(n8807), .ZN(n13505) );
  XNOR2_X1 U7281 ( .A(n10108), .B(n10107), .ZN(n11338) );
  INV_X1 U7282 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14177) );
  NAND2_X1 U7283 ( .A1(n7821), .A2(n7800), .ZN(n14172) );
  NOR2_X4 U7284 ( .A1(n8720), .A2(n10865), .ZN(n14916) );
  XNOR2_X2 U7285 ( .A(n12505), .B(n12506), .ZN(n13245) );
  NAND2_X2 U7286 ( .A1(n13598), .A2(n7153), .ZN(n13586) );
  OAI21_X2 U7287 ( .B1(n12261), .B2(n14621), .A(n12260), .ZN(n12731) );
  XNOR2_X1 U7288 ( .A(n10946), .B(n10962), .ZN(n15209) );
  NAND2_X2 U7289 ( .A1(n7270), .A2(n7268), .ZN(n12505) );
  NOR2_X2 U7290 ( .A1(n10840), .A2(n10839), .ZN(n11160) );
  INV_X4 U7292 ( .A(n11800), .ZN(n12485) );
  NOR2_X2 U7293 ( .A1(n15389), .A2(n8504), .ZN(n14538) );
  NOR2_X2 U7294 ( .A1(n15391), .A2(n15390), .ZN(n15389) );
  INV_X4 U7295 ( .A(n8898), .ZN(n9097) );
  INV_X2 U7296 ( .A(n8092), .ZN(n8364) );
  XNOR2_X2 U7297 ( .A(n7823), .B(n7822), .ZN(n8092) );
  BUF_X2 U7298 ( .A(n10669), .Z(n6477) );
  OAI211_X1 U7299 ( .C1(n9140), .C2(n10349), .A(n8866), .B(n8865), .ZN(n10669)
         );
  XNOR2_X2 U7300 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n8499) );
  INV_X1 U7301 ( .A(n6483), .ZN(n6478) );
  OAI22_X2 U7302 ( .A1(n14191), .A2(n14190), .B1(n14414), .B2(n14069), .ZN(
        n12427) );
  AOI21_X2 U7303 ( .B1(n14249), .B2(n7053), .A(n7050), .ZN(n14191) );
  XNOR2_X2 U7304 ( .A(n7826), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8422) );
  OAI21_X2 U7305 ( .B1(n7771), .B2(n7543), .A(n7542), .ZN(n7544) );
  NAND2_X2 U7306 ( .A1(n7174), .A2(n7173), .ZN(n7771) );
  BUF_X2 U7307 ( .A(n10058), .Z(n6480) );
  NAND2_X1 U7308 ( .A1(n10941), .A2(n9592), .ZN(n10058) );
  XNOR2_X2 U7309 ( .A(n8495), .B(n8494), .ZN(n8506) );
  XNOR2_X2 U7310 ( .A(n8455), .B(n8454), .ZN(n8495) );
  AOI21_X2 U7311 ( .B1(n12780), .B2(n12803), .A(n14587), .ZN(n12828) );
  NOR2_X2 U7312 ( .A1(n15228), .A2(n15227), .ZN(n15226) );
  NOR2_X2 U7313 ( .A1(n12849), .A2(n10254), .ZN(n12835) );
  NOR2_X2 U7314 ( .A1(n12850), .A2(n12852), .ZN(n12849) );
  XNOR2_X2 U7315 ( .A(n12089), .B(n11851), .ZN(n11497) );
  OAI22_X2 U7316 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13775), .B1(n10046), 
        .B2(n10045), .ZN(n10057) );
  AND2_X1 U7317 ( .A1(n13407), .A2(n13404), .ZN(n7146) );
  OR2_X1 U7318 ( .A1(n13887), .A2(n13997), .ZN(n13962) );
  AND2_X1 U7319 ( .A1(n8547), .A2(n8548), .ZN(n14531) );
  NAND2_X1 U7320 ( .A1(n14009), .A2(n14008), .ZN(n14007) );
  AND2_X1 U7321 ( .A1(n12513), .A2(n13183), .ZN(n13185) );
  AND2_X1 U7322 ( .A1(n10022), .A2(n10021), .ZN(n13071) );
  NAND2_X1 U7323 ( .A1(n14380), .A2(n7971), .ZN(n14361) );
  NAND2_X1 U7324 ( .A1(n12757), .A2(n12759), .ZN(n12797) );
  OAI21_X1 U7325 ( .B1(n7625), .B2(n6525), .A(n6638), .ZN(n6715) );
  NAND2_X1 U7326 ( .A1(n7129), .A2(n8980), .ZN(n11783) );
  OAI22_X1 U7327 ( .A1(n9307), .A2(n7339), .B1(n9308), .B2(n7340), .ZN(n9314)
         );
  OR2_X1 U7328 ( .A1(n15383), .A2(n15384), .ZN(n6896) );
  NOR2_X1 U7329 ( .A1(n14541), .A2(n8515), .ZN(n8517) );
  XNOR2_X2 U7330 ( .A(n14085), .B(n13916), .ZN(n11054) );
  INV_X1 U7331 ( .A(n14083), .ZN(n11854) );
  INV_X4 U7332 ( .A(n8341), .ZN(n6481) );
  INV_X2 U7333 ( .A(n13855), .ZN(n11847) );
  INV_X1 U7334 ( .A(n13935), .ZN(n13838) );
  INV_X2 U7335 ( .A(n6502), .ZN(n9477) );
  BUF_X2 U7336 ( .A(n9693), .Z(n10063) );
  INV_X1 U7337 ( .A(n6485), .ZN(n10323) );
  NOR2_X1 U7338 ( .A1(n10887), .A2(n8422), .ZN(n6485) );
  BUF_X2 U7339 ( .A(n7672), .Z(n8390) );
  CLKBUF_X2 U7340 ( .A(n8899), .Z(n9096) );
  OR2_X2 U7341 ( .A1(n11208), .A2(n9512), .ZN(n12548) );
  INV_X1 U7342 ( .A(n10512), .ZN(n7675) );
  INV_X4 U7343 ( .A(n7963), .ZN(n6482) );
  NAND2_X1 U7344 ( .A1(n8802), .A2(n8801), .ZN(n13379) );
  CLKBUF_X1 U7345 ( .A(n10206), .Z(n6501) );
  XNOR2_X1 U7346 ( .A(n6918), .B(n8815), .ZN(n9257) );
  INV_X4 U7348 ( .A(n7515), .ZN(n10344) );
  NAND2_X1 U7349 ( .A1(n7501), .A2(n7500), .ZN(n6713) );
  NAND2_X1 U7350 ( .A1(n9684), .A2(n9581), .ZN(n6973) );
  NAND2_X1 U7351 ( .A1(n7498), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6714) );
  NAND3_X1 U7352 ( .A1(n8154), .A2(n8097), .A3(n10322), .ZN(n8721) );
  OR2_X1 U7353 ( .A1(n14425), .A2(n14424), .ZN(n14492) );
  OAI21_X1 U7354 ( .B1(n13653), .B2(n13724), .A(n6734), .ZN(n13732) );
  OAI21_X1 U7355 ( .B1(n7146), .B2(n15145), .A(n9274), .ZN(n6706) );
  AND2_X1 U7356 ( .A1(n6490), .A2(n6491), .ZN(n13131) );
  NAND2_X1 U7357 ( .A1(n7128), .A2(n7126), .ZN(n13436) );
  OR2_X1 U7358 ( .A1(n12541), .A2(n12543), .ZN(n7275) );
  AND2_X1 U7359 ( .A1(n13999), .A2(n13998), .ZN(n14000) );
  NAND2_X1 U7360 ( .A1(n7309), .A2(n6553), .ZN(n14270) );
  NAND2_X1 U7361 ( .A1(n13464), .A2(n9167), .ZN(n13453) );
  NAND2_X1 U7362 ( .A1(n8393), .A2(n8392), .ZN(n8424) );
  NAND2_X1 U7363 ( .A1(n14303), .A2(n8133), .ZN(n14275) );
  OR2_X1 U7364 ( .A1(n13733), .A2(n13427), .ZN(n9204) );
  XNOR2_X1 U7365 ( .A(n13656), .B(n13441), .ZN(n13433) );
  NAND2_X1 U7366 ( .A1(n14007), .A2(n6554), .ZN(n13949) );
  NAND2_X1 U7367 ( .A1(n8751), .A2(n8750), .ZN(n13401) );
  XNOR2_X1 U7368 ( .A(n7606), .B(n7605), .ZN(n12425) );
  XNOR2_X1 U7369 ( .A(n14427), .B(n14070), .ZN(n14237) );
  NAND2_X1 U7370 ( .A1(n7612), .A2(n7578), .ZN(n7606) );
  NAND2_X2 U7371 ( .A1(n7820), .A2(n7819), .ZN(n14420) );
  NAND2_X1 U7372 ( .A1(n9156), .A2(n9155), .ZN(n13739) );
  NAND2_X1 U7373 ( .A1(n14037), .A2(n14038), .ZN(n14036) );
  OAI22_X1 U7374 ( .A1(n7818), .A2(n7575), .B1(n7816), .B2(n8689), .ZN(n7610)
         );
  AND2_X2 U7375 ( .A1(n9142), .A2(n9141), .ZN(n13490) );
  NAND2_X1 U7376 ( .A1(n13600), .A2(n13599), .ZN(n13598) );
  NAND2_X1 U7377 ( .A1(n7571), .A2(n7168), .ZN(n7166) );
  XOR2_X1 U7378 ( .A(n12798), .B(n12797), .Z(n12758) );
  AND2_X1 U7379 ( .A1(n12508), .A2(n12509), .ZN(n7277) );
  NAND2_X1 U7380 ( .A1(n7629), .A2(n7628), .ZN(n14438) );
  INV_X1 U7381 ( .A(n6715), .ZN(n7568) );
  NAND2_X1 U7382 ( .A1(n9085), .A2(n9084), .ZN(n13707) );
  NAND2_X1 U7383 ( .A1(n7802), .A2(n7801), .ZN(n14465) );
  NAND2_X1 U7384 ( .A1(n7810), .A2(n7809), .ZN(n7812) );
  OR2_X1 U7385 ( .A1(n14553), .A2(n14554), .ZN(n6902) );
  AOI21_X1 U7386 ( .B1(n7632), .B2(n7551), .A(n7550), .ZN(n7777) );
  NAND2_X1 U7387 ( .A1(n9015), .A2(n9014), .ZN(n12115) );
  NAND2_X1 U7388 ( .A1(n11420), .A2(n6584), .ZN(n11419) );
  NAND2_X1 U7389 ( .A1(n9001), .A2(n9000), .ZN(n14931) );
  AND2_X1 U7390 ( .A1(n11341), .A2(n10223), .ZN(n11420) );
  NAND2_X1 U7391 ( .A1(n8984), .A2(n8983), .ZN(n11902) );
  NAND2_X1 U7392 ( .A1(n7762), .A2(n7761), .ZN(n12319) );
  NAND2_X1 U7393 ( .A1(n14547), .A2(n14548), .ZN(n14544) );
  NAND2_X1 U7394 ( .A1(n6647), .A2(n6646), .ZN(n14546) );
  NAND2_X1 U7395 ( .A1(n6709), .A2(n11523), .ZN(n11524) );
  NAND2_X1 U7396 ( .A1(n7756), .A2(n7755), .ZN(n12200) );
  NAND2_X1 U7397 ( .A1(n8971), .A2(n8970), .ZN(n11620) );
  NAND2_X1 U7398 ( .A1(n7749), .A2(n7748), .ZN(n12153) );
  NAND2_X1 U7399 ( .A1(n6896), .A2(n6550), .ZN(n8519) );
  NAND2_X1 U7400 ( .A1(n8958), .A2(n8957), .ZN(n11701) );
  NAND2_X1 U7401 ( .A1(n7751), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U7402 ( .A1(n8942), .A2(n8941), .ZN(n11396) );
  XNOR2_X1 U7403 ( .A(n8517), .B(n8518), .ZN(n15383) );
  NAND2_X1 U7404 ( .A1(n7743), .A2(n7532), .ZN(n7751) );
  NAND2_X1 U7405 ( .A1(n10725), .A2(n10674), .ZN(n10698) );
  NOR2_X1 U7406 ( .A1(n8910), .A2(n7124), .ZN(n7123) );
  NAND2_X1 U7407 ( .A1(n8914), .A2(n8913), .ZN(n11183) );
  INV_X2 U7408 ( .A(n6481), .ZN(n8368) );
  AND2_X1 U7409 ( .A1(n10112), .A2(n10111), .ZN(n11024) );
  OAI211_X1 U7410 ( .C1(n8875), .C2(n13286), .A(n8895), .B(n8894), .ZN(n11268)
         );
  OAI211_X2 U7411 ( .C1(n7813), .C2(n10341), .A(n7690), .B(n7689), .ZN(n13916)
         );
  AND2_X1 U7412 ( .A1(n7709), .A2(n7708), .ZN(n10367) );
  AND3_X2 U7413 ( .A1(n7049), .A2(n7048), .A3(n7047), .ZN(n11704) );
  NAND4_X1 U7414 ( .A1(n8909), .A2(n8908), .A3(n8907), .A4(n8906), .ZN(n13266)
         );
  NAND2_X1 U7415 ( .A1(n8094), .A2(n8093), .ZN(n14384) );
  NAND2_X1 U7416 ( .A1(n6485), .A2(n14172), .ZN(n10846) );
  OR2_X1 U7417 ( .A1(n15376), .A2(n15377), .ZN(n6897) );
  INV_X1 U7418 ( .A(n7672), .ZN(n7813) );
  INV_X2 U7419 ( .A(n9140), .ZN(n9468) );
  NAND2_X1 U7420 ( .A1(n8166), .A2(n12379), .ZN(n10850) );
  AND2_X1 U7421 ( .A1(n9605), .A2(n13121), .ZN(n9695) );
  AND2_X1 U7422 ( .A1(n10512), .A2(n10344), .ZN(n7672) );
  OR2_X1 U7423 ( .A1(n8364), .A2(n8194), .ZN(n10887) );
  AND2_X1 U7424 ( .A1(n7841), .A2(n14513), .ZN(n7853) );
  NAND2_X1 U7425 ( .A1(n6876), .A2(n6873), .ZN(n10181) );
  INV_X4 U7426 ( .A(n10907), .ZN(n12823) );
  NAND2_X1 U7427 ( .A1(n12579), .A2(n8850), .ZN(n8869) );
  INV_X1 U7428 ( .A(n13768), .ZN(n8850) );
  NAND2_X1 U7429 ( .A1(n8800), .A2(n8799), .ZN(n8802) );
  XNOR2_X1 U7430 ( .A(n9601), .B(n13115), .ZN(n12578) );
  CLKBUF_X1 U7431 ( .A(n9216), .Z(n9529) );
  AND2_X1 U7432 ( .A1(n8165), .A2(n8159), .ZN(n12379) );
  XNOR2_X1 U7434 ( .A(n7835), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7840) );
  MUX2_X1 U7435 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10199), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n10201) );
  OAI21_X1 U7436 ( .B1(n10345), .B2(n6711), .A(n6710), .ZN(n7516) );
  CLKBUF_X1 U7437 ( .A(n9257), .Z(n9258) );
  NAND2_X2 U7438 ( .A1(n9592), .A2(P1_U3086), .ZN(n14527) );
  NAND2_X1 U7439 ( .A1(n9595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U7440 ( .A1(n7207), .A2(SI_5_), .ZN(n7518) );
  OR2_X1 U7441 ( .A1(n10193), .A2(n9589), .ZN(n9591) );
  NAND2_X1 U7442 ( .A1(n8818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8817) );
  AND2_X1 U7443 ( .A1(n8155), .A2(n6595), .ZN(n14506) );
  NAND2_X1 U7444 ( .A1(n8450), .A2(n6664), .ZN(n8451) );
  INV_X4 U7445 ( .A(n10344), .ZN(n9592) );
  NOR2_X2 U7446 ( .A1(n7787), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7797) );
  AND2_X1 U7447 ( .A1(n10195), .A2(n7422), .ZN(n10193) );
  OR2_X1 U7448 ( .A1(n8816), .A2(n8741), .ZN(n6918) );
  AND2_X1 U7449 ( .A1(n9622), .A2(n6542), .ZN(n6850) );
  NOR2_X1 U7450 ( .A1(n8747), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7233) );
  INV_X1 U7451 ( .A(n7668), .ZN(n6484) );
  NAND2_X1 U7452 ( .A1(n6506), .A2(n7089), .ZN(n7787) );
  AND2_X1 U7453 ( .A1(n9580), .A2(n6975), .ZN(n10188) );
  NAND2_X2 U7454 ( .A1(n6714), .A2(n6713), .ZN(n7515) );
  NOR2_X1 U7455 ( .A1(n9621), .A2(n6973), .ZN(n6970) );
  AND2_X1 U7456 ( .A1(n8911), .A2(n8770), .ZN(n8787) );
  AND2_X1 U7457 ( .A1(n8770), .A2(n8735), .ZN(n8736) );
  AND2_X1 U7458 ( .A1(n7350), .A2(n7598), .ZN(n7349) );
  NAND2_X1 U7459 ( .A1(n7598), .A2(n7463), .ZN(n7462) );
  AND2_X2 U7460 ( .A1(n6946), .A2(n6945), .ZN(n9684) );
  AND3_X1 U7461 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8770) );
  AND2_X1 U7462 ( .A1(n8738), .A2(n8752), .ZN(n8745) );
  NOR2_X1 U7463 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7593) );
  INV_X1 U7464 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8997) );
  NOR2_X1 U7465 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8728) );
  INV_X1 U7466 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8168) );
  INV_X4 U7467 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7468 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7798) );
  INV_X4 U7469 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7470 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6945) );
  INV_X1 U7471 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9727) );
  INV_X1 U7472 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9944) );
  INV_X1 U7473 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6946) );
  INV_X1 U7474 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7638) );
  INV_X1 U7475 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8793) );
  INV_X1 U7476 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7583) );
  INV_X1 U7477 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9582) );
  NOR2_X1 U7478 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n9581) );
  NOR2_X1 U7479 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n6658) );
  NOR2_X1 U7480 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n6657) );
  INV_X1 U7481 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9796) );
  INV_X1 U7482 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9927) );
  NOR2_X1 U7483 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9577) );
  INV_X4 U7484 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7485 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8879) );
  AND2_X2 U7486 ( .A1(n15278), .A2(n15272), .ZN(n15276) );
  NAND2_X1 U7487 ( .A1(n10910), .A2(n11015), .ZN(n10994) );
  NAND2_X1 U7488 ( .A1(n13180), .A2(n6489), .ZN(n6486) );
  AND2_X2 U7489 ( .A1(n6486), .A2(n6487), .ZN(n13222) );
  OR2_X1 U7490 ( .A1(n6488), .A2(n13183), .ZN(n6487) );
  INV_X1 U7491 ( .A(n12517), .ZN(n6488) );
  AND2_X1 U7492 ( .A1(n13182), .A2(n12517), .ZN(n6489) );
  NAND2_X1 U7493 ( .A1(n13171), .A2(n6493), .ZN(n6490) );
  OR2_X1 U7494 ( .A1(n6492), .A2(n6603), .ZN(n6491) );
  INV_X1 U7495 ( .A(n12558), .ZN(n6492) );
  AND2_X1 U7496 ( .A1(n13173), .A2(n12558), .ZN(n6493) );
  NAND2_X1 U7497 ( .A1(n8820), .A2(n13768), .ZN(n9453) );
  CLKBUF_X1 U7498 ( .A(n11714), .Z(n6494) );
  NAND2_X1 U7499 ( .A1(n14197), .A2(n7323), .ZN(n6495) );
  CLKBUF_X1 U7500 ( .A(n11680), .Z(n6496) );
  NAND2_X1 U7501 ( .A1(n8111), .A2(n8110), .ZN(n11714) );
  NAND2_X1 U7502 ( .A1(n14197), .A2(n7323), .ZN(n12438) );
  NAND2_X1 U7503 ( .A1(n11049), .A2(n8103), .ZN(n11680) );
  OAI21_X2 U7504 ( .B1(n11783), .B2(n8994), .A(n8995), .ZN(n11919) );
  NOR2_X2 U7505 ( .A1(n13581), .A2(n13702), .ZN(n6933) );
  AND2_X1 U7506 ( .A1(n12443), .A2(n7840), .ZN(n6497) );
  AOI21_X2 U7507 ( .B1(n14585), .B2(n12805), .A(n12806), .ZN(n12817) );
  NAND2_X1 U7508 ( .A1(n6714), .A2(n6713), .ZN(n6498) );
  INV_X1 U7509 ( .A(n10344), .ZN(n10345) );
  OR2_X1 U7510 ( .A1(n9217), .A2(n9216), .ZN(n11208) );
  NOR2_X1 U7511 ( .A1(n13379), .A2(n9217), .ZN(n9276) );
  BUF_X4 U7512 ( .A(n8870), .Z(n6499) );
  NAND2_X1 U7513 ( .A1(n8850), .A2(n8820), .ZN(n8870) );
  XNOR2_X1 U7514 ( .A(n9588), .B(n9587), .ZN(n10206) );
  AND4_X1 U7515 ( .A1(n7584), .A2(n7638), .A3(n7590), .A4(n7591), .ZN(n7089)
         );
  OAI222_X1 U7516 ( .A1(n14527), .A2(n12445), .B1(P1_U3086), .B2(n12443), .C1(
        n14521), .C2(n12580), .ZN(P1_U3325) );
  AOI21_X2 U7517 ( .B1(n12085), .B2(n12084), .A(n7476), .ZN(n12071) );
  OAI21_X2 U7518 ( .B1(n11844), .B2(n7135), .A(n7131), .ZN(n12085) );
  INV_X2 U7519 ( .A(n11600), .ZN(n11596) );
  AND2_X1 U7520 ( .A1(n10855), .A2(n10892), .ZN(n10893) );
  NAND4_X4 U7521 ( .A1(n7849), .A2(n7848), .A3(n7847), .A4(n7846), .ZN(n8099)
         );
  BUF_X8 U7522 ( .A(n9482), .Z(n6502) );
  NAND2_X1 U7523 ( .A1(n9275), .A2(n9276), .ZN(n9482) );
  NAND2_X1 U7524 ( .A1(n8116), .A2(n8115), .ZN(n11976) );
  AOI21_X2 U7525 ( .B1(n11374), .B2(n11373), .A(n11372), .ZN(n11376) );
  INV_X4 U7526 ( .A(n6483), .ZN(n12562) );
  NAND2_X1 U7527 ( .A1(n8120), .A2(n8119), .ZN(n12119) );
  NAND2_X2 U7528 ( .A1(n8128), .A2(n7314), .ZN(n14323) );
  NAND2_X2 U7529 ( .A1(n14378), .A2(n8123), .ZN(n8125) );
  NAND2_X2 U7530 ( .A1(n12231), .A2(n8122), .ZN(n14378) );
  AND2_X1 U7531 ( .A1(n8100), .A2(n11704), .ZN(n8201) );
  NAND2_X1 U7532 ( .A1(n8099), .A2(n10873), .ZN(n11036) );
  AND2_X1 U7533 ( .A1(n7841), .A2(n7840), .ZN(n7867) );
  XNOR2_X2 U7534 ( .A(n7599), .B(n7831), .ZN(n7828) );
  OAI222_X1 U7535 ( .A1(P3_U3151), .A2(n10959), .B1(n13125), .B2(n7504), .C1(
        n13123), .C2(n10399), .ZN(P3_U3294) );
  INV_X1 U7536 ( .A(n13112), .ZN(n13123) );
  NAND2_X1 U7537 ( .A1(n6752), .A2(n6545), .ZN(n6967) );
  NAND2_X1 U7538 ( .A1(n13453), .A2(n9179), .ZN(n7128) );
  AOI21_X1 U7539 ( .B1(n7015), .B2(n7018), .A(n6586), .ZN(n7014) );
  INV_X1 U7540 ( .A(n10155), .ZN(n7018) );
  AND4_X1 U7541 ( .A1(n9579), .A2(n10107), .A3(n9944), .A4(n9927), .ZN(n9580)
         );
  INV_X1 U7542 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8739) );
  AOI21_X1 U7543 ( .B1(n7189), .B2(n7191), .A(n7186), .ZN(n7185) );
  INV_X1 U7544 ( .A(n7557), .ZN(n7186) );
  NAND2_X1 U7545 ( .A1(n12483), .A2(n12636), .ZN(n12638) );
  AND2_X1 U7546 ( .A1(n11445), .A2(n11075), .ZN(n10939) );
  NAND2_X1 U7547 ( .A1(n6967), .A2(n6635), .ZN(n6962) );
  AOI21_X1 U7548 ( .B1(n7002), .B2(n7001), .A(n10150), .ZN(n7000) );
  INV_X1 U7549 ( .A(n6532), .ZN(n7001) );
  AOI21_X1 U7550 ( .B1(n7079), .B2(n6766), .A(n6644), .ZN(n6765) );
  INV_X1 U7551 ( .A(n7083), .ZN(n6766) );
  AOI21_X1 U7552 ( .B1(n13132), .B2(n12561), .A(n7244), .ZN(n7252) );
  INV_X1 U7553 ( .A(n12567), .ZN(n7244) );
  INV_X1 U7554 ( .A(n13733), .ZN(n9255) );
  NOR2_X1 U7555 ( .A1(n9190), .A2(n7127), .ZN(n7126) );
  INV_X1 U7556 ( .A(n9180), .ZN(n7127) );
  INV_X1 U7557 ( .A(n8356), .ZN(n8086) );
  AOI21_X1 U7558 ( .B1(n7296), .B2(n7295), .A(n6563), .ZN(n7294) );
  INV_X1 U7559 ( .A(n7300), .ZN(n7295) );
  AND2_X1 U7560 ( .A1(n8401), .A2(n7472), .ZN(n7471) );
  NAND2_X1 U7561 ( .A1(n7474), .A2(n7473), .ZN(n7472) );
  NOR2_X1 U7562 ( .A1(n8271), .A2(n7475), .ZN(n7474) );
  AOI21_X1 U7563 ( .B1(n6891), .B2(n12143), .A(n6890), .ZN(n6889) );
  INV_X1 U7564 ( .A(n12296), .ZN(n6890) );
  AOI21_X1 U7565 ( .B1(n6885), .B2(n6888), .A(n9906), .ZN(n6884) );
  INV_X1 U7566 ( .A(n6889), .ZN(n6888) );
  INV_X1 U7567 ( .A(n9567), .ZN(n7078) );
  INV_X1 U7568 ( .A(n13530), .ZN(n7212) );
  NOR2_X1 U7569 ( .A1(n9229), .A2(n6840), .ZN(n6839) );
  INV_X1 U7570 ( .A(n9228), .ZN(n6840) );
  NAND4_X1 U7571 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8997), .ZN(n8786)
         );
  NAND2_X1 U7572 ( .A1(n6721), .A2(n8453), .ZN(n8455) );
  NAND2_X1 U7573 ( .A1(n8496), .A2(n8452), .ZN(n6721) );
  OR2_X1 U7574 ( .A1(n10574), .A2(n7354), .ZN(n7353) );
  OR2_X1 U7575 ( .A1(n14615), .A2(n11285), .ZN(n10087) );
  AND2_X1 U7576 ( .A1(n6744), .A2(n6743), .ZN(n12791) );
  NAND2_X1 U7577 ( .A1(n12801), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6743) );
  AND2_X1 U7578 ( .A1(n10140), .A2(n9985), .ZN(n10176) );
  OR2_X1 U7579 ( .A1(n12683), .A2(n12991), .ZN(n10136) );
  NAND4_X1 U7580 ( .A1(n6658), .A2(n6657), .A3(n9727), .A4(n9582), .ZN(n6974)
         );
  NOR2_X1 U7581 ( .A1(n9551), .A2(n6783), .ZN(n6782) );
  AND2_X1 U7582 ( .A1(n10383), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9551) );
  INV_X1 U7583 ( .A(n9550), .ZN(n6783) );
  NAND2_X1 U7584 ( .A1(n13223), .A2(n7266), .ZN(n13153) );
  NOR2_X1 U7585 ( .A1(n13156), .A2(n7267), .ZN(n7266) );
  INV_X1 U7586 ( .A(n12523), .ZN(n7267) );
  AOI21_X1 U7587 ( .B1(n7484), .B2(n9106), .A(n6566), .ZN(n7120) );
  OR2_X1 U7588 ( .A1(n11178), .A2(n6838), .ZN(n6835) );
  INV_X1 U7589 ( .A(n6839), .ZN(n6838) );
  INV_X1 U7590 ( .A(n11225), .ZN(n8883) );
  NAND2_X1 U7591 ( .A1(n8745), .A2(n8739), .ZN(n8740) );
  INV_X1 U7592 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U7593 ( .A1(n8338), .A2(n7452), .ZN(n7451) );
  AND3_X1 U7594 ( .A1(n8418), .A2(n14212), .A3(n12439), .ZN(n7172) );
  NAND2_X1 U7595 ( .A1(n7051), .A2(n6552), .ZN(n7050) );
  AND2_X1 U7596 ( .A1(n7054), .A2(n14212), .ZN(n7053) );
  INV_X1 U7597 ( .A(n14267), .ZN(n8135) );
  NAND2_X1 U7598 ( .A1(n8349), .A2(n8348), .ZN(n8376) );
  INV_X1 U7599 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7463) );
  INV_X1 U7600 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7598) );
  INV_X1 U7601 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7350) );
  OAI211_X1 U7602 ( .C1(n7166), .C2(n7169), .A(n6666), .B(n6640), .ZN(n7818)
         );
  INV_X1 U7603 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7595) );
  AND2_X1 U7604 ( .A1(n7571), .A2(n7170), .ZN(n7169) );
  INV_X1 U7605 ( .A(n7619), .ZN(n7170) );
  NAND2_X1 U7606 ( .A1(n7812), .A2(n6618), .ZN(n7183) );
  INV_X1 U7607 ( .A(n7633), .ZN(n7550) );
  AND2_X1 U7608 ( .A1(n7631), .A2(n7634), .ZN(n7551) );
  INV_X1 U7609 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7093) );
  AND2_X1 U7610 ( .A1(n7631), .A2(n7547), .ZN(n7643) );
  XNOR2_X1 U7611 ( .A(n7540), .B(n10401), .ZN(n7763) );
  XNOR2_X1 U7612 ( .A(n7537), .B(SI_11_), .ZN(n7757) );
  INV_X1 U7613 ( .A(n7686), .ZN(n7584) );
  INV_X1 U7614 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9546) );
  OAI21_X1 U7615 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n8474), .A(n8473), .ZN(
        n8488) );
  NAND2_X1 U7616 ( .A1(n7358), .A2(n7361), .ZN(n7356) );
  INV_X1 U7617 ( .A(n12470), .ZN(n7377) );
  NAND2_X1 U7618 ( .A1(n14605), .A2(n10104), .ZN(n10161) );
  AND4_X1 U7619 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n12475)
         );
  CLKBUF_X2 U7620 ( .A(n9696), .Z(n10098) );
  AND2_X1 U7621 ( .A1(n9602), .A2(n9605), .ZN(n9693) );
  AND2_X1 U7622 ( .A1(n12578), .A2(n13121), .ZN(n9696) );
  XNOR2_X1 U7623 ( .A(n10961), .B(n10960), .ZN(n10988) );
  OR2_X1 U7624 ( .A1(n11009), .A2(n6747), .ZN(n6746) );
  AND2_X1 U7625 ( .A1(n9684), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6747) );
  OR2_X1 U7626 ( .A1(n15233), .A2(n10967), .ZN(n11096) );
  INV_X1 U7627 ( .A(n11517), .ZN(n6938) );
  AND2_X1 U7628 ( .A1(n11824), .A2(n11823), .ZN(n12000) );
  INV_X1 U7629 ( .A(n12004), .ZN(n6943) );
  OR2_X1 U7630 ( .A1(n12760), .A2(n12785), .ZN(n6966) );
  NOR2_X1 U7631 ( .A1(n12785), .A2(n12784), .ZN(n12787) );
  AND2_X1 U7632 ( .A1(n12753), .A2(n12760), .ZN(n12784) );
  XNOR2_X1 U7633 ( .A(n13003), .B(n12700), .ZN(n12842) );
  OR2_X1 U7634 ( .A1(n10038), .A2(n10061), .ZN(n12858) );
  NAND2_X1 U7635 ( .A1(n7412), .A2(n6557), .ZN(n12850) );
  INV_X1 U7636 ( .A(n10151), .ZN(n7004) );
  AOI21_X1 U7637 ( .B1(n7410), .B2(n7408), .A(n6567), .ZN(n7407) );
  INV_X1 U7638 ( .A(n10249), .ZN(n7408) );
  NAND2_X1 U7639 ( .A1(n12919), .A2(n10249), .ZN(n7411) );
  AOI21_X1 U7640 ( .B1(n7026), .B2(n12967), .A(n7024), .ZN(n7023) );
  INV_X1 U7641 ( .A(n10140), .ZN(n7024) );
  NAND2_X1 U7642 ( .A1(n7030), .A2(n7029), .ZN(n7028) );
  INV_X1 U7643 ( .A(n12968), .ZN(n7030) );
  OR2_X1 U7644 ( .A1(n12094), .A2(n10127), .ZN(n10129) );
  INV_X1 U7645 ( .A(n10181), .ZN(n11075) );
  OR2_X1 U7646 ( .A1(n11075), .A2(n11445), .ZN(n15357) );
  NAND2_X1 U7647 ( .A1(n6765), .A2(n6763), .ZN(n6762) );
  NAND2_X1 U7648 ( .A1(n6767), .A2(n10095), .ZN(n6763) );
  AND2_X1 U7649 ( .A1(n10195), .A2(n6594), .ZN(n9599) );
  AND2_X1 U7650 ( .A1(n9944), .A2(n10107), .ZN(n6878) );
  NAND2_X1 U7651 ( .A1(n6756), .A2(n7066), .ZN(n9824) );
  AOI21_X1 U7652 ( .B1(n7068), .B2(n7070), .A(n6623), .ZN(n7066) );
  NAND2_X1 U7653 ( .A1(n9795), .A2(n7068), .ZN(n6756) );
  XNOR2_X1 U7654 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9748) );
  AOI21_X1 U7655 ( .B1(n7063), .B2(n9658), .A(n6580), .ZN(n7062) );
  NOR2_X1 U7656 ( .A1(n10823), .A2(n7257), .ZN(n7256) );
  INV_X1 U7657 ( .A(n7263), .ZN(n7257) );
  NOR2_X1 U7658 ( .A1(n12424), .A2(n10344), .ZN(n7159) );
  OAI21_X1 U7659 ( .B1(n7273), .B2(n7271), .A(n12503), .ZN(n7269) );
  OR2_X1 U7660 ( .A1(n6499), .A2(n11237), .ZN(n8859) );
  NOR2_X1 U7661 ( .A1(n15040), .A2(n13366), .ZN(n13367) );
  NAND2_X1 U7662 ( .A1(n13427), .A2(n13614), .ZN(n6687) );
  AND2_X1 U7663 ( .A1(n9178), .A2(n9177), .ZN(n13461) );
  AND2_X1 U7664 ( .A1(n13577), .A2(n9081), .ZN(n7153) );
  AND2_X1 U7665 ( .A1(n13638), .A2(n9052), .ZN(n13619) );
  OAI21_X1 U7666 ( .B1(n13629), .B2(n9237), .A(n9238), .ZN(n13611) );
  NAND2_X1 U7667 ( .A1(n14657), .A2(n7150), .ZN(n13638) );
  NOR2_X1 U7668 ( .A1(n7152), .A2(n7151), .ZN(n7150) );
  INV_X1 U7669 ( .A(n9041), .ZN(n7151) );
  INV_X2 U7670 ( .A(n13379), .ZN(n11210) );
  NAND2_X1 U7671 ( .A1(n8835), .A2(n11273), .ZN(n7162) );
  NAND2_X1 U7673 ( .A1(n13415), .A2(n6735), .ZN(n13653) );
  NAND2_X1 U7674 ( .A1(n6733), .A2(n13408), .ZN(n6735) );
  INV_X1 U7675 ( .A(n13416), .ZN(n6733) );
  INV_X1 U7676 ( .A(n8748), .ZN(n7234) );
  XNOR2_X1 U7677 ( .A(n14420), .B(n14229), .ZN(n14212) );
  NAND2_X1 U7678 ( .A1(n8142), .A2(n8141), .ZN(n7313) );
  AND2_X1 U7679 ( .A1(n7156), .A2(n7155), .ZN(n7154) );
  INV_X1 U7680 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7155) );
  AND2_X1 U7681 ( .A1(n6908), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8500) );
  INV_X1 U7682 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6908) );
  INV_X1 U7683 ( .A(n6692), .ZN(n8527) );
  OR2_X1 U7684 ( .A1(n11825), .A2(n11955), .ZN(n6751) );
  XNOR2_X1 U7685 ( .A(n12000), .B(n12015), .ZN(n11825) );
  NAND2_X1 U7686 ( .A1(n10807), .A2(n10806), .ZN(n11424) );
  INV_X1 U7687 ( .A(n7247), .ZN(n7246) );
  OAI211_X1 U7688 ( .C1(n12569), .C2(n7250), .A(n7248), .B(n12568), .ZN(n7247)
         );
  NAND2_X1 U7689 ( .A1(n13132), .A2(n12561), .ZN(n7250) );
  NOR2_X1 U7690 ( .A1(n13375), .A2(n6698), .ZN(n6697) );
  OR2_X1 U7691 ( .A1(n15027), .A2(n13379), .ZN(n6698) );
  NAND2_X1 U7692 ( .A1(n13409), .A2(n13408), .ZN(n13411) );
  INV_X1 U7693 ( .A(n13409), .ZN(n7219) );
  NAND2_X1 U7694 ( .A1(n8072), .A2(n8071), .ZN(n14069) );
  NAND2_X1 U7695 ( .A1(n14733), .A2(n14997), .ZN(n14732) );
  AOI21_X1 U7696 ( .B1(n7441), .B2(n7439), .A(n7438), .ZN(n7437) );
  OR2_X1 U7697 ( .A1(n9319), .A2(n9320), .ZN(n7305) );
  NOR2_X1 U7698 ( .A1(n7308), .A2(n7307), .ZN(n7306) );
  INV_X1 U7699 ( .A(n9349), .ZN(n7344) );
  AND2_X1 U7700 ( .A1(n7468), .A2(n8278), .ZN(n7467) );
  NAND2_X1 U7701 ( .A1(n7471), .A2(n7469), .ZN(n7468) );
  INV_X1 U7702 ( .A(n7471), .ZN(n7470) );
  AOI21_X1 U7703 ( .B1(n9709), .B2(n6866), .A(n6865), .ZN(n6864) );
  INV_X1 U7704 ( .A(n9712), .ZN(n6865) );
  INV_X1 U7705 ( .A(n9714), .ZN(n6862) );
  INV_X1 U7706 ( .A(n10111), .ZN(n6863) );
  NAND2_X1 U7707 ( .A1(n8288), .A2(n8399), .ZN(n7458) );
  NOR2_X1 U7708 ( .A1(n7338), .A2(n7336), .ZN(n7335) );
  NOR2_X1 U7709 ( .A1(n9391), .A2(n9390), .ZN(n7336) );
  NOR2_X1 U7710 ( .A1(n6872), .A2(n6871), .ZN(n6870) );
  NAND2_X1 U7711 ( .A1(n11808), .A2(n6537), .ZN(n6871) );
  NOR2_X1 U7712 ( .A1(n9740), .A2(n10294), .ZN(n6872) );
  AND2_X1 U7713 ( .A1(n6894), .A2(n6892), .ZN(n6891) );
  INV_X1 U7714 ( .A(n9887), .ZN(n6894) );
  NAND2_X1 U7715 ( .A1(n6895), .A2(n6893), .ZN(n6892) );
  INV_X1 U7716 ( .A(n9419), .ZN(n7322) );
  INV_X1 U7717 ( .A(n8310), .ZN(n6683) );
  AOI21_X1 U7718 ( .B1(n6884), .B2(n6882), .A(n9908), .ZN(n6881) );
  INV_X1 U7719 ( .A(n6885), .ZN(n6882) );
  INV_X1 U7720 ( .A(n6884), .ZN(n6883) );
  AND2_X1 U7721 ( .A1(n8315), .A2(n8314), .ZN(n7445) );
  OR2_X1 U7722 ( .A1(n8315), .A2(n8314), .ZN(n7444) );
  INV_X1 U7723 ( .A(n8313), .ZN(n7448) );
  INV_X1 U7724 ( .A(n9432), .ZN(n7331) );
  NAND2_X1 U7725 ( .A1(n7327), .A2(n9434), .ZN(n7330) );
  OR2_X1 U7726 ( .A1(n8362), .A2(n11743), .ZN(n8196) );
  NAND2_X1 U7727 ( .A1(n8327), .A2(n7429), .ZN(n7428) );
  NOR2_X1 U7728 ( .A1(n7429), .A2(n8327), .ZN(n7430) );
  NOR2_X1 U7729 ( .A1(n6560), .A2(n7016), .ZN(n7015) );
  NAND2_X1 U7730 ( .A1(n6660), .A2(n10159), .ZN(n7016) );
  INV_X1 U7731 ( .A(n10154), .ZN(n7017) );
  NOR2_X1 U7732 ( .A1(n7072), .A2(n10152), .ZN(n7071) );
  NAND2_X1 U7733 ( .A1(n10178), .A2(n12868), .ZN(n7072) );
  NAND2_X1 U7734 ( .A1(n13071), .A2(n10252), .ZN(n10253) );
  NAND2_X1 U7735 ( .A1(n12722), .A2(n15309), .ZN(n9713) );
  INV_X1 U7736 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U7737 ( .A1(n9443), .A2(n6543), .ZN(n7290) );
  NAND2_X1 U7738 ( .A1(n7211), .A2(n7218), .ZN(n7210) );
  INV_X1 U7739 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8843) );
  INV_X1 U7740 ( .A(n7924), .ZN(n7036) );
  INV_X1 U7741 ( .A(n7192), .ZN(n7191) );
  NAND2_X1 U7742 ( .A1(n7552), .A2(n10797), .ZN(n7192) );
  INV_X1 U7743 ( .A(n7650), .ZN(n7198) );
  INV_X1 U7744 ( .A(n12171), .ZN(n7360) );
  NAND2_X1 U7745 ( .A1(n10211), .A2(n15326), .ZN(n10579) );
  NAND2_X1 U7746 ( .A1(n6853), .A2(n6852), .ZN(n10044) );
  AND2_X1 U7747 ( .A1(n10016), .A2(n10017), .ZN(n6852) );
  INV_X1 U7748 ( .A(n10970), .ZN(n6741) );
  NAND2_X1 U7749 ( .A1(n6738), .A2(n11099), .ZN(n6737) );
  XOR2_X1 U7750 ( .A(n12007), .B(n12006), .Z(n11833) );
  OR2_X1 U7751 ( .A1(n10300), .A2(n12837), .ZN(n10155) );
  NAND2_X1 U7752 ( .A1(n12479), .A2(n12865), .ZN(n7007) );
  INV_X1 U7753 ( .A(n10141), .ZN(n7021) );
  OR2_X1 U7754 ( .A1(n12625), .A2(n12944), .ZN(n10142) );
  INV_X1 U7755 ( .A(n11642), .ZN(n10226) );
  AND2_X1 U7756 ( .A1(n10114), .A2(n10113), .ZN(n6983) );
  NAND2_X1 U7757 ( .A1(n9652), .A2(n15304), .ZN(n10112) );
  NAND2_X1 U7758 ( .A1(n9713), .A2(n10110), .ZN(n10214) );
  OAI21_X1 U7759 ( .B1(n9611), .B2(n9610), .A(n7086), .ZN(n7085) );
  NAND2_X1 U7760 ( .A1(n12190), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7086) );
  NOR2_X1 U7761 ( .A1(n9988), .A2(n6788), .ZN(n6787) );
  INV_X1 U7762 ( .A(n9576), .ZN(n6788) );
  AOI21_X1 U7763 ( .B1(n7076), .B2(n7078), .A(n6624), .ZN(n7074) );
  NOR2_X1 U7764 ( .A1(n7077), .A2(n6774), .ZN(n6772) );
  NAND2_X1 U7765 ( .A1(n9563), .A2(n9562), .ZN(n9564) );
  NAND2_X1 U7766 ( .A1(n9824), .A2(n9822), .ZN(n9563) );
  INV_X1 U7767 ( .A(n9748), .ZN(n6778) );
  OR2_X1 U7768 ( .A1(n6942), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n9660) );
  XNOR2_X1 U7769 ( .A(n14656), .B(n12518), .ZN(n12500) );
  NAND2_X1 U7770 ( .A1(n12522), .A2(n12521), .ZN(n13223) );
  NAND2_X1 U7771 ( .A1(n6585), .A2(n7223), .ZN(n7221) );
  OR2_X1 U7772 ( .A1(n13433), .A2(n9254), .ZN(n7220) );
  NOR2_X1 U7773 ( .A1(n6568), .A2(n6828), .ZN(n6827) );
  INV_X1 U7774 ( .A(n9249), .ZN(n6828) );
  NOR2_X1 U7775 ( .A1(n13499), .A2(n7143), .ZN(n7142) );
  INV_X1 U7776 ( .A(n9139), .ZN(n7143) );
  NAND2_X1 U7777 ( .A1(n13671), .A2(n13460), .ZN(n9252) );
  AND2_X1 U7778 ( .A1(n9252), .A2(n7236), .ZN(n7235) );
  AND2_X1 U7779 ( .A1(n9153), .A2(n9251), .ZN(n7236) );
  AND2_X1 U7780 ( .A1(n8809), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9016) );
  INV_X1 U7781 ( .A(n9234), .ZN(n7228) );
  AND2_X1 U7782 ( .A1(n11899), .A2(n6928), .ZN(n6929) );
  INV_X1 U7783 ( .A(n6931), .ZN(n6928) );
  AOI21_X1 U7784 ( .B1(n6839), .B2(n6837), .A(n6562), .ZN(n6836) );
  OR2_X1 U7785 ( .A1(n11314), .A2(n11332), .ZN(n11313) );
  OAI21_X1 U7786 ( .B1(n7227), .B2(n7226), .A(n7224), .ZN(n11178) );
  INV_X1 U7787 ( .A(n9227), .ZN(n7225) );
  OAI22_X1 U7788 ( .A1(n12055), .A2(n7133), .B1(n12053), .B2(n12054), .ZN(
        n7132) );
  NAND2_X1 U7789 ( .A1(n7134), .A2(n7137), .ZN(n7133) );
  INV_X1 U7790 ( .A(n7138), .ZN(n7134) );
  NAND2_X1 U7791 ( .A1(n14001), .A2(n13998), .ZN(n13887) );
  NAND2_X1 U7792 ( .A1(n6680), .A2(n13880), .ZN(n13876) );
  INV_X1 U7793 ( .A(n13967), .ZN(n6680) );
  INV_X1 U7794 ( .A(n8419), .ZN(n8420) );
  XNOR2_X1 U7795 ( .A(n8424), .B(n14179), .ZN(n8430) );
  NAND2_X1 U7796 ( .A1(n12436), .A2(n6799), .ZN(n6798) );
  AND2_X1 U7797 ( .A1(n14237), .A2(n8041), .ZN(n7054) );
  XNOR2_X1 U7798 ( .A(n14688), .B(n14074), .ZN(n8401) );
  AND2_X1 U7799 ( .A1(n6811), .A2(n14556), .ZN(n6812) );
  INV_X1 U7800 ( .A(n6814), .ZN(n6811) );
  INV_X1 U7801 ( .A(n11868), .ZN(n6813) );
  INV_X1 U7802 ( .A(n8201), .ZN(n8098) );
  NAND2_X1 U7803 ( .A1(n8040), .A2(n14245), .ZN(n14249) );
  NOR2_X1 U7804 ( .A1(n8123), .A2(n7041), .ZN(n7038) );
  OAI21_X1 U7805 ( .B1(n7610), .B2(n7203), .A(n7201), .ZN(n8349) );
  INV_X1 U7806 ( .A(n7202), .ZN(n7201) );
  OAI21_X1 U7807 ( .B1(n7609), .B2(n7203), .A(n7581), .ZN(n7202) );
  NAND2_X1 U7808 ( .A1(n7181), .A2(SI_22_), .ZN(n7567) );
  INV_X1 U7809 ( .A(n7803), .ZN(n7560) );
  AND2_X1 U7810 ( .A1(n7592), .A2(n7798), .ZN(n7156) );
  NAND2_X1 U7811 ( .A1(n7188), .A2(n7192), .ZN(n7781) );
  NAND2_X1 U7812 ( .A1(n7777), .A2(n7193), .ZN(n7188) );
  AOI21_X1 U7813 ( .B1(n7176), .B2(n7178), .A(n6578), .ZN(n7173) );
  NAND2_X1 U7814 ( .A1(n7515), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U7815 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6665), .ZN(n6664) );
  INV_X1 U7816 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6665) );
  INV_X1 U7817 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n8454) );
  XNOR2_X1 U7818 ( .A(n8457), .B(n6899), .ZN(n8507) );
  INV_X1 U7819 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U7820 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15268), .A(n8467), .ZN(
        n8491) );
  NAND2_X1 U7821 ( .A1(n15159), .A2(n15158), .ZN(n15157) );
  INV_X1 U7822 ( .A(n12615), .ZN(n7381) );
  AND2_X1 U7823 ( .A1(n11939), .A2(n11938), .ZN(n11940) );
  AND2_X1 U7824 ( .A1(n12400), .A2(n7372), .ZN(n7371) );
  OR2_X1 U7825 ( .A1(n12366), .A2(n7373), .ZN(n7372) );
  INV_X1 U7826 ( .A(n12369), .ZN(n7373) );
  NAND2_X1 U7827 ( .A1(n12478), .A2(n12654), .ZN(n12634) );
  AND2_X1 U7828 ( .A1(n11161), .A2(n12721), .ZN(n11162) );
  NAND2_X1 U7829 ( .A1(n7389), .A2(n7388), .ZN(n7392) );
  INV_X1 U7830 ( .A(n15174), .ZN(n7388) );
  INV_X1 U7831 ( .A(n15173), .ZN(n7389) );
  INV_X1 U7832 ( .A(n11815), .ZN(n7383) );
  NAND2_X1 U7833 ( .A1(n7385), .A2(n12716), .ZN(n7384) );
  INV_X1 U7834 ( .A(n11813), .ZN(n7385) );
  AND2_X1 U7835 ( .A1(n12606), .A2(n7366), .ZN(n7365) );
  OR2_X1 U7836 ( .A1(n12680), .A2(n7367), .ZN(n7366) );
  INV_X1 U7837 ( .A(n12461), .ZN(n7367) );
  NAND2_X1 U7838 ( .A1(n7376), .A2(n12933), .ZN(n7375) );
  NAND2_X1 U7839 ( .A1(n12471), .A2(n12470), .ZN(n7379) );
  AND2_X1 U7840 ( .A1(n9978), .A2(n9977), .ZN(n9992) );
  AND3_X1 U7841 ( .A1(n9642), .A2(n9641), .A3(n9640), .ZN(n11801) );
  AND2_X1 U7842 ( .A1(n10182), .A2(n10575), .ZN(n10183) );
  AND2_X1 U7843 ( .A1(n9602), .A2(n12578), .ZN(n9694) );
  AND2_X1 U7844 ( .A1(n6748), .A2(n6746), .ZN(n10986) );
  NOR2_X1 U7845 ( .A1(n10986), .A2(n6745), .ZN(n10963) );
  AND2_X1 U7846 ( .A1(n11001), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U7847 ( .A1(n15240), .A2(n6536), .ZN(n6753) );
  NAND2_X1 U7848 ( .A1(n15240), .A2(n6755), .ZN(n6754) );
  NOR2_X1 U7849 ( .A1(n11509), .A2(n11510), .ZN(n15260) );
  NOR2_X1 U7850 ( .A1(n15271), .A2(n15270), .ZN(n15269) );
  OR2_X1 U7851 ( .A1(n14577), .A2(n14576), .ZN(n6744) );
  INV_X1 U7852 ( .A(n14594), .ZN(n6742) );
  OR2_X1 U7853 ( .A1(n12842), .A2(n12836), .ZN(n10254) );
  NAND2_X1 U7854 ( .A1(n6999), .A2(n6998), .ZN(n12851) );
  AOI21_X1 U7855 ( .B1(n7000), .B2(n7003), .A(n10152), .ZN(n6998) );
  AND4_X1 U7856 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n12866) );
  NAND2_X1 U7857 ( .A1(n12876), .A2(n7007), .ZN(n7006) );
  OR2_X1 U7858 ( .A1(n12898), .A2(n12475), .ZN(n7497) );
  INV_X1 U7859 ( .A(n7410), .ZN(n7409) );
  AND2_X1 U7860 ( .A1(n12907), .A2(n6535), .ZN(n7410) );
  NAND2_X1 U7861 ( .A1(n12929), .A2(n10248), .ZN(n12919) );
  NAND2_X1 U7862 ( .A1(n7419), .A2(n7417), .ZN(n12929) );
  NOR2_X1 U7863 ( .A1(n12936), .A2(n7418), .ZN(n7417) );
  INV_X1 U7864 ( .A(n10247), .ZN(n7418) );
  NAND2_X1 U7865 ( .A1(n12942), .A2(n12951), .ZN(n7419) );
  INV_X1 U7866 ( .A(n10139), .ZN(n7027) );
  INV_X1 U7867 ( .A(n10176), .ZN(n12951) );
  OR2_X1 U7868 ( .A1(n12981), .A2(n10243), .ZN(n10137) );
  AOI21_X1 U7869 ( .B1(n7401), .B2(n7403), .A(n6620), .ZN(n7398) );
  AND2_X1 U7870 ( .A1(n10133), .A2(n10134), .ZN(n12361) );
  CLKBUF_X1 U7871 ( .A(n12357), .Z(n12358) );
  NOR2_X1 U7872 ( .A1(n10131), .A2(n9851), .ZN(n6996) );
  AND2_X1 U7873 ( .A1(n6617), .A2(n10235), .ZN(n7421) );
  AOI21_X1 U7874 ( .B1(n11991), .B2(n6980), .A(n9836), .ZN(n6979) );
  NOR2_X1 U7875 ( .A1(n6981), .A2(n6978), .ZN(n6977) );
  AOI21_X1 U7876 ( .B1(n6988), .B2(n6990), .A(n6559), .ZN(n6987) );
  NAND2_X1 U7877 ( .A1(n11638), .A2(n11642), .ZN(n11637) );
  AND2_X1 U7878 ( .A1(n10119), .A2(n9786), .ZN(n11642) );
  NAND2_X1 U7879 ( .A1(n10259), .A2(n10308), .ZN(n15317) );
  AND2_X1 U7880 ( .A1(n10273), .A2(n10272), .ZN(n12912) );
  INV_X1 U7881 ( .A(n15317), .ZN(n15308) );
  AND2_X1 U7882 ( .A1(n10937), .A2(n15325), .ZN(n10799) );
  AND2_X1 U7883 ( .A1(n10306), .A2(n10291), .ZN(n10807) );
  NAND2_X1 U7884 ( .A1(n10035), .A2(n10034), .ZN(n12857) );
  OR2_X1 U7885 ( .A1(n6480), .A2(n12447), .ZN(n10034) );
  NAND2_X1 U7886 ( .A1(n9594), .A2(n9593), .ZN(n13019) );
  NAND2_X1 U7887 ( .A1(n9991), .A2(n9990), .ZN(n12675) );
  INV_X1 U7888 ( .A(n15357), .ZN(n15325) );
  NAND2_X1 U7889 ( .A1(n10260), .A2(n10939), .ZN(n15303) );
  AND2_X1 U7890 ( .A1(n10565), .A2(n10573), .ZN(n10937) );
  AND2_X1 U7891 ( .A1(n6765), .A2(n10095), .ZN(n6759) );
  INV_X1 U7892 ( .A(n10091), .ZN(n7080) );
  INV_X1 U7893 ( .A(n7424), .ZN(n7422) );
  AND2_X1 U7894 ( .A1(n14526), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U7895 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7396) );
  NAND2_X1 U7896 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n12589), .ZN(n9576) );
  NAND2_X1 U7897 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n6877) );
  XNOR2_X1 U7898 ( .A(n9573), .B(n11748), .ZN(n9960) );
  NAND2_X1 U7899 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U7900 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n11259), .ZN(n9569) );
  NAND2_X1 U7901 ( .A1(n6773), .A2(n9565), .ZN(n9854) );
  NAND2_X1 U7902 ( .A1(n9837), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6773) );
  XNOR2_X1 U7903 ( .A(n9564), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U7904 ( .A1(n9558), .A2(n9557), .ZN(n9795) );
  INV_X1 U7905 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9556) );
  OR2_X1 U7906 ( .A1(n9751), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9780) );
  AOI21_X1 U7907 ( .B1(n6782), .B2(n6780), .A(n6518), .ZN(n6779) );
  OR2_X1 U7908 ( .A1(n9638), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U7909 ( .A1(n9548), .A2(n9547), .ZN(n9644) );
  NAND2_X1 U7910 ( .A1(n9589), .A2(n9582), .ZN(n6940) );
  NAND2_X1 U7911 ( .A1(n11066), .A2(n11065), .ZN(n7263) );
  NAND2_X1 U7912 ( .A1(n11067), .A2(n10876), .ZN(n7260) );
  NAND2_X1 U7913 ( .A1(n7260), .A2(n7263), .ZN(n7259) );
  NAND2_X1 U7914 ( .A1(n6663), .A2(n10819), .ZN(n7255) );
  NAND2_X1 U7915 ( .A1(n8812), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9110) );
  OR2_X1 U7916 ( .A1(n9110), .A2(n9109), .ZN(n9118) );
  AND2_X1 U7917 ( .A1(n10668), .A2(n12548), .ZN(n10671) );
  INV_X1 U7918 ( .A(n6499), .ZN(n9183) );
  NAND2_X1 U7919 ( .A1(n13341), .A2(n6701), .ZN(n13360) );
  NOR2_X1 U7920 ( .A1(n6631), .A2(n6702), .ZN(n6701) );
  NOR2_X1 U7921 ( .A1(n13368), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U7922 ( .A1(n7223), .A2(n9504), .ZN(n13426) );
  NAND2_X1 U7923 ( .A1(n13469), .A2(n13451), .ZN(n13446) );
  XNOR2_X1 U7924 ( .A(n13739), .B(n13481), .ZN(n13458) );
  NAND2_X1 U7925 ( .A1(n13519), .A2(n13518), .ZN(n13517) );
  NOR2_X1 U7926 ( .A1(n13550), .A2(n13541), .ZN(n13540) );
  AOI21_X1 U7927 ( .B1(n7120), .B2(n7118), .A(n6564), .ZN(n7117) );
  INV_X1 U7928 ( .A(n7120), .ZN(n7119) );
  OAI22_X1 U7929 ( .A1(n13611), .A2(n9239), .B1(n13625), .B2(n13256), .ZN(
        n13594) );
  OR2_X1 U7930 ( .A1(n13594), .A2(n13599), .ZN(n13596) );
  NOR2_X1 U7931 ( .A1(n14661), .A2(n13721), .ZN(n13632) );
  OAI21_X1 U7932 ( .B1(n14649), .B2(n9235), .A(n9236), .ZN(n13629) );
  NAND2_X1 U7933 ( .A1(n6704), .A2(n14648), .ZN(n14657) );
  NAND2_X1 U7934 ( .A1(n6818), .A2(n6817), .ZN(n11920) );
  AOI21_X1 U7935 ( .B1(n6820), .B2(n6822), .A(n6555), .ZN(n6817) );
  INV_X1 U7936 ( .A(n11484), .ZN(n11480) );
  INV_X1 U7937 ( .A(n13539), .ZN(n13612) );
  AND2_X1 U7938 ( .A1(n9262), .A2(n9258), .ZN(n13614) );
  OR2_X1 U7939 ( .A1(n9140), .A2(n10351), .ZN(n8895) );
  CLKBUF_X1 U7940 ( .A(n11260), .Z(n11261) );
  NAND2_X1 U7941 ( .A1(n9226), .A2(n9225), .ZN(n11263) );
  NAND2_X1 U7942 ( .A1(n10638), .A2(n10639), .ZN(n8868) );
  INV_X1 U7943 ( .A(n13392), .ZN(n9271) );
  NAND2_X1 U7944 ( .A1(n9073), .A2(n9072), .ZN(n13712) );
  INV_X1 U7945 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8819) );
  AND2_X1 U7946 ( .A1(n8743), .A2(n8745), .ZN(n8746) );
  NOR2_X1 U7947 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8735) );
  INV_X1 U7948 ( .A(n9126), .ZN(n7566) );
  OR2_X1 U7949 ( .A1(n7564), .A2(n7184), .ZN(n7182) );
  NAND2_X1 U7950 ( .A1(n7102), .A2(n7106), .ZN(n7101) );
  INV_X1 U7951 ( .A(n14046), .ZN(n7102) );
  XNOR2_X1 U7952 ( .A(n13787), .B(n12151), .ZN(n13929) );
  OAI21_X1 U7953 ( .B1(n11704), .B2(n13855), .A(n7087), .ZN(n10897) );
  NAND2_X1 U7954 ( .A1(n13932), .A2(n7088), .ZN(n7087) );
  INV_X1 U7955 ( .A(n7110), .ZN(n7109) );
  OAI21_X1 U7956 ( .B1(n7112), .B2(n14054), .A(n7111), .ZN(n7110) );
  OR2_X1 U7957 ( .A1(n8445), .A2(n8185), .ZN(n10867) );
  OAI21_X1 U7958 ( .B1(n8339), .B2(n6534), .A(n6681), .ZN(n8346) );
  AND2_X1 U7959 ( .A1(n7451), .A2(n8345), .ZN(n6681) );
  AND4_X1 U7960 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n13833)
         );
  NAND2_X1 U7961 ( .A1(n7867), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7849) );
  INV_X1 U7962 ( .A(n6797), .ZN(n6794) );
  INV_X1 U7963 ( .A(n8424), .ZN(n6795) );
  NOR2_X1 U7964 ( .A1(n14184), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U7965 ( .A1(n8145), .A2(n14190), .ZN(n14197) );
  NAND2_X1 U7966 ( .A1(n8149), .A2(n8147), .ZN(n12439) );
  NOR2_X1 U7967 ( .A1(n14205), .A2(n14219), .ZN(n14188) );
  NOR2_X1 U7968 ( .A1(n6805), .A2(n6803), .ZN(n6802) );
  INV_X1 U7969 ( .A(n6804), .ZN(n6803) );
  NAND3_X1 U7970 ( .A1(n14277), .A2(n6802), .A3(n6801), .ZN(n14219) );
  NAND2_X1 U7971 ( .A1(n14249), .A2(n7054), .ZN(n14225) );
  NAND2_X1 U7972 ( .A1(n14277), .A2(n14266), .ZN(n14264) );
  NOR2_X1 U7973 ( .A1(n14444), .A2(n14296), .ZN(n14277) );
  NAND2_X1 U7974 ( .A1(n14291), .A2(n14306), .ZN(n14290) );
  NAND2_X1 U7975 ( .A1(n7988), .A2(n7987), .ZN(n14356) );
  NAND2_X1 U7976 ( .A1(n7649), .A2(n7648), .ZN(n13812) );
  OR2_X1 U7977 ( .A1(n14688), .A2(n12121), .ZN(n12232) );
  NAND2_X1 U7978 ( .A1(n11872), .A2(n7924), .ZN(n11881) );
  NAND2_X1 U7979 ( .A1(n14850), .A2(n11591), .ZN(n7285) );
  OR2_X1 U7980 ( .A1(n8099), .A2(n11860), .ZN(n8197) );
  NAND2_X1 U7981 ( .A1(n7309), .A2(n8134), .ZN(n14268) );
  AND2_X2 U7982 ( .A1(n14528), .A2(n10512), .ZN(n14444) );
  OR2_X1 U7983 ( .A1(n11574), .A2(n7813), .ZN(n7791) );
  INV_X1 U7984 ( .A(n10323), .ZN(n14883) );
  INV_X1 U7985 ( .A(n14888), .ZN(n14904) );
  NOR2_X1 U7986 ( .A1(n7462), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7461) );
  INV_X1 U7987 ( .A(n7462), .ZN(n7460) );
  XNOR2_X1 U7988 ( .A(n7818), .B(n7817), .ZN(n13776) );
  XNOR2_X1 U7989 ( .A(n7636), .B(n7635), .ZN(n11256) );
  NAND2_X1 U7990 ( .A1(n6615), .A2(n7584), .ZN(n7091) );
  NAND2_X1 U7991 ( .A1(n7536), .A2(n7179), .ZN(n7175) );
  INV_X1 U7992 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7325) );
  INV_X1 U7993 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U7994 ( .A1(n7505), .A2(n7504), .ZN(n6842) );
  INV_X1 U7995 ( .A(n8500), .ZN(n6907) );
  XNOR2_X1 U7996 ( .A(n8507), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U7997 ( .A1(n6903), .A2(n6549), .ZN(n8547) );
  OR2_X1 U7998 ( .A1(n8538), .A2(n6904), .ZN(n6903) );
  OR2_X1 U7999 ( .A1(n14746), .A2(n6598), .ZN(n6904) );
  AND3_X1 U8000 ( .A1(n9755), .A2(n9754), .A3(n9753), .ZN(n15162) );
  AND2_X1 U8001 ( .A1(n12278), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U8002 ( .A1(n9613), .A2(n9612), .ZN(n12603) );
  INV_X1 U8003 ( .A(n7392), .ZN(n15171) );
  AND4_X1 U8004 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n12991)
         );
  NAND2_X1 U8005 ( .A1(n10060), .A2(n10059), .ZN(n13003) );
  INV_X1 U8006 ( .A(n12961), .ZN(n12934) );
  AND4_X1 U8007 ( .A1(n9886), .A2(n9885), .A3(n9884), .A4(n9883), .ZN(n12408)
         );
  AND4_X1 U8008 ( .A1(n9809), .A2(n9808), .A3(n9807), .A4(n9806), .ZN(n12352)
         );
  AOI21_X1 U8009 ( .B1(n10105), .B2(n10161), .A(n10156), .ZN(n10186) );
  INV_X1 U8010 ( .A(n10164), .ZN(n10156) );
  INV_X1 U8011 ( .A(n12866), .ZN(n12701) );
  NAND2_X1 U8012 ( .A1(n6751), .A2(n6548), .ZN(n6944) );
  AND2_X1 U8013 ( .A1(n6962), .A2(n6959), .ZN(n12786) );
  AND2_X1 U8014 ( .A1(n6966), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6961) );
  INV_X1 U8015 ( .A(n13092), .ZN(n12950) );
  AND3_X1 U8016 ( .A1(n9815), .A2(n9814), .A3(n9813), .ZN(n12331) );
  NAND2_X1 U8017 ( .A1(n10355), .A2(n10278), .ZN(n10280) );
  INV_X1 U8018 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9598) );
  INV_X1 U8019 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13115) );
  XNOR2_X1 U8020 ( .A(n9625), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11445) );
  OAI21_X1 U8021 ( .B1(n9626), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9625) );
  INV_X1 U8022 ( .A(n7252), .ZN(n7251) );
  AND2_X1 U8023 ( .A1(n10344), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7158) );
  NOR2_X1 U8024 ( .A1(n14924), .A2(n12104), .ZN(n7276) );
  OR2_X1 U8025 ( .A1(n8875), .A2(n8863), .ZN(n7265) );
  OR2_X1 U8026 ( .A1(n11574), .A2(n9140), .ZN(n9085) );
  INV_X1 U8027 ( .A(n13451), .ZN(n13661) );
  AND2_X1 U8028 ( .A1(n10689), .A2(n13419), .ZN(n13252) );
  OR2_X1 U8029 ( .A1(n9536), .A2(n9535), .ZN(n9537) );
  INV_X1 U8030 ( .A(n13536), .ZN(n13168) );
  NAND2_X1 U8031 ( .A1(n13376), .A2(n15033), .ZN(n6699) );
  NAND2_X1 U8032 ( .A1(n7128), .A2(n9180), .ZN(n13434) );
  OR2_X1 U8033 ( .A1(n12381), .A2(n9140), .ZN(n9142) );
  OR2_X1 U8034 ( .A1(n14668), .A2(n11210), .ZN(n13525) );
  INV_X1 U8035 ( .A(n13641), .ZN(n14665) );
  INV_X1 U8036 ( .A(n13636), .ZN(n14655) );
  OAI21_X1 U8037 ( .B1(n13398), .B2(n7145), .A(n7147), .ZN(n6729) );
  NAND2_X1 U8038 ( .A1(n15147), .A2(n15137), .ZN(n7145) );
  INV_X1 U8039 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U8040 ( .A1(n13733), .A2(n13749), .ZN(n7242) );
  AND2_X1 U8041 ( .A1(n13414), .A2(n7238), .ZN(n6734) );
  AND2_X1 U8042 ( .A1(n13651), .A2(n13413), .ZN(n7238) );
  NAND2_X1 U8043 ( .A1(n8798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8799) );
  INV_X1 U8044 ( .A(n8797), .ZN(n8800) );
  INV_X1 U8045 ( .A(n14235), .ZN(n6805) );
  NAND2_X1 U8046 ( .A1(n8062), .A2(n8061), .ZN(n14229) );
  AOI21_X1 U8047 ( .B1(n8096), .B2(n14384), .A(n8095), .ZN(n10322) );
  NOR2_X1 U8048 ( .A1(n13899), .A2(n14353), .ZN(n8095) );
  INV_X1 U8049 ( .A(n7313), .ZN(n7312) );
  OR2_X1 U8050 ( .A1(n11747), .A2(n7813), .ZN(n7808) );
  NOR2_X1 U8051 ( .A1(n15386), .A2(n15387), .ZN(n15385) );
  XNOR2_X1 U8052 ( .A(n8506), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15376) );
  NAND2_X1 U8053 ( .A1(n8519), .A2(n8520), .ZN(n14547) );
  INV_X1 U8054 ( .A(n8520), .ZN(n6646) );
  INV_X1 U8055 ( .A(n8519), .ZN(n6647) );
  XNOR2_X1 U8056 ( .A(n8531), .B(n8530), .ZN(n14733) );
  OAI21_X1 U8057 ( .B1(n14735), .B2(n14736), .A(n6708), .ZN(n6707) );
  INV_X1 U8058 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8059 ( .A1(n7440), .A2(n8232), .ZN(n7439) );
  NOR2_X1 U8060 ( .A1(n8232), .A2(n7440), .ZN(n7441) );
  INV_X1 U8061 ( .A(n9306), .ZN(n7340) );
  AOI21_X1 U8062 ( .B1(n7306), .B2(n7305), .A(n7303), .ZN(n7302) );
  INV_X1 U8063 ( .A(n9329), .ZN(n7303) );
  NAND2_X1 U8064 ( .A1(n8242), .A2(n8244), .ZN(n7432) );
  AND2_X1 U8065 ( .A1(n9333), .A2(n9334), .ZN(n7351) );
  NAND2_X1 U8066 ( .A1(n8253), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U8067 ( .A1(n6533), .A2(n7344), .ZN(n7343) );
  INV_X1 U8068 ( .A(n8272), .ZN(n7475) );
  NAND2_X1 U8069 ( .A1(n8271), .A2(n7475), .ZN(n7473) );
  INV_X1 U8070 ( .A(n7473), .ZN(n7469) );
  INV_X1 U8071 ( .A(n8281), .ZN(n7466) );
  NAND2_X1 U8072 ( .A1(n9391), .A2(n9390), .ZN(n7337) );
  NAND2_X1 U8073 ( .A1(n9400), .A2(n9389), .ZN(n7338) );
  AND2_X1 U8074 ( .A1(n6861), .A2(n6859), .ZN(n9734) );
  NOR2_X1 U8075 ( .A1(n10221), .A2(n6860), .ZN(n6859) );
  AND2_X1 U8076 ( .A1(n8289), .A2(n7457), .ZN(n7456) );
  OR2_X1 U8077 ( .A1(n8288), .A2(n8398), .ZN(n7457) );
  INV_X1 U8078 ( .A(n9871), .ZN(n6893) );
  AND2_X1 U8079 ( .A1(n9405), .A2(n9406), .ZN(n7352) );
  OR2_X1 U8080 ( .A1(n6869), .A2(n6868), .ZN(n9805) );
  OAI21_X1 U8081 ( .B1(n6870), .B2(n6507), .A(n6619), .ZN(n6868) );
  NOR3_X1 U8082 ( .A1(n9739), .A2(n10939), .A3(n6507), .ZN(n6869) );
  AOI21_X1 U8083 ( .B1(n6889), .B2(n6887), .A(n6886), .ZN(n6885) );
  INV_X1 U8084 ( .A(n9905), .ZN(n6886) );
  INV_X1 U8085 ( .A(n6891), .ZN(n6887) );
  NOR2_X1 U8086 ( .A1(n7320), .A2(n6569), .ZN(n7315) );
  NOR2_X1 U8087 ( .A1(n9424), .A2(n9423), .ZN(n7320) );
  INV_X1 U8088 ( .A(n9420), .ZN(n7321) );
  OAI21_X1 U8089 ( .B1(n9423), .B2(n6530), .A(n9424), .ZN(n7318) );
  NAND2_X1 U8090 ( .A1(n7319), .A2(n7316), .ZN(n9427) );
  AND2_X1 U8091 ( .A1(n7318), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U8092 ( .A1(n9421), .A2(n7315), .ZN(n7319) );
  NAND2_X1 U8093 ( .A1(n9423), .A2(n6530), .ZN(n7317) );
  AOI21_X1 U8094 ( .B1(n6881), .B2(n6883), .A(n6625), .ZN(n6880) );
  NAND2_X1 U8095 ( .A1(n8316), .A2(n7447), .ZN(n7446) );
  INV_X1 U8096 ( .A(n8317), .ZN(n7447) );
  NAND2_X1 U8097 ( .A1(n7326), .A2(n7328), .ZN(n9437) );
  AND2_X1 U8098 ( .A1(n6540), .A2(n7329), .ZN(n7328) );
  NOR2_X1 U8099 ( .A1(n12907), .A2(n6858), .ZN(n6857) );
  INV_X1 U8100 ( .A(n10000), .ZN(n6858) );
  OAI21_X1 U8101 ( .B1(n6856), .B2(n12892), .A(n6854), .ZN(n6853) );
  NOR2_X1 U8102 ( .A1(n6855), .A2(n12876), .ZN(n6854) );
  AOI21_X1 U8103 ( .B1(n10001), .B2(n6857), .A(n10002), .ZN(n6856) );
  NOR2_X1 U8104 ( .A1(n10003), .A2(n10147), .ZN(n6855) );
  INV_X1 U8105 ( .A(n15326), .ZN(n10212) );
  INV_X1 U8106 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U8107 ( .A1(n9444), .A2(n7293), .ZN(n7291) );
  AOI21_X1 U8108 ( .B1(n7430), .B2(n7428), .A(n8334), .ZN(n7426) );
  NAND2_X1 U8109 ( .A1(n6497), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U8110 ( .A1(n14212), .A2(n7052), .ZN(n7051) );
  INV_X1 U8111 ( .A(n8053), .ZN(n7052) );
  NAND2_X1 U8112 ( .A1(n7042), .A2(n8280), .ZN(n7041) );
  NAND2_X1 U8113 ( .A1(n12228), .A2(n7043), .ZN(n7042) );
  INV_X1 U8114 ( .A(n8274), .ZN(n7043) );
  NAND2_X1 U8115 ( .A1(n7578), .A2(n7204), .ZN(n7203) );
  INV_X1 U8116 ( .A(n7605), .ZN(n7204) );
  INV_X1 U8117 ( .A(n7190), .ZN(n7189) );
  OAI21_X1 U8118 ( .B1(n7193), .B2(n7191), .A(n7553), .ZN(n7190) );
  OR2_X1 U8119 ( .A1(n7552), .A2(n10797), .ZN(n7193) );
  INV_X1 U8120 ( .A(n7177), .ZN(n7176) );
  OAI21_X1 U8121 ( .B1(n7179), .B2(n7178), .A(n7763), .ZN(n7177) );
  INV_X1 U8122 ( .A(n7539), .ZN(n7178) );
  OR2_X1 U8123 ( .A1(n7013), .A2(n12841), .ZN(n6659) );
  NAND2_X1 U8124 ( .A1(n7014), .A2(n12822), .ZN(n7013) );
  NAND2_X1 U8125 ( .A1(n7012), .A2(n12822), .ZN(n7011) );
  INV_X1 U8126 ( .A(n10179), .ZN(n7073) );
  NAND2_X1 U8127 ( .A1(n10981), .A2(n6551), .ZN(n10946) );
  NAND2_X1 U8128 ( .A1(n11096), .A2(n10969), .ZN(n11097) );
  NAND2_X1 U8129 ( .A1(n11832), .A2(n11831), .ZN(n12006) );
  INV_X1 U8130 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12012) );
  NOR2_X1 U8131 ( .A1(n7416), .A2(n10149), .ZN(n7413) );
  INV_X1 U8132 ( .A(n10253), .ZN(n7416) );
  NAND2_X1 U8133 ( .A1(n10253), .A2(n7415), .ZN(n7414) );
  INV_X1 U8134 ( .A(n10250), .ZN(n7415) );
  OR2_X1 U8135 ( .A1(n12675), .A2(n12933), .ZN(n10145) );
  OR2_X1 U8136 ( .A1(n9949), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9963) );
  INV_X1 U8137 ( .A(n7402), .ZN(n7401) );
  OAI21_X1 U8138 ( .B1(n10241), .B2(n7403), .A(n12988), .ZN(n7402) );
  INV_X1 U8139 ( .A(n10242), .ZN(n7403) );
  INV_X1 U8140 ( .A(n6989), .ZN(n6988) );
  OAI21_X1 U8141 ( .B1(n11642), .B2(n6990), .A(n10120), .ZN(n6989) );
  INV_X1 U8142 ( .A(n10119), .ZN(n6990) );
  INV_X1 U8143 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U8144 ( .A1(n9586), .A2(n7395), .ZN(n7424) );
  NOR2_X1 U8145 ( .A1(n9621), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U8146 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n11746), .ZN(n9572) );
  INV_X1 U8147 ( .A(n7069), .ZN(n7068) );
  OAI21_X1 U8148 ( .B1(n9794), .B2(n7070), .A(n9810), .ZN(n7069) );
  INV_X1 U8149 ( .A(n9560), .ZN(n7070) );
  NOR2_X1 U8150 ( .A1(n7064), .A2(n7061), .ZN(n7060) );
  INV_X1 U8151 ( .A(n9549), .ZN(n7063) );
  NAND2_X1 U8152 ( .A1(n9684), .A2(n9582), .ZN(n6942) );
  INV_X2 U8153 ( .A(n10879), .ZN(n12547) );
  INV_X1 U8154 ( .A(n12112), .ZN(n7271) );
  INV_X1 U8155 ( .A(n7273), .ZN(n7272) );
  NAND2_X1 U8156 ( .A1(n7290), .A2(n7288), .ZN(n7292) );
  NOR2_X1 U8157 ( .A1(n9461), .A2(n7289), .ZN(n7288) );
  INV_X1 U8158 ( .A(n7291), .ZN(n7289) );
  OR2_X1 U8159 ( .A1(n6499), .A2(n14942), .ZN(n8829) );
  NAND2_X1 U8160 ( .A1(n7209), .A2(n6515), .ZN(n9246) );
  INV_X1 U8161 ( .A(n7484), .ZN(n7118) );
  AND2_X1 U8162 ( .A1(n7216), .A2(n9243), .ZN(n7215) );
  NAND2_X1 U8163 ( .A1(n9241), .A2(n7217), .ZN(n7216) );
  INV_X1 U8164 ( .A(n9240), .ZN(n7217) );
  NOR2_X1 U8165 ( .A1(n13621), .A2(n13712), .ZN(n6935) );
  INV_X1 U8166 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8986) );
  AND2_X1 U8167 ( .A1(n11785), .A2(n6821), .ZN(n6820) );
  NAND2_X1 U8168 ( .A1(n8979), .A2(n9232), .ZN(n6821) );
  INV_X1 U8169 ( .A(n9232), .ZN(n6822) );
  NAND2_X1 U8170 ( .A1(n15141), .A2(n6932), .ZN(n6931) );
  INV_X1 U8171 ( .A(n11387), .ZN(n6834) );
  INV_X1 U8172 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8730) );
  INV_X1 U8173 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U8174 ( .A1(n8790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8791) );
  INV_X1 U8175 ( .A(n8786), .ZN(n8795) );
  NAND2_X1 U8176 ( .A1(n7113), .A2(n13814), .ZN(n7111) );
  NOR2_X1 U8177 ( .A1(n13814), .A2(n7113), .ZN(n7112) );
  AOI21_X1 U8178 ( .B1(n6534), .B2(n7451), .A(n8345), .ZN(n7450) );
  NOR2_X1 U8179 ( .A1(n14433), .A2(n14438), .ZN(n6804) );
  INV_X1 U8180 ( .A(n8399), .ZN(n7298) );
  NOR2_X1 U8181 ( .A1(n14470), .A2(n6808), .ZN(n6806) );
  OR2_X1 U8182 ( .A1(n14688), .A2(n14058), .ZN(n8274) );
  OAI21_X1 U8183 ( .B1(n11871), .B2(n7035), .A(n6576), .ZN(n11979) );
  NAND2_X1 U8184 ( .A1(n7034), .A2(n7036), .ZN(n7033) );
  NAND2_X1 U8185 ( .A1(n14716), .A2(n6815), .ZN(n6814) );
  NAND2_X1 U8186 ( .A1(n7287), .A2(n7285), .ZN(n7283) );
  INV_X1 U8187 ( .A(n7285), .ZN(n7284) );
  NOR2_X1 U8188 ( .A1(n11567), .A2(n13916), .ZN(n6800) );
  NAND2_X1 U8189 ( .A1(n12117), .A2(n6547), .ZN(n7039) );
  INV_X1 U8190 ( .A(n7041), .ZN(n7037) );
  NAND2_X1 U8191 ( .A1(n7549), .A2(SI_16_), .ZN(n7633) );
  NAND2_X1 U8192 ( .A1(n7196), .A2(n7195), .ZN(n7194) );
  NOR2_X1 U8193 ( .A1(n7198), .A2(n7197), .ZN(n7196) );
  NAND2_X1 U8194 ( .A1(n7198), .A2(n7197), .ZN(n7195) );
  OR2_X1 U8195 ( .A1(n7759), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7765) );
  NOR2_X1 U8196 ( .A1(n7757), .A2(n7180), .ZN(n7179) );
  INV_X1 U8197 ( .A(n7535), .ZN(n7180) );
  AND2_X1 U8198 ( .A1(n7698), .A2(n7652), .ZN(n7718) );
  INV_X1 U8199 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U8200 ( .A1(n10345), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8201 ( .A1(n7516), .A2(SI_4_), .ZN(n7703) );
  INV_X1 U8202 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U8203 ( .A1(n6691), .A2(n8456), .ZN(n8457) );
  OAI21_X1 U8204 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n8462), .A(n8461), .ZN(
        n8463) );
  OAI21_X1 U8205 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15297), .A(n8468), .ZN(
        n8470) );
  INV_X1 U8206 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U8207 ( .A1(n15181), .A2(n6649), .ZN(n15159) );
  NAND2_X1 U8208 ( .A1(n11807), .A2(n12717), .ZN(n6649) );
  NAND2_X1 U8209 ( .A1(n7375), .A2(n7379), .ZN(n12473) );
  NAND2_X1 U8210 ( .A1(n10838), .A2(n10581), .ZN(n10584) );
  NOR2_X1 U8211 ( .A1(n9963), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9978) );
  AND2_X1 U8212 ( .A1(n12635), .A2(n12477), .ZN(n12654) );
  NAND2_X1 U8213 ( .A1(n12473), .A2(n12472), .ZN(n12653) );
  NAND2_X1 U8214 ( .A1(n9994), .A2(n9614), .ZN(n9615) );
  NOR2_X1 U8215 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9615), .ZN(n10010) );
  NAND2_X1 U8216 ( .A1(n12616), .A2(n12615), .ZN(n12614) );
  AND2_X1 U8217 ( .A1(n9757), .A2(n9756), .ZN(n9772) );
  NAND2_X1 U8218 ( .A1(n9772), .A2(n8586), .ZN(n9788) );
  INV_X1 U8219 ( .A(n7481), .ZN(n7361) );
  AND2_X1 U8220 ( .A1(n7359), .A2(n12178), .ZN(n7358) );
  NAND2_X1 U8221 ( .A1(n7481), .A2(n7360), .ZN(n7359) );
  AND2_X1 U8222 ( .A1(n9992), .A2(n12674), .ZN(n9994) );
  NAND2_X1 U8223 ( .A1(n12172), .A2(n12171), .ZN(n12342) );
  MUX2_X1 U8224 ( .A(n10580), .B(n10579), .S(n10585), .Z(n10838) );
  AND2_X1 U8225 ( .A1(n9915), .A2(n9914), .ZN(n9933) );
  NAND2_X1 U8226 ( .A1(n9933), .A2(n9932), .ZN(n9949) );
  NAND2_X1 U8227 ( .A1(n14610), .A2(n14603), .ZN(n10164) );
  AND3_X1 U8228 ( .A1(n10085), .A2(n10084), .A3(n10083), .ZN(n10088) );
  AND4_X1 U8229 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(n11025)
         );
  AOI21_X1 U8230 ( .B1(n11015), .B2(n11364), .A(n10944), .ZN(n11006) );
  NAND2_X1 U8231 ( .A1(n11096), .A2(n6510), .ZN(n6736) );
  NAND2_X1 U8232 ( .A1(n11520), .A2(n6741), .ZN(n6740) );
  OR2_X1 U8233 ( .A1(n15269), .A2(n11515), .ZN(n6939) );
  AND2_X1 U8234 ( .A1(n12256), .A2(n12255), .ZN(n12724) );
  OR2_X1 U8235 ( .A1(n12258), .A2(n12259), .ZN(n6752) );
  NAND2_X1 U8236 ( .A1(n12799), .A2(n12800), .ZN(n14568) );
  XNOR2_X1 U8237 ( .A(n12804), .B(n14583), .ZN(n14586) );
  XNOR2_X1 U8238 ( .A(n12791), .B(n14583), .ZN(n14594) );
  NAND2_X1 U8239 ( .A1(n14586), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14585) );
  AND2_X1 U8240 ( .A1(n10157), .A2(n10155), .ZN(n10266) );
  AND2_X1 U8241 ( .A1(n13003), .A2(n12700), .ZN(n10255) );
  NOR2_X1 U8242 ( .A1(n10037), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10061) );
  AND2_X1 U8243 ( .A1(n10061), .A2(n8562), .ZN(n14604) );
  NAND2_X1 U8244 ( .A1(n12894), .A2(n10148), .ZN(n12874) );
  AND2_X1 U8245 ( .A1(n12892), .A2(n7405), .ZN(n7404) );
  NAND2_X1 U8246 ( .A1(n7407), .A2(n7409), .ZN(n7405) );
  AND2_X1 U8247 ( .A1(n10145), .A2(n10144), .ZN(n12923) );
  OAI21_X1 U8248 ( .B1(n12968), .B2(n7022), .A(n7020), .ZN(n10143) );
  INV_X1 U8249 ( .A(n7023), .ZN(n7022) );
  AOI21_X1 U8250 ( .B1(n7023), .B2(n7025), .A(n7021), .ZN(n7020) );
  AND3_X1 U8251 ( .A1(n9984), .A2(n9983), .A3(n9982), .ZN(n12944) );
  NAND2_X1 U8252 ( .A1(n12974), .A2(n10245), .ZN(n12958) );
  AND2_X1 U8253 ( .A1(n12967), .A2(n10245), .ZN(n7425) );
  INV_X1 U8254 ( .A(n12707), .ZN(n12978) );
  OR2_X1 U8255 ( .A1(n9881), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9896) );
  NOR2_X1 U8256 ( .A1(n9896), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9915) );
  AOI21_X1 U8257 ( .B1(n6505), .B2(n6995), .A(n6993), .ZN(n6992) );
  INV_X1 U8258 ( .A(n10132), .ZN(n6993) );
  INV_X1 U8259 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U8260 ( .A1(n9865), .A2(n9864), .ZN(n9881) );
  AND3_X1 U8261 ( .A1(n9785), .A2(n9784), .A3(n9783), .ZN(n11799) );
  AND4_X1 U8262 ( .A1(n9747), .A2(n9746), .A3(n9745), .A4(n9744), .ZN(n11809)
         );
  NAND2_X1 U8263 ( .A1(n11405), .A2(n10225), .ZN(n11641) );
  AND2_X1 U8264 ( .A1(n10118), .A2(n9770), .ZN(n11808) );
  AOI21_X1 U8265 ( .B1(n10168), .B2(n10114), .A(n6584), .ZN(n6985) );
  NAND2_X1 U8266 ( .A1(n11077), .A2(n10113), .ZN(n11340) );
  NOR2_X1 U8267 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9717) );
  INV_X1 U8268 ( .A(n11024), .ZN(n10217) );
  CLKBUF_X1 U8269 ( .A(n10210), .Z(n15323) );
  NAND2_X1 U8270 ( .A1(n10009), .A2(n10008), .ZN(n12479) );
  NAND2_X1 U8271 ( .A1(n9976), .A2(n9975), .ZN(n12625) );
  INV_X1 U8272 ( .A(n12331), .ZN(n14622) );
  AND2_X1 U8273 ( .A1(n12912), .A2(n15359), .ZN(n14623) );
  INV_X1 U8274 ( .A(n10219), .ZN(n9652) );
  INV_X1 U8275 ( .A(n10047), .ZN(n7082) );
  NOR2_X1 U8276 ( .A1(n10074), .A2(n7084), .ZN(n7083) );
  INV_X1 U8277 ( .A(n10048), .ZN(n7084) );
  AND2_X1 U8278 ( .A1(n12426), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U8279 ( .A1(n7424), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7423) );
  OAI21_X1 U8280 ( .B1(n10004), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n10006), 
        .ZN(n10020) );
  INV_X1 U8281 ( .A(n7085), .ZN(n10005) );
  XNOR2_X1 U8282 ( .A(n7085), .B(n12377), .ZN(n10004) );
  NAND2_X1 U8283 ( .A1(n6786), .A2(n6636), .ZN(n9611) );
  INV_X1 U8284 ( .A(n6639), .ZN(n6785) );
  INV_X1 U8285 ( .A(n9621), .ZN(n9622) );
  NAND2_X1 U8286 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n7058), .ZN(n7057) );
  AOI21_X1 U8287 ( .B1(n6769), .B2(n7076), .A(n6768), .ZN(n6770) );
  INV_X1 U8288 ( .A(n7074), .ZN(n6768) );
  NAND2_X1 U8289 ( .A1(n9620), .A2(n9796), .ZN(n10187) );
  AOI21_X1 U8290 ( .B1(n6779), .B2(n6781), .A(n6778), .ZN(n6777) );
  XNOR2_X1 U8291 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9763) );
  AND2_X1 U8292 ( .A1(n9664), .A2(n9726), .ZN(n10965) );
  XNOR2_X1 U8293 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9682) );
  AND2_X1 U8294 ( .A1(n9542), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9681) );
  INV_X1 U8295 ( .A(n12561), .ZN(n7249) );
  NAND2_X1 U8296 ( .A1(n7252), .A2(n7249), .ZN(n7248) );
  OR2_X1 U8297 ( .A1(n9059), .A2(n8810), .ZN(n9075) );
  CLKBUF_X1 U8298 ( .A(n13180), .Z(n13181) );
  CLKBUF_X1 U8299 ( .A(n13143), .Z(n13144) );
  INV_X1 U8300 ( .A(n13193), .ZN(n7274) );
  XNOR2_X1 U8301 ( .A(n11231), .B(n10879), .ZN(n10694) );
  NAND2_X1 U8302 ( .A1(n12527), .A2(n13203), .ZN(n13201) );
  CLKBUF_X1 U8303 ( .A(n13153), .Z(n13154) );
  CLKBUF_X1 U8304 ( .A(n13223), .Z(n13224) );
  NAND2_X1 U8305 ( .A1(n8811), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9087) );
  INV_X1 U8306 ( .A(n9075), .ZN(n8811) );
  OR2_X1 U8307 ( .A1(n9087), .A2(n9086), .ZN(n9101) );
  AOI21_X1 U8308 ( .B1(n14965), .B2(n13279), .A(n13278), .ZN(n13294) );
  INV_X1 U8309 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11438) );
  OR2_X1 U8311 ( .A1(n9053), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9068) );
  OAI21_X1 U8312 ( .B1(n9074), .B2(n13363), .A(n15032), .ZN(n13364) );
  AOI21_X1 U8313 ( .B1(n6831), .B2(n13408), .A(n6830), .ZN(n6829) );
  INV_X1 U8314 ( .A(n7220), .ZN(n6831) );
  AND2_X1 U8315 ( .A1(n9255), .A2(n13427), .ZN(n6830) );
  NAND2_X1 U8316 ( .A1(n7221), .A2(n7220), .ZN(n13409) );
  AND2_X1 U8317 ( .A1(n9196), .A2(n9172), .ZN(n13449) );
  AND2_X1 U8318 ( .A1(n9505), .A2(n9504), .ZN(n13452) );
  INV_X1 U8319 ( .A(n6827), .ZN(n6824) );
  NAND2_X1 U8320 ( .A1(n13503), .A2(n13490), .ZN(n13487) );
  AOI21_X1 U8321 ( .B1(n7142), .B2(n13511), .A(n6582), .ZN(n7140) );
  INV_X1 U8322 ( .A(n7142), .ZN(n7141) );
  NAND2_X1 U8323 ( .A1(n8813), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U8324 ( .A1(n6933), .A2(n13554), .ZN(n13550) );
  OR2_X1 U8325 ( .A1(n13571), .A2(n9244), .ZN(n7484) );
  NAND2_X1 U8326 ( .A1(n13586), .A2(n9095), .ZN(n13573) );
  NAND2_X1 U8327 ( .A1(n7213), .A2(n7215), .ZN(n13563) );
  NAND2_X1 U8328 ( .A1(n7214), .A2(n9241), .ZN(n7213) );
  INV_X1 U8329 ( .A(n13596), .ZN(n7214) );
  NAND2_X1 U8330 ( .A1(n6935), .A2(n6934), .ZN(n13581) );
  INV_X1 U8331 ( .A(n6935), .ZN(n13601) );
  NAND2_X1 U8332 ( .A1(n6632), .A2(n6678), .ZN(n14661) );
  NAND2_X1 U8333 ( .A1(n9016), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9059) );
  OAI21_X1 U8334 ( .B1(n6843), .B2(n6583), .A(n9508), .ZN(n14649) );
  INV_X1 U8335 ( .A(n7229), .ZN(n6843) );
  INV_X1 U8336 ( .A(n9507), .ZN(n7230) );
  NOR2_X1 U8337 ( .A1(n11488), .A2(n14931), .ZN(n6927) );
  NOR2_X1 U8338 ( .A1(n8987), .A2(n8986), .ZN(n9002) );
  NAND2_X1 U8339 ( .A1(n11608), .A2(n9232), .ZN(n11786) );
  NAND2_X1 U8340 ( .A1(n6819), .A2(n6820), .ZN(n11784) );
  OR2_X1 U8341 ( .A1(n11609), .A2(n6822), .ZN(n6819) );
  INV_X1 U8342 ( .A(n11488), .ZN(n6930) );
  NOR2_X1 U8343 ( .A1(n11488), .A2(n6931), .ZN(n11792) );
  NAND2_X1 U8344 ( .A1(n11609), .A2(n11613), .ZN(n11608) );
  AND2_X1 U8345 ( .A1(n9231), .A2(n8965), .ZN(n11484) );
  NOR2_X1 U8346 ( .A1(n11488), .A2(n11701), .ZN(n11615) );
  NAND2_X1 U8347 ( .A1(n6835), .A2(n6836), .ZN(n11386) );
  NAND2_X1 U8348 ( .A1(n11304), .A2(n11291), .ZN(n11314) );
  AND2_X1 U8349 ( .A1(n15127), .A2(n11303), .ZN(n11304) );
  NOR2_X1 U8350 ( .A1(n11267), .A2(n11268), .ZN(n11303) );
  NAND2_X1 U8351 ( .A1(n6922), .A2(n6921), .ZN(n11267) );
  INV_X1 U8352 ( .A(n10639), .ZN(n10637) );
  NAND2_X1 U8353 ( .A1(n11278), .A2(n9222), .ZN(n7208) );
  AND2_X1 U8354 ( .A1(n8853), .A2(n8852), .ZN(n10715) );
  NAND2_X1 U8355 ( .A1(n9450), .A2(n9449), .ZN(n13384) );
  INV_X1 U8356 ( .A(n13490), .ZN(n13671) );
  NAND2_X1 U8357 ( .A1(n9116), .A2(n9115), .ZN(n13541) );
  NAND2_X1 U8358 ( .A1(n9046), .A2(n9045), .ZN(n13721) );
  INV_X1 U8359 ( .A(n15140), .ZN(n15100) );
  NAND2_X1 U8360 ( .A1(n6841), .A2(n9228), .ZN(n11319) );
  NAND2_X1 U8361 ( .A1(n11175), .A2(n11178), .ZN(n6841) );
  CLKBUF_X1 U8362 ( .A(n10662), .Z(n9219) );
  OR2_X1 U8363 ( .A1(n9217), .A2(n9220), .ZN(n15123) );
  AND2_X1 U8364 ( .A1(n10682), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10336) );
  NAND2_X1 U8365 ( .A1(n6919), .A2(n8749), .ZN(n9263) );
  NAND2_X1 U8366 ( .A1(n6920), .A2(n8744), .ZN(n6919) );
  NAND2_X1 U8367 ( .A1(n8743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8744) );
  AND2_X1 U8368 ( .A1(n8757), .A2(n8756), .ZN(n8769) );
  AOI21_X1 U8369 ( .B1(n8796), .B2(P2_IR_REG_31__SCAN_IN), .A(n8798), .ZN(
        n8797) );
  NAND2_X1 U8370 ( .A1(n8998), .A2(n8795), .ZN(n8796) );
  OR2_X1 U8371 ( .A1(n8937), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8939) );
  OR2_X1 U8372 ( .A1(n8939), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U8373 ( .A1(n7136), .A2(n7137), .ZN(n7135) );
  INV_X1 U8374 ( .A(n7132), .ZN(n7131) );
  INV_X1 U8375 ( .A(n12055), .ZN(n7136) );
  INV_X1 U8376 ( .A(n7101), .ZN(n7099) );
  NOR2_X1 U8377 ( .A1(n6531), .A2(n7098), .ZN(n7097) );
  INV_X1 U8378 ( .A(n13875), .ZN(n7098) );
  INV_X1 U8379 ( .A(n13929), .ZN(n7105) );
  INV_X1 U8380 ( .A(n13952), .ZN(n13850) );
  INV_X1 U8381 ( .A(n13887), .ZN(n13881) );
  XNOR2_X1 U8382 ( .A(n13868), .B(n12151), .ZN(n13877) );
  OR2_X1 U8383 ( .A1(n7993), .A2(n7992), .ZN(n8001) );
  OR2_X1 U8384 ( .A1(n8010), .A2(n13953), .ZN(n8016) );
  NAND2_X1 U8385 ( .A1(n7972), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7993) );
  INV_X1 U8386 ( .A(n7974), .ZN(n7972) );
  NAND2_X1 U8387 ( .A1(n7139), .A2(n11846), .ZN(n7138) );
  NAND2_X1 U8388 ( .A1(n11843), .A2(n11845), .ZN(n7137) );
  NOR2_X1 U8389 ( .A1(n7874), .A2(n7873), .ZN(n7882) );
  INV_X1 U8390 ( .A(n13876), .ZN(n13890) );
  NAND2_X1 U8391 ( .A1(n8194), .A2(n8364), .ZN(n10861) );
  INV_X1 U8392 ( .A(n13932), .ZN(n13854) );
  NAND2_X1 U8393 ( .A1(n14686), .A2(n7112), .ZN(n7116) );
  NAND2_X1 U8394 ( .A1(n14686), .A2(n13811), .ZN(n7108) );
  XNOR2_X1 U8395 ( .A(n7171), .B(n14172), .ZN(n8423) );
  OR2_X1 U8396 ( .A1(n8442), .A2(n6596), .ZN(n7482) );
  AND4_X1 U8397 ( .A1(n7962), .A2(n7961), .A3(n7960), .A4(n7959), .ZN(n13977)
         );
  NAND2_X1 U8398 ( .A1(n14118), .A2(n14117), .ZN(n14761) );
  AOI21_X1 U8399 ( .B1(n10628), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10627), .ZN(
        n10764) );
  AOI21_X1 U8400 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10652), .A(n10733), .ZN(
        n10655) );
  AOI21_X1 U8401 ( .B1(n10785), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10778), .ZN(
        n10757) );
  NAND2_X1 U8402 ( .A1(n11125), .A2(n6661), .ZN(n14785) );
  OR2_X1 U8403 ( .A1(n11126), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U8404 ( .A1(n14785), .A2(n14786), .ZN(n14784) );
  AOI21_X1 U8405 ( .B1(n11775), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11774), .ZN(
        n14148) );
  AOI21_X1 U8406 ( .B1(n12239), .B2(P1_REG1_REG_17__SCAN_IN), .A(n12238), .ZN(
        n14157) );
  INV_X1 U8407 ( .A(n6798), .ZN(n6796) );
  XNOR2_X1 U8408 ( .A(n8342), .B(n13944), .ZN(n8419) );
  AND2_X1 U8409 ( .A1(n10327), .A2(n8074), .ZN(n13942) );
  OR2_X1 U8410 ( .A1(n8055), .A2(n8054), .ZN(n8066) );
  AND2_X1 U8411 ( .A1(n14249), .A2(n8041), .ZN(n14226) );
  OR2_X1 U8412 ( .A1(n8016), .A2(n14028), .ZN(n8032) );
  INV_X1 U8413 ( .A(n6703), .ZN(n7044) );
  OAI21_X1 U8414 ( .B1(n7046), .B2(n14306), .A(n8020), .ZN(n6703) );
  NAND2_X1 U8415 ( .A1(n14336), .A2(n8293), .ZN(n14311) );
  NAND2_X1 U8416 ( .A1(n14389), .A2(n6807), .ZN(n14367) );
  NAND2_X1 U8417 ( .A1(n14389), .A2(n14395), .ZN(n14390) );
  NOR2_X1 U8418 ( .A1(n13812), .A2(n12232), .ZN(n14389) );
  INV_X1 U8419 ( .A(n7957), .ZN(n7955) );
  NAND2_X1 U8420 ( .A1(n7040), .A2(n8274), .ZN(n12224) );
  NAND2_X1 U8421 ( .A1(n12117), .A2(n8401), .ZN(n7040) );
  NAND2_X1 U8422 ( .A1(n6813), .A2(n6514), .ZN(n12121) );
  AND2_X1 U8423 ( .A1(n7932), .A2(n7931), .ZN(n7940) );
  NAND2_X1 U8424 ( .A1(n6813), .A2(n6812), .ZN(n12037) );
  NOR2_X1 U8425 ( .A1(n11868), .A2(n6814), .ZN(n11974) );
  INV_X1 U8426 ( .A(n8407), .ZN(n11886) );
  NAND2_X1 U8427 ( .A1(n7923), .A2(n7922), .ZN(n11872) );
  NOR2_X1 U8428 ( .A1(n11868), .A2(n12200), .ZN(n11887) );
  OR2_X1 U8429 ( .A1(n11721), .A2(n12153), .ZN(n11868) );
  OAI21_X1 U8430 ( .B1(n11496), .B2(n7899), .A(n7898), .ZN(n11654) );
  NOR2_X1 U8431 ( .A1(n11503), .A2(n12089), .ZN(n11657) );
  NAND2_X1 U8432 ( .A1(n6800), .A2(n14850), .ZN(n11681) );
  NOR2_X1 U8433 ( .A1(n13916), .A2(n11567), .ZN(n11682) );
  NAND2_X1 U8434 ( .A1(n11568), .A2(n14845), .ZN(n11567) );
  AND2_X1 U8435 ( .A1(n11704), .A2(n11860), .ZN(n11568) );
  OR2_X1 U8436 ( .A1(n10867), .A2(n10318), .ZN(n10325) );
  INV_X1 U8437 ( .A(n8202), .ZN(n7347) );
  OR2_X1 U8438 ( .A1(n10861), .A2(n14101), .ZN(n14351) );
  NAND2_X1 U8439 ( .A1(n7642), .A2(n7641), .ZN(n14480) );
  INV_X1 U8440 ( .A(n13812), .ZN(n14697) );
  OR2_X1 U8441 ( .A1(n10867), .A2(n8187), .ZN(n8720) );
  OR2_X1 U8442 ( .A1(n10887), .A2(n7827), .ZN(n14875) );
  AND2_X1 U8443 ( .A1(n10319), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10335) );
  NAND2_X1 U8444 ( .A1(n8174), .A2(n8188), .ZN(n10407) );
  XNOR2_X1 U8445 ( .A(n8353), .B(n8352), .ZN(n12444) );
  AND2_X1 U8446 ( .A1(n7611), .A2(n7612), .ZN(n13773) );
  OR2_X1 U8447 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  AND2_X1 U8448 ( .A1(n7597), .A2(n7349), .ZN(n7348) );
  INV_X1 U8449 ( .A(n8155), .ZN(n8161) );
  XNOR2_X1 U8450 ( .A(n7796), .B(n7795), .ZN(n11745) );
  INV_X1 U8451 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7585) );
  OR2_X1 U8452 ( .A1(n7544), .A2(SI_14_), .ZN(n7200) );
  NAND2_X1 U8453 ( .A1(n7536), .A2(n7535), .ZN(n7758) );
  NOR2_X1 U8454 ( .A1(n7744), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7752) );
  OR2_X1 U8455 ( .A1(n7727), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7735) );
  OR2_X1 U8456 ( .A1(n7735), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7744) );
  NOR2_X1 U8457 ( .A1(n7679), .A2(n7511), .ZN(n7512) );
  INV_X1 U8458 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U8459 ( .A1(n7584), .A2(n7583), .ZN(n7696) );
  NAND2_X1 U8460 ( .A1(n6679), .A2(n6484), .ZN(n7682) );
  INV_X1 U8461 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11366) );
  NAND2_X1 U8462 ( .A1(n8449), .A2(n6719), .ZN(n8498) );
  NAND2_X1 U8463 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6720), .ZN(n6719) );
  INV_X1 U8464 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6720) );
  XNOR2_X1 U8465 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n8497) );
  XNOR2_X1 U8466 ( .A(n8451), .B(n6693), .ZN(n8496) );
  INV_X1 U8467 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U8468 ( .A1(n8510), .A2(n15378), .ZN(n8514) );
  NAND2_X1 U8469 ( .A1(n6902), .A2(n6900), .ZN(n6692) );
  NAND2_X1 U8470 ( .A1(n6901), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8471 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n8476), .A(n8475), .ZN(
        n8485) );
  NAND2_X1 U8472 ( .A1(n14740), .A2(n6915), .ZN(n6912) );
  NAND2_X1 U8473 ( .A1(n6914), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6913) );
  INV_X1 U8474 ( .A(n14740), .ZN(n6914) );
  NOR2_X1 U8475 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14747), .ZN(n8538) );
  NAND2_X1 U8476 ( .A1(n6655), .A2(n12653), .ZN(n12599) );
  OR2_X1 U8477 ( .A1(n12473), .A2(n12472), .ZN(n6655) );
  AOI21_X1 U8478 ( .B1(n6654), .B2(n7382), .A(n6653), .ZN(n11943) );
  INV_X1 U8479 ( .A(n7380), .ZN(n6653) );
  AOI21_X1 U8480 ( .B1(n7381), .B2(n7382), .A(n11940), .ZN(n7380) );
  AND3_X1 U8481 ( .A1(n9801), .A2(n9800), .A3(n9799), .ZN(n11947) );
  NAND2_X1 U8482 ( .A1(n7364), .A2(n12461), .ZN(n12607) );
  NAND2_X1 U8483 ( .A1(n12681), .A2(n12680), .ZN(n7364) );
  AOI21_X1 U8484 ( .B1(n7371), .B2(n7373), .A(n6575), .ZN(n7369) );
  AOI21_X1 U8485 ( .B1(n7390), .B2(n15174), .A(n6581), .ZN(n7386) );
  NAND2_X1 U8486 ( .A1(n7392), .A2(n7390), .ZN(n11245) );
  AND2_X1 U8487 ( .A1(n12614), .A2(n7382), .ZN(n11941) );
  NAND2_X1 U8488 ( .A1(n12614), .A2(n7384), .ZN(n11814) );
  AOI21_X1 U8489 ( .B1(n7365), .B2(n7367), .A(n6579), .ZN(n7362) );
  INV_X1 U8490 ( .A(n7375), .ZN(n7374) );
  NAND2_X1 U8491 ( .A1(n7376), .A2(n7379), .ZN(n12673) );
  AND4_X1 U8492 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(n12334)
         );
  AND2_X1 U8493 ( .A1(n10600), .A2(n10799), .ZN(n15186) );
  NAND2_X1 U8494 ( .A1(n7370), .A2(n12369), .ZN(n12401) );
  NAND2_X1 U8495 ( .A1(n12367), .A2(n12366), .ZN(n7370) );
  INV_X1 U8496 ( .A(n15193), .ZN(n12696) );
  INV_X1 U8497 ( .A(n15180), .ZN(n15172) );
  INV_X1 U8498 ( .A(n12944), .ZN(n12705) );
  INV_X1 U8499 ( .A(n12979), .ZN(n12706) );
  INV_X1 U8500 ( .A(n12991), .ZN(n12964) );
  INV_X1 U8501 ( .A(n12408), .ZN(n12709) );
  INV_X1 U8502 ( .A(n11809), .ZN(n11810) );
  INV_X1 U8503 ( .A(n11025), .ZN(n12722) );
  AND4_X1 U8504 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n10209)
         );
  NAND2_X1 U8505 ( .A1(n10982), .A2(n10983), .ZN(n10981) );
  OAI21_X1 U8506 ( .B1(n10961), .B2(P3_REG1_REG_2__SCAN_IN), .A(n6727), .ZN(
        n10983) );
  NAND2_X1 U8507 ( .A1(n10961), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6727) );
  INV_X1 U8508 ( .A(n6746), .ZN(n10987) );
  AOI21_X1 U8509 ( .B1(n15206), .B2(n10964), .A(n15195), .ZN(n15215) );
  INV_X1 U8510 ( .A(n15259), .ZN(n6749) );
  INV_X1 U8511 ( .A(n6939), .ZN(n11518) );
  XNOR2_X1 U8512 ( .A(n12724), .B(n12257), .ZN(n12258) );
  INV_X1 U8513 ( .A(n6752), .ZN(n12725) );
  INV_X1 U8514 ( .A(n6967), .ZN(n12730) );
  NAND2_X1 U8515 ( .A1(n12753), .A2(n6964), .ZN(n6963) );
  INV_X1 U8516 ( .A(n6744), .ZN(n14578) );
  NOR2_X1 U8517 ( .A1(n10974), .A2(n10973), .ZN(n14593) );
  OAI21_X1 U8518 ( .B1(n12792), .B2(n6958), .A(n12815), .ZN(n6957) );
  NAND2_X1 U8519 ( .A1(n6948), .A2(n6642), .ZN(n6952) );
  NAND2_X1 U8520 ( .A1(n12792), .A2(n12815), .ZN(n6948) );
  NAND2_X1 U8521 ( .A1(n6958), .A2(n12815), .ZN(n6947) );
  NAND2_X1 U8522 ( .A1(n6539), .A2(n6725), .ZN(n6724) );
  INV_X1 U8523 ( .A(n12832), .ZN(n6725) );
  NOR2_X1 U8524 ( .A1(n6955), .A2(n6958), .ZN(n6950) );
  INV_X1 U8525 ( .A(n14610), .ZN(n14605) );
  NAND2_X1 U8526 ( .A1(n10078), .A2(n10077), .ZN(n14615) );
  AOI21_X1 U8527 ( .B1(n12840), .B2(n12839), .A(n12838), .ZN(n13006) );
  NAND2_X1 U8528 ( .A1(n6997), .A2(n7000), .ZN(n12853) );
  OR2_X1 U8529 ( .A1(n12894), .A2(n7003), .ZN(n6997) );
  OAI21_X1 U8530 ( .B1(n12864), .B2(n15308), .A(n6731), .ZN(n13011) );
  INV_X1 U8531 ( .A(n6732), .ZN(n6731) );
  OAI22_X1 U8532 ( .A1(n12866), .A2(n15303), .B1(n15302), .B2(n12865), .ZN(
        n6732) );
  NAND2_X1 U8533 ( .A1(n7005), .A2(n7006), .ZN(n12867) );
  NAND2_X1 U8534 ( .A1(n12894), .A2(n6532), .ZN(n7005) );
  NAND2_X1 U8535 ( .A1(n7411), .A2(n7410), .ZN(n12906) );
  NAND2_X1 U8536 ( .A1(n7419), .A2(n10247), .ZN(n12931) );
  NAND2_X1 U8537 ( .A1(n7019), .A2(n7023), .ZN(n12935) );
  NAND2_X1 U8538 ( .A1(n12968), .A2(n7026), .ZN(n7019) );
  NAND2_X1 U8539 ( .A1(n7028), .A2(n7026), .ZN(n12954) );
  NAND2_X1 U8540 ( .A1(n7028), .A2(n10139), .ZN(n12952) );
  NAND2_X1 U8541 ( .A1(n12358), .A2(n10241), .ZN(n7400) );
  NAND2_X1 U8542 ( .A1(n6994), .A2(n10130), .ZN(n12297) );
  OAI21_X1 U8543 ( .B1(n10129), .B2(n6995), .A(n6505), .ZN(n12295) );
  NAND2_X1 U8544 ( .A1(n10129), .A2(n6996), .ZN(n6994) );
  NAND2_X1 U8545 ( .A1(n10129), .A2(n10128), .ZN(n12144) );
  NAND2_X1 U8546 ( .A1(n10236), .A2(n10235), .ZN(n12091) );
  AND3_X1 U8547 ( .A1(n9829), .A2(n9828), .A3(n9827), .ZN(n14617) );
  NAND2_X1 U8548 ( .A1(n11992), .A2(n11991), .ZN(n11990) );
  NAND2_X1 U8549 ( .A1(n6982), .A2(n10124), .ZN(n11992) );
  NAND2_X1 U8550 ( .A1(n11951), .A2(n10172), .ZN(n6982) );
  NAND2_X1 U8551 ( .A1(n11637), .A2(n10119), .ZN(n11728) );
  NAND2_X1 U8552 ( .A1(n11082), .A2(n10222), .ZN(n11343) );
  INV_X1 U8553 ( .A(n15331), .ZN(n12946) );
  OR2_X1 U8554 ( .A1(n11424), .A2(n10811), .ZN(n12997) );
  NAND2_X1 U8555 ( .A1(n12946), .A2(n11424), .ZN(n15334) );
  AND2_X2 U8556 ( .A1(n10807), .A2(n10299), .ZN(n15374) );
  AND2_X1 U8557 ( .A1(n14612), .A2(n14611), .ZN(n14629) );
  NOR2_X1 U8558 ( .A1(n13011), .A2(n6730), .ZN(n13068) );
  AND2_X1 U8559 ( .A1(n13012), .A2(n15339), .ZN(n6730) );
  OR3_X1 U8560 ( .A1(n13023), .A2(n13022), .A3(n13021), .ZN(n13076) );
  AND2_X1 U8561 ( .A1(n9962), .A2(n9961), .ZN(n13092) );
  NAND2_X1 U8562 ( .A1(n9948), .A2(n9947), .ZN(n13095) );
  AOI21_X1 U8563 ( .B1(n10796), .B2(n10076), .A(n9913), .ZN(n13105) );
  NAND2_X1 U8564 ( .A1(n9863), .A2(n9862), .ZN(n12330) );
  NAND2_X1 U8565 ( .A1(n9842), .A2(n9841), .ZN(n12222) );
  INV_X1 U8566 ( .A(n15162), .ZN(n11674) );
  NAND2_X1 U8567 ( .A1(n15365), .A2(n15325), .ZN(n13110) );
  AND2_X2 U8568 ( .A1(n10312), .A2(n10937), .ZN(n15365) );
  NOR2_X1 U8569 ( .A1(n10355), .A2(n10354), .ZN(n10419) );
  INV_X1 U8570 ( .A(n10573), .ZN(n10354) );
  NAND2_X1 U8571 ( .A1(n7079), .A2(n10096), .ZN(n6764) );
  OAI21_X1 U8572 ( .B1(n6765), .B2(n10096), .A(n6762), .ZN(n6761) );
  XNOR2_X1 U8573 ( .A(n10092), .B(n10091), .ZN(n12575) );
  AOI21_X1 U8574 ( .B1(n10057), .B2(n7083), .A(n7081), .ZN(n10092) );
  NAND2_X1 U8575 ( .A1(n13114), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U8576 ( .A1(n9600), .A2(n13114), .ZN(n13121) );
  NOR2_X1 U8577 ( .A1(n10193), .A2(n7394), .ZN(n7393) );
  AND2_X1 U8578 ( .A1(n9589), .A2(n7395), .ZN(n7394) );
  NAND2_X1 U8579 ( .A1(n6789), .A2(n9576), .ZN(n9989) );
  NAND2_X1 U8580 ( .A1(n9974), .A2(n9972), .ZN(n6789) );
  OR2_X1 U8581 ( .A1(n9624), .A2(n6877), .ZN(n6876) );
  AND2_X1 U8582 ( .A1(n6878), .A2(n9627), .ZN(n6875) );
  INV_X1 U8583 ( .A(SI_20_), .ZN(n11336) );
  INV_X1 U8584 ( .A(SI_16_), .ZN(n10546) );
  NAND2_X1 U8585 ( .A1(n7075), .A2(n9567), .ZN(n9876) );
  NAND2_X1 U8586 ( .A1(n9854), .A2(n9853), .ZN(n7075) );
  INV_X1 U8587 ( .A(SI_15_), .ZN(n10522) );
  INV_X1 U8588 ( .A(SI_12_), .ZN(n10401) );
  NAND2_X1 U8589 ( .A1(n7067), .A2(n9560), .ZN(n9811) );
  NAND2_X1 U8590 ( .A1(n9795), .A2(n9794), .ZN(n7067) );
  XNOR2_X1 U8591 ( .A(n9767), .B(n9766), .ZN(n15256) );
  NAND2_X1 U8592 ( .A1(n6776), .A2(n6779), .ZN(n9749) );
  OR2_X1 U8593 ( .A1(n9725), .A2(n6781), .ZN(n6776) );
  NAND2_X1 U8594 ( .A1(n6784), .A2(n9550), .ZN(n9634) );
  NAND2_X1 U8595 ( .A1(n7065), .A2(n9549), .ZN(n9659) );
  NAND2_X1 U8596 ( .A1(n9644), .A2(n9643), .ZN(n7065) );
  NAND2_X1 U8597 ( .A1(n9686), .A2(n9685), .ZN(n10959) );
  INV_X1 U8598 ( .A(n7258), .ZN(n11189) );
  OR2_X1 U8599 ( .A1(n12130), .A2(n7273), .ZN(n12504) );
  NAND2_X1 U8600 ( .A1(n11186), .A2(n7262), .ZN(n7261) );
  INV_X1 U8601 ( .A(n11187), .ZN(n7262) );
  AND3_X1 U8602 ( .A1(n9114), .A2(n9113), .A3(n9112), .ZN(n13538) );
  NAND2_X1 U8603 ( .A1(n12106), .A2(n12105), .ZN(n14925) );
  NAND2_X1 U8604 ( .A1(n9056), .A2(n9055), .ZN(n14644) );
  NOR2_X1 U8605 ( .A1(n10824), .A2(n10823), .ZN(n10878) );
  INV_X1 U8606 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11379) );
  AOI21_X1 U8607 ( .B1(n11276), .B2(n6483), .A(n11279), .ZN(n10709) );
  OR2_X1 U8609 ( .A1(n12109), .A2(n12108), .ZN(n12110) );
  NOR2_X1 U8610 ( .A1(n12111), .A2(n12112), .ZN(n12130) );
  AND2_X1 U8611 ( .A1(n9131), .A2(n9130), .ZN(n13521) );
  OR2_X1 U8612 ( .A1(n12136), .A2(n9140), .ZN(n9131) );
  INV_X1 U8613 ( .A(n13261), .ZN(n11788) );
  NAND2_X1 U8614 ( .A1(n10664), .A2(n10666), .ZN(n10667) );
  INV_X1 U8615 ( .A(n10665), .ZN(n10666) );
  NAND2_X1 U8616 ( .A1(n13172), .A2(n12552), .ZN(n13230) );
  INV_X1 U8617 ( .A(n13252), .ZN(n14930) );
  CLKBUF_X1 U8618 ( .A(n13241), .Z(n13242) );
  INV_X1 U8619 ( .A(n14926), .ZN(n13243) );
  NAND2_X2 U8620 ( .A1(n6528), .A2(n8874), .ZN(n13268) );
  OR2_X1 U8621 ( .A1(n8869), .A2(n10462), .ZN(n8858) );
  OR2_X1 U8622 ( .A1(n8904), .A2(n8855), .ZN(n8860) );
  CLKBUF_X1 U8623 ( .A(n9221), .Z(n13269) );
  OAI21_X1 U8624 ( .B1(n13294), .B2(n13293), .A(n13292), .ZN(n13309) );
  AND2_X1 U8625 ( .A1(n14985), .A2(n13326), .ZN(n13328) );
  NAND2_X1 U8626 ( .A1(n6695), .A2(n6694), .ZN(n14999) );
  OR2_X1 U8627 ( .A1(n13354), .A2(n13353), .ZN(n13370) );
  NAND2_X1 U8628 ( .A1(n13360), .A2(n6634), .ZN(n15034) );
  INV_X1 U8629 ( .A(n13405), .ZN(n6669) );
  NAND2_X1 U8630 ( .A1(n6687), .A2(n6686), .ZN(n6685) );
  XNOR2_X1 U8631 ( .A(n13426), .B(n9190), .ZN(n6688) );
  NAND2_X1 U8632 ( .A1(n13428), .A2(n13612), .ZN(n6686) );
  AND2_X1 U8633 ( .A1(n9169), .A2(n9168), .ZN(n13451) );
  NAND2_X1 U8634 ( .A1(n13517), .A2(n9139), .ZN(n13500) );
  NAND2_X1 U8635 ( .A1(n13598), .A2(n9081), .ZN(n13588) );
  NAND2_X1 U8636 ( .A1(n13596), .A2(n9240), .ZN(n13578) );
  NAND2_X1 U8637 ( .A1(n14657), .A2(n9041), .ZN(n13640) );
  NAND2_X1 U8638 ( .A1(n7229), .A2(n9234), .ZN(n11905) );
  NAND2_X1 U8639 ( .A1(n8897), .A2(n7125), .ZN(n11297) );
  NAND2_X1 U8640 ( .A1(n11261), .A2(n8896), .ZN(n7125) );
  NAND2_X1 U8641 ( .A1(n7227), .A2(n9227), .ZN(n11299) );
  OR2_X1 U8642 ( .A1(n14668), .A2(n11229), .ZN(n13636) );
  INV_X1 U8643 ( .A(n7162), .ZN(n7161) );
  NAND2_X1 U8644 ( .A1(n10688), .A2(n15090), .ZN(n13419) );
  AND2_X1 U8645 ( .A1(n15156), .A2(n13648), .ZN(n6925) );
  OR2_X1 U8646 ( .A1(n10382), .A2(n9140), .ZN(n8914) );
  INV_X1 U8647 ( .A(n13384), .ZN(n13728) );
  AND2_X1 U8648 ( .A1(n15147), .A2(n13648), .ZN(n6926) );
  INV_X1 U8649 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7241) );
  INV_X1 U8650 ( .A(n13521), .ZN(n13748) );
  INV_X1 U8651 ( .A(n13541), .ZN(n13755) );
  AND2_X1 U8652 ( .A1(n10683), .A2(n10336), .ZN(n15090) );
  NOR2_X1 U8653 ( .A1(n8747), .A2(n7232), .ZN(n7231) );
  NAND2_X1 U8654 ( .A1(n8815), .A2(n8819), .ZN(n7232) );
  CLKBUF_X1 U8655 ( .A(n9263), .Z(n13774) );
  INV_X1 U8656 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11748) );
  INV_X1 U8657 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10383) );
  INV_X1 U8658 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10370) );
  INV_X1 U8659 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10343) );
  INV_X1 U8660 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U8661 ( .A1(n7103), .A2(n7107), .ZN(n7100) );
  NAND2_X1 U8662 ( .A1(n12204), .A2(n12203), .ZN(n12308) );
  AND2_X1 U8663 ( .A1(n12205), .A2(n12202), .ZN(n12203) );
  AOI21_X1 U8664 ( .B1(n11584), .B2(n11583), .A(n7486), .ZN(n13915) );
  NAND2_X1 U8665 ( .A1(n14036), .A2(n7094), .ZN(n13923) );
  NOR2_X1 U8666 ( .A1(n13921), .A2(n7095), .ZN(n7094) );
  INV_X1 U8667 ( .A(n13837), .ZN(n7095) );
  NAND2_X1 U8668 ( .A1(n14036), .A2(n13837), .ZN(n13922) );
  NAND2_X1 U8669 ( .A1(n14007), .A2(n13848), .ZN(n13951) );
  NAND2_X1 U8670 ( .A1(n7815), .A2(n7814), .ZN(n14449) );
  OR2_X1 U8671 ( .A1(n12588), .A2(n7813), .ZN(n7815) );
  XNOR2_X1 U8672 ( .A(n13877), .B(n13878), .ZN(n14001) );
  NAND2_X1 U8673 ( .A1(n11599), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14696) );
  INV_X1 U8674 ( .A(n14078), .ZN(n12317) );
  NAND2_X1 U8675 ( .A1(n12308), .A2(n12307), .ZN(n12311) );
  NAND2_X1 U8676 ( .A1(n7130), .A2(n7137), .ZN(n12056) );
  NAND2_X1 U8677 ( .A1(n11844), .A2(n7138), .ZN(n7130) );
  OR2_X1 U8678 ( .A1(n10867), .A2(n10866), .ZN(n14049) );
  AND2_X1 U8679 ( .A1(n12148), .A2(n14882), .ZN(n14687) );
  NAND2_X1 U8680 ( .A1(n7115), .A2(n7116), .ZN(n14053) );
  NAND2_X1 U8681 ( .A1(n8051), .A2(n8050), .ZN(n14070) );
  INV_X1 U8682 ( .A(n11591), .ZN(n14084) );
  NAND3_X2 U8683 ( .A1(n7864), .A2(n7863), .A3(n7862), .ZN(n14085) );
  NOR2_X1 U8684 ( .A1(n10850), .A2(n10413), .ZN(n14102) );
  AOI21_X1 U8685 ( .B1(n10650), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10649), .ZN(
        n10735) );
  AOI21_X1 U8686 ( .B1(n11965), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11960), .ZN(
        n11962) );
  NAND2_X1 U8687 ( .A1(n6794), .A2(n8424), .ZN(n6793) );
  AND2_X1 U8688 ( .A1(n8148), .A2(n8146), .ZN(n7323) );
  NAND2_X1 U8689 ( .A1(n14197), .A2(n8146), .ZN(n12440) );
  AOI21_X1 U8690 ( .B1(n12431), .B2(n14384), .A(n12430), .ZN(n14412) );
  OR2_X1 U8691 ( .A1(n14189), .A2(n14188), .ZN(n14415) );
  NAND2_X1 U8692 ( .A1(n14277), .A2(n6802), .ZN(n14217) );
  NAND2_X1 U8693 ( .A1(n14225), .A2(n8053), .ZN(n14213) );
  NAND2_X1 U8694 ( .A1(n14290), .A2(n7045), .ZN(n14282) );
  INV_X1 U8695 ( .A(n14444), .ZN(n14281) );
  AND2_X1 U8696 ( .A1(n14310), .A2(n8127), .ZN(n7314) );
  NAND2_X1 U8697 ( .A1(n8128), .A2(n8127), .ZN(n14324) );
  AND2_X1 U8698 ( .A1(n14356), .A2(n7989), .ZN(n7492) );
  NAND2_X1 U8699 ( .A1(n8125), .A2(n7300), .ZN(n7299) );
  NAND2_X1 U8700 ( .A1(n7341), .A2(n8121), .ZN(n12229) );
  NAND2_X1 U8701 ( .A1(n7768), .A2(n7767), .ZN(n12387) );
  INV_X1 U8702 ( .A(n14394), .ZN(n14322) );
  INV_X1 U8703 ( .A(n14172), .ZN(n11874) );
  NAND2_X1 U8704 ( .A1(n7281), .A2(n7285), .ZN(n11455) );
  NAND2_X1 U8705 ( .A1(n6496), .A2(n7286), .ZN(n7281) );
  NAND2_X1 U8706 ( .A1(n8197), .A2(n8193), .ZN(n11865) );
  INV_X1 U8707 ( .A(n14400), .ZN(n14325) );
  OR2_X1 U8708 ( .A1(n14432), .A2(n14431), .ZN(n14493) );
  OR2_X1 U8709 ( .A1(n14443), .A2(n14442), .ZN(n14495) );
  INV_X1 U8710 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7459) );
  NAND2_X1 U8711 ( .A1(n6790), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7599) );
  INV_X1 U8712 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U8713 ( .A1(n7621), .A2(n7622), .ZN(n12381) );
  XNOR2_X1 U8714 ( .A(n7630), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14528) );
  NAND2_X1 U8715 ( .A1(n7824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U8716 ( .A1(n7205), .A2(n7561), .ZN(n7806) );
  NAND2_X1 U8717 ( .A1(n7561), .A2(n7559), .ZN(n7804) );
  NAND2_X1 U8718 ( .A1(n7793), .A2(n7786), .ZN(n11574) );
  AND2_X1 U8719 ( .A1(n7647), .A2(n7646), .ZN(n14803) );
  INV_X1 U8720 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10518) );
  INV_X1 U8721 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10417) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10403) );
  INV_X1 U8723 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U8724 ( .A1(n7325), .A2(n7324), .ZN(n7673) );
  NAND2_X1 U8725 ( .A1(n7509), .A2(n6842), .ZN(n7661) );
  XNOR2_X1 U8726 ( .A(n7665), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U8727 ( .A1(n14537), .A2(n6916), .ZN(n15386) );
  OAI21_X1 U8728 ( .B1(n14538), .B2(n14539), .A(n6917), .ZN(n6916) );
  INV_X1 U8729 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6917) );
  XNOR2_X1 U8730 ( .A(n6898), .B(n8508), .ZN(n15380) );
  INV_X1 U8731 ( .A(n8509), .ZN(n6898) );
  NAND2_X1 U8732 ( .A1(n15380), .A2(n15379), .ZN(n15378) );
  XNOR2_X1 U8733 ( .A(n6692), .B(n8526), .ZN(n14731) );
  NAND2_X1 U8734 ( .A1(n14732), .A2(n8532), .ZN(n14735) );
  AND2_X1 U8735 ( .A1(n6911), .A2(n6909), .ZN(n14742) );
  NOR2_X1 U8736 ( .A1(n14744), .A2(n6910), .ZN(n6909) );
  INV_X1 U8737 ( .A(n6912), .ZN(n6910) );
  INV_X1 U8738 ( .A(n14563), .ZN(n6905) );
  AND2_X1 U8739 ( .A1(n12597), .A2(n6651), .ZN(n6650) );
  NOR2_X1 U8740 ( .A1(n6616), .A2(n6523), .ZN(n6651) );
  NAND2_X1 U8741 ( .A1(n6849), .A2(n10936), .ZN(n6848) );
  INV_X1 U8742 ( .A(n6751), .ZN(n12001) );
  INV_X1 U8743 ( .A(n6944), .ZN(n12003) );
  NAND2_X1 U8744 ( .A1(n7246), .A2(n7251), .ZN(n7245) );
  AOI21_X1 U8745 ( .B1(n9538), .B2(n7493), .A(n9537), .ZN(n9539) );
  NAND2_X1 U8746 ( .A1(n6700), .A2(n6696), .ZN(n13382) );
  NAND2_X1 U8747 ( .A1(n6699), .A2(n6697), .ZN(n6696) );
  NAND2_X1 U8748 ( .A1(n13380), .A2(n13379), .ZN(n6700) );
  NAND2_X1 U8749 ( .A1(n6670), .A2(n6667), .ZN(P2_U3236) );
  INV_X1 U8750 ( .A(n6668), .ZN(n6667) );
  NAND2_X1 U8751 ( .A1(n13406), .A2(n14665), .ZN(n6670) );
  OAI21_X1 U8752 ( .B1(n13407), .B2(n14668), .A(n6669), .ZN(n6668) );
  AND2_X1 U8753 ( .A1(n13414), .A2(n13413), .ZN(n13652) );
  AOI21_X1 U8754 ( .B1(n13396), .B2(n13688), .A(n6673), .ZN(n6672) );
  NOR2_X1 U8755 ( .A1(n15156), .A2(n13650), .ZN(n6673) );
  OR2_X1 U8756 ( .A1(n15156), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8757 ( .A1(n6718), .A2(n6717), .ZN(n6716) );
  AOI21_X1 U8758 ( .B1(n13396), .B2(n13749), .A(n6676), .ZN(n6675) );
  NOR2_X1 U8759 ( .A1(n15147), .A2(n13730), .ZN(n6676) );
  INV_X1 U8760 ( .A(n6729), .ZN(n6728) );
  AOI21_X1 U8761 ( .B1(n13732), .B2(n15147), .A(n7239), .ZN(n13734) );
  NAND2_X1 U8762 ( .A1(n7242), .A2(n7240), .ZN(n7239) );
  OR2_X1 U8763 ( .A1(n15147), .A2(n7241), .ZN(n7240) );
  CLKBUF_X2 U8764 ( .A(n14102), .Z(P1_U4016) );
  MUX2_X1 U8765 ( .A(n14174), .B(n14173), .S(n14172), .Z(n14176) );
  NAND2_X1 U8766 ( .A1(n8721), .A2(n14504), .ZN(n8192) );
  INV_X1 U8767 ( .A(n6897), .ZN(n15375) );
  INV_X1 U8768 ( .A(n6896), .ZN(n15382) );
  INV_X1 U8769 ( .A(n14546), .ZN(n14545) );
  INV_X1 U8770 ( .A(n6902), .ZN(n14552) );
  NAND2_X1 U8771 ( .A1(n14739), .A2(n14740), .ZN(n14738) );
  OR2_X1 U8772 ( .A1(n14532), .A2(n8549), .ZN(n7487) );
  AND2_X1 U8773 ( .A1(n12296), .A2(n6511), .ZN(n6505) );
  INV_X1 U8774 ( .A(n7867), .ZN(n7963) );
  INV_X1 U8775 ( .A(n8340), .ZN(n7452) );
  CLKBUF_X3 U8776 ( .A(n11847), .Z(n13933) );
  NAND2_X1 U8777 ( .A1(n7108), .A2(n13814), .ZN(n7115) );
  NOR2_X1 U8778 ( .A1(n6973), .A2(n6974), .ZN(n9620) );
  NAND2_X1 U8779 ( .A1(n8854), .A2(n8835), .ZN(n9509) );
  AND4_X1 U8780 ( .A1(n7588), .A2(n7589), .A3(n7583), .A4(n7093), .ZN(n6506)
         );
  INV_X2 U8781 ( .A(n9895), .ZN(n10036) );
  NAND2_X1 U8782 ( .A1(n9771), .A2(n11642), .ZN(n6507) );
  NAND2_X1 U8783 ( .A1(n9620), .A2(n6542), .ZN(n6508) );
  INV_X1 U8784 ( .A(n7003), .ZN(n7002) );
  NAND2_X1 U8785 ( .A1(n7006), .A2(n7004), .ZN(n7003) );
  INV_X1 U8786 ( .A(n13811), .ZN(n7113) );
  AND4_X1 U8787 ( .A1(n10161), .A2(n7073), .A3(n6587), .A4(n10164), .ZN(n6509)
         );
  INV_X1 U8788 ( .A(n11231), .ZN(n6921) );
  NAND2_X1 U8789 ( .A1(n7604), .A2(n7603), .ZN(n8342) );
  INV_X1 U8790 ( .A(n8342), .ZN(n6799) );
  AND2_X1 U8791 ( .A1(n10969), .A2(n11520), .ZN(n6510) );
  INV_X1 U8792 ( .A(n10168), .ZN(n11344) );
  OR2_X1 U8793 ( .A1(n6996), .A2(n6995), .ZN(n6511) );
  AND2_X1 U8794 ( .A1(n7597), .A2(n7350), .ZN(n6512) );
  AND2_X1 U8795 ( .A1(n7383), .A2(n7384), .ZN(n7382) );
  OR2_X2 U8796 ( .A1(n7103), .A2(n6531), .ZN(n6513) );
  AND2_X1 U8797 ( .A1(n6812), .A2(n6816), .ZN(n6514) );
  AND2_X1 U8798 ( .A1(n6577), .A2(n7210), .ZN(n6515) );
  NAND2_X1 U8799 ( .A1(n6742), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n14592) );
  AND2_X1 U8800 ( .A1(n6626), .A2(n7115), .ZN(n6516) );
  AND2_X1 U8801 ( .A1(n9470), .A2(n9469), .ZN(n13731) );
  INV_X1 U8802 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7397) );
  INV_X1 U8803 ( .A(n7035), .ZN(n7034) );
  OAI21_X1 U8804 ( .B1(n7922), .B2(n7036), .A(n8407), .ZN(n7035) );
  OR2_X1 U8805 ( .A1(n8423), .A2(n8428), .ZN(n6517) );
  AND2_X1 U8806 ( .A1(n10380), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6518) );
  AND2_X1 U8807 ( .A1(n7015), .A2(n10576), .ZN(n6519) );
  INV_X1 U8808 ( .A(n11248), .ZN(n12719) );
  AND4_X1 U8809 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n11248)
         );
  AND2_X1 U8810 ( .A1(n12309), .A2(n12307), .ZN(n6520) );
  AND2_X1 U8811 ( .A1(n10226), .A2(n10225), .ZN(n6521) );
  AND2_X1 U8812 ( .A1(n6737), .A2(n6740), .ZN(n6522) );
  INV_X1 U8813 ( .A(n10172), .ZN(n6978) );
  XNOR2_X1 U8814 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9658) );
  INV_X1 U8815 ( .A(n9658), .ZN(n7064) );
  AND2_X1 U8816 ( .A1(n12696), .A2(n12858), .ZN(n6523) );
  AND2_X1 U8817 ( .A1(n13054), .A2(n12990), .ZN(n9906) );
  INV_X1 U8818 ( .A(n9906), .ZN(n10134) );
  AND2_X1 U8819 ( .A1(n12143), .A2(n6622), .ZN(n6524) );
  AND2_X1 U8820 ( .A1(n7626), .A2(SI_23_), .ZN(n6525) );
  OAI21_X1 U8821 ( .B1(n6965), .B2(n12742), .A(n6961), .ZN(n6960) );
  OR2_X1 U8822 ( .A1(n15147), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6526) );
  OR2_X1 U8823 ( .A1(n15156), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6527) );
  NOR2_X2 U8824 ( .A1(n7841), .A2(n7840), .ZN(n7852) );
  AND3_X1 U8825 ( .A1(n8873), .A2(n8872), .A3(n8871), .ZN(n6528) );
  OR2_X1 U8826 ( .A1(n8538), .A2(n14746), .ZN(n6906) );
  AND2_X1 U8827 ( .A1(n14277), .A2(n6804), .ZN(n6529) );
  NAND2_X1 U8828 ( .A1(n7639), .A2(n7597), .ZN(n8159) );
  AND2_X1 U8829 ( .A1(n9419), .A2(n9420), .ZN(n6530) );
  OR2_X1 U8830 ( .A1(n13930), .A2(n7099), .ZN(n6531) );
  AND2_X1 U8831 ( .A1(n7007), .A2(n10148), .ZN(n6532) );
  NOR2_X1 U8832 ( .A1(n8748), .A2(n8747), .ZN(n8816) );
  INV_X1 U8833 ( .A(n14931), .ZN(n14676) );
  AND2_X1 U8834 ( .A1(n9348), .A2(n9347), .ZN(n6533) );
  NOR2_X1 U8835 ( .A1(n7452), .A2(n8338), .ZN(n6534) );
  INV_X1 U8836 ( .A(n8290), .ZN(n14337) );
  OR2_X1 U8837 ( .A1(n12675), .A2(n12909), .ZN(n6535) );
  AND2_X1 U8838 ( .A1(n15223), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8839 ( .A1(n7400), .A2(n10242), .ZN(n12987) );
  OR2_X1 U8840 ( .A1(n10115), .A2(n10294), .ZN(n6537) );
  AND2_X1 U8841 ( .A1(n9250), .A2(n9249), .ZN(n6538) );
  OR2_X1 U8842 ( .A1(n12831), .A2(n15241), .ZN(n6539) );
  OR2_X1 U8843 ( .A1(n7327), .A2(n9434), .ZN(n6540) );
  AND3_X1 U8844 ( .A1(n12494), .A2(n12490), .A3(n15180), .ZN(n6541) );
  INV_X1 U8845 ( .A(n14054), .ZN(n7114) );
  AND2_X1 U8846 ( .A1(n9796), .A2(n6851), .ZN(n6542) );
  XNOR2_X1 U8847 ( .A(n12479), .B(n12865), .ZN(n12876) );
  INV_X1 U8848 ( .A(n8254), .ZN(n7435) );
  NAND2_X1 U8849 ( .A1(n13201), .A2(n12531), .ZN(n13161) );
  NAND2_X1 U8850 ( .A1(n13144), .A2(n7275), .ZN(n13192) );
  INV_X1 U8851 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7653) );
  INV_X1 U8852 ( .A(n8329), .ZN(n7429) );
  OR2_X1 U8853 ( .A1(n7293), .A2(n9444), .ZN(n6543) );
  OR2_X1 U8854 ( .A1(n12569), .A2(n7249), .ZN(n6544) );
  OR2_X1 U8855 ( .A1(n12257), .A2(n12724), .ZN(n6545) );
  OR2_X1 U8856 ( .A1(n12581), .A2(n14623), .ZN(n6546) );
  INV_X1 U8857 ( .A(n12967), .ZN(n7029) );
  AND2_X1 U8858 ( .A1(n12228), .A2(n8401), .ZN(n6547) );
  OR2_X1 U8859 ( .A1(n12015), .A2(n12000), .ZN(n6548) );
  AND4_X1 U8860 ( .A1(n9762), .A2(n9761), .A3(n9760), .A4(n9759), .ZN(n11816)
         );
  INV_X1 U8861 ( .A(n10152), .ZN(n12852) );
  INV_X1 U8862 ( .A(n13554), .ZN(n13697) );
  AND2_X1 U8863 ( .A1(n9108), .A2(n9107), .ZN(n13554) );
  OR2_X1 U8864 ( .A1(n6905), .A2(n15038), .ZN(n6549) );
  INV_X1 U8865 ( .A(n8238), .ZN(n7438) );
  OR2_X1 U8866 ( .A1(n8517), .A2(n8518), .ZN(n6550) );
  OR2_X1 U8867 ( .A1(n10961), .A2(n10945), .ZN(n6551) );
  AND2_X1 U8868 ( .A1(n8355), .A2(n8354), .ZN(n14407) );
  INV_X1 U8869 ( .A(n14407), .ZN(n14184) );
  INV_X1 U8870 ( .A(n8234), .ZN(n7440) );
  NAND2_X1 U8871 ( .A1(n14420), .A2(n8063), .ZN(n6552) );
  AND2_X1 U8872 ( .A1(n8135), .A2(n8134), .ZN(n6553) );
  AND2_X1 U8873 ( .A1(n13850), .A2(n13848), .ZN(n6554) );
  AND2_X1 U8874 ( .A1(n11902), .A2(n14922), .ZN(n6555) );
  AND2_X1 U8875 ( .A1(n10703), .A2(n11306), .ZN(n6556) );
  INV_X1 U8876 ( .A(n10214), .ZN(n15300) );
  AND2_X1 U8877 ( .A1(n7485), .A2(n7414), .ZN(n6557) );
  NOR2_X1 U8878 ( .A1(n15214), .A2(n6536), .ZN(n6558) );
  AND2_X1 U8879 ( .A1(n11939), .A2(n11799), .ZN(n6559) );
  INV_X1 U8880 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7395) );
  AND2_X1 U8881 ( .A1(n7017), .A2(n10155), .ZN(n6560) );
  NOR2_X1 U8882 ( .A1(n13814), .A2(n7114), .ZN(n6561) );
  OR2_X1 U8883 ( .A1(n13812), .A2(n13977), .ZN(n8280) );
  AND2_X1 U8884 ( .A1(n10142), .A2(n10141), .ZN(n12936) );
  NOR2_X1 U8885 ( .A1(n11332), .A2(n9325), .ZN(n6562) );
  NOR2_X1 U8886 ( .A1(n14470), .A2(n14363), .ZN(n6563) );
  NOR2_X1 U8887 ( .A1(n13554), .A2(n13538), .ZN(n6564) );
  AND2_X1 U8888 ( .A1(n7374), .A2(n7379), .ZN(n6565) );
  AND2_X1 U8889 ( .A1(n13554), .A2(n13538), .ZN(n6566) );
  INV_X1 U8890 ( .A(n9241), .ZN(n7218) );
  AND2_X1 U8891 ( .A1(n12603), .A2(n12704), .ZN(n6567) );
  INV_X1 U8892 ( .A(n10130), .ZN(n6995) );
  AND2_X1 U8893 ( .A1(n13505), .A2(n13483), .ZN(n6568) );
  AND2_X1 U8894 ( .A1(n7322), .A2(n7321), .ZN(n6569) );
  AND2_X1 U8895 ( .A1(n11854), .A2(n11596), .ZN(n6570) );
  OR2_X1 U8896 ( .A1(n10194), .A2(n9589), .ZN(n6571) );
  NAND2_X1 U8897 ( .A1(n14242), .A2(n8141), .ZN(n6572) );
  NAND2_X1 U8898 ( .A1(n7797), .A2(n7592), .ZN(n6573) );
  INV_X1 U8899 ( .A(n6808), .ZN(n6807) );
  NAND2_X1 U8900 ( .A1(n14395), .A2(n6809), .ZN(n6808) );
  AND2_X1 U8901 ( .A1(n11804), .A2(n11803), .ZN(n6574) );
  INV_X1 U8902 ( .A(n7046), .ZN(n7045) );
  NAND2_X1 U8903 ( .A1(n14283), .A2(n8015), .ZN(n7046) );
  AND2_X1 U8904 ( .A1(n9232), .A2(n8978), .ZN(n11613) );
  AND2_X1 U8905 ( .A1(n12403), .A2(n12709), .ZN(n6575) );
  AND2_X1 U8906 ( .A1(n7033), .A2(n7930), .ZN(n6576) );
  AND2_X1 U8907 ( .A1(n13532), .A2(n13531), .ZN(n6577) );
  INV_X1 U8908 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9590) );
  INV_X1 U8909 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7831) );
  AND2_X1 U8910 ( .A1(n7541), .A2(n10401), .ZN(n6578) );
  AND2_X1 U8911 ( .A1(n12463), .A2(n12706), .ZN(n6579) );
  XNOR2_X1 U8912 ( .A(n8791), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9216) );
  AND2_X1 U8913 ( .A1(n10343), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6580) );
  AND2_X1 U8914 ( .A1(n11244), .A2(n11248), .ZN(n6581) );
  NOR2_X1 U8915 ( .A1(n13505), .A2(n13512), .ZN(n6582) );
  INV_X1 U8916 ( .A(n7297), .ZN(n7296) );
  OR2_X1 U8917 ( .A1(n8126), .A2(n7298), .ZN(n7297) );
  OR2_X1 U8918 ( .A1(n7230), .A2(n7228), .ZN(n6583) );
  NAND2_X1 U8919 ( .A1(n10116), .A2(n10115), .ZN(n6584) );
  AND2_X1 U8920 ( .A1(n7222), .A2(n9504), .ZN(n6585) );
  INV_X1 U8921 ( .A(n7287), .ZN(n7286) );
  NOR2_X1 U8922 ( .A1(n14850), .A2(n11591), .ZN(n7287) );
  NAND2_X1 U8923 ( .A1(n10161), .A2(n10163), .ZN(n6586) );
  AND3_X1 U8924 ( .A1(n10266), .A2(n12842), .A3(n7071), .ZN(n6587) );
  NAND2_X1 U8925 ( .A1(n9221), .A2(n12548), .ZN(n10664) );
  OR2_X1 U8926 ( .A1(n8443), .A2(n7482), .ZN(n6588) );
  INV_X1 U8927 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8815) );
  XNOR2_X1 U8928 ( .A(n8833), .B(P2_IR_REG_1__SCAN_IN), .ZN(n14944) );
  AND3_X1 U8929 ( .A1(n8420), .A2(n7172), .A3(n8430), .ZN(n6589) );
  INV_X1 U8930 ( .A(n9319), .ZN(n7308) );
  AND2_X1 U8931 ( .A1(n6797), .A2(n6795), .ZN(n6590) );
  AND2_X1 U8932 ( .A1(n7331), .A2(n9430), .ZN(n6591) );
  AND2_X1 U8933 ( .A1(n12223), .A2(n8121), .ZN(n6592) );
  AND2_X1 U8934 ( .A1(n11306), .A2(n13266), .ZN(n6593) );
  AND2_X1 U8935 ( .A1(n7423), .A2(n9587), .ZN(n6594) );
  AND2_X1 U8936 ( .A1(n7461), .A2(n7459), .ZN(n6595) );
  AND2_X1 U8937 ( .A1(n8441), .A2(n8440), .ZN(n6596) );
  AND2_X1 U8938 ( .A1(n11097), .A2(n10970), .ZN(n6597) );
  AND2_X1 U8939 ( .A1(n6905), .A2(n15038), .ZN(n6598) );
  NAND2_X1 U8940 ( .A1(n8506), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n6599) );
  OAI22_X1 U8941 ( .A1(n6878), .A2(n6877), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_21__SCAN_IN), .ZN(n6874) );
  AND2_X1 U8942 ( .A1(n14290), .A2(n8015), .ZN(n6600) );
  AND2_X1 U8943 ( .A1(n12532), .A2(n12531), .ZN(n6601) );
  AND2_X1 U8944 ( .A1(n6906), .A2(n6905), .ZN(n6602) );
  AND2_X1 U8945 ( .A1(n12553), .A2(n12552), .ZN(n6603) );
  OR2_X1 U8946 ( .A1(n7435), .A2(n8253), .ZN(n6604) );
  OR2_X1 U8947 ( .A1(n8244), .A2(n8242), .ZN(n6605) );
  AND2_X1 U8948 ( .A1(n14337), .A2(n7989), .ZN(n6606) );
  AND2_X1 U8949 ( .A1(n7246), .A2(n6544), .ZN(n6607) );
  AND2_X1 U8950 ( .A1(n7397), .A2(n6851), .ZN(n6608) );
  AND2_X1 U8951 ( .A1(n7411), .A2(n6535), .ZN(n6609) );
  AND2_X1 U8952 ( .A1(n7194), .A2(n7643), .ZN(n6610) );
  AND2_X1 U8953 ( .A1(n6506), .A2(n7460), .ZN(n6611) );
  INV_X1 U8954 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n10107) );
  OR2_X1 U8955 ( .A1(n6533), .A2(n7344), .ZN(n6612) );
  INV_X1 U8956 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8743) );
  AND2_X1 U8957 ( .A1(n7215), .A2(n7212), .ZN(n7211) );
  NAND2_X1 U8958 ( .A1(n7332), .A2(n9432), .ZN(n6613) );
  NAND2_X1 U8959 ( .A1(n7105), .A2(n13928), .ZN(n6614) );
  INV_X1 U8960 ( .A(n6739), .ZN(n6738) );
  NAND2_X1 U8961 ( .A1(n11534), .A2(n10970), .ZN(n6739) );
  AND2_X1 U8962 ( .A1(n10126), .A2(n10125), .ZN(n11991) );
  INV_X1 U8963 ( .A(n11991), .ZN(n6981) );
  INV_X1 U8964 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7058) );
  OAI21_X1 U8965 ( .B1(n9853), .B2(n7078), .A(n9874), .ZN(n7077) );
  INV_X1 U8966 ( .A(n12143), .ZN(n6895) );
  NAND2_X1 U8967 ( .A1(n7299), .A2(n8399), .ZN(n14344) );
  XNOR2_X1 U8968 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9643) );
  INV_X1 U8969 ( .A(n9643), .ZN(n7061) );
  XNOR2_X1 U8970 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9724) );
  INV_X1 U8971 ( .A(n9724), .ZN(n6780) );
  INV_X1 U8972 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n6851) );
  INV_X1 U8973 ( .A(n10124), .ZN(n6980) );
  NAND2_X1 U8974 ( .A1(n7591), .A2(n7590), .ZN(n7092) );
  NAND2_X1 U8975 ( .A1(n13224), .A2(n12523), .ZN(n13152) );
  NAND2_X1 U8976 ( .A1(n12508), .A2(n13242), .ZN(n14638) );
  INV_X1 U8977 ( .A(n14420), .ZN(n6801) );
  AND3_X1 U8978 ( .A1(n7588), .A2(n7589), .A3(n7583), .ZN(n6615) );
  AND2_X1 U8979 ( .A1(n12857), .A2(n15186), .ZN(n6616) );
  INV_X1 U8980 ( .A(n7026), .ZN(n7025) );
  NOR2_X1 U8981 ( .A1(n12951), .A2(n7027), .ZN(n7026) );
  OR2_X1 U8982 ( .A1(n12222), .A2(n12179), .ZN(n6617) );
  AND2_X1 U8983 ( .A1(n7564), .A2(n7184), .ZN(n6618) );
  INV_X1 U8984 ( .A(n6933), .ZN(n13567) );
  INV_X1 U8985 ( .A(n12933), .ZN(n12909) );
  AND3_X1 U8986 ( .A1(n9997), .A2(n9996), .A3(n9995), .ZN(n12933) );
  NAND2_X1 U8987 ( .A1(n14389), .A2(n6806), .ZN(n6810) );
  INV_X1 U8988 ( .A(n7077), .ZN(n7076) );
  AND2_X1 U8989 ( .A1(n9787), .A2(n10228), .ZN(n6619) );
  AND2_X1 U8990 ( .A1(n12650), .A2(n12707), .ZN(n6620) );
  OR2_X1 U8991 ( .A1(n7091), .A2(n7092), .ZN(n6621) );
  NAND2_X1 U8992 ( .A1(n12222), .A2(n12179), .ZN(n6622) );
  AND2_X1 U8993 ( .A1(n10518), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6623) );
  AND2_X1 U8994 ( .A1(n9568), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6624) );
  NOR2_X1 U8995 ( .A1(n10133), .A2(n10294), .ZN(n6625) );
  AND2_X1 U8996 ( .A1(n7116), .A2(n7114), .ZN(n6626) );
  NOR2_X1 U8997 ( .A1(n12130), .A2(n12129), .ZN(n6627) );
  INV_X1 U8998 ( .A(n12659), .ZN(n12704) );
  AND3_X1 U8999 ( .A1(n9619), .A2(n9618), .A3(n9617), .ZN(n12659) );
  AND2_X1 U9000 ( .A1(n7420), .A2(n6622), .ZN(n6628) );
  AND2_X1 U9001 ( .A1(n7039), .A2(n7037), .ZN(n6629) );
  AND2_X1 U9002 ( .A1(n7182), .A2(n7566), .ZN(n6630) );
  INV_X1 U9003 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8863) );
  INV_X1 U9004 ( .A(n12785), .ZN(n12798) );
  INV_X1 U9005 ( .A(n9518), .ZN(n7152) );
  OAI21_X1 U9006 ( .B1(n12172), .B2(n7361), .A(n7358), .ZN(n12279) );
  NAND2_X1 U9007 ( .A1(n7780), .A2(n7779), .ZN(n14475) );
  INV_X1 U9008 ( .A(n14475), .ZN(n6809) );
  BUF_X1 U9009 ( .A(n9215), .Z(n8803) );
  AND2_X1 U9010 ( .A1(n13368), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6631) );
  INV_X1 U9011 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7056) );
  NOR2_X1 U9012 ( .A1(n11925), .A2(n12115), .ZN(n6632) );
  NAND2_X1 U9013 ( .A1(n12760), .A2(n12785), .ZN(n6965) );
  INV_X1 U9014 ( .A(n13707), .ZN(n6934) );
  NAND2_X1 U9015 ( .A1(n15157), .A2(n11812), .ZN(n12616) );
  NAND2_X1 U9016 ( .A1(n7774), .A2(n7773), .ZN(n14710) );
  INV_X1 U9017 ( .A(n14710), .ZN(n6816) );
  NAND2_X1 U9018 ( .A1(n12131), .A2(n12128), .ZN(n7273) );
  NOR2_X1 U9019 ( .A1(n8748), .A2(n8740), .ZN(n8755) );
  INV_X1 U9020 ( .A(n7354), .ZN(n10575) );
  AND2_X1 U9021 ( .A1(n6929), .A2(n6930), .ZN(n6633) );
  OR2_X1 U9022 ( .A1(n13361), .A2(n13362), .ZN(n6634) );
  AND2_X1 U9023 ( .A1(n12742), .A2(n12798), .ZN(n6635) );
  OR2_X1 U9024 ( .A1(n6787), .A2(n6785), .ZN(n6636) );
  NAND2_X1 U9025 ( .A1(n10189), .A2(n10188), .ZN(n6637) );
  OR2_X1 U9026 ( .A1(n7626), .A2(SI_23_), .ZN(n6638) );
  NAND2_X1 U9027 ( .A1(n12138), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U9028 ( .A1(n7573), .A2(n12169), .ZN(n6640) );
  INV_X1 U9029 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11573) );
  INV_X1 U9030 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11357) );
  AND2_X1 U9031 ( .A1(n6639), .A2(n9972), .ZN(n6641) );
  INV_X1 U9032 ( .A(n6965), .ZN(n6964) );
  INV_X1 U9033 ( .A(n10896), .ZN(n7088) );
  INV_X1 U9034 ( .A(n11701), .ZN(n6932) );
  AND2_X1 U9035 ( .A1(n7391), .A2(n11164), .ZN(n7390) );
  AND2_X2 U9036 ( .A1(n9273), .A2(n15089), .ZN(n15147) );
  INV_X1 U9037 ( .A(n14583), .ZN(n12803) );
  OAI21_X1 U9038 ( .B1(n11260), .B2(n7122), .A(n7121), .ZN(n11174) );
  INV_X1 U9039 ( .A(n12200), .ZN(n6815) );
  INV_X1 U9040 ( .A(n11228), .ZN(n6922) );
  AND2_X1 U9041 ( .A1(n15147), .A2(n15100), .ZN(n13749) );
  INV_X1 U9042 ( .A(n10668), .ZN(n6671) );
  AND2_X1 U9043 ( .A1(n6947), .A2(n6955), .ZN(n6642) );
  AND2_X1 U9044 ( .A1(n7161), .A2(n8854), .ZN(n6643) );
  AND2_X1 U9045 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n10093), .ZN(n6644) );
  OAI21_X1 U9046 ( .B1(n10074), .B2(n7082), .A(n10073), .ZN(n7081) );
  INV_X1 U9047 ( .A(n7079), .ZN(n6767) );
  NOR2_X1 U9048 ( .A1(n7081), .A2(n7080), .ZN(n7079) );
  OR2_X1 U9049 ( .A1(n10208), .A2(n10207), .ZN(n6645) );
  INV_X1 U9050 ( .A(n12794), .ZN(n6958) );
  AND2_X1 U9051 ( .A1(n11338), .A2(n10576), .ZN(n15311) );
  INV_X1 U9052 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7503) );
  INV_X1 U9053 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6723) );
  INV_X1 U9054 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6711) );
  INV_X1 U9055 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6774) );
  AOI21_X1 U9056 ( .B1(n6688), .B2(n9268), .A(n6685), .ZN(n13657) );
  OAI21_X1 U9057 ( .B1(n6498), .B2(n7503), .A(n7502), .ZN(n7506) );
  NAND2_X1 U9058 ( .A1(n7683), .A2(n7514), .ZN(n7691) );
  NAND2_X1 U9059 ( .A1(n7206), .A2(n7561), .ZN(n7810) );
  NAND2_X1 U9060 ( .A1(n6648), .A2(n6610), .ZN(n7632) );
  NAND2_X1 U9061 ( .A1(n7544), .A2(n7195), .ZN(n6648) );
  INV_X1 U9062 ( .A(n6706), .ZN(n6705) );
  NAND2_X1 U9063 ( .A1(n6707), .A2(n14734), .ZN(n14739) );
  NAND2_X1 U9064 ( .A1(n14729), .A2(n8528), .ZN(n8531) );
  NAND2_X1 U9065 ( .A1(n10280), .A2(n10279), .ZN(n10574) );
  AOI21_X1 U9066 ( .B1(n12667), .B2(n12666), .A(n12466), .ZN(n12627) );
  INV_X1 U9067 ( .A(n12616), .ZN(n6654) );
  AOI21_X1 U9068 ( .B1(n10583), .B2(n10582), .A(n10584), .ZN(n10840) );
  NAND2_X1 U9069 ( .A1(n6969), .A2(n9584), .ZN(n6968) );
  OAI22_X1 U9070 ( .A1(n11160), .A2(n11159), .B1(n12722), .B2(n11158), .ZN(
        n15173) );
  NAND2_X2 U9071 ( .A1(n12458), .A2(n12457), .ZN(n12681) );
  NAND2_X2 U9072 ( .A1(n12282), .A2(n12281), .ZN(n12367) );
  AOI21_X2 U9073 ( .B1(n11806), .B2(n11805), .A(n6574), .ZN(n15183) );
  NAND2_X1 U9074 ( .A1(n6652), .A2(n6650), .ZN(P3_U3154) );
  NAND2_X1 U9075 ( .A1(n6656), .A2(n15180), .ZN(n6652) );
  NAND2_X1 U9076 ( .A1(n11943), .A2(n11942), .ZN(n12172) );
  NAND2_X1 U9077 ( .A1(n6689), .A2(n12659), .ZN(n12598) );
  NAND2_X1 U9078 ( .A1(n12594), .A2(n12595), .ZN(n6656) );
  NAND2_X1 U9079 ( .A1(n7363), .A2(n7362), .ZN(n12667) );
  NAND3_X1 U9080 ( .A1(n7009), .A2(n7008), .A3(n6659), .ZN(n10184) );
  NAND2_X1 U9081 ( .A1(n9575), .A2(n9574), .ZN(n9974) );
  NAND2_X1 U9082 ( .A1(n6944), .A2(n6943), .ZN(n12256) );
  NAND2_X1 U9083 ( .A1(n6939), .A2(n6938), .ZN(n11824) );
  NAND2_X1 U9084 ( .A1(n6757), .A2(n9572), .ZN(n9573) );
  NAND2_X1 U9085 ( .A1(n15262), .A2(n11512), .ZN(n11514) );
  XNOR2_X1 U9086 ( .A(n11514), .B(n15284), .ZN(n15271) );
  OAI21_X1 U9087 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(n14519), .A(n10031), 
        .ZN(n10045) );
  INV_X1 U9088 ( .A(n10988), .ZN(n6748) );
  NOR2_X1 U9089 ( .A1(n10972), .A2(n10971), .ZN(n11509) );
  NAND2_X1 U9090 ( .A1(n9705), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n6941) );
  INV_X1 U9091 ( .A(n7015), .ZN(n7012) );
  XNOR2_X1 U9092 ( .A(n10963), .B(n10962), .ZN(n15196) );
  NAND2_X1 U9093 ( .A1(n9555), .A2(n9554), .ZN(n9779) );
  INV_X1 U9094 ( .A(n9565), .ZN(n6769) );
  NAND2_X1 U9095 ( .A1(n9570), .A2(n9569), .ZN(n9910) );
  NAND2_X1 U9096 ( .A1(n6758), .A2(n7055), .ZN(n9942) );
  NAND2_X1 U9097 ( .A1(n9571), .A2(n7057), .ZN(n9925) );
  AOI21_X1 U9098 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10030) );
  NAND2_X1 U9099 ( .A1(n6771), .A2(n6770), .ZN(n9890) );
  NAND2_X1 U9100 ( .A1(n6558), .A2(n10966), .ZN(n6936) );
  NAND2_X1 U9101 ( .A1(n6937), .A2(n6936), .ZN(n15234) );
  AOI21_X1 U9102 ( .B1(n10185), .B2(n15327), .A(n11741), .ZN(n6846) );
  INV_X1 U9103 ( .A(n10160), .ZN(n6660) );
  NAND2_X1 U9104 ( .A1(n13619), .A2(n13618), .ZN(n13617) );
  NAND2_X1 U9105 ( .A1(n13416), .A2(n6832), .ZN(n13415) );
  OAI21_X2 U9106 ( .B1(n13573), .B2(n7119), .A(n7117), .ZN(n13529) );
  OAI21_X1 U9107 ( .B1(n11914), .B2(n9026), .A(n9025), .ZN(n14659) );
  AOI21_X1 U9108 ( .B1(n7704), .B2(n7520), .A(n7519), .ZN(n7715) );
  AND2_X2 U9109 ( .A1(n8787), .A2(n8788), .ZN(n8792) );
  NAND2_X1 U9110 ( .A1(n11437), .A2(n11436), .ZN(n11664) );
  NAND2_X1 U9111 ( .A1(n6662), .A2(n7261), .ZN(n11374) );
  NAND3_X1 U9112 ( .A1(n7254), .A2(n7259), .A3(n7253), .ZN(n6662) );
  XNOR2_X2 U9113 ( .A(n10879), .B(n10663), .ZN(n10665) );
  NAND4_X2 U9114 ( .A1(n8725), .A2(n8863), .A3(n8879), .A4(n8724), .ZN(n8892)
         );
  INV_X1 U9115 ( .A(n7255), .ZN(n10824) );
  INV_X1 U9116 ( .A(n10820), .ZN(n6663) );
  NAND3_X1 U9117 ( .A1(n8101), .A2(n7346), .A3(n7345), .ZN(n11562) );
  NAND2_X1 U9118 ( .A1(n8415), .A2(n14275), .ZN(n7309) );
  NAND2_X1 U9119 ( .A1(n7544), .A2(SI_14_), .ZN(n7199) );
  NAND2_X1 U9120 ( .A1(n7167), .A2(n7165), .ZN(n6666) );
  NAND3_X1 U9121 ( .A1(n6513), .A2(n7096), .A3(n6614), .ZN(n13939) );
  NAND2_X1 U9122 ( .A1(n13773), .A2(n9468), .ZN(n9182) );
  NAND2_X1 U9123 ( .A1(n7517), .A2(n7691), .ZN(n7704) );
  NAND2_X1 U9124 ( .A1(n13915), .A2(n13914), .ZN(n13913) );
  NAND2_X2 U9125 ( .A1(n13810), .A2(n13809), .ZN(n14686) );
  OAI21_X2 U9126 ( .B1(n14686), .B2(n6561), .A(n7109), .ZN(n13974) );
  NAND2_X2 U9127 ( .A1(n13466), .A2(n13465), .ZN(n13464) );
  NOR2_X1 U9128 ( .A1(n10341), .A2(n9140), .ZN(n8882) );
  INV_X1 U9129 ( .A(n7669), .ZN(n6679) );
  XNOR2_X2 U9130 ( .A(n11231), .B(n13268), .ZN(n11225) );
  OAI211_X1 U9131 ( .C1(n13398), .C2(n13724), .A(n7146), .B(n15156), .ZN(n6845) );
  NOR2_X2 U9132 ( .A1(n9125), .A2(n7480), .ZN(n13519) );
  NAND3_X2 U9133 ( .A1(n8771), .A2(n8736), .A3(n8737), .ZN(n8748) );
  NAND2_X1 U9134 ( .A1(n9584), .A2(n6608), .ZN(n6972) );
  NAND2_X1 U9135 ( .A1(n10244), .A2(n10243), .ZN(n12974) );
  NAND2_X1 U9136 ( .A1(n10236), .A2(n7421), .ZN(n7420) );
  AOI21_X1 U9137 ( .B1(n10264), .B2(n15317), .A(n10263), .ZN(n12587) );
  NOR2_X2 U9138 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8725) );
  INV_X1 U9139 ( .A(n8898), .ZN(n8861) );
  XNOR2_X2 U9140 ( .A(n6477), .B(n6671), .ZN(n10639) );
  NOR2_X1 U9141 ( .A1(n13529), .A2(n13534), .ZN(n9125) );
  OAI21_X1 U9142 ( .B1(n13519), .B2(n7141), .A(n7140), .ZN(n7144) );
  NAND2_X2 U9143 ( .A1(n8875), .A2(n10344), .ZN(n8898) );
  NAND2_X1 U9144 ( .A1(n7175), .A2(n7539), .ZN(n7764) );
  NAND2_X1 U9145 ( .A1(n6674), .A2(n6672), .ZN(P2_U3529) );
  OR2_X1 U9146 ( .A1(n13729), .A2(n15154), .ZN(n6674) );
  NAND2_X1 U9147 ( .A1(n6677), .A2(n6675), .ZN(P2_U3497) );
  OR2_X1 U9148 ( .A1(n13729), .A2(n15145), .ZN(n6677) );
  NOR2_X2 U9149 ( .A1(n13656), .A2(n13446), .ZN(n13429) );
  INV_X1 U9150 ( .A(n14656), .ZN(n6678) );
  OAI21_X2 U9151 ( .B1(n7667), .B2(n7513), .A(n7512), .ZN(n7683) );
  NAND3_X1 U9152 ( .A1(n6842), .A2(n7659), .A3(n7509), .ZN(n7663) );
  NAND2_X1 U9153 ( .A1(n8421), .A2(n6589), .ZN(n7171) );
  OAI21_X1 U9154 ( .B1(n8312), .B2(n8311), .A(n6682), .ZN(n8315) );
  NAND2_X1 U9155 ( .A1(n6684), .A2(n6683), .ZN(n6682) );
  NAND2_X1 U9156 ( .A1(n8312), .A2(n8311), .ZN(n6684) );
  AOI21_X1 U9157 ( .B1(n7467), .B2(n7470), .A(n7466), .ZN(n7465) );
  NAND4_X1 U9158 ( .A1(n6588), .A2(n6517), .A3(n8439), .A4(n7164), .ZN(n6712)
         );
  NAND3_X1 U9159 ( .A1(n6825), .A2(n9252), .A3(n6823), .ZN(n13459) );
  NOR2_X1 U9160 ( .A1(n6972), .A2(n6974), .ZN(n6971) );
  NAND2_X1 U9161 ( .A1(n7378), .A2(n7377), .ZN(n7376) );
  NAND2_X1 U9162 ( .A1(n12598), .A2(n12653), .ZN(n12478) );
  INV_X1 U9163 ( .A(n12599), .ZN(n6689) );
  NAND2_X1 U9164 ( .A1(n15183), .A2(n15182), .ZN(n15181) );
  NAND2_X1 U9165 ( .A1(n7387), .A2(n7386), .ZN(n11806) );
  AND3_X2 U9166 ( .A1(n6971), .A2(n6970), .A3(n9580), .ZN(n10195) );
  NAND3_X1 U9167 ( .A1(n11082), .A2(n10168), .A3(n10222), .ZN(n11341) );
  NAND2_X1 U9168 ( .A1(n11079), .A2(n10221), .ZN(n11082) );
  OAI211_X2 U9169 ( .C1(n10058), .C2(n10394), .A(n9676), .B(n9675), .ZN(n10812) );
  NAND2_X1 U9170 ( .A1(n13171), .A2(n13173), .ZN(n13172) );
  INV_X1 U9171 ( .A(n13408), .ZN(n6832) );
  OAI21_X1 U9172 ( .B1(n7221), .B2(n6832), .A(n6829), .ZN(n6833) );
  NAND2_X1 U9173 ( .A1(n7406), .A2(n7404), .ZN(n12886) );
  NAND2_X1 U9174 ( .A1(n6728), .A2(n6705), .ZN(P2_U3496) );
  NAND2_X1 U9175 ( .A1(n7200), .A2(n7199), .ZN(n7651) );
  NAND2_X1 U9176 ( .A1(n8287), .A2(n8286), .ZN(n7454) );
  NAND2_X1 U9177 ( .A1(n8321), .A2(n8322), .ZN(n8320) );
  NAND2_X1 U9178 ( .A1(n7442), .A2(n7446), .ZN(n8321) );
  NAND2_X1 U9179 ( .A1(n7427), .A2(n7426), .ZN(n8331) );
  NAND2_X1 U9180 ( .A1(n6712), .A2(n8444), .ZN(n7163) );
  INV_X1 U9181 ( .A(n7206), .ZN(n7205) );
  NAND2_X1 U9182 ( .A1(n6690), .A2(n9272), .ZN(P2_U3528) );
  NAND2_X1 U9183 ( .A1(n6845), .A2(n6844), .ZN(n6690) );
  NAND2_X1 U9184 ( .A1(n9129), .A2(n7567), .ZN(n7625) );
  NAND2_X1 U9185 ( .A1(n7559), .A2(n7560), .ZN(n7206) );
  AOI21_X1 U9186 ( .B1(n7123), .B2(n11262), .A(n6593), .ZN(n7121) );
  NAND2_X1 U9187 ( .A1(n14743), .A2(n14744), .ZN(n8533) );
  NAND2_X1 U9188 ( .A1(n6911), .A2(n6912), .ZN(n14743) );
  NAND2_X1 U9189 ( .A1(n8495), .A2(n8494), .ZN(n6691) );
  NOR2_X1 U9190 ( .A1(n14549), .A2(n8523), .ZN(n14553) );
  NOR2_X1 U9191 ( .A1(n14999), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14998) );
  NAND2_X1 U9192 ( .A1(n13335), .A2(n13349), .ZN(n6694) );
  INV_X1 U9193 ( .A(n13336), .ZN(n6695) );
  NAND2_X1 U9194 ( .A1(n7812), .A2(n7564), .ZN(n7181) );
  NAND2_X1 U9195 ( .A1(n7183), .A2(n7567), .ZN(n9127) );
  NAND2_X1 U9196 ( .A1(n7663), .A2(n7509), .ZN(n7667) );
  NAND2_X2 U9197 ( .A1(n7568), .A2(SI_24_), .ZN(n7571) );
  INV_X1 U9198 ( .A(n7166), .ZN(n7167) );
  INV_X1 U9199 ( .A(n11175), .ZN(n6837) );
  INV_X1 U9200 ( .A(n14659), .ZN(n6704) );
  OR2_X1 U9201 ( .A1(n8755), .A2(n8741), .ZN(n8742) );
  INV_X1 U9202 ( .A(n7123), .ZN(n7122) );
  NAND2_X1 U9203 ( .A1(n13476), .A2(n13478), .ZN(n13475) );
  OR2_X1 U9204 ( .A1(n13267), .A2(n11268), .ZN(n8897) );
  NAND2_X1 U9205 ( .A1(n8936), .A2(n8935), .ZN(n11383) );
  NAND2_X1 U9206 ( .A1(n8967), .A2(n8966), .ZN(n11614) );
  NAND2_X1 U9207 ( .A1(n8498), .A2(n8497), .ZN(n8450) );
  NAND2_X1 U9208 ( .A1(n7280), .A2(n7279), .ZN(n11469) );
  NAND2_X1 U9209 ( .A1(n14553), .A2(n14554), .ZN(n6901) );
  NOR2_X1 U9210 ( .A1(n14543), .A2(n14542), .ZN(n14541) );
  AND2_X2 U9211 ( .A1(n6512), .A2(n7639), .ZN(n8155) );
  AND2_X1 U9212 ( .A1(n11459), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U9213 ( .A1(n15173), .A2(n7390), .ZN(n7387) );
  NAND2_X1 U9214 ( .A1(n12627), .A2(n12628), .ZN(n12626) );
  NAND2_X1 U9215 ( .A1(n7368), .A2(n7369), .ZN(n12452) );
  NAND2_X1 U9216 ( .A1(n10181), .A2(n10180), .ZN(n7354) );
  NAND2_X1 U9217 ( .A1(n9624), .A2(n9944), .ZN(n10106) );
  NAND2_X1 U9218 ( .A1(n12595), .A2(n6541), .ZN(n12498) );
  NAND2_X1 U9219 ( .A1(n12758), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U9220 ( .A1(n12736), .A2(n12741), .ZN(n12757) );
  NAND2_X1 U9221 ( .A1(n15254), .A2(n15255), .ZN(n6709) );
  NAND2_X1 U9222 ( .A1(n13142), .A2(n13145), .ZN(n13143) );
  NAND2_X1 U9223 ( .A1(n8443), .A2(n7483), .ZN(n8439) );
  NAND2_X1 U9224 ( .A1(n8346), .A2(n8347), .ZN(n8443) );
  NAND2_X1 U9225 ( .A1(n7726), .A2(n7526), .ZN(n7732) );
  NOR2_X1 U9226 ( .A1(n7508), .A2(n10394), .ZN(n7659) );
  INV_X1 U9227 ( .A(n7570), .ZN(n7165) );
  NAND2_X1 U9228 ( .A1(n7187), .A2(n7185), .ZN(n7558) );
  AOI21_X1 U9229 ( .B1(n13732), .B2(n15156), .A(n6716), .ZN(n13654) );
  OR2_X1 U9230 ( .A1(n15156), .A2(n9200), .ZN(n6717) );
  NAND2_X1 U9231 ( .A1(n13733), .A2(n13688), .ZN(n6718) );
  INV_X1 U9232 ( .A(n6973), .ZN(n6969) );
  INV_X1 U9233 ( .A(n13891), .ZN(n7104) );
  NOR2_X1 U9234 ( .A1(n6968), .A2(n6974), .ZN(n9585) );
  NAND2_X1 U9235 ( .A1(n7357), .A2(n7355), .ZN(n12282) );
  AOI21_X2 U9236 ( .B1(n10274), .B2(n12167), .A(n12254), .ZN(n10355) );
  AND2_X1 U9237 ( .A1(n8536), .A2(n8537), .ZN(n14746) );
  NAND2_X4 U9238 ( .A1(n7624), .A2(n7623), .ZN(n14433) );
  OAI21_X1 U9239 ( .B1(n7515), .B2(n6723), .A(n6722), .ZN(n7510) );
  NAND2_X1 U9240 ( .A1(n7100), .A2(n7101), .ZN(n13931) );
  NAND2_X1 U9241 ( .A1(n14739), .A2(n6913), .ZN(n6911) );
  NOR2_X1 U9242 ( .A1(n13898), .A2(n7104), .ZN(n7103) );
  AOI21_X1 U9243 ( .B1(n6726), .B2(n15287), .A(n6724), .ZN(n12833) );
  XNOR2_X1 U9244 ( .A(n12819), .B(n12824), .ZN(n6726) );
  NAND2_X1 U9245 ( .A1(n12733), .A2(n12734), .ZN(n12736) );
  XNOR2_X1 U9246 ( .A(n6833), .B(n9214), .ZN(n9269) );
  INV_X1 U9247 ( .A(n12802), .ZN(n12804) );
  NAND2_X4 U9248 ( .A1(n10205), .A2(n10206), .ZN(n10941) );
  XNOR2_X2 U9249 ( .A(n9591), .B(n9590), .ZN(n10205) );
  NAND2_X2 U9250 ( .A1(n11407), .A2(n11406), .ZN(n11405) );
  NAND2_X1 U9251 ( .A1(n10233), .A2(n10232), .ZN(n11988) );
  NAND2_X1 U9252 ( .A1(n7399), .A2(n7398), .ZN(n12976) );
  NAND2_X1 U9253 ( .A1(n12875), .A2(n10250), .ZN(n12863) );
  NAND2_X1 U9254 ( .A1(n8742), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6920) );
  INV_X1 U9255 ( .A(n8897), .ZN(n7124) );
  XNOR2_X2 U9256 ( .A(n8817), .B(n8819), .ZN(n13768) );
  NAND2_X1 U9257 ( .A1(n11614), .A2(n8979), .ZN(n7129) );
  NAND2_X1 U9258 ( .A1(n7715), .A2(n7714), .ZN(n7717) );
  XNOR2_X2 U9259 ( .A(n7651), .B(n7650), .ZN(n10890) );
  INV_X1 U9260 ( .A(n7269), .ZN(n7268) );
  OAI211_X1 U9261 ( .C1(n11096), .C2(n6739), .A(n6522), .B(n6736), .ZN(n10972)
         );
  NAND2_X1 U9262 ( .A1(n6750), .A2(n6749), .ZN(n15262) );
  INV_X1 U9263 ( .A(n15260), .ZN(n6750) );
  OAI21_X1 U9264 ( .B1(n15215), .B2(n6754), .A(n6753), .ZN(n10967) );
  INV_X1 U9265 ( .A(n15216), .ZN(n6755) );
  NOR2_X1 U9266 ( .A1(n15215), .A2(n15216), .ZN(n15214) );
  NAND2_X1 U9267 ( .A1(n9942), .A2(n9940), .ZN(n6757) );
  NAND2_X1 U9268 ( .A1(n9925), .A2(n9923), .ZN(n6758) );
  NAND2_X1 U9269 ( .A1(n10057), .A2(n6759), .ZN(n6760) );
  OAI211_X1 U9270 ( .C1(n10057), .C2(n6764), .A(n6761), .B(n6760), .ZN(n13113)
         );
  NAND2_X1 U9271 ( .A1(n9837), .A2(n6772), .ZN(n6771) );
  NAND2_X1 U9272 ( .A1(n6775), .A2(n6777), .ZN(n9553) );
  NAND2_X1 U9273 ( .A1(n9725), .A2(n6779), .ZN(n6775) );
  NAND2_X1 U9274 ( .A1(n9725), .A2(n9724), .ZN(n6784) );
  INV_X1 U9275 ( .A(n6782), .ZN(n6781) );
  NAND2_X1 U9276 ( .A1(n9974), .A2(n6641), .ZN(n6786) );
  NAND3_X1 U9277 ( .A1(n6611), .A2(n6512), .A3(n6476), .ZN(n6790) );
  AND2_X2 U9278 ( .A1(n7090), .A2(n6506), .ZN(n7639) );
  AND2_X1 U9279 ( .A1(n14188), .A2(n6796), .ZN(n14182) );
  NAND2_X1 U9280 ( .A1(n14188), .A2(n6797), .ZN(n14403) );
  NAND3_X1 U9281 ( .A1(n6792), .A2(n6791), .A3(n6793), .ZN(n14402) );
  NAND2_X1 U9282 ( .A1(n14188), .A2(n6590), .ZN(n6791) );
  OR2_X1 U9283 ( .A1(n14188), .A2(n6795), .ZN(n6792) );
  NAND2_X1 U9284 ( .A1(n14188), .A2(n12436), .ZN(n12432) );
  NAND3_X1 U9285 ( .A1(n6800), .A2(n14850), .A3(n11596), .ZN(n11473) );
  NAND3_X1 U9286 ( .A1(n14335), .A2(n6806), .A3(n14389), .ZN(n14331) );
  INV_X1 U9287 ( .A(n6810), .ZN(n14330) );
  NAND2_X1 U9288 ( .A1(n11609), .A2(n6820), .ZN(n6818) );
  INV_X1 U9289 ( .A(n9250), .ZN(n6826) );
  NAND2_X1 U9290 ( .A1(n7235), .A2(n6824), .ZN(n6823) );
  NAND2_X1 U9291 ( .A1(n6826), .A2(n7235), .ZN(n6825) );
  NAND2_X1 U9292 ( .A1(n7237), .A2(n7235), .ZN(n13480) );
  NAND2_X1 U9293 ( .A1(n9250), .A2(n6827), .ZN(n7237) );
  NAND3_X1 U9294 ( .A1(n6835), .A2(n6836), .A3(n6834), .ZN(n11384) );
  NAND2_X1 U9295 ( .A1(n7506), .A2(SI_1_), .ZN(n7509) );
  NAND2_X1 U9296 ( .A1(n10186), .A2(n6846), .ZN(n6847) );
  OAI211_X1 U9297 ( .C1(n10186), .C2(n6848), .A(n6847), .B(n6645), .ZN(
        P3_U3296) );
  NAND2_X1 U9298 ( .A1(n10185), .A2(n10296), .ZN(n6849) );
  NAND2_X1 U9299 ( .A1(n9620), .A2(n6850), .ZN(n9926) );
  INV_X1 U9300 ( .A(n9926), .ZN(n9623) );
  AND2_X1 U9301 ( .A1(n9715), .A2(n10939), .ZN(n6860) );
  OAI21_X1 U9302 ( .B1(n6864), .B2(n6863), .A(n6862), .ZN(n6861) );
  NOR2_X1 U9303 ( .A1(n6867), .A2(n10214), .ZN(n6866) );
  INV_X1 U9304 ( .A(n9710), .ZN(n6867) );
  AOI21_X1 U9305 ( .B1(n9624), .B2(n6875), .A(n6874), .ZN(n6873) );
  NAND2_X1 U9306 ( .A1(n9624), .A2(n6878), .ZN(n9626) );
  NAND2_X1 U9307 ( .A1(n6879), .A2(n6880), .ZN(n9922) );
  NAND2_X1 U9308 ( .A1(n9872), .A2(n6881), .ZN(n6879) );
  AND2_X2 U9309 ( .A1(n6897), .A2(n6599), .ZN(n8508) );
  INV_X1 U9310 ( .A(n6906), .ZN(n14564) );
  XNOR2_X1 U9311 ( .A(n8499), .B(n6907), .ZN(n8502) );
  AOI21_X1 U9312 ( .B1(n8533), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n14742), .ZN(
        n8536) );
  INV_X1 U9313 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6915) );
  NAND2_X2 U9314 ( .A1(n9263), .A2(n9257), .ZN(n8875) );
  NOR2_X2 U9315 ( .A1(n13487), .A2(n13739), .ZN(n13469) );
  NOR2_X2 U9316 ( .A1(n13520), .A2(n13505), .ZN(n13503) );
  NAND2_X1 U9317 ( .A1(n6923), .A2(n6527), .ZN(n13647) );
  NAND2_X1 U9318 ( .A1(n13645), .A2(n6925), .ZN(n6923) );
  NAND2_X1 U9319 ( .A1(n6924), .A2(n6526), .ZN(n13727) );
  NAND2_X1 U9320 ( .A1(n13645), .A2(n6926), .ZN(n6924) );
  NAND2_X1 U9321 ( .A1(n6929), .A2(n6927), .ZN(n11925) );
  INV_X1 U9322 ( .A(n10967), .ZN(n6937) );
  AND3_X2 U9323 ( .A1(n6942), .A2(n6941), .A3(n6940), .ZN(n10961) );
  NAND2_X1 U9324 ( .A1(n14592), .A2(n12792), .ZN(n12793) );
  NAND2_X1 U9325 ( .A1(n14596), .A2(n6950), .ZN(n6949) );
  NAND2_X1 U9326 ( .A1(n12793), .A2(n12794), .ZN(n12816) );
  NAND3_X1 U9327 ( .A1(n6954), .A2(n6951), .A3(n6949), .ZN(n12834) );
  OAI21_X1 U9328 ( .B1(n6957), .B2(n6953), .A(n6952), .ZN(n6951) );
  NOR2_X1 U9329 ( .A1(n12794), .A2(n12825), .ZN(n6953) );
  NAND3_X1 U9330 ( .A1(n6956), .A2(n14592), .A3(n6955), .ZN(n6954) );
  INV_X1 U9331 ( .A(n12825), .ZN(n6955) );
  INV_X1 U9332 ( .A(n6957), .ZN(n6956) );
  NAND2_X1 U9333 ( .A1(n6967), .A2(n12742), .ZN(n12753) );
  AOI21_X1 U9334 ( .B1(n12730), .B2(n6964), .A(n6960), .ZN(n6959) );
  NAND3_X1 U9335 ( .A1(n6963), .A2(n6966), .A3(n6962), .ZN(n12754) );
  NAND4_X1 U9336 ( .A1(n9578), .A2(n9577), .A3(n9838), .A4(n9857), .ZN(n9621)
         );
  NAND2_X1 U9337 ( .A1(n11951), .A2(n6977), .ZN(n6976) );
  NAND2_X1 U9338 ( .A1(n6976), .A2(n6979), .ZN(n12094) );
  NAND2_X1 U9339 ( .A1(n11077), .A2(n6983), .ZN(n6984) );
  NAND2_X1 U9340 ( .A1(n6984), .A2(n6985), .ZN(n10117) );
  NAND2_X1 U9341 ( .A1(n11339), .A2(n10114), .ZN(n11418) );
  NAND2_X1 U9342 ( .A1(n11340), .A2(n11344), .ZN(n11339) );
  NAND2_X1 U9343 ( .A1(n11638), .A2(n6988), .ZN(n6986) );
  NAND2_X1 U9344 ( .A1(n6986), .A2(n6987), .ZN(n11753) );
  NAND2_X1 U9345 ( .A1(n10129), .A2(n6505), .ZN(n6991) );
  NAND2_X1 U9346 ( .A1(n6991), .A2(n6992), .ZN(n12362) );
  NAND2_X1 U9347 ( .A1(n12894), .A2(n7000), .ZN(n6999) );
  NAND2_X1 U9348 ( .A1(n12841), .A2(n10154), .ZN(n10265) );
  NAND2_X1 U9349 ( .A1(n12841), .A2(n6519), .ZN(n7008) );
  OAI21_X1 U9350 ( .B1(n7014), .B2(n10576), .A(n7010), .ZN(n7009) );
  NAND2_X1 U9351 ( .A1(n7014), .A2(n7011), .ZN(n7010) );
  NAND2_X1 U9352 ( .A1(n7039), .A2(n7038), .ZN(n14380) );
  OAI21_X2 U9353 ( .B1(n14291), .B2(n7046), .A(n7044), .ZN(n14258) );
  OAI21_X1 U9354 ( .B1(n7850), .B2(n8202), .A(n8098), .ZN(n11559) );
  NAND2_X1 U9355 ( .A1(n7675), .A2(n14090), .ZN(n7047) );
  NAND2_X1 U9356 ( .A1(n7685), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U9357 ( .A1(n7672), .A2(n7664), .ZN(n7049) );
  NAND2_X1 U9358 ( .A1(n14356), .A2(n6606), .ZN(n14336) );
  INV_X1 U9359 ( .A(n14311), .ZN(n8008) );
  NAND2_X1 U9360 ( .A1(n11471), .A2(n7888), .ZN(n7890) );
  NAND2_X1 U9361 ( .A1(n11456), .A2(n7881), .ZN(n11471) );
  OR2_X1 U9362 ( .A1(n11458), .A2(n11459), .ZN(n11456) );
  OAI22_X1 U9363 ( .A1(n11687), .A2(n7872), .B1(n11591), .B2(n11684), .ZN(
        n11458) );
  NAND2_X1 U9364 ( .A1(n9644), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U9365 ( .A1(n7059), .A2(n7062), .ZN(n9725) );
  AOI21_X1 U9366 ( .B1(n10057), .B2(n10048), .A(n10047), .ZN(n10075) );
  NAND2_X1 U9367 ( .A1(n9910), .A2(n9909), .ZN(n9571) );
  NAND2_X1 U9368 ( .A1(n9888), .A2(n9890), .ZN(n9570) );
  NAND2_X1 U9369 ( .A1(n13960), .A2(n13875), .ZN(n7107) );
  NAND2_X1 U9370 ( .A1(n13960), .A2(n7097), .ZN(n7096) );
  NAND2_X1 U9371 ( .A1(n7107), .A2(n13891), .ZN(n14045) );
  INV_X1 U9372 ( .A(n13898), .ZN(n7106) );
  OAI21_X1 U9373 ( .B1(n13573), .B2(n9106), .A(n7484), .ZN(n13549) );
  NAND2_X1 U9374 ( .A1(n11174), .A2(n6837), .ZN(n8922) );
  NAND2_X1 U9375 ( .A1(n12308), .A2(n6520), .ZN(n12391) );
  INV_X1 U9376 ( .A(n11843), .ZN(n7139) );
  INV_X1 U9377 ( .A(n7144), .ZN(n13476) );
  XNOR2_X2 U9378 ( .A(n7149), .B(n9214), .ZN(n13398) );
  NAND2_X1 U9379 ( .A1(n13415), .A2(n9205), .ZN(n7149) );
  OR2_X1 U9380 ( .A1(n15147), .A2(n7148), .ZN(n7147) );
  NAND2_X1 U9381 ( .A1(n7797), .A2(n7156), .ZN(n7821) );
  NAND2_X1 U9382 ( .A1(n7797), .A2(n7154), .ZN(n7824) );
  OAI21_X1 U9383 ( .B1(n7159), .B2(n7158), .A(n8875), .ZN(n7157) );
  NAND2_X2 U9384 ( .A1(n7157), .A2(n7160), .ZN(n10663) );
  NAND3_X1 U9385 ( .A1(n13774), .A2(n9258), .A3(n14944), .ZN(n7160) );
  NAND2_X2 U9386 ( .A1(n8875), .A2(n9592), .ZN(n9140) );
  INV_X1 U9387 ( .A(n8875), .ZN(n8899) );
  NAND2_X1 U9388 ( .A1(n8854), .A2(n7162), .ZN(n10638) );
  NAND2_X1 U9389 ( .A1(n7163), .A2(n8448), .ZN(P1_U3242) );
  INV_X1 U9390 ( .A(n8438), .ZN(n7164) );
  NAND2_X1 U9391 ( .A1(n7169), .A2(n7570), .ZN(n7622) );
  NAND2_X1 U9392 ( .A1(n7570), .A2(n7571), .ZN(n7620) );
  NAND2_X1 U9393 ( .A1(n7622), .A2(n7571), .ZN(n7616) );
  INV_X1 U9394 ( .A(n7615), .ZN(n7168) );
  NAND2_X1 U9395 ( .A1(n7536), .A2(n7176), .ZN(n7174) );
  OAI211_X1 U9396 ( .C1(n7812), .C2(n7184), .A(n7183), .B(n6630), .ZN(n9129)
         );
  INV_X1 U9397 ( .A(SI_22_), .ZN(n7184) );
  NAND2_X1 U9398 ( .A1(n7777), .A2(n7189), .ZN(n7187) );
  OAI21_X1 U9399 ( .B1(n7544), .B2(n7196), .A(n7195), .ZN(n7644) );
  INV_X1 U9400 ( .A(SI_14_), .ZN(n7197) );
  NAND2_X1 U9401 ( .A1(n7610), .A2(n7609), .ZN(n7612) );
  OAI21_X1 U9402 ( .B1(n7207), .B2(SI_5_), .A(n7518), .ZN(n7705) );
  MUX2_X1 U9403 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n10344), .Z(n7207) );
  NAND2_X1 U9404 ( .A1(n7208), .A2(n10637), .ZN(n9224) );
  XNOR2_X1 U9405 ( .A(n7208), .B(n10639), .ZN(n10640) );
  NAND2_X1 U9406 ( .A1(n13596), .A2(n7211), .ZN(n7209) );
  NAND4_X1 U9407 ( .A1(n8832), .A2(n8831), .A3(n8829), .A4(n8830), .ZN(n9221)
         );
  NAND2_X1 U9408 ( .A1(n7219), .A2(n6832), .ZN(n13410) );
  NAND2_X1 U9409 ( .A1(n13440), .A2(n9505), .ZN(n7223) );
  INV_X1 U9410 ( .A(n9254), .ZN(n7222) );
  AOI21_X1 U9411 ( .B1(n11298), .B2(n7225), .A(n6556), .ZN(n7224) );
  INV_X1 U9412 ( .A(n11298), .ZN(n7226) );
  NAND2_X1 U9413 ( .A1(n11263), .A2(n11262), .ZN(n7227) );
  NAND2_X1 U9414 ( .A1(n11920), .A2(n9233), .ZN(n7229) );
  NAND2_X1 U9415 ( .A1(n7234), .A2(n7233), .ZN(n8818) );
  NAND2_X1 U9416 ( .A1(n7234), .A2(n7231), .ZN(n13763) );
  NAND2_X1 U9417 ( .A1(n9252), .A2(n9153), .ZN(n13478) );
  NAND2_X1 U9418 ( .A1(n7237), .A2(n9251), .ZN(n13477) );
  NAND2_X1 U9419 ( .A1(n13131), .A2(n6607), .ZN(n7243) );
  OAI211_X1 U9420 ( .C1(n13131), .C2(n7245), .A(n7243), .B(n12574), .ZN(
        P2_U3192) );
  OR2_X1 U9421 ( .A1(n13131), .A2(n13132), .ZN(n13133) );
  INV_X1 U9422 ( .A(n11188), .ZN(n7253) );
  NAND2_X1 U9423 ( .A1(n7255), .A2(n7256), .ZN(n7254) );
  OAI21_X1 U9424 ( .B1(n10878), .B2(n7260), .A(n7263), .ZN(n7258) );
  NOR2_X1 U9425 ( .A1(n10878), .A2(n10877), .ZN(n11068) );
  AND2_X1 U9426 ( .A1(n10715), .A2(n11276), .ZN(n11279) );
  NAND2_X2 U9427 ( .A1(n7265), .A2(n7264), .ZN(n11276) );
  NAND2_X1 U9428 ( .A1(n8875), .A2(n13784), .ZN(n7264) );
  NAND2_X1 U9429 ( .A1(n12111), .A2(n7272), .ZN(n7270) );
  NAND3_X1 U9430 ( .A1(n13143), .A2(n7275), .A3(n7274), .ZN(n13194) );
  NAND2_X1 U9431 ( .A1(n12106), .A2(n7276), .ZN(n14923) );
  NAND2_X2 U9432 ( .A1(n11668), .A2(n11667), .ZN(n12106) );
  NAND2_X1 U9434 ( .A1(n13241), .A2(n7277), .ZN(n13180) );
  NAND2_X1 U9435 ( .A1(n13180), .A2(n13182), .ZN(n12513) );
  OAI22_X1 U9436 ( .A1(n9288), .A2(n9289), .B1(n9292), .B2(n7278), .ZN(n9294)
         );
  AOI22_X1 U9437 ( .A1(n9296), .A2(n9297), .B1(n9292), .B2(n7278), .ZN(n9293)
         );
  NAND2_X1 U9438 ( .A1(n9286), .A2(n9287), .ZN(n7278) );
  NAND2_X1 U9439 ( .A1(n11680), .A2(n7282), .ZN(n7280) );
  AOI21_X1 U9440 ( .B1(n7282), .B2(n7284), .A(n6570), .ZN(n7279) );
  NAND2_X1 U9441 ( .A1(n7290), .A2(n7291), .ZN(n9462) );
  NAND2_X1 U9442 ( .A1(n7292), .A2(n9445), .ZN(n9464) );
  INV_X1 U9443 ( .A(n9442), .ZN(n7293) );
  OAI21_X2 U9444 ( .B1(n8125), .B2(n7297), .A(n7294), .ZN(n14329) );
  NAND2_X1 U9445 ( .A1(n8125), .A2(n8124), .ZN(n14372) );
  NOR2_X1 U9446 ( .A1(n7301), .A2(n8398), .ZN(n7300) );
  INV_X1 U9447 ( .A(n8124), .ZN(n7301) );
  OAI21_X1 U9448 ( .B1(n9321), .B2(n7306), .A(n7305), .ZN(n9330) );
  NAND2_X1 U9449 ( .A1(n7304), .A2(n7302), .ZN(n9327) );
  NAND2_X1 U9450 ( .A1(n9321), .A2(n7305), .ZN(n7304) );
  INV_X1 U9451 ( .A(n9320), .ZN(n7307) );
  OAI211_X2 U9452 ( .C1(n14242), .C2(n7311), .A(n7310), .B(n14208), .ZN(n14211) );
  NAND2_X1 U9453 ( .A1(n7313), .A2(n8143), .ZN(n7310) );
  INV_X1 U9454 ( .A(n8143), .ZN(n7311) );
  NAND2_X1 U9455 ( .A1(n14238), .A2(n8143), .ZN(n14209) );
  NAND2_X1 U9456 ( .A1(n7312), .A2(n14242), .ZN(n14238) );
  NAND3_X1 U9459 ( .A1(n7325), .A2(n7324), .A3(n7582), .ZN(n7686) );
  NAND3_X1 U9460 ( .A1(n9431), .A2(n6613), .A3(n7330), .ZN(n7326) );
  INV_X1 U9461 ( .A(n9433), .ZN(n7327) );
  NAND2_X1 U9462 ( .A1(n7330), .A2(n6591), .ZN(n7329) );
  INV_X1 U9463 ( .A(n9430), .ZN(n7332) );
  NAND2_X1 U9464 ( .A1(n7333), .A2(n7335), .ZN(n9402) );
  NAND3_X1 U9465 ( .A1(n9373), .A2(n7337), .A3(n7334), .ZN(n7333) );
  OR2_X1 U9466 ( .A1(n9375), .A2(n9374), .ZN(n7334) );
  NOR2_X1 U9467 ( .A1(n9309), .A2(n9306), .ZN(n7339) );
  AOI21_X1 U9468 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9316) );
  NAND2_X1 U9469 ( .A1(n7341), .A2(n6592), .ZN(n12231) );
  OR2_X2 U9470 ( .A1(n12119), .A2(n8401), .ZN(n7341) );
  NAND3_X1 U9471 ( .A1(n9345), .A2(n9346), .A3(n6612), .ZN(n7342) );
  NAND2_X1 U9472 ( .A1(n7342), .A2(n7343), .ZN(n9355) );
  NAND2_X1 U9473 ( .A1(n11036), .A2(n8202), .ZN(n7345) );
  NAND2_X1 U9474 ( .A1(n8201), .A2(n11036), .ZN(n7346) );
  NAND2_X1 U9475 ( .A1(n11039), .A2(n11036), .ZN(n11035) );
  NAND2_X1 U9476 ( .A1(n7347), .A2(n8098), .ZN(n11039) );
  NAND2_X1 U9477 ( .A1(n7639), .A2(n7348), .ZN(n8157) );
  OAI22_X1 U9478 ( .A1(n9335), .A2(n7351), .B1(n9333), .B2(n9334), .ZN(n9341)
         );
  NAND2_X1 U9479 ( .A1(n9341), .A2(n9340), .ZN(n9344) );
  OAI22_X1 U9480 ( .A1(n9407), .A2(n7352), .B1(n9405), .B2(n9406), .ZN(n9413)
         );
  NAND2_X1 U9481 ( .A1(n9413), .A2(n9414), .ZN(n9412) );
  NAND2_X2 U9482 ( .A1(n7353), .A2(n10578), .ZN(n10585) );
  INV_X2 U9483 ( .A(n10585), .ZN(n11800) );
  NAND2_X1 U9484 ( .A1(n12172), .A2(n7358), .ZN(n7357) );
  NAND2_X1 U9485 ( .A1(n12681), .A2(n7365), .ZN(n7363) );
  NAND2_X1 U9486 ( .A1(n12367), .A2(n7371), .ZN(n7368) );
  INV_X1 U9487 ( .A(n12471), .ZN(n7378) );
  INV_X1 U9488 ( .A(n11162), .ZN(n7391) );
  NOR2_X1 U9489 ( .A1(n15171), .A2(n11162), .ZN(n11163) );
  OAI21_X2 U9490 ( .B1(n6571), .B2(n7395), .A(n7393), .ZN(n12254) );
  NAND3_X1 U9491 ( .A1(n9585), .A2(n7396), .A3(n10188), .ZN(n10192) );
  NAND2_X1 U9492 ( .A1(n9585), .A2(n10188), .ZN(n10198) );
  INV_X1 U9493 ( .A(n10837), .ZN(n15309) );
  NAND2_X1 U9494 ( .A1(n12357), .A2(n7401), .ZN(n7399) );
  NAND2_X1 U9495 ( .A1(n12919), .A2(n7407), .ZN(n7406) );
  OAI21_X1 U9496 ( .B1(n12919), .B2(n7409), .A(n7407), .ZN(n12887) );
  NAND2_X1 U9497 ( .A1(n12877), .A2(n12876), .ZN(n12875) );
  NAND2_X1 U9498 ( .A1(n12877), .A2(n7413), .ZN(n7412) );
  NAND2_X1 U9499 ( .A1(n7420), .A2(n6524), .ZN(n12139) );
  AND2_X2 U9500 ( .A1(n11639), .A2(n10227), .ZN(n11731) );
  NAND2_X1 U9501 ( .A1(n11405), .A2(n6521), .ZN(n11639) );
  NAND2_X1 U9502 ( .A1(n10195), .A2(n7423), .ZN(n9595) );
  NAND2_X1 U9503 ( .A1(n12974), .A2(n7425), .ZN(n12960) );
  XNOR2_X2 U9504 ( .A(n7833), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7841) );
  OAI21_X1 U9505 ( .B1(n8328), .B2(n7430), .A(n7428), .ZN(n8332) );
  NAND2_X1 U9506 ( .A1(n8328), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U9507 ( .A1(n7431), .A2(n7432), .ZN(n8247) );
  NAND3_X1 U9508 ( .A1(n8241), .A2(n6605), .A3(n8240), .ZN(n7431) );
  NAND2_X1 U9509 ( .A1(n7433), .A2(n7434), .ZN(n8257) );
  NAND3_X1 U9510 ( .A1(n8252), .A2(n6604), .A3(n8251), .ZN(n7433) );
  OAI21_X1 U9511 ( .B1(n8233), .B2(n7441), .A(n7439), .ZN(n8237) );
  NAND2_X1 U9512 ( .A1(n7436), .A2(n7437), .ZN(n8236) );
  NAND2_X1 U9513 ( .A1(n8233), .A2(n7439), .ZN(n7436) );
  OAI211_X1 U9514 ( .C1(n7445), .C2(n7448), .A(n7444), .B(n7443), .ZN(n7442)
         );
  NAND2_X1 U9515 ( .A1(n8318), .A2(n8317), .ZN(n7443) );
  NAND2_X1 U9516 ( .A1(n8339), .A2(n7451), .ZN(n7449) );
  NAND2_X1 U9517 ( .A1(n7449), .A2(n7450), .ZN(n8344) );
  NAND2_X1 U9518 ( .A1(n8283), .A2(n8282), .ZN(n7455) );
  NAND2_X1 U9519 ( .A1(n7453), .A2(n7456), .ZN(n8299) );
  NAND3_X1 U9520 ( .A1(n7455), .A2(n7454), .A3(n7458), .ZN(n7453) );
  NAND2_X1 U9521 ( .A1(n8155), .A2(n7461), .ZN(n7834) );
  NAND2_X1 U9522 ( .A1(n8273), .A2(n7467), .ZN(n7464) );
  NAND2_X1 U9523 ( .A1(n7464), .A2(n7465), .ZN(n8284) );
  NAND2_X1 U9524 ( .A1(n13401), .A2(n13749), .ZN(n9274) );
  NAND2_X1 U9525 ( .A1(n13401), .A2(n13688), .ZN(n9272) );
  XNOR2_X1 U9526 ( .A(n11594), .B(n11590), .ZN(n11626) );
  NAND2_X1 U9527 ( .A1(n13913), .A2(n11588), .ZN(n11594) );
  CLKBUF_X1 U9528 ( .A(n11584), .Z(n10901) );
  NAND2_X1 U9529 ( .A1(n8792), .A2(n8793), .ZN(n8790) );
  OAI21_X1 U9530 ( .B1(n7515), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7507), .ZN(
        n7508) );
  NAND2_X1 U9531 ( .A1(n7515), .A2(n9542), .ZN(n7507) );
  NAND2_X1 U9532 ( .A1(n6498), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7502) );
  NAND2_X2 U9533 ( .A1(n7879), .A2(n7478), .ZN(n14083) );
  NOR2_X1 U9534 ( .A1(n9429), .A2(n9428), .ZN(n9431) );
  OAI21_X1 U9535 ( .B1(n10322), .B2(n14377), .A(n10332), .ZN(n10333) );
  INV_X1 U9536 ( .A(n10211), .ZN(n12723) );
  XNOR2_X2 U9537 ( .A(n7825), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U9538 ( .A1(n7851), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U9539 ( .A1(n8208), .A2(n8201), .ZN(n8204) );
  AND2_X2 U9540 ( .A1(n12443), .A2(n7840), .ZN(n7851) );
  NAND2_X1 U9541 ( .A1(n9599), .A2(n9598), .ZN(n13114) );
  INV_X1 U9542 ( .A(n9599), .ZN(n9596) );
  NOR2_X1 U9543 ( .A1(n9502), .A2(n9503), .ZN(n9540) );
  OAI22_X1 U9544 ( .A1(n10698), .A2(n10697), .B1(n10696), .B2(n10695), .ZN(
        n10702) );
  AND2_X1 U9545 ( .A1(n10671), .A2(n10670), .ZN(n10672) );
  NOR2_X1 U9546 ( .A1(n10671), .A2(n10670), .ZN(n10673) );
  XNOR2_X1 U9547 ( .A(n8349), .B(n8348), .ZN(n13766) );
  NAND2_X1 U9548 ( .A1(n11216), .A2(n8834), .ZN(n8854) );
  INV_X1 U9549 ( .A(n8820), .ZN(n12579) );
  INV_X1 U9550 ( .A(n10192), .ZN(n10194) );
  AND2_X1 U9551 ( .A1(n12062), .A2(n12061), .ZN(n7476) );
  NOR2_X1 U9552 ( .A1(n15365), .A2(n10315), .ZN(n7477) );
  NOR2_X1 U9553 ( .A1(n12583), .A2(n13110), .ZN(n10314) );
  AND2_X1 U9554 ( .A1(n15334), .A2(n11076), .ZN(n12999) );
  NOR2_X1 U9555 ( .A1(n12583), .A2(n13062), .ZN(n10301) );
  INV_X1 U9556 ( .A(n8792), .ZN(n8801) );
  INV_X1 U9557 ( .A(n12479), .ZN(n13075) );
  AND3_X1 U9558 ( .A1(n7878), .A2(n7877), .A3(n7876), .ZN(n7478) );
  OR2_X1 U9559 ( .A1(n14504), .A2(n8191), .ZN(n7479) );
  AND2_X1 U9560 ( .A1(n13755), .A2(n13514), .ZN(n7480) );
  AND2_X1 U9561 ( .A1(n12343), .A2(n12174), .ZN(n7481) );
  AND2_X1 U9562 ( .A1(n7489), .A2(n7494), .ZN(n7483) );
  OR2_X1 U9563 ( .A1(n13071), .A2(n10252), .ZN(n7485) );
  AND2_X1 U9564 ( .A1(n11582), .A2(n11581), .ZN(n7486) );
  INV_X1 U9565 ( .A(n14310), .ZN(n8007) );
  INV_X1 U9566 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11257) );
  AND2_X1 U9567 ( .A1(n9473), .A2(n9256), .ZN(n13593) );
  INV_X1 U9568 ( .A(n13593), .ZN(n9268) );
  INV_X1 U9569 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9561) );
  INV_X1 U9570 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12421) );
  INV_X1 U9571 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11259) );
  INV_X1 U9572 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10563) );
  AND2_X1 U9573 ( .A1(n8151), .A2(n10848), .ZN(n7488) );
  INV_X1 U9574 ( .A(n14916), .ZN(n14917) );
  INV_X1 U9575 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7500) );
  NAND2_X1 U9576 ( .A1(n8371), .A2(n8370), .ZN(n7489) );
  INV_X1 U9577 ( .A(n14353), .ZN(n14364) );
  NAND2_X2 U9578 ( .A1(n13419), .A2(n11205), .ZN(n7490) );
  INV_X2 U9579 ( .A(n7490), .ZN(n14668) );
  AND2_X1 U9580 ( .A1(n7916), .A2(n10786), .ZN(n7491) );
  INV_X1 U9581 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11880) );
  INV_X1 U9582 ( .A(n14349), .ZN(n7987) );
  INV_X1 U9583 ( .A(n15284), .ZN(n11544) );
  AND4_X1 U9584 ( .A1(n9530), .A2(n11210), .A3(n9534), .A4(n11879), .ZN(n7493)
         );
  AND2_X1 U9585 ( .A1(n8430), .A2(n8397), .ZN(n7494) );
  AND2_X1 U9586 ( .A1(n8383), .A2(n8380), .ZN(n7495) );
  OR2_X1 U9587 ( .A1(n10321), .A2(n14400), .ZN(n7496) );
  AND4_X1 U9588 ( .A1(n10015), .A2(n10014), .A3(n10013), .A4(n10012), .ZN(
        n12865) );
  NAND2_X1 U9589 ( .A1(n8202), .A2(n8223), .ZN(n8203) );
  OAI22_X1 U9590 ( .A1(n8201), .A2(n8208), .B1(n8223), .B2(n8202), .ZN(n8199)
         );
  NOR2_X1 U9591 ( .A1(n8205), .A2(n11561), .ZN(n8206) );
  MUX2_X1 U9592 ( .A(n8211), .B(n8210), .S(n8209), .Z(n8212) );
  AOI21_X1 U9593 ( .B1(n10668), .B2(n9477), .A(n9285), .ZN(n9292) );
  INV_X1 U9594 ( .A(n9356), .ZN(n9357) );
  INV_X1 U9595 ( .A(n10112), .ZN(n9715) );
  OAI21_X1 U9596 ( .B1(n8307), .B2(n8306), .A(n8305), .ZN(n8309) );
  INV_X1 U9597 ( .A(n9410), .ZN(n9411) );
  NOR2_X1 U9598 ( .A1(n9427), .A2(n9426), .ZN(n9429) );
  NAND2_X1 U9599 ( .A1(n8362), .A2(n8092), .ZN(n8195) );
  OAI21_X1 U9600 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9438) );
  INV_X2 U9601 ( .A(n8208), .ZN(n8223) );
  INV_X1 U9602 ( .A(n12341), .ZN(n12173) );
  INV_X1 U9603 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U9604 ( .A1(n12352), .A2(n12173), .ZN(n12174) );
  NAND2_X1 U9605 ( .A1(n10162), .A2(n14605), .ZN(n10163) );
  INV_X1 U9606 ( .A(n12702), .ZN(n10252) );
  INV_X1 U9607 ( .A(n14640), .ZN(n12509) );
  XNOR2_X1 U9608 ( .A(n14184), .B(n14067), .ZN(n8421) );
  INV_X1 U9609 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7592) );
  AND2_X1 U9610 ( .A1(n9583), .A2(n9796), .ZN(n9584) );
  INV_X1 U9611 ( .A(n13226), .ZN(n12521) );
  NAND2_X1 U9612 ( .A1(n12479), .A2(n12703), .ZN(n10250) );
  INV_X1 U9613 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10093) );
  INV_X1 U9614 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9586) );
  INV_X1 U9615 ( .A(n9101), .ZN(n8812) );
  INV_X1 U9616 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8724) );
  OAI22_X1 U9617 ( .A1(n10896), .A2(n13855), .B1(n11704), .B2(n13838), .ZN(
        n10895) );
  INV_X1 U9618 ( .A(n8001), .ZN(n7999) );
  OR2_X1 U9619 ( .A1(n12280), .A2(n12711), .ZN(n12278) );
  INV_X1 U9620 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9716) );
  INV_X1 U9621 ( .A(n15240), .ZN(n10966) );
  INV_X1 U9622 ( .A(n11514), .ZN(n11513) );
  OR2_X1 U9623 ( .A1(n12791), .A2(n14583), .ZN(n12792) );
  INV_X1 U9624 ( .A(n12822), .ZN(n10576) );
  NAND2_X1 U9625 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n9561), .ZN(n9562) );
  INV_X1 U9626 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9559) );
  INV_X1 U9627 ( .A(n9118), .ZN(n8813) );
  AND2_X1 U9628 ( .A1(n9486), .A2(n9485), .ZN(n9487) );
  OR2_X1 U9629 ( .A1(n9171), .A2(n9170), .ZN(n9196) );
  OR3_X1 U9630 ( .A1(n9132), .A2(n13214), .A3(n13147), .ZN(n9145) );
  OR2_X1 U9631 ( .A1(n8972), .A2(n11438), .ZN(n8987) );
  INV_X1 U9632 ( .A(n8803), .ZN(n9512) );
  NAND2_X1 U9633 ( .A1(n13436), .A2(n9191), .ZN(n13416) );
  OR2_X1 U9634 ( .A1(n8959), .A2(n11379), .ZN(n8972) );
  AND3_X1 U9635 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8915) );
  INV_X1 U9636 ( .A(n10663), .ZN(n8834) );
  INV_X1 U9637 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8798) );
  INV_X1 U9638 ( .A(n12312), .ZN(n12309) );
  INV_X1 U9639 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7873) );
  OR2_X1 U9640 ( .A1(n11587), .A2(n11586), .ZN(n11588) );
  INV_X1 U9641 ( .A(n13789), .ZN(n13790) );
  OR2_X1 U9642 ( .A1(n8073), .A2(n13940), .ZN(n10327) );
  INV_X1 U9643 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10786) );
  INV_X1 U9644 ( .A(n14245), .ZN(n8137) );
  NAND2_X1 U9645 ( .A1(n7999), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U9646 ( .A1(n14883), .A2(n11874), .ZN(n10869) );
  NAND2_X1 U9647 ( .A1(n7545), .A2(n10522), .ZN(n7631) );
  NAND2_X1 U9648 ( .A1(n7533), .A2(SI_10_), .ZN(n7535) );
  AND2_X1 U9649 ( .A1(n7518), .A2(n7705), .ZN(n7519) );
  NAND2_X1 U9650 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  OR2_X1 U9651 ( .A1(n9816), .A2(n9603), .ZN(n9843) );
  NOR2_X1 U9652 ( .A1(n9843), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9865) );
  OR2_X1 U9653 ( .A1(n9788), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9816) );
  OR2_X1 U9654 ( .A1(n10023), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10037) );
  OR2_X1 U9655 ( .A1(n10598), .A2(n10597), .ZN(n15189) );
  OR2_X1 U9656 ( .A1(n14604), .A2(n10062), .ZN(n12844) );
  INV_X1 U9657 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n11008) );
  INV_X1 U9658 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10985) );
  INV_X1 U9659 ( .A(n11520), .ZN(n11534) );
  INV_X1 U9660 ( .A(n12732), .ZN(n12257) );
  OR2_X1 U9661 ( .A1(n6501), .A2(n12823), .ZN(n10973) );
  INV_X1 U9662 ( .A(n10266), .ZN(n10256) );
  INV_X1 U9663 ( .A(n10243), .ZN(n12980) );
  INV_X1 U9664 ( .A(n12708), .ZN(n12990) );
  AND2_X1 U9665 ( .A1(n9903), .A2(n10132), .ZN(n12296) );
  AND2_X1 U9666 ( .A1(n10124), .A2(n9833), .ZN(n10172) );
  INV_X1 U9667 ( .A(n15311), .ZN(n15327) );
  OR2_X1 U9668 ( .A1(n10801), .A2(n10574), .ZN(n10306) );
  INV_X1 U9669 ( .A(n10095), .ZN(n10096) );
  OR2_X1 U9670 ( .A1(n9891), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U9671 ( .A1(n9553), .A2(n9552), .ZN(n9765) );
  NAND2_X1 U9672 ( .A1(n11431), .A2(n11430), .ZN(n11432) );
  NAND2_X1 U9673 ( .A1(n13268), .A2(n6478), .ZN(n10695) );
  INV_X1 U9674 ( .A(n13512), .ZN(n13483) );
  INV_X1 U9675 ( .A(n9498), .ZN(n9499) );
  INV_X1 U9676 ( .A(n9453), .ZN(n9207) );
  OR2_X1 U9677 ( .A1(n14983), .A2(n14982), .ZN(n14985) );
  AND2_X1 U9678 ( .A1(n15001), .A2(n15000), .ZN(n15002) );
  AND2_X1 U9679 ( .A1(n15023), .A2(n15022), .ZN(n15029) );
  AND2_X1 U9680 ( .A1(n9138), .A2(n9137), .ZN(n13536) );
  INV_X1 U9681 ( .A(n13259), .ZN(n11787) );
  OR2_X1 U9682 ( .A1(n10677), .A2(n9258), .ZN(n13539) );
  NOR2_X1 U9683 ( .A1(n10663), .A2(n11276), .ZN(n11275) );
  OR2_X1 U9684 ( .A1(n11208), .A2(n10679), .ZN(n15140) );
  NAND2_X1 U9685 ( .A1(n6483), .A2(n11210), .ZN(n10687) );
  NOR2_X1 U9686 ( .A1(n7916), .A2(n10786), .ZN(n7932) );
  OR2_X1 U9687 ( .A1(n7892), .A2(n7891), .ZN(n7908) );
  AND2_X1 U9688 ( .A1(n12392), .A2(n12389), .ZN(n12390) );
  OR2_X1 U9689 ( .A1(n7965), .A2(n7964), .ZN(n7974) );
  OR2_X1 U9690 ( .A1(n13865), .A2(n13907), .ZN(n13998) );
  INV_X1 U9691 ( .A(n11593), .ZN(n11590) );
  NAND2_X1 U9692 ( .A1(n7940), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U9693 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  NAND2_X1 U9694 ( .A1(n12306), .A2(n12305), .ZN(n12307) );
  NAND2_X1 U9695 ( .A1(n7955), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7965) );
  AND2_X1 U9696 ( .A1(n8066), .A2(n8056), .ZN(n14220) );
  NAND2_X1 U9697 ( .A1(n14069), .A2(n14364), .ZN(n12428) );
  INV_X1 U9698 ( .A(n8409), .ZN(n12036) );
  INV_X1 U9699 ( .A(n10869), .ZN(n10320) );
  INV_X1 U9700 ( .A(n10407), .ZN(n8190) );
  OAI21_X1 U9701 ( .B1(n7533), .B2(SI_10_), .A(n7535), .ZN(n7750) );
  INV_X1 U9702 ( .A(n7691), .ZN(n7693) );
  OAI21_X1 U9703 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n8481), .A(n8480), .ZN(
        n8535) );
  NOR2_X1 U9704 ( .A1(n9741), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9757) );
  OR2_X1 U9705 ( .A1(n9719), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9741) );
  AND2_X1 U9706 ( .A1(n10592), .A2(n10937), .ZN(n15180) );
  AND4_X1 U9707 ( .A1(n10103), .A2(n10053), .A3(n10052), .A4(n10051), .ZN(
        n12837) );
  AND4_X1 U9708 ( .A1(n9954), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(n12979)
         );
  INV_X1 U9709 ( .A(n15241), .ZN(n15280) );
  INV_X1 U9710 ( .A(n14592), .ZN(n14596) );
  AND2_X1 U9711 ( .A1(n12954), .A2(n12953), .ZN(n13037) );
  INV_X1 U9712 ( .A(n15302), .ZN(n12963) );
  AND2_X1 U9713 ( .A1(n14603), .A2(n14602), .ZN(n14614) );
  INV_X1 U9714 ( .A(n14623), .ZN(n15339) );
  AND2_X1 U9715 ( .A1(n10938), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10573) );
  INV_X1 U9716 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9838) );
  AND2_X1 U9717 ( .A1(n9152), .A2(n9151), .ZN(n13460) );
  OR2_X1 U9718 ( .A1(n10475), .A2(n10474), .ZN(n15042) );
  INV_X1 U9719 ( .A(n15042), .ZN(n15021) );
  AND2_X1 U9720 ( .A1(n10455), .A2(n10454), .ZN(n15027) );
  INV_X1 U9721 ( .A(n15039), .ZN(n15051) );
  INV_X1 U9722 ( .A(n13731), .ZN(n13396) );
  INV_X1 U9723 ( .A(n9266), .ZN(n9267) );
  INV_X1 U9724 ( .A(n13525), .ZN(n14664) );
  AND2_X1 U9725 ( .A1(n15156), .A2(n15100), .ZN(n13688) );
  AND2_X1 U9726 ( .A1(n9219), .A2(n15123), .ZN(n13724) );
  INV_X1 U9727 ( .A(n13724), .ZN(n15137) );
  AND3_X1 U9728 ( .A1(n15091), .A2(n8804), .A3(n10687), .ZN(n9273) );
  AND2_X1 U9729 ( .A1(n8769), .A2(n8765), .ZN(n15055) );
  AND2_X1 U9730 ( .A1(n8767), .A2(n8766), .ZN(n11202) );
  OR2_X1 U9731 ( .A1(n8748), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8762) );
  NOR2_X1 U9732 ( .A1(n8999), .A2(n9028), .ZN(n14994) );
  OR2_X1 U9733 ( .A1(n7949), .A2(n7948), .ZN(n7957) );
  INV_X1 U9734 ( .A(n14875), .ZN(n14882) );
  INV_X1 U9735 ( .A(n14065), .ZN(n14689) );
  INV_X1 U9736 ( .A(n14696), .ZN(n14063) );
  OR2_X1 U9737 ( .A1(n14203), .A2(n7963), .ZN(n8072) );
  AND4_X1 U9738 ( .A1(n7998), .A2(n7997), .A3(n7996), .A4(n7995), .ZN(n14352)
         );
  INV_X1 U9739 ( .A(n14775), .ZN(n14804) );
  OR2_X1 U9740 ( .A1(n14760), .A2(n14749), .ZN(n14168) );
  INV_X1 U9741 ( .A(n8415), .ZN(n14283) );
  NAND2_X1 U9742 ( .A1(n10320), .A2(n10406), .ZN(n14386) );
  NAND2_X1 U9743 ( .A1(n10325), .A2(n14386), .ZN(n14393) );
  INV_X1 U9744 ( .A(n10859), .ZN(n10865) );
  AND2_X1 U9745 ( .A1(n14860), .A2(n8153), .ZN(n14888) );
  INV_X1 U9746 ( .A(n14860), .ZN(n14879) );
  AOI21_X1 U9747 ( .B1(n8190), .B2(n8189), .A(n10408), .ZN(n10859) );
  INV_X1 U9748 ( .A(n10860), .ZN(n10406) );
  INV_X1 U9749 ( .A(n10335), .ZN(n10413) );
  XNOR2_X1 U9750 ( .A(n7656), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14151) );
  AND2_X1 U9751 ( .A1(n10955), .A2(n10954), .ZN(n15245) );
  AND2_X1 U9752 ( .A1(n11155), .A2(n11741), .ZN(n15193) );
  AND4_X1 U9753 ( .A1(n10103), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n11285) );
  OR2_X1 U9754 ( .A1(n10565), .A2(n10354), .ZN(n12720) );
  INV_X1 U9755 ( .A(n15245), .ZN(n15296) );
  INV_X1 U9756 ( .A(n14593), .ZN(n15291) );
  AND2_X1 U9757 ( .A1(n12966), .A2(n12965), .ZN(n13042) );
  AND2_X1 U9758 ( .A1(n12142), .A2(n12285), .ZN(n12324) );
  NOR2_X1 U9759 ( .A1(n10301), .A2(n10303), .ZN(n10304) );
  NAND2_X1 U9760 ( .A1(n15374), .A2(n15325), .ZN(n13062) );
  INV_X1 U9761 ( .A(n15374), .ZN(n15371) );
  INV_X1 U9762 ( .A(n11947), .ZN(n11936) );
  INV_X1 U9763 ( .A(n15365), .ZN(n15363) );
  INV_X1 U9764 ( .A(SI_17_), .ZN(n10797) );
  INV_X1 U9765 ( .A(SI_11_), .ZN(n10378) );
  NAND2_X1 U9766 ( .A1(n10712), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14934) );
  OR2_X1 U9767 ( .A1(n10686), .A2(n10678), .ZN(n14926) );
  OR2_X1 U9768 ( .A1(n9094), .A2(n9093), .ZN(n13564) );
  INV_X1 U9769 ( .A(n15027), .ZN(n15048) );
  INV_X1 U9770 ( .A(n15033), .ZN(n15053) );
  OR2_X1 U9771 ( .A1(n10455), .A2(P2_U3088), .ZN(n15039) );
  OR2_X1 U9772 ( .A1(n14668), .A2(n11227), .ZN(n13641) );
  INV_X1 U9773 ( .A(n15156), .ZN(n15154) );
  AND2_X2 U9774 ( .A1(n9273), .A2(n10675), .ZN(n15156) );
  INV_X1 U9775 ( .A(n13749), .ZN(n13754) );
  INV_X1 U9776 ( .A(n15147), .ZN(n15145) );
  INV_X1 U9777 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12138) );
  INV_X1 U9778 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11200) );
  INV_X1 U9779 ( .A(n14465), .ZN(n14335) );
  NAND2_X1 U9780 ( .A1(n10863), .A2(n10862), .ZN(n14065) );
  NAND2_X1 U9781 ( .A1(n8080), .A2(n8079), .ZN(n14193) );
  INV_X1 U9782 ( .A(n13833), .ZN(n14363) );
  OR2_X1 U9783 ( .A1(n10604), .A2(n10603), .ZN(n14760) );
  OR2_X1 U9784 ( .A1(n14760), .A2(n14101), .ZN(n14775) );
  INV_X1 U9785 ( .A(n14771), .ZN(n14807) );
  AND2_X1 U9786 ( .A1(n12227), .A2(n12226), .ZN(n14702) );
  NAND2_X1 U9787 ( .A1(n14393), .A2(n14879), .ZN(n14400) );
  NAND2_X1 U9788 ( .A1(n14393), .A2(n10324), .ZN(n14394) );
  AND2_X1 U9789 ( .A1(n14702), .A2(n14701), .ZN(n14722) );
  OR2_X1 U9790 ( .A1(n8720), .A2(n10859), .ZN(n14905) );
  INV_X1 U9791 ( .A(n7840), .ZN(n14513) );
  INV_X1 U9792 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10795) );
  INV_X1 U9793 ( .A(n12720), .ZN(P3_U3897) );
  NAND2_X1 U9794 ( .A1(n7496), .A2(n10334), .ZN(P1_U3356) );
  NAND2_X1 U9795 ( .A1(n8723), .A2(n8722), .ZN(P1_U3557) );
  NAND2_X1 U9796 ( .A1(n8192), .A2(n7479), .ZN(P1_U3525) );
  XNOR2_X1 U9797 ( .A(n7487), .B(n8719), .ZN(SUB_1596_U4) );
  INV_X2 U9798 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13383) );
  INV_X2 U9799 ( .A(P1_RD_REG_SCAN_IN), .ZN(n14536) );
  NAND3_X1 U9800 ( .A1(n14177), .A2(n13383), .A3(n14536), .ZN(n7498) );
  INV_X2 U9801 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7499) );
  NAND3_X1 U9802 ( .A1(n7499), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7501) );
  INV_X1 U9803 ( .A(n7506), .ZN(n7505) );
  INV_X1 U9804 ( .A(SI_1_), .ZN(n7504) );
  INV_X1 U9805 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9672) );
  INV_X1 U9806 ( .A(SI_0_), .ZN(n10394) );
  INV_X1 U9807 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10350) );
  MUX2_X1 U9808 ( .A(n10350), .B(n9546), .S(n6498), .Z(n7668) );
  INV_X1 U9809 ( .A(SI_2_), .ZN(n10389) );
  NOR2_X1 U9810 ( .A1(n7668), .A2(n10389), .ZN(n7513) );
  NAND2_X1 U9811 ( .A1(n7510), .A2(SI_3_), .ZN(n7514) );
  OAI21_X1 U9812 ( .B1(n7510), .B2(SI_3_), .A(n7514), .ZN(n7679) );
  NOR2_X1 U9813 ( .A1(n6484), .A2(SI_2_), .ZN(n7511) );
  OAI21_X1 U9814 ( .B1(n7516), .B2(SI_4_), .A(n7703), .ZN(n7692) );
  INV_X1 U9815 ( .A(n7692), .ZN(n7517) );
  AND2_X1 U9816 ( .A1(n7703), .A2(n7518), .ZN(n7520) );
  MUX2_X1 U9817 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9592), .Z(n7521) );
  NAND2_X1 U9818 ( .A1(n7521), .A2(SI_6_), .ZN(n7523) );
  OAI21_X1 U9819 ( .B1(SI_6_), .B2(n7521), .A(n7523), .ZN(n7522) );
  INV_X1 U9820 ( .A(n7522), .ZN(n7714) );
  NAND2_X1 U9821 ( .A1(n7717), .A2(n7523), .ZN(n7724) );
  MUX2_X1 U9822 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9592), .Z(n7524) );
  NAND2_X1 U9823 ( .A1(n7524), .A2(SI_7_), .ZN(n7526) );
  OAI21_X1 U9824 ( .B1(n7524), .B2(SI_7_), .A(n7526), .ZN(n7525) );
  INV_X1 U9825 ( .A(n7525), .ZN(n7723) );
  NAND2_X1 U9826 ( .A1(n7724), .A2(n7723), .ZN(n7726) );
  MUX2_X1 U9827 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9592), .Z(n7527) );
  NAND2_X1 U9828 ( .A1(n7527), .A2(SI_8_), .ZN(n7529) );
  OAI21_X1 U9829 ( .B1(SI_8_), .B2(n7527), .A(n7529), .ZN(n7528) );
  INV_X1 U9830 ( .A(n7528), .ZN(n7731) );
  NAND2_X1 U9831 ( .A1(n7732), .A2(n7731), .ZN(n7734) );
  NAND2_X1 U9832 ( .A1(n7734), .A2(n7529), .ZN(n7741) );
  MUX2_X1 U9833 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9592), .Z(n7530) );
  NAND2_X1 U9834 ( .A1(n7530), .A2(SI_9_), .ZN(n7532) );
  OAI21_X1 U9835 ( .B1(SI_9_), .B2(n7530), .A(n7532), .ZN(n7531) );
  INV_X1 U9836 ( .A(n7531), .ZN(n7740) );
  NAND2_X1 U9837 ( .A1(n7741), .A2(n7740), .ZN(n7743) );
  MUX2_X1 U9838 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9592), .Z(n7533) );
  INV_X1 U9839 ( .A(n7750), .ZN(n7534) );
  MUX2_X1 U9840 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9592), .Z(n7537) );
  INV_X1 U9841 ( .A(n7537), .ZN(n7538) );
  NAND2_X1 U9842 ( .A1(n7538), .A2(n10378), .ZN(n7539) );
  MUX2_X1 U9843 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n9592), .Z(n7540) );
  INV_X1 U9844 ( .A(n7540), .ZN(n7541) );
  MUX2_X1 U9845 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9592), .Z(n7769) );
  NOR2_X1 U9846 ( .A1(n7769), .A2(SI_13_), .ZN(n7543) );
  NAND2_X1 U9847 ( .A1(n7769), .A2(SI_13_), .ZN(n7542) );
  MUX2_X1 U9848 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9592), .Z(n7650) );
  MUX2_X1 U9849 ( .A(n9568), .B(n11200), .S(n9592), .Z(n7545) );
  INV_X1 U9850 ( .A(n7545), .ZN(n7546) );
  NAND2_X1 U9851 ( .A1(n7546), .A2(SI_15_), .ZN(n7547) );
  MUX2_X1 U9852 ( .A(n11259), .B(n11257), .S(n9592), .Z(n7548) );
  NAND2_X1 U9853 ( .A1(n7548), .A2(n10546), .ZN(n7634) );
  INV_X1 U9854 ( .A(n7548), .ZN(n7549) );
  MUX2_X1 U9855 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n9592), .Z(n7775) );
  INV_X1 U9856 ( .A(n7775), .ZN(n7552) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9592), .Z(n7782) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9592), .Z(n7794) );
  AOI22_X1 U9859 ( .A1(SI_18_), .A2(n7782), .B1(n7794), .B2(SI_19_), .ZN(n7553) );
  OAI21_X1 U9860 ( .B1(n7782), .B2(SI_18_), .A(SI_19_), .ZN(n7556) );
  INV_X1 U9861 ( .A(n7794), .ZN(n7555) );
  NOR2_X1 U9862 ( .A1(SI_18_), .A2(SI_19_), .ZN(n7554) );
  INV_X1 U9863 ( .A(n7782), .ZN(n7784) );
  AOI22_X1 U9864 ( .A1(n7556), .A2(n7555), .B1(n7554), .B2(n7784), .ZN(n7557)
         );
  NAND2_X1 U9865 ( .A1(n7558), .A2(n11336), .ZN(n7559) );
  INV_X1 U9866 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11744) );
  MUX2_X1 U9867 ( .A(n11744), .B(n11748), .S(n9592), .Z(n7803) );
  MUX2_X1 U9868 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9592), .Z(n7562) );
  NAND2_X1 U9869 ( .A1(n7562), .A2(SI_21_), .ZN(n7564) );
  OAI21_X1 U9870 ( .B1(SI_21_), .B2(n7562), .A(n7564), .ZN(n7563) );
  INV_X1 U9871 ( .A(n7563), .ZN(n7809) );
  INV_X1 U9872 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7565) );
  MUX2_X1 U9873 ( .A(n7565), .B(n12138), .S(n9592), .Z(n9126) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9592), .Z(n7626) );
  INV_X1 U9875 ( .A(SI_24_), .ZN(n7569) );
  NAND2_X1 U9876 ( .A1(n6715), .A2(n7569), .ZN(n7570) );
  INV_X1 U9877 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12380) );
  INV_X1 U9878 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12377) );
  MUX2_X1 U9879 ( .A(n12380), .B(n12377), .S(n9592), .Z(n7619) );
  MUX2_X1 U9880 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9592), .Z(n7572) );
  XNOR2_X1 U9881 ( .A(n7572), .B(SI_25_), .ZN(n7615) );
  INV_X1 U9882 ( .A(n7572), .ZN(n7573) );
  INV_X1 U9883 ( .A(SI_25_), .ZN(n12169) );
  INV_X1 U9884 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13777) );
  MUX2_X1 U9885 ( .A(n14519), .B(n13777), .S(n9592), .Z(n7816) );
  INV_X1 U9886 ( .A(n7816), .ZN(n7574) );
  NOR2_X1 U9887 ( .A1(n7574), .A2(SI_26_), .ZN(n7575) );
  INV_X1 U9888 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14518) );
  INV_X1 U9889 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13775) );
  MUX2_X1 U9890 ( .A(n14518), .B(n13775), .S(n9592), .Z(n7576) );
  XNOR2_X1 U9891 ( .A(n7576), .B(SI_27_), .ZN(n7609) );
  INV_X1 U9892 ( .A(n7576), .ZN(n7577) );
  NAND2_X1 U9893 ( .A1(n7577), .A2(SI_27_), .ZN(n7578) );
  MUX2_X1 U9894 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9592), .Z(n7579) );
  XNOR2_X1 U9895 ( .A(n7579), .B(SI_28_), .ZN(n7605) );
  INV_X1 U9896 ( .A(n7579), .ZN(n7580) );
  INV_X1 U9897 ( .A(SI_28_), .ZN(n13128) );
  NAND2_X1 U9898 ( .A1(n7580), .A2(n13128), .ZN(n7581) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9592), .Z(n8350) );
  INV_X1 U9900 ( .A(SI_29_), .ZN(n13124) );
  XNOR2_X1 U9901 ( .A(n8350), .B(n13124), .ZN(n8348) );
  INV_X1 U9902 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7587) );
  INV_X1 U9903 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7586) );
  NOR2_X1 U9904 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7589) );
  NOR2_X1 U9905 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n7588) );
  NOR2_X1 U9906 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7594) );
  NAND4_X1 U9907 ( .A1(n7594), .A2(n7593), .A3(n7798), .A4(n7592), .ZN(n8163)
         );
  NAND3_X1 U9908 ( .A1(n7638), .A2(n8168), .A3(n7595), .ZN(n7596) );
  NAND2_X1 U9909 ( .A1(n8157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U9910 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7600), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n7602) );
  NAND2_X2 U9911 ( .A1(n7602), .A2(n6790), .ZN(n14516) );
  NAND2_X2 U9912 ( .A1(n7828), .A2(n14516), .ZN(n10512) );
  NAND2_X1 U9913 ( .A1(n13766), .A2(n8390), .ZN(n7604) );
  BUF_X4 U9914 ( .A(n7685), .Z(n8391) );
  NAND2_X1 U9915 ( .A1(n8391), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9916 ( .A1(n12425), .A2(n8390), .ZN(n7608) );
  NAND2_X1 U9917 ( .A1(n8391), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7607) );
  NAND2_X2 U9918 ( .A1(n7608), .A2(n7607), .ZN(n14409) );
  INV_X1 U9919 ( .A(n14409), .ZN(n12436) );
  NAND2_X1 U9920 ( .A1(n13773), .A2(n8390), .ZN(n7614) );
  NAND2_X1 U9921 ( .A1(n8391), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7613) );
  XNOR2_X1 U9922 ( .A(n7616), .B(n7615), .ZN(n13779) );
  NAND2_X1 U9923 ( .A1(n13779), .A2(n8390), .ZN(n7618) );
  NAND2_X1 U9924 ( .A1(n8391), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7617) );
  NAND2_X2 U9925 ( .A1(n7618), .A2(n7617), .ZN(n14427) );
  INV_X1 U9926 ( .A(n14427), .ZN(n14235) );
  NAND2_X1 U9927 ( .A1(n7620), .A2(n7619), .ZN(n7621) );
  OR2_X2 U9928 ( .A1(n12381), .A2(n7813), .ZN(n7624) );
  NAND2_X1 U9929 ( .A1(n8391), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7623) );
  XNOR2_X1 U9930 ( .A(n7626), .B(SI_23_), .ZN(n7627) );
  XNOR2_X1 U9931 ( .A(n7625), .B(n7627), .ZN(n12192) );
  NAND2_X1 U9932 ( .A1(n12192), .A2(n8390), .ZN(n7629) );
  NAND2_X1 U9933 ( .A1(n8391), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7628) );
  INV_X1 U9934 ( .A(n14438), .ZN(n14266) );
  OR2_X1 U9935 ( .A1(n9127), .A2(n9592), .ZN(n7630) );
  NAND2_X1 U9936 ( .A1(n7632), .A2(n7631), .ZN(n7636) );
  AND2_X1 U9937 ( .A1(n7634), .A2(n7633), .ZN(n7635) );
  NAND2_X1 U9938 ( .A1(n11256), .A2(n8390), .ZN(n7642) );
  INV_X1 U9939 ( .A(n7639), .ZN(n7646) );
  NAND2_X1 U9940 ( .A1(n7646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7637) );
  MUX2_X1 U9941 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7637), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n7640) );
  NAND2_X1 U9942 ( .A1(n7640), .A2(n7787), .ZN(n11772) );
  INV_X1 U9943 ( .A(n11772), .ZN(n11965) );
  AOI22_X1 U9944 ( .A1(n8391), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6504), .B2(
        n11965), .ZN(n7641) );
  INV_X1 U9945 ( .A(n14480), .ZN(n14395) );
  XNOR2_X1 U9946 ( .A(n7644), .B(n7643), .ZN(n11172) );
  NAND2_X1 U9947 ( .A1(n11172), .A2(n8390), .ZN(n7649) );
  NAND2_X1 U9948 ( .A1(n6621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7645) );
  MUX2_X1 U9949 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7645), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n7647) );
  AOI22_X1 U9950 ( .A1(n8391), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6503), .B2(
        n14803), .ZN(n7648) );
  NAND2_X1 U9951 ( .A1(n10890), .A2(n8390), .ZN(n7658) );
  NOR2_X1 U9952 ( .A1(n7696), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U9953 ( .A1(n7718), .A2(n7653), .ZN(n7727) );
  INV_X1 U9954 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U9955 ( .A1(n7752), .A2(n7654), .ZN(n7759) );
  OAI21_X1 U9956 ( .B1(n7765), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U9957 ( .A1(n7772), .A2(n7585), .ZN(n7655) );
  NAND2_X1 U9958 ( .A1(n7655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7656) );
  AOI22_X1 U9959 ( .A1(n14151), .A2(n6504), .B1(n8391), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7657) );
  NAND2_X2 U9960 ( .A1(n7658), .A2(n7657), .ZN(n14688) );
  INV_X1 U9961 ( .A(n7659), .ZN(n7660) );
  NAND2_X1 U9962 ( .A1(n7661), .A2(n7660), .ZN(n7662) );
  NAND2_X1 U9963 ( .A1(n7663), .A2(n7662), .ZN(n12424) );
  INV_X1 U9964 ( .A(n12424), .ZN(n7664) );
  NAND2_X1 U9965 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7665) );
  INV_X1 U9966 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14752) );
  NOR2_X1 U9967 ( .A1(n9592), .A2(n10394), .ZN(n7666) );
  XNOR2_X1 U9968 ( .A(n7666), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14529) );
  MUX2_X1 U9969 ( .A(n14752), .B(n14529), .S(n10512), .Z(n11860) );
  NAND2_X1 U9970 ( .A1(n7667), .A2(SI_2_), .ZN(n7680) );
  OAI21_X1 U9971 ( .B1(n7667), .B2(SI_2_), .A(n7680), .ZN(n7669) );
  NAND2_X1 U9972 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  NAND2_X1 U9973 ( .A1(n7682), .A2(n7670), .ZN(n10349) );
  INV_X1 U9974 ( .A(n10349), .ZN(n7671) );
  NAND2_X1 U9975 ( .A1(n7672), .A2(n7671), .ZN(n7678) );
  NAND2_X1 U9976 ( .A1(n7685), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U9977 ( .A1(n7673), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7674) );
  XNOR2_X1 U9978 ( .A(n7674), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U9979 ( .A1(n6503), .A2(n14113), .ZN(n7676) );
  AND3_X2 U9980 ( .A1(n7678), .A2(n7677), .A3(n7676), .ZN(n14845) );
  AND2_X1 U9981 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  NAND2_X1 U9982 ( .A1(n7682), .A2(n7681), .ZN(n7684) );
  NAND2_X1 U9983 ( .A1(n7683), .A2(n7684), .ZN(n10341) );
  NAND2_X1 U9984 ( .A1(n7685), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U9985 ( .A1(n7686), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7687) );
  MUX2_X1 U9986 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7687), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n7688) );
  AND2_X1 U9987 ( .A1(n7688), .A2(n7696), .ZN(n14120) );
  NAND2_X1 U9988 ( .A1(n6504), .A2(n14120), .ZN(n7689) );
  NAND2_X1 U9989 ( .A1(n7693), .A2(n7692), .ZN(n7694) );
  NAND2_X1 U9990 ( .A1(n7694), .A2(n7704), .ZN(n10351) );
  INV_X1 U9991 ( .A(n10351), .ZN(n7695) );
  NAND2_X1 U9992 ( .A1(n7695), .A2(n8390), .ZN(n7702) );
  NAND2_X1 U9993 ( .A1(n7696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7697) );
  MUX2_X1 U9994 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7697), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7699) );
  INV_X1 U9995 ( .A(n7698), .ZN(n7710) );
  NAND2_X1 U9996 ( .A1(n7699), .A2(n7710), .ZN(n14774) );
  INV_X1 U9997 ( .A(n14774), .ZN(n10628) );
  NAND2_X1 U9998 ( .A1(n6503), .A2(n10628), .ZN(n7701) );
  NAND2_X1 U9999 ( .A1(n8391), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U10000 ( .A1(n7704), .A2(n7703), .ZN(n7707) );
  INV_X1 U10001 ( .A(n7705), .ZN(n7706) );
  NAND2_X1 U10002 ( .A1(n7707), .A2(n7706), .ZN(n7709) );
  OR2_X1 U10003 ( .A1(n7707), .A2(n7706), .ZN(n7708) );
  NAND2_X1 U10004 ( .A1(n10367), .A2(n8390), .ZN(n7713) );
  NAND2_X1 U10005 ( .A1(n7710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7711) );
  XNOR2_X1 U10006 ( .A(n7711), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U10007 ( .A1(n8391), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6503), .B2(
        n10629), .ZN(n7712) );
  OR2_X1 U10008 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  NAND2_X1 U10009 ( .A1(n7717), .A2(n7716), .ZN(n10382) );
  OR2_X1 U10010 ( .A1(n10382), .A2(n7813), .ZN(n7722) );
  INV_X1 U10011 ( .A(n7718), .ZN(n7719) );
  NAND2_X1 U10012 ( .A1(n7719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7720) );
  XNOR2_X1 U10013 ( .A(n7720), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U10014 ( .A1(n8391), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6504), .B2(
        n10650), .ZN(n7721) );
  NAND2_X1 U10015 ( .A1(n7722), .A2(n7721), .ZN(n14864) );
  OR2_X1 U10016 ( .A1(n11473), .A2(n14864), .ZN(n11503) );
  OR2_X1 U10017 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  NAND2_X1 U10018 ( .A1(n7726), .A2(n7725), .ZN(n10404) );
  OR2_X1 U10019 ( .A1(n10404), .A2(n7813), .ZN(n7730) );
  NAND2_X1 U10020 ( .A1(n7727), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7728) );
  XNOR2_X1 U10021 ( .A(n7728), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U10022 ( .A1(n8391), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6503), .B2(
        n10652), .ZN(n7729) );
  NAND2_X1 U10023 ( .A1(n7730), .A2(n7729), .ZN(n12089) );
  OR2_X1 U10024 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U10025 ( .A1(n7734), .A2(n7733), .ZN(n10416) );
  OR2_X1 U10026 ( .A1(n10416), .A2(n7813), .ZN(n7739) );
  NAND2_X1 U10027 ( .A1(n7735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7736) );
  MUX2_X1 U10028 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7736), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n7737) );
  NAND2_X1 U10029 ( .A1(n7737), .A2(n7744), .ZN(n10748) );
  INV_X1 U10030 ( .A(n10748), .ZN(n10753) );
  AOI22_X1 U10031 ( .A1(n8391), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6504), .B2(
        n10753), .ZN(n7738) );
  NAND2_X1 U10032 ( .A1(n7739), .A2(n7738), .ZN(n14881) );
  INV_X1 U10033 ( .A(n14881), .ZN(n12079) );
  NAND2_X1 U10034 ( .A1(n11657), .A2(n12079), .ZN(n11721) );
  OR2_X1 U10035 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  NAND2_X1 U10036 ( .A1(n7743), .A2(n7742), .ZN(n10442) );
  OR2_X1 U10037 ( .A1(n10442), .A2(n7813), .ZN(n7749) );
  NAND2_X1 U10038 ( .A1(n7744), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7745) );
  MUX2_X1 U10039 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7745), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n7746) );
  INV_X1 U10040 ( .A(n7746), .ZN(n7747) );
  NOR2_X1 U10041 ( .A1(n7747), .A2(n7752), .ZN(n14138) );
  AOI22_X1 U10042 ( .A1(n8391), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6504), .B2(
        n14138), .ZN(n7748) );
  XNOR2_X1 U10043 ( .A(n7751), .B(n7750), .ZN(n10509) );
  NAND2_X1 U10044 ( .A1(n10509), .A2(n8390), .ZN(n7756) );
  INV_X1 U10045 ( .A(n7752), .ZN(n7753) );
  NAND2_X1 U10046 ( .A1(n7753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7754) );
  XNOR2_X1 U10047 ( .A(n7754), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U10048 ( .A1(n8391), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6503), 
        .B2(n10785), .ZN(n7755) );
  XNOR2_X1 U10049 ( .A(n7758), .B(n7757), .ZN(n10517) );
  NAND2_X1 U10050 ( .A1(n10517), .A2(n8390), .ZN(n7762) );
  NAND2_X1 U10051 ( .A1(n7759), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7760) );
  XNOR2_X1 U10052 ( .A(n7760), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U10053 ( .A1(n8391), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6503), 
        .B2(n11126), .ZN(n7761) );
  INV_X1 U10054 ( .A(n12319), .ZN(n14716) );
  XNOR2_X1 U10055 ( .A(n7764), .B(n7763), .ZN(n10561) );
  NAND2_X1 U10056 ( .A1(n10561), .A2(n8390), .ZN(n7768) );
  NAND2_X1 U10057 ( .A1(n7765), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7766) );
  XNOR2_X1 U10058 ( .A(n7766), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14788) );
  AOI22_X1 U10059 ( .A1(n8391), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n14788), 
        .B2(n6504), .ZN(n7767) );
  INV_X1 U10060 ( .A(n12387), .ZN(n14556) );
  INV_X1 U10061 ( .A(SI_13_), .ZN(n10440) );
  XNOR2_X1 U10062 ( .A(n7769), .B(n10440), .ZN(n7770) );
  XNOR2_X1 U10063 ( .A(n7771), .B(n7770), .ZN(n10792) );
  NAND2_X1 U10064 ( .A1(n10792), .A2(n8390), .ZN(n7774) );
  XNOR2_X1 U10065 ( .A(n7772), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U10066 ( .A1(n11775), .A2(n6503), .B1(n8391), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n7773) );
  XNOR2_X1 U10067 ( .A(n7775), .B(n10797), .ZN(n7776) );
  XNOR2_X1 U10068 ( .A(n7777), .B(n7776), .ZN(n11355) );
  NAND2_X1 U10069 ( .A1(n11355), .A2(n8390), .ZN(n7780) );
  NAND2_X1 U10070 ( .A1(n7787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7778) );
  XNOR2_X1 U10071 ( .A(n7778), .B(P1_IR_REG_17__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U10072 ( .A1(n8391), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6503), 
        .B2(n12239), .ZN(n7779) );
  XNOR2_X1 U10073 ( .A(n7781), .B(SI_18_), .ZN(n7783) );
  NAND2_X1 U10074 ( .A1(n7783), .A2(n7782), .ZN(n7793) );
  INV_X1 U10075 ( .A(n7783), .ZN(n7785) );
  NAND2_X1 U10076 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  INV_X1 U10077 ( .A(n7797), .ZN(n7788) );
  NAND2_X1 U10078 ( .A1(n7788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7789) );
  XNOR2_X1 U10079 ( .A(n7789), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U10080 ( .A1(n8391), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6504), 
        .B2(n14162), .ZN(n7790) );
  NAND2_X2 U10081 ( .A1(n7791), .A2(n7790), .ZN(n14470) );
  INV_X1 U10082 ( .A(SI_18_), .ZN(n10832) );
  OR2_X1 U10083 ( .A1(n7781), .A2(n10832), .ZN(n7792) );
  NAND2_X1 U10084 ( .A1(n7793), .A2(n7792), .ZN(n7796) );
  XNOR2_X1 U10085 ( .A(n7794), .B(SI_19_), .ZN(n7795) );
  NAND2_X1 U10086 ( .A1(n11745), .A2(n8390), .ZN(n7802) );
  NAND2_X1 U10087 ( .A1(n6573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7799) );
  MUX2_X1 U10088 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7799), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n7800) );
  AOI22_X1 U10089 ( .A1(n8391), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6503), 
        .B2(n11874), .ZN(n7801) );
  NAND2_X1 U10090 ( .A1(n7804), .A2(n7803), .ZN(n7805) );
  NAND2_X1 U10091 ( .A1(n7806), .A2(n7805), .ZN(n11747) );
  NAND2_X1 U10092 ( .A1(n8391), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7807) );
  NAND2_X2 U10093 ( .A1(n7808), .A2(n7807), .ZN(n14455) );
  NOR2_X1 U10094 ( .A1(n14331), .A2(n14455), .ZN(n14456) );
  OR2_X1 U10095 ( .A1(n7810), .A2(n7809), .ZN(n7811) );
  NAND2_X1 U10096 ( .A1(n7812), .A2(n7811), .ZN(n12588) );
  NAND2_X1 U10097 ( .A1(n8391), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7814) );
  INV_X1 U10098 ( .A(n14449), .ZN(n14302) );
  NAND2_X1 U10099 ( .A1(n14456), .A2(n14302), .ZN(n14296) );
  XNOR2_X1 U10100 ( .A(n7816), .B(SI_26_), .ZN(n7817) );
  NAND2_X1 U10101 ( .A1(n13776), .A2(n8390), .ZN(n7820) );
  NAND2_X1 U10102 ( .A1(n8391), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7819) );
  AOI21_X1 U10103 ( .B1(n8342), .B2(n12432), .A(n14182), .ZN(n10331) );
  INV_X1 U10104 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7822) );
  OAI21_X2 U10105 ( .B1(n7824), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7825) );
  INV_X2 U10106 ( .A(n8422), .ZN(n11743) );
  NAND2_X1 U10107 ( .A1(n11743), .A2(n14172), .ZN(n8171) );
  INV_X1 U10108 ( .A(n8171), .ZN(n7827) );
  INV_X1 U10109 ( .A(n7828), .ZN(n14101) );
  INV_X1 U10110 ( .A(P1_B_REG_SCAN_IN), .ZN(n7829) );
  NOR2_X1 U10111 ( .A1(n14516), .A2(n7829), .ZN(n7830) );
  NOR2_X1 U10112 ( .A1(n14351), .A2(n7830), .ZN(n14178) );
  INV_X1 U10113 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7832) );
  OR2_X2 U10114 ( .A1(n14506), .A2(n7832), .ZN(n7833) );
  INV_X1 U10115 ( .A(n7841), .ZN(n12443) );
  NAND2_X1 U10116 ( .A1(n7834), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7835) );
  INV_X1 U10117 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10118 ( .A1(n8083), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10119 ( .A1(n8358), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7836) );
  OAI211_X1 U10120 ( .C1(n8086), .C2(n7838), .A(n7837), .B(n7836), .ZN(n14067)
         );
  NAND2_X1 U10121 ( .A1(n14178), .A2(n14067), .ZN(n10326) );
  OAI21_X1 U10122 ( .B1(n6799), .B2(n14875), .A(n10326), .ZN(n7839) );
  AOI21_X1 U10123 ( .B1(n10331), .B2(n14883), .A(n7839), .ZN(n8097) );
  NAND2_X1 U10124 ( .A1(n7867), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10125 ( .A1(n7853), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10126 ( .A1(n7852), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U10128 ( .A1(n7853), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10129 ( .A1(n7852), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7846) );
  INV_X1 U10130 ( .A(n8197), .ZN(n7850) );
  NAND2_X1 U10131 ( .A1(n7851), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7857) );
  NAND2_X1 U10132 ( .A1(n7852), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10133 ( .A1(n7867), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10134 ( .A1(n7853), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7854) );
  XNOR2_X2 U10135 ( .A(n14086), .B(n14845), .ZN(n11561) );
  INV_X1 U10136 ( .A(n14086), .ZN(n11117) );
  INV_X1 U10137 ( .A(n14845), .ZN(n8209) );
  NAND2_X1 U10138 ( .A1(n11117), .A2(n8209), .ZN(n7858) );
  OAI21_X1 U10139 ( .B1(n11559), .B2(n11561), .A(n7858), .ZN(n11053) );
  NAND2_X1 U10140 ( .A1(n8357), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10141 ( .A1(n7851), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10142 ( .A1(n7852), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7861) );
  INV_X1 U10143 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10144 ( .A1(n7867), .A2(n7859), .ZN(n7860) );
  AND2_X1 U10145 ( .A1(n7861), .A2(n7860), .ZN(n7862) );
  NAND2_X1 U10146 ( .A1(n11053), .A2(n11054), .ZN(n7866) );
  INV_X1 U10147 ( .A(n14085), .ZN(n11629) );
  NAND2_X1 U10148 ( .A1(n11629), .A2(n13916), .ZN(n7865) );
  NAND2_X1 U10149 ( .A1(n7866), .A2(n7865), .ZN(n11687) );
  NAND2_X1 U10150 ( .A1(n8357), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10151 ( .A1(n7852), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10152 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7874) );
  OAI21_X1 U10153 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7874), .ZN(n11630) );
  INV_X1 U10154 ( .A(n11630), .ZN(n11683) );
  NAND2_X1 U10155 ( .A1(n6482), .A2(n11683), .ZN(n7869) );
  NAND2_X1 U10156 ( .A1(n8356), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7868) );
  AND4_X2 U10157 ( .A1(n7871), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n11591)
         );
  INV_X1 U10158 ( .A(n14850), .ZN(n11684) );
  AND2_X1 U10159 ( .A1(n11591), .A2(n11684), .ZN(n7872) );
  NAND2_X1 U10160 ( .A1(n8357), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10161 ( .A1(n7851), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7878) );
  AND2_X1 U10162 ( .A1(n7874), .A2(n7873), .ZN(n7875) );
  NOR2_X1 U10163 ( .A1(n7882), .A2(n7875), .ZN(n11605) );
  NAND2_X1 U10164 ( .A1(n7867), .A2(n11605), .ZN(n7877) );
  NAND2_X1 U10165 ( .A1(n7852), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10166 ( .A1(n11854), .A2(n11600), .ZN(n7881) );
  NAND2_X1 U10167 ( .A1(n14083), .A2(n11596), .ZN(n7880) );
  NAND2_X1 U10168 ( .A1(n7881), .A2(n7880), .ZN(n11459) );
  INV_X1 U10169 ( .A(n14864), .ZN(n11476) );
  NAND2_X1 U10170 ( .A1(n8358), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10171 ( .A1(n8357), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10172 ( .A1(n7882), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7892) );
  OR2_X1 U10173 ( .A1(n7882), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7883) );
  AND2_X1 U10174 ( .A1(n7892), .A2(n7883), .ZN(n11856) );
  NAND2_X1 U10175 ( .A1(n6482), .A2(n11856), .ZN(n7885) );
  NAND2_X1 U10176 ( .A1(n8356), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7884) );
  NAND4_X1 U10177 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n14082) );
  NAND2_X1 U10178 ( .A1(n11476), .A2(n14082), .ZN(n7888) );
  INV_X1 U10179 ( .A(n14082), .ZN(n8105) );
  NAND2_X1 U10180 ( .A1(n14864), .A2(n8105), .ZN(n7889) );
  NAND2_X1 U10181 ( .A1(n7890), .A2(n7889), .ZN(n11496) );
  NAND2_X1 U10182 ( .A1(n8083), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10183 ( .A1(n8358), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7896) );
  INV_X1 U10184 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10185 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  AND2_X1 U10186 ( .A1(n7908), .A2(n7893), .ZN(n11505) );
  NAND2_X1 U10187 ( .A1(n6482), .A2(n11505), .ZN(n7895) );
  NAND2_X1 U10188 ( .A1(n8356), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7894) );
  NAND4_X1 U10189 ( .A1(n7897), .A2(n7896), .A3(n7895), .A4(n7894), .ZN(n14081) );
  INV_X1 U10190 ( .A(n14081), .ZN(n11851) );
  AND2_X1 U10191 ( .A1(n12089), .A2(n11851), .ZN(n7899) );
  OR2_X1 U10192 ( .A1(n12089), .A2(n11851), .ZN(n7898) );
  NAND2_X1 U10193 ( .A1(n8357), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10194 ( .A1(n8358), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7902) );
  XNOR2_X1 U10195 ( .A(n7908), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n12076) );
  NAND2_X1 U10196 ( .A1(n6482), .A2(n12076), .ZN(n7901) );
  NAND2_X1 U10197 ( .A1(n8356), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7900) );
  NAND4_X1 U10198 ( .A1(n7903), .A2(n7902), .A3(n7901), .A4(n7900), .ZN(n14080) );
  XNOR2_X1 U10199 ( .A(n14881), .B(n14080), .ZN(n11652) );
  INV_X1 U10200 ( .A(n14080), .ZN(n12161) );
  NOR2_X1 U10201 ( .A1(n14881), .A2(n12161), .ZN(n7904) );
  AOI21_X1 U10202 ( .B1(n11654), .B2(n11652), .A(n7904), .ZN(n11716) );
  NAND2_X1 U10203 ( .A1(n8083), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10204 ( .A1(n8358), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U10205 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n7905) );
  OR2_X1 U10206 ( .A1(n7908), .A2(n7905), .ZN(n7916) );
  INV_X1 U10207 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7907) );
  INV_X1 U10208 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7906) );
  OAI21_X1 U10209 ( .B1(n7908), .B2(n7907), .A(n7906), .ZN(n7909) );
  AND2_X1 U10210 ( .A1(n7916), .A2(n7909), .ZN(n12163) );
  NAND2_X1 U10211 ( .A1(n6482), .A2(n12163), .ZN(n7911) );
  NAND2_X1 U10212 ( .A1(n8356), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7910) );
  NAND4_X1 U10213 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n14079) );
  XNOR2_X1 U10214 ( .A(n12153), .B(n14079), .ZN(n11717) );
  NAND2_X1 U10215 ( .A1(n11716), .A2(n11717), .ZN(n7915) );
  INV_X1 U10216 ( .A(n14079), .ZN(n12209) );
  NAND2_X1 U10217 ( .A1(n12153), .A2(n12209), .ZN(n7914) );
  NAND2_X1 U10218 ( .A1(n7915), .A2(n7914), .ZN(n11871) );
  INV_X1 U10219 ( .A(n11871), .ZN(n7923) );
  NAND2_X1 U10220 ( .A1(n8358), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10221 ( .A1(n8357), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7919) );
  NOR2_X1 U10222 ( .A1(n7932), .A2(n7491), .ZN(n12211) );
  NAND2_X1 U10223 ( .A1(n6482), .A2(n12211), .ZN(n7918) );
  NAND2_X1 U10224 ( .A1(n8356), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7917) );
  NAND4_X1 U10225 ( .A1(n7920), .A2(n7919), .A3(n7918), .A4(n7917), .ZN(n14078) );
  OR2_X1 U10226 ( .A1(n12200), .A2(n12317), .ZN(n7924) );
  NAND2_X1 U10227 ( .A1(n12200), .A2(n12317), .ZN(n7921) );
  NAND2_X1 U10228 ( .A1(n7924), .A2(n7921), .ZN(n11870) );
  INV_X1 U10229 ( .A(n11870), .ZN(n7922) );
  NAND2_X1 U10230 ( .A1(n8358), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7929) );
  INV_X1 U10231 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7925) );
  XNOR2_X1 U10232 ( .A(n7932), .B(n7925), .ZN(n12314) );
  NAND2_X1 U10233 ( .A1(n6482), .A2(n12314), .ZN(n7928) );
  NAND2_X1 U10234 ( .A1(n8356), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U10235 ( .A1(n8357), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7926) );
  NAND4_X1 U10236 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n14077) );
  XNOR2_X1 U10237 ( .A(n12319), .B(n14077), .ZN(n8407) );
  INV_X1 U10238 ( .A(n14077), .ZN(n12395) );
  OR2_X1 U10239 ( .A1(n12319), .A2(n12395), .ZN(n7930) );
  NAND2_X1 U10240 ( .A1(n8358), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U10241 ( .A1(n8357), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7936) );
  AND2_X1 U10242 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n7931) );
  AOI21_X1 U10243 ( .B1(n7932), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n7933) );
  OR2_X1 U10244 ( .A1(n7940), .A2(n7933), .ZN(n11984) );
  INV_X1 U10245 ( .A(n11984), .ZN(n12397) );
  NAND2_X1 U10246 ( .A1(n6482), .A2(n12397), .ZN(n7935) );
  NAND2_X1 U10247 ( .A1(n8356), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7934) );
  NAND4_X1 U10248 ( .A1(n7937), .A2(n7936), .A3(n7935), .A4(n7934), .ZN(n14076) );
  XNOR2_X1 U10249 ( .A(n12387), .B(n14076), .ZN(n11977) );
  NAND2_X1 U10250 ( .A1(n11979), .A2(n11977), .ZN(n7939) );
  INV_X1 U10251 ( .A(n14076), .ZN(n12385) );
  OR2_X1 U10252 ( .A1(n12387), .A2(n12385), .ZN(n7938) );
  NAND2_X1 U10253 ( .A1(n7939), .A2(n7938), .ZN(n12030) );
  NAND2_X1 U10254 ( .A1(n8083), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10255 ( .A1(n8358), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7944) );
  OR2_X1 U10256 ( .A1(n7940), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7941) );
  AND2_X1 U10257 ( .A1(n7941), .A2(n7949), .ZN(n14021) );
  NAND2_X1 U10258 ( .A1(n6482), .A2(n14021), .ZN(n7943) );
  NAND2_X1 U10259 ( .A1(n8356), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7942) );
  NAND4_X1 U10260 ( .A1(n7945), .A2(n7944), .A3(n7943), .A4(n7942), .ZN(n14075) );
  XNOR2_X1 U10261 ( .A(n14710), .B(n14075), .ZN(n8409) );
  NAND2_X1 U10262 ( .A1(n12030), .A2(n8409), .ZN(n7947) );
  INV_X1 U10263 ( .A(n14075), .ZN(n13794) );
  OR2_X1 U10264 ( .A1(n14710), .A2(n13794), .ZN(n7946) );
  NAND2_X1 U10265 ( .A1(n7947), .A2(n7946), .ZN(n12117) );
  NAND2_X1 U10266 ( .A1(n8358), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7954) );
  INV_X1 U10267 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10268 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  NAND2_X1 U10269 ( .A1(n7957), .A2(n7950), .ZN(n14695) );
  INV_X1 U10270 ( .A(n14695), .ZN(n12123) );
  NAND2_X1 U10271 ( .A1(n6482), .A2(n12123), .ZN(n7953) );
  NAND2_X1 U10272 ( .A1(n8356), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10273 ( .A1(n8083), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7951) );
  NAND4_X1 U10274 ( .A1(n7954), .A2(n7953), .A3(n7952), .A4(n7951), .ZN(n14074) );
  INV_X1 U10275 ( .A(n14074), .ZN(n14058) );
  NAND2_X1 U10276 ( .A1(n8083), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10277 ( .A1(n8358), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7961) );
  INV_X1 U10278 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10279 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  AND2_X1 U10280 ( .A1(n7965), .A2(n7958), .ZN(n14062) );
  NAND2_X1 U10281 ( .A1(n6482), .A2(n14062), .ZN(n7960) );
  NAND2_X1 U10282 ( .A1(n8356), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10283 ( .A1(n13812), .A2(n13977), .ZN(n8279) );
  NAND2_X1 U10284 ( .A1(n8280), .A2(n8279), .ZN(n12223) );
  INV_X1 U10285 ( .A(n12223), .ZN(n12228) );
  NAND2_X1 U10286 ( .A1(n8357), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10287 ( .A1(n8358), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7969) );
  INV_X1 U10288 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10289 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  AND2_X1 U10290 ( .A1(n7974), .A2(n7966), .ZN(n14379) );
  NAND2_X1 U10291 ( .A1(n6482), .A2(n14379), .ZN(n7968) );
  NAND2_X1 U10292 ( .A1(n8356), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7967) );
  NAND4_X1 U10293 ( .A1(n7970), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n14365) );
  XNOR2_X1 U10294 ( .A(n14480), .B(n14365), .ZN(n14381) );
  INV_X1 U10295 ( .A(n14381), .ZN(n8123) );
  INV_X1 U10296 ( .A(n14365), .ZN(n13993) );
  NAND2_X1 U10297 ( .A1(n14480), .A2(n13993), .ZN(n7971) );
  NAND2_X1 U10298 ( .A1(n8083), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U10299 ( .A1(n8358), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7978) );
  INV_X1 U10300 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U10301 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  AND2_X1 U10302 ( .A1(n7993), .A2(n7975), .ZN(n14370) );
  NAND2_X1 U10303 ( .A1(n6482), .A2(n14370), .ZN(n7977) );
  NAND2_X1 U10304 ( .A1(n8356), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7976) );
  NAND4_X1 U10305 ( .A1(n7979), .A2(n7978), .A3(n7977), .A4(n7976), .ZN(n14072) );
  INV_X1 U10306 ( .A(n14072), .ZN(n14354) );
  OR2_X1 U10307 ( .A1(n14475), .A2(n14354), .ZN(n7980) );
  NAND2_X1 U10308 ( .A1(n14361), .A2(n7980), .ZN(n7982) );
  NAND2_X1 U10309 ( .A1(n14475), .A2(n14354), .ZN(n7981) );
  NAND2_X1 U10310 ( .A1(n7982), .A2(n7981), .ZN(n14350) );
  INV_X1 U10311 ( .A(n14350), .ZN(n7988) );
  NAND2_X1 U10312 ( .A1(n8357), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10313 ( .A1(n8358), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7985) );
  XNOR2_X1 U10314 ( .A(n7993), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U10315 ( .A1(n6482), .A2(n14345), .ZN(n7984) );
  NAND2_X1 U10316 ( .A1(n8356), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7983) );
  XNOR2_X1 U10317 ( .A(n14470), .B(n13833), .ZN(n14349) );
  OR2_X1 U10318 ( .A1(n14470), .A2(n13833), .ZN(n7989) );
  NAND2_X1 U10319 ( .A1(n8083), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10320 ( .A1(n8358), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7997) );
  INV_X1 U10321 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7991) );
  INV_X1 U10322 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7990) );
  OAI21_X1 U10323 ( .B1(n7993), .B2(n7991), .A(n7990), .ZN(n7994) );
  NAND2_X1 U10324 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7992) );
  AND2_X1 U10325 ( .A1(n7994), .A2(n8001), .ZN(n14333) );
  NAND2_X1 U10326 ( .A1(n6482), .A2(n14333), .ZN(n7996) );
  NAND2_X1 U10327 ( .A1(n8356), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7995) );
  OR2_X1 U10328 ( .A1(n14465), .A2(n14352), .ZN(n8295) );
  NAND2_X1 U10329 ( .A1(n14465), .A2(n14352), .ZN(n8293) );
  NAND2_X1 U10330 ( .A1(n8295), .A2(n8293), .ZN(n8290) );
  INV_X1 U10331 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10332 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  NAND2_X1 U10333 ( .A1(n8010), .A2(n8002), .ZN(n14317) );
  OR2_X1 U10334 ( .A1(n14317), .A2(n7963), .ZN(n8006) );
  NAND2_X1 U10335 ( .A1(n8357), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U10336 ( .A1(n8358), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U10337 ( .A1(n8356), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8003) );
  NAND4_X1 U10338 ( .A1(n8006), .A2(n8005), .A3(n8004), .A4(n8003), .ZN(n14292) );
  INV_X1 U10339 ( .A(n14292), .ZN(n13843) );
  XNOR2_X1 U10340 ( .A(n14455), .B(n13843), .ZN(n14310) );
  NAND2_X1 U10341 ( .A1(n8008), .A2(n8007), .ZN(n14313) );
  OR2_X1 U10342 ( .A1(n14455), .A2(n13843), .ZN(n8009) );
  NAND2_X1 U10343 ( .A1(n14313), .A2(n8009), .ZN(n14291) );
  INV_X1 U10344 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8014) );
  INV_X1 U10345 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13953) );
  NAND2_X1 U10346 ( .A1(n8010), .A2(n13953), .ZN(n8011) );
  NAND2_X1 U10347 ( .A1(n8016), .A2(n8011), .ZN(n14299) );
  OR2_X1 U10348 ( .A1(n14299), .A2(n7963), .ZN(n8013) );
  AOI22_X1 U10349 ( .A1(n8083), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n8358), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n8012) );
  OAI211_X1 U10350 ( .C1(n8086), .C2(n8014), .A(n8013), .B(n8012), .ZN(n14285)
         );
  XNOR2_X1 U10351 ( .A(n14449), .B(n14285), .ZN(n14306) );
  NAND2_X1 U10352 ( .A1(n14302), .A2(n14285), .ZN(n8015) );
  INV_X1 U10353 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U10354 ( .A1(n8016), .A2(n14028), .ZN(n8017) );
  NAND2_X1 U10355 ( .A1(n8032), .A2(n8017), .ZN(n14278) );
  AOI22_X1 U10356 ( .A1(n8083), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n8358), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10357 ( .A1(n8356), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8018) );
  OAI211_X1 U10358 ( .C1(n14278), .C2(n7963), .A(n8019), .B(n8018), .ZN(n14293) );
  XNOR2_X1 U10359 ( .A(n14281), .B(n14293), .ZN(n8415) );
  INV_X1 U10360 ( .A(n14293), .ZN(n13954) );
  NAND2_X1 U10361 ( .A1(n14444), .A2(n13954), .ZN(n8020) );
  XNOR2_X1 U10362 ( .A(n8032), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U10363 ( .A1(n14262), .A2(n6482), .ZN(n8026) );
  INV_X1 U10364 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8023) );
  NAND2_X1 U10365 ( .A1(n8357), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10366 ( .A1(n8358), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8021) );
  OAI211_X1 U10367 ( .C1(n8023), .C2(n8086), .A(n8022), .B(n8021), .ZN(n8024)
         );
  INV_X1 U10368 ( .A(n8024), .ZN(n8025) );
  NAND2_X1 U10369 ( .A1(n8026), .A2(n8025), .ZN(n14284) );
  XNOR2_X1 U10370 ( .A(n14438), .B(n14284), .ZN(n14267) );
  NAND2_X1 U10371 ( .A1(n14258), .A2(n14267), .ZN(n8028) );
  INV_X1 U10372 ( .A(n14284), .ZN(n14029) );
  NAND2_X1 U10373 ( .A1(n14438), .A2(n14029), .ZN(n8027) );
  NAND2_X1 U10374 ( .A1(n8028), .A2(n8027), .ZN(n14246) );
  INV_X1 U10375 ( .A(n14246), .ZN(n8040) );
  INV_X1 U10376 ( .A(n8032), .ZN(n8030) );
  AND2_X1 U10377 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n8029) );
  NAND2_X1 U10378 ( .A1(n8030), .A2(n8029), .ZN(n8044) );
  INV_X1 U10379 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13908) );
  INV_X1 U10380 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8031) );
  OAI21_X1 U10381 ( .B1(n8032), .B2(n13908), .A(n8031), .ZN(n8033) );
  NAND2_X1 U10382 ( .A1(n8044), .A2(n8033), .ZN(n14253) );
  OR2_X1 U10383 ( .A1(n14253), .A2(n7963), .ZN(n8039) );
  INV_X1 U10384 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10385 ( .A1(n8358), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10386 ( .A1(n8083), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8034) );
  OAI211_X1 U10387 ( .C1(n8036), .C2(n8086), .A(n8035), .B(n8034), .ZN(n8037)
         );
  INV_X1 U10388 ( .A(n8037), .ZN(n8038) );
  NAND2_X1 U10389 ( .A1(n8039), .A2(n8038), .ZN(n14228) );
  XNOR2_X1 U10390 ( .A(n14433), .B(n14228), .ZN(n14245) );
  INV_X1 U10391 ( .A(n14433), .ZN(n8140) );
  NAND2_X1 U10392 ( .A1(n8140), .A2(n14228), .ZN(n8041) );
  INV_X1 U10393 ( .A(n8044), .ZN(n8042) );
  NAND2_X1 U10394 ( .A1(n8042), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8055) );
  INV_X1 U10395 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U10396 ( .A1(n8044), .A2(n8043), .ZN(n8045) );
  NAND2_X1 U10397 ( .A1(n8055), .A2(n8045), .ZN(n14232) );
  OR2_X1 U10398 ( .A1(n14232), .A2(n7963), .ZN(n8051) );
  INV_X1 U10399 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10400 ( .A1(n8357), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10401 ( .A1(n8358), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U10402 ( .C1(n8048), .C2(n8086), .A(n8047), .B(n8046), .ZN(n8049)
         );
  INV_X1 U10403 ( .A(n8049), .ZN(n8050) );
  INV_X1 U10404 ( .A(n14070), .ZN(n8052) );
  NAND2_X1 U10405 ( .A1(n14427), .A2(n8052), .ZN(n8053) );
  INV_X1 U10406 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10407 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  NAND2_X1 U10408 ( .A1(n14220), .A2(n6482), .ZN(n8062) );
  INV_X1 U10409 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10410 ( .A1(n8083), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10411 ( .A1(n8358), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8057) );
  OAI211_X1 U10412 ( .C1(n8059), .C2(n8086), .A(n8058), .B(n8057), .ZN(n8060)
         );
  INV_X1 U10413 ( .A(n8060), .ZN(n8061) );
  INV_X1 U10414 ( .A(n14229), .ZN(n8063) );
  INV_X1 U10415 ( .A(n8066), .ZN(n8064) );
  NAND2_X1 U10416 ( .A1(n8064), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8073) );
  INV_X1 U10417 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10418 ( .A1(n8066), .A2(n8065), .ZN(n8067) );
  NAND2_X1 U10419 ( .A1(n8073), .A2(n8067), .ZN(n14203) );
  INV_X1 U10420 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14418) );
  NAND2_X1 U10421 ( .A1(n8357), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10422 ( .A1(n8358), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8068) );
  OAI211_X1 U10423 ( .C1(n14418), .C2(n8086), .A(n8069), .B(n8068), .ZN(n8070)
         );
  INV_X1 U10424 ( .A(n8070), .ZN(n8071) );
  INV_X1 U10425 ( .A(n14069), .ZN(n13941) );
  XNOR2_X1 U10426 ( .A(n14205), .B(n13941), .ZN(n14190) );
  INV_X1 U10427 ( .A(n14205), .ZN(n14414) );
  INV_X1 U10428 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13940) );
  NAND2_X1 U10429 ( .A1(n8073), .A2(n13940), .ZN(n8074) );
  NAND2_X1 U10430 ( .A1(n13942), .A2(n6482), .ZN(n8080) );
  INV_X1 U10431 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10432 ( .A1(n8083), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10433 ( .A1(n8358), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8075) );
  OAI211_X1 U10434 ( .C1(n8077), .C2(n8086), .A(n8076), .B(n8075), .ZN(n8078)
         );
  INV_X1 U10435 ( .A(n8078), .ZN(n8079) );
  NOR2_X1 U10436 ( .A1(n12436), .A2(n14193), .ZN(n8081) );
  INV_X1 U10437 ( .A(n14193), .ZN(n13899) );
  OAI22_X1 U10438 ( .A1(n12427), .A2(n8081), .B1(n13899), .B2(n14409), .ZN(
        n8091) );
  INV_X1 U10439 ( .A(n10327), .ZN(n8082) );
  NAND2_X1 U10440 ( .A1(n8082), .A2(n6482), .ZN(n8090) );
  INV_X1 U10441 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10442 ( .A1(n8083), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U10443 ( .A1(n8358), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8084) );
  OAI211_X1 U10444 ( .C1(n8087), .C2(n8086), .A(n8085), .B(n8084), .ZN(n8088)
         );
  INV_X1 U10445 ( .A(n8088), .ZN(n8089) );
  NAND2_X1 U10446 ( .A1(n8090), .A2(n8089), .ZN(n14068) );
  INV_X1 U10447 ( .A(n14068), .ZN(n13944) );
  XNOR2_X1 U10448 ( .A(n8091), .B(n8419), .ZN(n8096) );
  NAND2_X1 U10449 ( .A1(n8194), .A2(n11874), .ZN(n8094) );
  OR2_X1 U10450 ( .A1(n8092), .A2(n11743), .ZN(n8093) );
  OR2_X1 U10451 ( .A1(n10861), .A2(n7828), .ZN(n14353) );
  INV_X1 U10452 ( .A(n11860), .ZN(n10873) );
  INV_X1 U10453 ( .A(n8100), .ZN(n10896) );
  NAND2_X1 U10454 ( .A1(n10896), .A2(n11704), .ZN(n8101) );
  NAND2_X1 U10455 ( .A1(n11562), .A2(n11561), .ZN(n11560) );
  NAND2_X1 U10456 ( .A1(n11117), .A2(n14845), .ZN(n8102) );
  INV_X1 U10457 ( .A(n11054), .ZN(n11051) );
  NAND2_X1 U10458 ( .A1(n11050), .A2(n11051), .ZN(n11049) );
  INV_X1 U10459 ( .A(n13916), .ZN(n12414) );
  NAND2_X1 U10460 ( .A1(n11629), .A2(n12414), .ZN(n8103) );
  XNOR2_X1 U10461 ( .A(n14864), .B(n14082), .ZN(n11470) );
  INV_X1 U10462 ( .A(n11470), .ZN(n8104) );
  NAND2_X1 U10463 ( .A1(n11469), .A2(n8104), .ZN(n8107) );
  NAND2_X1 U10464 ( .A1(n11476), .A2(n8105), .ZN(n8106) );
  NAND2_X1 U10465 ( .A1(n8107), .A2(n8106), .ZN(n11495) );
  NAND2_X1 U10466 ( .A1(n11495), .A2(n11497), .ZN(n8109) );
  OR2_X1 U10467 ( .A1(n12089), .A2(n14081), .ZN(n8108) );
  NAND2_X1 U10468 ( .A1(n8109), .A2(n8108), .ZN(n11651) );
  INV_X1 U10469 ( .A(n11652), .ZN(n11653) );
  NAND2_X1 U10470 ( .A1(n11651), .A2(n11653), .ZN(n8111) );
  OR2_X1 U10471 ( .A1(n14881), .A2(n14080), .ZN(n8110) );
  INV_X1 U10472 ( .A(n11717), .ZN(n11715) );
  NAND2_X1 U10473 ( .A1(n11714), .A2(n11715), .ZN(n8113) );
  OR2_X1 U10474 ( .A1(n12153), .A2(n14079), .ZN(n8112) );
  NAND2_X1 U10475 ( .A1(n8113), .A2(n8112), .ZN(n11867) );
  OR2_X1 U10476 ( .A1(n12200), .A2(n14078), .ZN(n8114) );
  NAND2_X1 U10477 ( .A1(n11885), .A2(n11886), .ZN(n8116) );
  OR2_X1 U10478 ( .A1(n12319), .A2(n14077), .ZN(n8115) );
  INV_X1 U10479 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U10480 ( .A1(n11976), .A2(n11978), .ZN(n8118) );
  OR2_X1 U10481 ( .A1(n12387), .A2(n14076), .ZN(n8117) );
  NAND2_X1 U10482 ( .A1(n8118), .A2(n8117), .ZN(n12035) );
  NAND2_X1 U10483 ( .A1(n12035), .A2(n12036), .ZN(n8120) );
  OR2_X1 U10484 ( .A1(n14710), .A2(n14075), .ZN(n8119) );
  NAND2_X1 U10485 ( .A1(n14688), .A2(n14074), .ZN(n8121) );
  INV_X1 U10486 ( .A(n13977), .ZN(n14073) );
  OR2_X1 U10487 ( .A1(n13812), .A2(n14073), .ZN(n8122) );
  OR2_X1 U10488 ( .A1(n14480), .A2(n14365), .ZN(n8124) );
  NOR2_X1 U10489 ( .A1(n14475), .A2(n14072), .ZN(n8398) );
  NAND2_X1 U10490 ( .A1(n14475), .A2(n14072), .ZN(n8399) );
  AND2_X1 U10491 ( .A1(n14470), .A2(n14363), .ZN(n8126) );
  NAND2_X1 U10492 ( .A1(n14329), .A2(n8290), .ZN(n8128) );
  INV_X1 U10493 ( .A(n14352), .ZN(n14071) );
  OR2_X1 U10494 ( .A1(n14465), .A2(n14071), .ZN(n8127) );
  NAND2_X1 U10495 ( .A1(n14455), .A2(n14292), .ZN(n8129) );
  INV_X1 U10496 ( .A(n14306), .ZN(n8130) );
  NAND2_X1 U10497 ( .A1(n15401), .A2(n8130), .ZN(n14303) );
  INV_X1 U10498 ( .A(n14285), .ZN(n8132) );
  NAND2_X1 U10499 ( .A1(n14302), .A2(n8132), .ZN(n8133) );
  OR2_X1 U10500 ( .A1(n14444), .A2(n14293), .ZN(n8134) );
  NAND2_X1 U10501 ( .A1(n14438), .A2(n14284), .ZN(n8136) );
  NAND2_X1 U10502 ( .A1(n14270), .A2(n8136), .ZN(n14244) );
  INV_X1 U10503 ( .A(n14244), .ZN(n8138) );
  NAND2_X1 U10504 ( .A1(n8138), .A2(n8137), .ZN(n14242) );
  INV_X1 U10505 ( .A(n14228), .ZN(n8139) );
  NAND2_X1 U10506 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  INV_X1 U10507 ( .A(n14237), .ZN(n8142) );
  NAND2_X1 U10508 ( .A1(n14427), .A2(n14070), .ZN(n8143) );
  INV_X1 U10509 ( .A(n14212), .ZN(n14208) );
  NAND2_X1 U10510 ( .A1(n14420), .A2(n14229), .ZN(n8144) );
  NAND2_X1 U10511 ( .A1(n14211), .A2(n8144), .ZN(n14194) );
  INV_X1 U10512 ( .A(n14194), .ZN(n8145) );
  INV_X1 U10513 ( .A(n14190), .ZN(n14195) );
  OR2_X1 U10514 ( .A1(n14205), .A2(n14069), .ZN(n8146) );
  NAND2_X1 U10515 ( .A1(n14409), .A2(n14193), .ZN(n8149) );
  OR2_X1 U10516 ( .A1(n14409), .A2(n14193), .ZN(n8147) );
  INV_X1 U10517 ( .A(n12439), .ZN(n8148) );
  NAND2_X1 U10518 ( .A1(n12438), .A2(n8149), .ZN(n8150) );
  XNOR2_X1 U10519 ( .A(n8150), .B(n8419), .ZN(n10321) );
  NAND2_X1 U10520 ( .A1(n8194), .A2(n14172), .ZN(n8151) );
  NAND2_X2 U10521 ( .A1(n8364), .A2(n11743), .ZN(n10848) );
  NAND2_X1 U10522 ( .A1(n12151), .A2(n10861), .ZN(n14860) );
  INV_X1 U10523 ( .A(n8194), .ZN(n8152) );
  NAND2_X1 U10524 ( .A1(n8152), .A2(n11743), .ZN(n8394) );
  OR2_X1 U10525 ( .A1(n8394), .A2(n14172), .ZN(n8153) );
  OR2_X2 U10526 ( .A1(n10321), .A2(n14888), .ZN(n8154) );
  INV_X1 U10527 ( .A(n10861), .ZN(n8172) );
  NAND2_X1 U10528 ( .A1(n8161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8156) );
  MUX2_X1 U10529 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8156), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8158) );
  NAND2_X1 U10530 ( .A1(n8158), .A2(n8157), .ZN(n14522) );
  NAND2_X1 U10531 ( .A1(n8159), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8160) );
  MUX2_X1 U10532 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8160), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8162) );
  NAND2_X1 U10533 ( .A1(n8162), .A2(n8161), .ZN(n14523) );
  NOR2_X1 U10534 ( .A1(n14522), .A2(n14523), .ZN(n8166) );
  OR2_X1 U10535 ( .A1(n7787), .A2(n8163), .ZN(n8167) );
  OAI21_X1 U10536 ( .B1(n8167), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8164) );
  MUX2_X1 U10537 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8164), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8165) );
  NAND2_X1 U10538 ( .A1(n8167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8169) );
  XNOR2_X1 U10539 ( .A(n8169), .B(n8168), .ZN(n10319) );
  NAND2_X1 U10540 ( .A1(n10850), .A2(n10319), .ZN(n8170) );
  AOI21_X1 U10541 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n10871) );
  NAND2_X1 U10542 ( .A1(n10871), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10543 ( .A1(n14523), .A2(P1_B_REG_SCAN_IN), .ZN(n8173) );
  MUX2_X1 U10544 ( .A(n8173), .B(P1_B_REG_SCAN_IN), .S(n12379), .Z(n8174) );
  INV_X1 U10545 ( .A(n14522), .ZN(n8188) );
  NOR4_X1 U10546 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8183) );
  NOR4_X1 U10547 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8182) );
  INV_X1 U10548 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14843) );
  INV_X1 U10549 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14842) );
  INV_X1 U10550 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14841) );
  INV_X1 U10551 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14840) );
  NAND4_X1 U10552 ( .A1(n14843), .A2(n14842), .A3(n14841), .A4(n14840), .ZN(
        n8180) );
  NOR4_X1 U10553 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8178) );
  NOR4_X1 U10554 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8177) );
  NOR4_X1 U10555 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8176) );
  NOR4_X1 U10556 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8175) );
  NAND4_X1 U10557 ( .A1(n8178), .A2(n8177), .A3(n8176), .A4(n8175), .ZN(n8179)
         );
  NOR4_X1 U10558 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8180), .A4(n8179), .ZN(n8181) );
  NAND3_X1 U10559 ( .A1(n8183), .A2(n8182), .A3(n8181), .ZN(n8184) );
  NAND2_X1 U10560 ( .A1(n8190), .A2(n8184), .ZN(n10857) );
  INV_X1 U10561 ( .A(n10857), .ZN(n8185) );
  INV_X1 U10562 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8186) );
  AND2_X1 U10563 ( .A1(n14522), .A2(n14523), .ZN(n10411) );
  AOI21_X1 U10564 ( .B1(n8190), .B2(n8186), .A(n10411), .ZN(n10858) );
  INV_X1 U10565 ( .A(n10858), .ZN(n10864) );
  NAND2_X1 U10566 ( .A1(n10869), .A2(n10864), .ZN(n8187) );
  INV_X1 U10567 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8189) );
  NOR2_X1 U10568 ( .A1(n12379), .A2(n8188), .ZN(n10408) );
  INV_X2 U10569 ( .A(n14905), .ZN(n14504) );
  INV_X1 U10570 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U10571 ( .A1(n8099), .A2(n11860), .ZN(n8193) );
  XNOR2_X1 U10572 ( .A(n8194), .B(n14172), .ZN(n8362) );
  NAND2_X2 U10573 ( .A1(n8196), .A2(n8195), .ZN(n8208) );
  XNOR2_X1 U10574 ( .A(n8197), .B(n8223), .ZN(n8198) );
  OAI21_X1 U10575 ( .B1(n11865), .B2(n10848), .A(n8198), .ZN(n8200) );
  NAND2_X1 U10576 ( .A1(n8200), .A2(n8199), .ZN(n8207) );
  NAND2_X1 U10577 ( .A1(n8204), .A2(n8203), .ZN(n8205) );
  NAND2_X1 U10578 ( .A1(n8207), .A2(n8206), .ZN(n8213) );
  NAND2_X1 U10579 ( .A1(n8223), .A2(n14086), .ZN(n8211) );
  NAND2_X1 U10580 ( .A1(n8208), .A2(n11117), .ZN(n8210) );
  NAND3_X1 U10581 ( .A1(n8213), .A2(n8212), .A3(n11054), .ZN(n8217) );
  NAND2_X1 U10582 ( .A1(n8223), .A2(n13916), .ZN(n8215) );
  NAND2_X1 U10583 ( .A1(n8208), .A2(n12414), .ZN(n8214) );
  MUX2_X1 U10584 ( .A(n8215), .B(n8214), .S(n14085), .Z(n8216) );
  NAND2_X1 U10585 ( .A1(n8217), .A2(n8216), .ZN(n8220) );
  MUX2_X1 U10586 ( .A(n11591), .B(n14850), .S(n8208), .Z(n8219) );
  MUX2_X1 U10587 ( .A(n11684), .B(n14084), .S(n8341), .Z(n8218) );
  OAI21_X1 U10588 ( .B1(n8220), .B2(n8219), .A(n8218), .ZN(n8222) );
  NAND2_X1 U10589 ( .A1(n8220), .A2(n8219), .ZN(n8221) );
  NAND2_X1 U10590 ( .A1(n8222), .A2(n8221), .ZN(n8226) );
  INV_X2 U10591 ( .A(n8223), .ZN(n8341) );
  MUX2_X1 U10592 ( .A(n11600), .B(n14083), .S(n8341), .Z(n8227) );
  NAND2_X1 U10593 ( .A1(n8226), .A2(n8227), .ZN(n8225) );
  MUX2_X1 U10594 ( .A(n14083), .B(n11600), .S(n8341), .Z(n8224) );
  NAND2_X1 U10595 ( .A1(n8225), .A2(n8224), .ZN(n8231) );
  INV_X1 U10596 ( .A(n8226), .ZN(n8229) );
  INV_X1 U10597 ( .A(n8227), .ZN(n8228) );
  NAND2_X1 U10598 ( .A1(n8229), .A2(n8228), .ZN(n8230) );
  NAND2_X1 U10599 ( .A1(n8231), .A2(n8230), .ZN(n8233) );
  MUX2_X1 U10600 ( .A(n14864), .B(n14082), .S(n6481), .Z(n8234) );
  MUX2_X1 U10601 ( .A(n14864), .B(n14082), .S(n8341), .Z(n8232) );
  MUX2_X1 U10602 ( .A(n12089), .B(n14081), .S(n8341), .Z(n8238) );
  MUX2_X1 U10603 ( .A(n14081), .B(n12089), .S(n8341), .Z(n8235) );
  NAND2_X1 U10604 ( .A1(n8236), .A2(n8235), .ZN(n8241) );
  INV_X1 U10605 ( .A(n8237), .ZN(n8239) );
  NAND2_X1 U10606 ( .A1(n8239), .A2(n7438), .ZN(n8240) );
  MUX2_X1 U10607 ( .A(n14080), .B(n14881), .S(n8341), .Z(n8243) );
  MUX2_X1 U10608 ( .A(n14080), .B(n14881), .S(n6481), .Z(n8242) );
  INV_X1 U10609 ( .A(n8243), .ZN(n8244) );
  MUX2_X1 U10610 ( .A(n14079), .B(n12153), .S(n6481), .Z(n8248) );
  NAND2_X1 U10611 ( .A1(n8247), .A2(n8248), .ZN(n8246) );
  MUX2_X1 U10612 ( .A(n14079), .B(n12153), .S(n8368), .Z(n8245) );
  NAND2_X1 U10613 ( .A1(n8246), .A2(n8245), .ZN(n8252) );
  INV_X1 U10614 ( .A(n8247), .ZN(n8250) );
  INV_X1 U10615 ( .A(n8248), .ZN(n8249) );
  NAND2_X1 U10616 ( .A1(n8250), .A2(n8249), .ZN(n8251) );
  MUX2_X1 U10617 ( .A(n14078), .B(n12200), .S(n8368), .Z(n8254) );
  MUX2_X1 U10618 ( .A(n14078), .B(n12200), .S(n6481), .Z(n8253) );
  MUX2_X1 U10619 ( .A(n14077), .B(n12319), .S(n6481), .Z(n8258) );
  NAND2_X1 U10620 ( .A1(n8257), .A2(n8258), .ZN(n8256) );
  MUX2_X1 U10621 ( .A(n14077), .B(n12319), .S(n8368), .Z(n8255) );
  NAND2_X1 U10622 ( .A1(n8256), .A2(n8255), .ZN(n8262) );
  INV_X1 U10623 ( .A(n8257), .ZN(n8260) );
  INV_X1 U10624 ( .A(n8258), .ZN(n8259) );
  NAND2_X1 U10625 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  NAND2_X1 U10626 ( .A1(n8262), .A2(n8261), .ZN(n8265) );
  MUX2_X1 U10627 ( .A(n14076), .B(n12387), .S(n8368), .Z(n8266) );
  NAND2_X1 U10628 ( .A1(n8265), .A2(n8266), .ZN(n8264) );
  MUX2_X1 U10629 ( .A(n14076), .B(n12387), .S(n6481), .Z(n8263) );
  NAND2_X1 U10630 ( .A1(n8264), .A2(n8263), .ZN(n8270) );
  INV_X1 U10631 ( .A(n8265), .ZN(n8268) );
  INV_X1 U10632 ( .A(n8266), .ZN(n8267) );
  NAND2_X1 U10633 ( .A1(n8268), .A2(n8267), .ZN(n8269) );
  NAND2_X1 U10634 ( .A1(n8270), .A2(n8269), .ZN(n8273) );
  MUX2_X1 U10635 ( .A(n14075), .B(n14710), .S(n6481), .Z(n8272) );
  MUX2_X1 U10636 ( .A(n14075), .B(n14710), .S(n8368), .Z(n8271) );
  NAND2_X1 U10637 ( .A1(n8280), .A2(n8274), .ZN(n8276) );
  INV_X1 U10638 ( .A(n14688), .ZN(n14703) );
  OAI21_X1 U10639 ( .B1(n14703), .B2(n14074), .A(n8279), .ZN(n8275) );
  MUX2_X1 U10640 ( .A(n8276), .B(n8275), .S(n8368), .Z(n8277) );
  INV_X1 U10641 ( .A(n8277), .ZN(n8278) );
  MUX2_X1 U10642 ( .A(n8280), .B(n8279), .S(n6481), .Z(n8281) );
  MUX2_X1 U10643 ( .A(n14365), .B(n14480), .S(n6481), .Z(n8285) );
  NAND2_X1 U10644 ( .A1(n8284), .A2(n8285), .ZN(n8283) );
  MUX2_X1 U10645 ( .A(n14365), .B(n14480), .S(n8368), .Z(n8282) );
  INV_X1 U10646 ( .A(n8284), .ZN(n8287) );
  INV_X1 U10647 ( .A(n8285), .ZN(n8286) );
  MUX2_X1 U10648 ( .A(n14072), .B(n14475), .S(n8368), .Z(n8288) );
  NOR2_X1 U10649 ( .A1(n8290), .A2(n14349), .ZN(n8289) );
  NAND3_X1 U10650 ( .A1(n14470), .A2(n8368), .A3(n13833), .ZN(n8292) );
  OR3_X1 U10651 ( .A1(n14470), .A2(n8368), .A3(n13833), .ZN(n8291) );
  NAND2_X1 U10652 ( .A1(n8292), .A2(n8291), .ZN(n8297) );
  OR2_X1 U10653 ( .A1(n8293), .A2(n6481), .ZN(n8294) );
  OAI211_X1 U10654 ( .C1(n8295), .C2(n8368), .A(n8294), .B(n8007), .ZN(n8296)
         );
  AOI21_X1 U10655 ( .B1(n14337), .B2(n8297), .A(n8296), .ZN(n8298) );
  NAND2_X1 U10656 ( .A1(n8299), .A2(n8298), .ZN(n8303) );
  AND2_X1 U10657 ( .A1(n8341), .A2(n14292), .ZN(n8301) );
  OAI21_X1 U10658 ( .B1(n8368), .B2(n14292), .A(n14455), .ZN(n8300) );
  OAI21_X1 U10659 ( .B1(n8301), .B2(n14455), .A(n8300), .ZN(n8302) );
  NAND2_X1 U10660 ( .A1(n8303), .A2(n8302), .ZN(n8307) );
  MUX2_X1 U10661 ( .A(n14449), .B(n14285), .S(n6481), .Z(n8304) );
  INV_X1 U10662 ( .A(n8304), .ZN(n8306) );
  MUX2_X1 U10663 ( .A(n14449), .B(n14285), .S(n8368), .Z(n8305) );
  NAND2_X1 U10664 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  NAND2_X1 U10665 ( .A1(n8309), .A2(n8308), .ZN(n8312) );
  MUX2_X1 U10666 ( .A(n14444), .B(n14293), .S(n8341), .Z(n8311) );
  MUX2_X1 U10667 ( .A(n14281), .B(n13954), .S(n6481), .Z(n8310) );
  MUX2_X1 U10668 ( .A(n14284), .B(n14438), .S(n8368), .Z(n8314) );
  MUX2_X1 U10669 ( .A(n14284), .B(n14438), .S(n6481), .Z(n8313) );
  MUX2_X1 U10670 ( .A(n14228), .B(n14433), .S(n8341), .Z(n8316) );
  INV_X1 U10671 ( .A(n8316), .ZN(n8318) );
  MUX2_X1 U10672 ( .A(n14433), .B(n14228), .S(n8368), .Z(n8317) );
  MUX2_X1 U10673 ( .A(n14070), .B(n14427), .S(n8341), .Z(n8322) );
  MUX2_X1 U10674 ( .A(n14070), .B(n14427), .S(n6481), .Z(n8319) );
  NAND2_X1 U10675 ( .A1(n8320), .A2(n8319), .ZN(n8326) );
  INV_X1 U10676 ( .A(n8321), .ZN(n8324) );
  INV_X1 U10677 ( .A(n8322), .ZN(n8323) );
  NAND2_X1 U10678 ( .A1(n8324), .A2(n8323), .ZN(n8325) );
  NAND2_X1 U10679 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  MUX2_X1 U10680 ( .A(n14229), .B(n14420), .S(n6481), .Z(n8329) );
  MUX2_X1 U10681 ( .A(n14229), .B(n14420), .S(n8368), .Z(n8327) );
  MUX2_X1 U10682 ( .A(n14205), .B(n14069), .S(n6481), .Z(n8333) );
  MUX2_X1 U10683 ( .A(n14205), .B(n14069), .S(n8341), .Z(n8330) );
  NAND2_X1 U10684 ( .A1(n8331), .A2(n8330), .ZN(n8337) );
  INV_X1 U10685 ( .A(n8332), .ZN(n8335) );
  INV_X1 U10686 ( .A(n8333), .ZN(n8334) );
  NAND2_X1 U10687 ( .A1(n8335), .A2(n8334), .ZN(n8336) );
  NAND2_X1 U10688 ( .A1(n8337), .A2(n8336), .ZN(n8339) );
  MUX2_X1 U10689 ( .A(n14193), .B(n14409), .S(n6481), .Z(n8340) );
  MUX2_X1 U10690 ( .A(n14193), .B(n14409), .S(n8341), .Z(n8338) );
  MUX2_X1 U10691 ( .A(n14068), .B(n8342), .S(n6481), .Z(n8345) );
  MUX2_X1 U10692 ( .A(n13944), .B(n6799), .S(n8368), .Z(n8343) );
  NAND2_X1 U10693 ( .A1(n8344), .A2(n8343), .ZN(n8347) );
  INV_X1 U10694 ( .A(n8350), .ZN(n8351) );
  NAND2_X1 U10695 ( .A1(n8351), .A2(n13124), .ZN(n8381) );
  NAND2_X1 U10696 ( .A1(n8376), .A2(n8381), .ZN(n8353) );
  MUX2_X1 U10697 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10345), .Z(n8377) );
  INV_X1 U10698 ( .A(n8377), .ZN(n8378) );
  XNOR2_X1 U10699 ( .A(n8378), .B(SI_30_), .ZN(n8352) );
  NAND2_X1 U10700 ( .A1(n12444), .A2(n8390), .ZN(n8355) );
  NAND2_X1 U10701 ( .A1(n8391), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10702 ( .A1(n14184), .A2(n6481), .ZN(n8367) );
  NAND2_X1 U10703 ( .A1(n8356), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10704 ( .A1(n8357), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10705 ( .A1(n8358), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8359) );
  AND3_X1 U10706 ( .A1(n8361), .A2(n8360), .A3(n8359), .ZN(n8425) );
  INV_X1 U10707 ( .A(n8362), .ZN(n8363) );
  OAI22_X1 U10708 ( .A1(n6481), .A2(n8425), .B1(n8364), .B2(n8363), .ZN(n8365)
         );
  NAND2_X1 U10709 ( .A1(n8365), .A2(n14067), .ZN(n8366) );
  NAND2_X1 U10710 ( .A1(n8367), .A2(n8366), .ZN(n8440) );
  INV_X1 U10711 ( .A(n8440), .ZN(n8371) );
  INV_X1 U10712 ( .A(n8425), .ZN(n14179) );
  OAI21_X1 U10713 ( .B1(n14179), .B2(n11743), .A(n14067), .ZN(n8369) );
  MUX2_X1 U10714 ( .A(n8369), .B(n14407), .S(n8368), .Z(n8441) );
  INV_X1 U10715 ( .A(n8441), .ZN(n8370) );
  INV_X1 U10716 ( .A(n8376), .ZN(n8373) );
  MUX2_X1 U10717 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9592), .Z(n8372) );
  INV_X1 U10718 ( .A(SI_31_), .ZN(n13119) );
  XNOR2_X1 U10719 ( .A(n8372), .B(n13119), .ZN(n8383) );
  NAND2_X1 U10720 ( .A1(n8377), .A2(SI_30_), .ZN(n8380) );
  NAND2_X1 U10721 ( .A1(n8373), .A2(n7495), .ZN(n8389) );
  OAI21_X1 U10722 ( .B1(SI_30_), .B2(n8377), .A(n8381), .ZN(n8374) );
  NOR2_X1 U10723 ( .A1(n8374), .A2(n8383), .ZN(n8375) );
  NAND2_X1 U10724 ( .A1(n8376), .A2(n8375), .ZN(n8388) );
  INV_X1 U10725 ( .A(SI_30_), .ZN(n12576) );
  OAI21_X1 U10726 ( .B1(n8383), .B2(n12576), .A(n8377), .ZN(n8386) );
  INV_X1 U10727 ( .A(n8383), .ZN(n8379) );
  OAI21_X1 U10728 ( .B1(n8379), .B2(SI_30_), .A(n8378), .ZN(n8385) );
  INV_X1 U10729 ( .A(n8380), .ZN(n8382) );
  NOR2_X1 U10730 ( .A1(n8382), .A2(n8381), .ZN(n8384) );
  AOI22_X1 U10731 ( .A1(n8386), .A2(n8385), .B1(n8384), .B2(n8383), .ZN(n8387)
         );
  NAND3_X1 U10732 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n13762) );
  NAND2_X1 U10733 ( .A1(n13762), .A2(n8390), .ZN(n8393) );
  NAND2_X1 U10734 ( .A1(n8391), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10735 ( .A1(n10861), .A2(n8394), .ZN(n8396) );
  OR2_X1 U10736 ( .A1(n10848), .A2(n14172), .ZN(n8395) );
  NAND2_X1 U10737 ( .A1(n8396), .A2(n8395), .ZN(n8434) );
  INV_X1 U10738 ( .A(n8434), .ZN(n8397) );
  INV_X1 U10739 ( .A(n8398), .ZN(n8400) );
  NAND2_X1 U10740 ( .A1(n8400), .A2(n8399), .ZN(n14373) );
  INV_X1 U10741 ( .A(n8401), .ZN(n12120) );
  INV_X1 U10742 ( .A(n11561), .ZN(n11558) );
  XNOR2_X1 U10743 ( .A(n14084), .B(n11684), .ZN(n11686) );
  AND2_X1 U10744 ( .A1(n11558), .A2(n11686), .ZN(n8403) );
  NOR3_X1 U10745 ( .A1(n11459), .A2(n11039), .A3(n11865), .ZN(n8402) );
  NAND4_X1 U10746 ( .A1(n11054), .A2(n8403), .A3(n8402), .A4(n11470), .ZN(
        n8404) );
  NOR2_X1 U10747 ( .A1(n8404), .A2(n11497), .ZN(n8405) );
  NAND3_X1 U10748 ( .A1(n11717), .A2(n8405), .A3(n11652), .ZN(n8406) );
  NOR2_X1 U10749 ( .A1(n11870), .A2(n8406), .ZN(n8408) );
  NAND4_X1 U10750 ( .A1(n8409), .A2(n8408), .A3(n11977), .A4(n8407), .ZN(n8410) );
  NOR3_X1 U10751 ( .A1(n12223), .A2(n12120), .A3(n8410), .ZN(n8411) );
  NAND3_X1 U10752 ( .A1(n14373), .A2(n8411), .A3(n14381), .ZN(n8412) );
  NOR2_X1 U10753 ( .A1(n14310), .A2(n8412), .ZN(n8413) );
  NAND4_X1 U10754 ( .A1(n14306), .A2(n14337), .A3(n8413), .A4(n7987), .ZN(
        n8414) );
  NOR2_X1 U10755 ( .A1(n8415), .A2(n8414), .ZN(n8416) );
  NAND4_X1 U10756 ( .A1(n14237), .A2(n8416), .A3(n14245), .A4(n14267), .ZN(
        n8417) );
  NOR2_X1 U10757 ( .A1(n14190), .A2(n8417), .ZN(n8418) );
  NAND2_X1 U10758 ( .A1(n8092), .A2(n8422), .ZN(n8428) );
  AND2_X1 U10759 ( .A1(n8424), .A2(n8425), .ZN(n8427) );
  NOR2_X1 U10760 ( .A1(n8424), .A2(n8425), .ZN(n8426) );
  MUX2_X1 U10761 ( .A(n8427), .B(n8426), .S(n6481), .Z(n8433) );
  INV_X1 U10762 ( .A(n8433), .ZN(n8429) );
  AND2_X1 U10763 ( .A1(n8434), .A2(n8428), .ZN(n8431) );
  NAND2_X1 U10764 ( .A1(n8429), .A2(n8431), .ZN(n8442) );
  INV_X1 U10765 ( .A(n8430), .ZN(n8432) );
  NAND2_X1 U10766 ( .A1(n8432), .A2(n8431), .ZN(n8435) );
  MUX2_X1 U10767 ( .A(n8435), .B(n8434), .S(n8433), .Z(n8437) );
  NAND3_X1 U10768 ( .A1(n7494), .A2(n8440), .A3(n8441), .ZN(n8436) );
  OAI211_X1 U10769 ( .C1(n8442), .C2(n7489), .A(n8437), .B(n8436), .ZN(n8438)
         );
  INV_X1 U10770 ( .A(n10319), .ZN(n10511) );
  NAND2_X1 U10771 ( .A1(n10511), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12193) );
  INV_X1 U10772 ( .A(n12193), .ZN(n8444) );
  NOR3_X1 U10773 ( .A1(n8445), .A2(n14516), .A3(n14353), .ZN(n8447) );
  OAI21_X1 U10774 ( .B1(n8194), .B2(n12193), .A(P1_B_REG_SCAN_IN), .ZN(n8446)
         );
  OR2_X1 U10775 ( .A1(n8447), .A2(n8446), .ZN(n8448) );
  INV_X1 U10776 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15038) );
  XNOR2_X1 U10777 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n8482) );
  INV_X1 U10778 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8481) );
  XNOR2_X1 U10779 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8484) );
  INV_X1 U10780 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8479) );
  INV_X1 U10781 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n8476) );
  XNOR2_X1 U10782 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n8487) );
  INV_X1 U10783 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n8474) );
  XNOR2_X1 U10784 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .ZN(n8524) );
  INV_X1 U10785 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n8469) );
  INV_X1 U10786 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15297) );
  XNOR2_X1 U10787 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n8490) );
  INV_X1 U10788 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15268) );
  XNOR2_X1 U10789 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n8492) );
  INV_X1 U10790 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10791 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n8511) );
  NAND2_X1 U10792 ( .A1(n8500), .A2(n8499), .ZN(n8449) );
  NAND2_X1 U10793 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8451), .ZN(n8453) );
  INV_X1 U10794 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10795 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8455), .ZN(n8456) );
  NAND2_X1 U10796 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8457), .ZN(n8460) );
  INV_X1 U10797 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10798 ( .A1(n8507), .A2(n8458), .ZN(n8459) );
  NAND2_X1 U10799 ( .A1(n8460), .A2(n8459), .ZN(n8512) );
  NAND2_X1 U10800 ( .A1(n8511), .A2(n8512), .ZN(n8461) );
  NAND2_X1 U10801 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n8463), .ZN(n8466) );
  XOR2_X1 U10802 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8463), .Z(n8516) );
  INV_X1 U10803 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10804 ( .A1(n8516), .A2(n8464), .ZN(n8465) );
  NAND2_X1 U10805 ( .A1(n8466), .A2(n8465), .ZN(n8493) );
  NAND2_X1 U10806 ( .A1(n8492), .A2(n8493), .ZN(n8467) );
  NAND2_X1 U10807 ( .A1(n8490), .A2(n8491), .ZN(n8468) );
  NAND2_X1 U10808 ( .A1(n8469), .A2(n8470), .ZN(n8472) );
  XNOR2_X1 U10809 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n8470), .ZN(n8489) );
  NAND2_X1 U10810 ( .A1(n8489), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10811 ( .A1(n8472), .A2(n8471), .ZN(n8525) );
  NAND2_X1 U10812 ( .A1(n8524), .A2(n8525), .ZN(n8473) );
  NAND2_X1 U10813 ( .A1(n8487), .A2(n8488), .ZN(n8475) );
  INV_X1 U10814 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U10815 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8477), .ZN(n8478) );
  AOI22_X1 U10816 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n8479), .B1(n8485), .B2(
        n8478), .ZN(n8483) );
  NAND2_X1 U10817 ( .A1(n8484), .A2(n8483), .ZN(n8480) );
  XNOR2_X1 U10818 ( .A(n8482), .B(n8535), .ZN(n14744) );
  XNOR2_X1 U10819 ( .A(n8484), .B(n8483), .ZN(n14740) );
  XNOR2_X1 U10820 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n8486) );
  XOR2_X1 U10821 ( .A(n8486), .B(n8485), .Z(n14736) );
  XOR2_X1 U10822 ( .A(n8488), .B(n8487), .Z(n8529) );
  XOR2_X1 U10823 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n8489), .Z(n14554) );
  XOR2_X1 U10824 ( .A(n8491), .B(n8490), .Z(n8521) );
  XNOR2_X1 U10825 ( .A(n8493), .B(n8492), .ZN(n8520) );
  INV_X1 U10826 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8494) );
  XNOR2_X1 U10827 ( .A(n8496), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15387) );
  XOR2_X1 U10828 ( .A(n8498), .B(n8497), .Z(n14539) );
  INV_X1 U10829 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8503) );
  NOR2_X1 U10830 ( .A1(n8502), .A2(n8503), .ZN(n8504) );
  AOI21_X1 U10831 ( .B1(n11366), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n8500), .ZN(
        n8501) );
  INV_X1 U10832 ( .A(n8501), .ZN(n15381) );
  NAND2_X1 U10833 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15381), .ZN(n15391) );
  XNOR2_X1 U10834 ( .A(n8503), .B(n8502), .ZN(n15390) );
  NAND2_X1 U10835 ( .A1(n14539), .A2(n14538), .ZN(n14537) );
  NAND2_X1 U10836 ( .A1(n15387), .A2(n15386), .ZN(n8505) );
  AOI21_X1 U10837 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n8505), .A(n15385), .ZN(
        n15377) );
  NAND2_X1 U10838 ( .A1(n8508), .A2(n8509), .ZN(n8510) );
  INV_X1 U10839 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15379) );
  INV_X1 U10840 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8513) );
  NOR2_X1 U10841 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  XOR2_X1 U10842 ( .A(n8512), .B(n8511), .Z(n14543) );
  XNOR2_X1 U10843 ( .A(n8514), .B(n8513), .ZN(n14542) );
  INV_X1 U10844 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8518) );
  XNOR2_X1 U10845 ( .A(n8516), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15384) );
  INV_X1 U10846 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14548) );
  NAND2_X1 U10847 ( .A1(n14546), .A2(n14544), .ZN(n8522) );
  NOR2_X1 U10848 ( .A1(n8521), .A2(n8522), .ZN(n8523) );
  XNOR2_X1 U10849 ( .A(n8522), .B(n8521), .ZN(n14551) );
  INV_X1 U10850 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14550) );
  NOR2_X1 U10851 ( .A1(n14551), .A2(n14550), .ZN(n14549) );
  XOR2_X1 U10852 ( .A(n8525), .B(n8524), .Z(n8526) );
  INV_X1 U10853 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14730) );
  NAND2_X1 U10854 ( .A1(n14731), .A2(n14730), .ZN(n14729) );
  NAND2_X1 U10855 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  NAND2_X1 U10856 ( .A1(n8529), .A2(n8531), .ZN(n8532) );
  INV_X1 U10857 ( .A(n8529), .ZN(n8530) );
  INV_X1 U10858 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U10859 ( .A1(n14736), .A2(n14735), .ZN(n14734) );
  INV_X1 U10860 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8542) );
  XNOR2_X1 U10861 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n8542), .ZN(n8540) );
  INV_X1 U10862 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14813) );
  NOR2_X1 U10863 ( .A1(n14813), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n8534) );
  INV_X1 U10864 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12766) );
  OAI22_X1 U10865 ( .A1(n8535), .A2(n8534), .B1(n12766), .B2(
        P1_ADDR_REG_15__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10866 ( .A(n8540), .B(n8539), .ZN(n8537) );
  NOR2_X1 U10867 ( .A1(n8536), .A2(n8537), .ZN(n14747) );
  OR2_X1 U10868 ( .A1(n8540), .A2(n8539), .ZN(n8541) );
  OAI21_X1 U10869 ( .B1(n8542), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n8541), .ZN(
        n8543) );
  XOR2_X1 U10870 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8543), .Z(n8544) );
  XNOR2_X1 U10871 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8544), .ZN(n14563) );
  NOR2_X1 U10872 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8543), .ZN(n8546) );
  AND2_X1 U10873 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n8544), .ZN(n8545) );
  NOR2_X1 U10874 ( .A1(n8546), .A2(n8545), .ZN(n8550) );
  XOR2_X1 U10875 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n8551) );
  XNOR2_X1 U10876 ( .A(n8550), .B(n8551), .ZN(n8548) );
  NOR2_X1 U10877 ( .A1(n8547), .A2(n8548), .ZN(n14532) );
  NOR2_X1 U10878 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14531), .ZN(n8549) );
  INV_X1 U10879 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n8553) );
  OR2_X1 U10880 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  OAI21_X1 U10881 ( .B1(n8553), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n8552), .ZN(
        n8556) );
  XNOR2_X1 U10882 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n8554) );
  XNOR2_X1 U10883 ( .A(n8554), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8555) );
  XNOR2_X1 U10884 ( .A(n8556), .B(n8555), .ZN(n8718) );
  AOI22_X1 U10885 ( .A1(n11336), .A2(keyinput_g12), .B1(n10394), .B2(
        keyinput_g32), .ZN(n8557) );
  OAI221_X1 U10886 ( .B1(n11336), .B2(keyinput_g12), .C1(n10394), .C2(
        keyinput_g32), .A(n8557), .ZN(n8567) );
  INV_X1 U10887 ( .A(SI_6_), .ZN(n10387) );
  INV_X1 U10888 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14535) );
  AOI22_X1 U10889 ( .A1(n10387), .A2(keyinput_g26), .B1(keyinput_g33), .B2(
        n14535), .ZN(n8558) );
  OAI221_X1 U10890 ( .B1(n10387), .B2(keyinput_g26), .C1(n14535), .C2(
        keyinput_g33), .A(n8558), .ZN(n8566) );
  INV_X1 U10891 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9977) );
  INV_X1 U10892 ( .A(SI_23_), .ZN(n8560) );
  AOI22_X1 U10893 ( .A1(n9977), .A2(keyinput_g45), .B1(keyinput_g9), .B2(n8560), .ZN(n8559) );
  OAI221_X1 U10894 ( .B1(n9977), .B2(keyinput_g45), .C1(n8560), .C2(
        keyinput_g9), .A(n8559), .ZN(n8565) );
  INV_X1 U10895 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8563) );
  INV_X1 U10896 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8562) );
  AOI22_X1 U10897 ( .A1(n8563), .A2(keyinput_g36), .B1(n8562), .B2(
        keyinput_g42), .ZN(n8561) );
  OAI221_X1 U10898 ( .B1(n8563), .B2(keyinput_g36), .C1(n8562), .C2(
        keyinput_g42), .A(n8561), .ZN(n8564) );
  NOR4_X1 U10899 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n8597)
         );
  AOI22_X1 U10900 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n8568) );
  OAI221_X1 U10901 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n8568), .ZN(n8575) );
  AOI22_X1 U10902 ( .A1(SI_4_), .A2(keyinput_g28), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n8569) );
  OAI221_X1 U10903 ( .B1(SI_4_), .B2(keyinput_g28), .C1(SI_22_), .C2(
        keyinput_g10), .A(n8569), .ZN(n8574) );
  INV_X1 U10904 ( .A(SI_5_), .ZN(n10396) );
  INV_X1 U10905 ( .A(P3_WR_REG_SCAN_IN), .ZN(n8664) );
  AOI22_X1 U10906 ( .A1(n10396), .A2(keyinput_g27), .B1(keyinput_g0), .B2(
        n8664), .ZN(n8570) );
  OAI221_X1 U10907 ( .B1(n10396), .B2(keyinput_g27), .C1(n8664), .C2(
        keyinput_g0), .A(n8570), .ZN(n8573) );
  INV_X1 U10908 ( .A(SI_21_), .ZN(n11402) );
  INV_X1 U10909 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15220) );
  AOI22_X1 U10910 ( .A1(n11402), .A2(keyinput_g11), .B1(n15220), .B2(
        keyinput_g52), .ZN(n8571) );
  OAI221_X1 U10911 ( .B1(n11402), .B2(keyinput_g11), .C1(n15220), .C2(
        keyinput_g52), .A(n8571), .ZN(n8572) );
  NOR4_X1 U10912 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n8596)
         );
  AOI22_X1 U10913 ( .A1(n10832), .A2(keyinput_g14), .B1(keyinput_g16), .B2(
        n10546), .ZN(n8576) );
  OAI221_X1 U10914 ( .B1(n10832), .B2(keyinput_g14), .C1(n10546), .C2(
        keyinput_g16), .A(n8576), .ZN(n8583) );
  INV_X1 U10915 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U10916 ( .A1(n10797), .A2(keyinput_g15), .B1(n12608), .B2(
        keyinput_g41), .ZN(n8577) );
  OAI221_X1 U10917 ( .B1(n10797), .B2(keyinput_g15), .C1(n12608), .C2(
        keyinput_g41), .A(n8577), .ZN(n8582) );
  INV_X1 U10918 ( .A(SI_19_), .ZN(n11032) );
  AOI22_X1 U10919 ( .A1(n10440), .A2(keyinput_g19), .B1(n11032), .B2(
        keyinput_g13), .ZN(n8578) );
  OAI221_X1 U10920 ( .B1(n10440), .B2(keyinput_g19), .C1(n11032), .C2(
        keyinput_g13), .A(n8578), .ZN(n8581) );
  AOI22_X1 U10921 ( .A1(n7197), .A2(keyinput_g18), .B1(n10522), .B2(
        keyinput_g17), .ZN(n8579) );
  OAI221_X1 U10922 ( .B1(n7197), .B2(keyinput_g18), .C1(n10522), .C2(
        keyinput_g17), .A(n8579), .ZN(n8580) );
  NOR4_X1 U10923 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n8595)
         );
  INV_X1 U10924 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15203) );
  AOI22_X1 U10925 ( .A1(n15203), .A2(keyinput_g40), .B1(n9756), .B2(
        keyinput_g43), .ZN(n8584) );
  OAI221_X1 U10926 ( .B1(n15203), .B2(keyinput_g40), .C1(n9756), .C2(
        keyinput_g43), .A(n8584), .ZN(n8593) );
  INV_X1 U10927 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8586) );
  AOI22_X1 U10928 ( .A1(n7504), .A2(keyinput_g31), .B1(n8586), .B2(
        keyinput_g53), .ZN(n8585) );
  OAI221_X1 U10929 ( .B1(n7504), .B2(keyinput_g31), .C1(n8586), .C2(
        keyinput_g53), .A(n8585), .ZN(n8592) );
  AOI22_X1 U10930 ( .A1(n13128), .A2(keyinput_g4), .B1(keyinput_g2), .B2(
        n12576), .ZN(n8587) );
  OAI221_X1 U10931 ( .B1(n13128), .B2(keyinput_g4), .C1(n12576), .C2(
        keyinput_g2), .A(n8587), .ZN(n8591) );
  INV_X1 U10932 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8589) );
  AOI22_X1 U10933 ( .A1(n7569), .A2(keyinput_g8), .B1(n8589), .B2(keyinput_g55), .ZN(n8588) );
  OAI221_X1 U10934 ( .B1(n7569), .B2(keyinput_g8), .C1(n8589), .C2(
        keyinput_g55), .A(n8588), .ZN(n8590) );
  NOR4_X1 U10935 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), .ZN(n8594)
         );
  AND4_X1 U10936 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n8716)
         );
  OAI22_X1 U10937 ( .A1(SI_29_), .A2(keyinput_g3), .B1(keyinput_g24), .B2(
        SI_8_), .ZN(n8598) );
  AOI221_X1 U10938 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_8_), .C2(
        keyinput_g24), .A(n8598), .ZN(n8605) );
  OAI22_X1 U10939 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .ZN(n8599) );
  AOI221_X1 U10940 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g49), .C2(P3_REG3_REG_5__SCAN_IN), .A(n8599), .ZN(n8604) );
  OAI22_X1 U10941 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n8600) );
  AOI221_X1 U10942 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g39), .C2(P3_REG3_REG_10__SCAN_IN), .A(n8600), .ZN(n8603) );
  OAI22_X1 U10943 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .ZN(n8601) );
  AOI221_X1 U10944 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        keyinput_g54), .C2(P3_REG3_REG_0__SCAN_IN), .A(n8601), .ZN(n8602) );
  NAND4_X1 U10945 ( .A1(n8605), .A2(n8604), .A3(n8603), .A4(n8602), .ZN(n8632)
         );
  OAI22_X1 U10946 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        keyinput_g25), .B2(SI_7_), .ZN(n8606) );
  AOI221_X1 U10947 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        SI_7_), .C2(keyinput_g25), .A(n8606), .ZN(n8612) );
  OAI22_X1 U10948 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        keyinput_g59), .B2(P3_REG3_REG_2__SCAN_IN), .ZN(n8607) );
  AOI221_X1 U10949 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput_g59), .A(n8607), .ZN(n8611) );
  OAI22_X1 U10950 ( .A1(SI_11_), .A2(keyinput_g21), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n8608) );
  AOI221_X1 U10951 ( .B1(SI_11_), .B2(keyinput_g21), .C1(keyinput_g22), .C2(
        SI_10_), .A(n8608), .ZN(n8610) );
  XNOR2_X1 U10952 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_g46), .ZN(n8609)
         );
  NAND4_X1 U10953 ( .A1(n8612), .A2(n8611), .A3(n8610), .A4(n8609), .ZN(n8631)
         );
  OAI22_X1 U10954 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g62), .B2(P3_REG3_REG_26__SCAN_IN), .ZN(n8613) );
  AOI221_X1 U10955 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n8613), .ZN(n8620) );
  OAI22_X1 U10956 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n8614) );
  AOI221_X1 U10957 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        keyinput_g63), .C2(P3_REG3_REG_15__SCAN_IN), .A(n8614), .ZN(n8619) );
  OAI22_X1 U10958 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(SI_3_), 
        .B2(keyinput_g29), .ZN(n8615) );
  AOI221_X1 U10959 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        keyinput_g29), .C2(SI_3_), .A(n8615), .ZN(n8618) );
  OAI22_X1 U10960 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        keyinput_g38), .B2(P3_REG3_REG_23__SCAN_IN), .ZN(n8616) );
  AOI221_X1 U10961 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n8616), .ZN(n8617) );
  NAND4_X1 U10962 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n8630)
         );
  OAI22_X1 U10963 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g44), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n8621) );
  AOI221_X1 U10964 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P3_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n8621), .ZN(n8628) );
  OAI22_X1 U10965 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        SI_26_), .B2(keyinput_g6), .ZN(n8622) );
  AOI221_X1 U10966 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g6), .C2(SI_26_), .A(n8622), .ZN(n8627) );
  OAI22_X1 U10967 ( .A1(SI_9_), .A2(keyinput_g23), .B1(keyinput_g20), .B2(
        SI_12_), .ZN(n8623) );
  AOI221_X1 U10968 ( .B1(SI_9_), .B2(keyinput_g23), .C1(SI_12_), .C2(
        keyinput_g20), .A(n8623), .ZN(n8626) );
  OAI22_X1 U10969 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g5), .B2(SI_27_), .ZN(n8624) );
  AOI221_X1 U10970 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        SI_27_), .C2(keyinput_g5), .A(n8624), .ZN(n8625) );
  NAND4_X1 U10971 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n8629)
         );
  NOR4_X1 U10972 ( .A1(n8632), .A2(n8631), .A3(n8630), .A4(n8629), .ZN(n8715)
         );
  AOI22_X1 U10973 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n8633) );
  OAI221_X1 U10974 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n8633), .ZN(n8640) );
  AOI22_X1 U10975 ( .A1(SI_18_), .A2(keyinput_f14), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n8634) );
  OAI221_X1 U10976 ( .B1(SI_18_), .B2(keyinput_f14), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n8634), .ZN(n8639) );
  AOI22_X1 U10977 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n8635) );
  OAI221_X1 U10978 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n8635), .ZN(n8638) );
  AOI22_X1 U10979 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_19_), .B2(
        keyinput_f13), .ZN(n8636) );
  OAI221_X1 U10980 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_19_), .C2(
        keyinput_f13), .A(n8636), .ZN(n8637) );
  NOR4_X1 U10981 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n8709)
         );
  AOI22_X1 U10982 ( .A1(SI_21_), .A2(keyinput_f11), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n8641) );
  OAI221_X1 U10983 ( .B1(SI_21_), .B2(keyinput_f11), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n8641), .ZN(n8648) );
  AOI22_X1 U10984 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n8642) );
  OAI221_X1 U10985 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n8642), .ZN(n8647) );
  AOI22_X1 U10986 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n8643) );
  OAI221_X1 U10987 ( .B1(SI_28_), .B2(keyinput_f4), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n8643), .ZN(n8646) );
  AOI22_X1 U10988 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n8644) );
  OAI221_X1 U10989 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n8644), .ZN(n8645) );
  NOR4_X1 U10990 ( .A1(n8648), .A2(n8647), .A3(n8646), .A4(n8645), .ZN(n8708)
         );
  AOI22_X1 U10991 ( .A1(SI_0_), .A2(keyinput_f32), .B1(SI_4_), .B2(
        keyinput_f28), .ZN(n8649) );
  OAI221_X1 U10992 ( .B1(SI_0_), .B2(keyinput_f32), .C1(SI_4_), .C2(
        keyinput_f28), .A(n8649), .ZN(n8706) );
  AOI22_X1 U10993 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n8650) );
  OAI221_X1 U10994 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n8650), .ZN(n8705) );
  AOI22_X1 U10995 ( .A1(SI_17_), .A2(keyinput_f15), .B1(n7184), .B2(
        keyinput_f10), .ZN(n8651) );
  OAI221_X1 U10996 ( .B1(SI_17_), .B2(keyinput_f15), .C1(n7184), .C2(
        keyinput_f10), .A(n8651), .ZN(n8661) );
  OAI22_X1 U10997 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n8652) );
  AOI221_X1 U10998 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        keyinput_f58), .C2(P3_REG3_REG_11__SCAN_IN), .A(n8652), .ZN(n8659) );
  OAI22_X1 U10999 ( .A1(SI_15_), .A2(keyinput_f17), .B1(SI_16_), .B2(
        keyinput_f16), .ZN(n8653) );
  AOI221_X1 U11000 ( .B1(SI_15_), .B2(keyinput_f17), .C1(keyinput_f16), .C2(
        SI_16_), .A(n8653), .ZN(n8658) );
  OAI22_X1 U11001 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P3_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n8654) );
  AOI221_X1 U11002 ( .B1(SI_23_), .B2(keyinput_f9), .C1(keyinput_f33), .C2(
        P3_RD_REG_SCAN_IN), .A(n8654), .ZN(n8657) );
  OAI22_X1 U11003 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(
        keyinput_f19), .B2(SI_13_), .ZN(n8655) );
  AOI221_X1 U11004 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        SI_13_), .C2(keyinput_f19), .A(n8655), .ZN(n8656) );
  NAND4_X1 U11005 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n8660)
         );
  AOI211_X1 U11006 ( .C1(keyinput_f51), .C2(P3_REG3_REG_24__SCAN_IN), .A(n8661), .B(n8660), .ZN(n8662) );
  OAI21_X1 U11007 ( .B1(keyinput_f51), .B2(P3_REG3_REG_24__SCAN_IN), .A(n8662), 
        .ZN(n8704) );
  AOI22_X1 U11008 ( .A1(n9864), .A2(keyinput_f37), .B1(keyinput_f0), .B2(n8664), .ZN(n8663) );
  OAI221_X1 U11009 ( .B1(n9864), .B2(keyinput_f37), .C1(n8664), .C2(
        keyinput_f0), .A(n8663), .ZN(n8671) );
  INV_X1 U11010 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15160) );
  INV_X1 U11011 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U11012 ( .A1(n15160), .A2(keyinput_f35), .B1(n9914), .B2(
        keyinput_f50), .ZN(n8665) );
  OAI221_X1 U11013 ( .B1(n15160), .B2(keyinput_f35), .C1(n9914), .C2(
        keyinput_f50), .A(n8665), .ZN(n8670) );
  INV_X1 U11014 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U11015 ( .A1(n12270), .A2(keyinput_f56), .B1(keyinput_f52), .B2(
        n15220), .ZN(n8666) );
  OAI221_X1 U11016 ( .B1(n12270), .B2(keyinput_f56), .C1(n15220), .C2(
        keyinput_f52), .A(n8666), .ZN(n8669) );
  INV_X1 U11017 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9614) );
  AOI22_X1 U11018 ( .A1(n12169), .A2(keyinput_f7), .B1(n9614), .B2(
        keyinput_f38), .ZN(n8667) );
  OAI221_X1 U11019 ( .B1(n12169), .B2(keyinput_f7), .C1(n9614), .C2(
        keyinput_f38), .A(n8667), .ZN(n8668) );
  NOR4_X1 U11020 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n8702)
         );
  AOI22_X1 U11021 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n8672) );
  OAI221_X1 U11022 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n8672), .ZN(n8679) );
  AOI22_X1 U11023 ( .A1(SI_20_), .A2(keyinput_f12), .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n8673) );
  OAI221_X1 U11024 ( .B1(SI_20_), .B2(keyinput_f12), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n8673), .ZN(n8678) );
  INV_X1 U11025 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U11026 ( .A1(n12765), .A2(keyinput_f63), .B1(keyinput_f26), .B2(
        n10387), .ZN(n8674) );
  OAI221_X1 U11027 ( .B1(n12765), .B2(keyinput_f63), .C1(n10387), .C2(
        keyinput_f26), .A(n8674), .ZN(n8677) );
  AOI22_X1 U11028 ( .A1(SI_10_), .A2(keyinput_f22), .B1(n10378), .B2(
        keyinput_f21), .ZN(n8675) );
  OAI221_X1 U11029 ( .B1(SI_10_), .B2(keyinput_f22), .C1(n10378), .C2(
        keyinput_f21), .A(n8675), .ZN(n8676) );
  NOR4_X1 U11030 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n8701)
         );
  INV_X1 U11031 ( .A(SI_8_), .ZN(n10372) );
  INV_X1 U11032 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U11033 ( .A1(n10372), .A2(keyinput_f24), .B1(keyinput_f54), .B2(
        n11365), .ZN(n8680) );
  OAI221_X1 U11034 ( .B1(n10372), .B2(keyinput_f24), .C1(n11365), .C2(
        keyinput_f54), .A(n8680), .ZN(n8687) );
  AOI22_X1 U11035 ( .A1(n13124), .A2(keyinput_f3), .B1(keyinput_f31), .B2(
        n7504), .ZN(n8681) );
  OAI221_X1 U11036 ( .B1(n13124), .B2(keyinput_f3), .C1(n7504), .C2(
        keyinput_f31), .A(n8681), .ZN(n8686) );
  AOI22_X1 U11037 ( .A1(n13119), .A2(keyinput_f1), .B1(n7197), .B2(
        keyinput_f18), .ZN(n8682) );
  OAI221_X1 U11038 ( .B1(n13119), .B2(keyinput_f1), .C1(n7197), .C2(
        keyinput_f18), .A(n8682), .ZN(n8685) );
  INV_X1 U11039 ( .A(SI_27_), .ZN(n12447) );
  AOI22_X1 U11040 ( .A1(n9977), .A2(keyinput_f45), .B1(keyinput_f5), .B2(
        n12447), .ZN(n8683) );
  OAI221_X1 U11041 ( .B1(n9977), .B2(keyinput_f45), .C1(n12447), .C2(
        keyinput_f5), .A(n8683), .ZN(n8684) );
  NOR4_X1 U11042 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n8700)
         );
  INV_X1 U11043 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10984) );
  INV_X1 U11044 ( .A(SI_26_), .ZN(n8689) );
  AOI22_X1 U11045 ( .A1(n10984), .A2(keyinput_f59), .B1(keyinput_f6), .B2(
        n8689), .ZN(n8688) );
  OAI221_X1 U11046 ( .B1(n10984), .B2(keyinput_f59), .C1(n8689), .C2(
        keyinput_f6), .A(n8688), .ZN(n8698) );
  INV_X1 U11047 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8691) );
  AOI22_X1 U11048 ( .A1(n15203), .A2(keyinput_f40), .B1(n8691), .B2(
        keyinput_f48), .ZN(n8690) );
  OAI221_X1 U11049 ( .B1(n15203), .B2(keyinput_f40), .C1(n8691), .C2(
        keyinput_f48), .A(n8690), .ZN(n8697) );
  INV_X1 U11050 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n8693) );
  AOI22_X1 U11051 ( .A1(n8693), .A2(keyinput_f61), .B1(n12012), .B2(
        keyinput_f46), .ZN(n8692) );
  OAI221_X1 U11052 ( .B1(n8693), .B2(keyinput_f61), .C1(n12012), .C2(
        keyinput_f46), .A(n8692), .ZN(n8696) );
  INV_X1 U11053 ( .A(SI_9_), .ZN(n10346) );
  AOI22_X1 U11054 ( .A1(n7569), .A2(keyinput_f8), .B1(keyinput_f23), .B2(
        n10346), .ZN(n8694) );
  OAI221_X1 U11055 ( .B1(n7569), .B2(keyinput_f8), .C1(n10346), .C2(
        keyinput_f23), .A(n8694), .ZN(n8695) );
  NOR4_X1 U11056 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(n8699)
         );
  NAND4_X1 U11057 ( .A1(n8702), .A2(n8701), .A3(n8700), .A4(n8699), .ZN(n8703)
         );
  NOR4_X1 U11058 ( .A1(n8706), .A2(n8705), .A3(n8704), .A4(n8703), .ZN(n8707)
         );
  NAND3_X1 U11059 ( .A1(n8709), .A2(n8708), .A3(n8707), .ZN(n8711) );
  AOI21_X1 U11060 ( .B1(keyinput_f30), .B2(n8711), .A(SI_2_), .ZN(n8713) );
  INV_X1 U11061 ( .A(keyinput_f30), .ZN(n8710) );
  AOI21_X1 U11062 ( .B1(n8711), .B2(n8710), .A(keyinput_g30), .ZN(n8712) );
  AOI22_X1 U11063 ( .A1(keyinput_g30), .A2(n8713), .B1(SI_2_), .B2(n8712), 
        .ZN(n8714) );
  AOI21_X1 U11064 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8717) );
  XNOR2_X1 U11065 ( .A(n8718), .B(n8717), .ZN(n8719) );
  NAND2_X1 U11066 ( .A1(n8721), .A2(n14916), .ZN(n8723) );
  NAND2_X1 U11067 ( .A1(n14917), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8722) );
  INV_X1 U11068 ( .A(n8892), .ZN(n8737) );
  NOR2_X2 U11069 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8727) );
  NOR2_X2 U11070 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n8726) );
  NAND4_X1 U11071 ( .A1(n8793), .A2(n8798), .A3(n8730), .A4(n8729), .ZN(n8731)
         );
  NOR2_X2 U11072 ( .A1(n8786), .A2(n8731), .ZN(n8771) );
  NOR2_X1 U11073 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8734) );
  NOR2_X1 U11074 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8733) );
  NOR2_X1 U11075 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8732) );
  INV_X1 U11076 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11077 ( .A1(n8746), .A2(n8739), .ZN(n8747) );
  INV_X1 U11078 ( .A(n8816), .ZN(n8749) );
  NAND2_X1 U11079 ( .A1(n13766), .A2(n9468), .ZN(n8751) );
  NAND2_X1 U11080 ( .A1(n9097), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8750) );
  INV_X1 U11081 ( .A(n8762), .ZN(n8753) );
  NAND2_X1 U11082 ( .A1(n8753), .A2(n8752), .ZN(n8759) );
  NAND2_X1 U11083 ( .A1(n8759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U11084 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8754), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8757) );
  INV_X1 U11085 ( .A(n8755), .ZN(n8756) );
  NAND2_X1 U11086 ( .A1(n8762), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8758) );
  MUX2_X1 U11087 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8758), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8760) );
  NAND2_X1 U11088 ( .A1(n8760), .A2(n8759), .ZN(n13780) );
  NAND2_X1 U11089 ( .A1(n8748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8761) );
  MUX2_X1 U11090 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8761), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8763) );
  NAND2_X1 U11091 ( .A1(n8763), .A2(n8762), .ZN(n12378) );
  XNOR2_X1 U11092 ( .A(n12378), .B(P2_B_REG_SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11093 ( .A1(n13780), .A2(n8764), .ZN(n8765) );
  INV_X1 U11094 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15092) );
  NAND2_X1 U11095 ( .A1(n15055), .A2(n15092), .ZN(n8767) );
  INV_X1 U11096 ( .A(n8769), .ZN(n13778) );
  NAND2_X1 U11097 ( .A1(n13778), .A2(n13780), .ZN(n8766) );
  NOR2_X1 U11098 ( .A1(n13780), .A2(n12378), .ZN(n8768) );
  NAND2_X1 U11099 ( .A1(n8769), .A2(n8768), .ZN(n10683) );
  NOR2_X2 U11100 ( .A1(n8892), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8911) );
  INV_X1 U11101 ( .A(n8998), .ZN(n8773) );
  INV_X1 U11102 ( .A(n8771), .ZN(n8772) );
  OAI21_X1 U11103 ( .B1(n8773), .B2(n8772), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8775) );
  INV_X1 U11104 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8774) );
  XNOR2_X1 U11105 ( .A(n8775), .B(n8774), .ZN(n10682) );
  INV_X1 U11106 ( .A(n15090), .ZN(n15093) );
  NOR2_X1 U11107 ( .A1(n11202), .A2(n15093), .ZN(n15091) );
  NOR4_X1 U11108 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8779) );
  NOR4_X1 U11109 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8778) );
  NOR4_X1 U11110 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8777) );
  NOR4_X1 U11111 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8776) );
  NAND4_X1 U11112 ( .A1(n8779), .A2(n8778), .A3(n8777), .A4(n8776), .ZN(n8785)
         );
  NOR2_X1 U11113 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8783) );
  NOR4_X1 U11114 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8782) );
  NOR4_X1 U11115 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8781) );
  NOR4_X1 U11116 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8780) );
  NAND4_X1 U11117 ( .A1(n8783), .A2(n8782), .A3(n8781), .A4(n8780), .ZN(n8784)
         );
  OAI21_X1 U11118 ( .B1(n8785), .B2(n8784), .A(n15055), .ZN(n11203) );
  AND2_X1 U11119 ( .A1(n8795), .A2(n8798), .ZN(n8788) );
  OAI21_X2 U11120 ( .B1(n8790), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8789) );
  XNOR2_X2 U11121 ( .A(n8789), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11122 ( .A1(n9217), .A2(n9529), .ZN(n10677) );
  NAND2_X1 U11123 ( .A1(n8801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8794) );
  XNOR2_X1 U11124 ( .A(n8794), .B(n8793), .ZN(n9215) );
  NAND2_X1 U11125 ( .A1(n8803), .A2(n13379), .ZN(n9531) );
  INV_X1 U11126 ( .A(n9531), .ZN(n10679) );
  OR2_X1 U11127 ( .A1(n10677), .A2(n10679), .ZN(n11201) );
  AND2_X1 U11128 ( .A1(n11203), .A2(n11201), .ZN(n8804) );
  INV_X1 U11129 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U11130 ( .A1(n15055), .A2(n15088), .ZN(n8806) );
  NAND2_X1 U11131 ( .A1(n13778), .A2(n12378), .ZN(n8805) );
  NAND2_X1 U11132 ( .A1(n8806), .A2(n8805), .ZN(n15089) );
  INV_X1 U11133 ( .A(n15089), .ZN(n10675) );
  NAND2_X1 U11134 ( .A1(n12192), .A2(n9468), .ZN(n8808) );
  NAND2_X1 U11135 ( .A1(n9097), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11136 ( .A1(n8915), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8928) );
  INV_X1 U11137 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8927) );
  NOR2_X1 U11138 ( .A1(n8928), .A2(n8927), .ZN(n8943) );
  NAND2_X1 U11139 ( .A1(n8943), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11140 ( .A1(n9002), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9018) );
  INV_X1 U11141 ( .A(n9018), .ZN(n8809) );
  NAND2_X1 U11142 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8810) );
  INV_X1 U11143 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9086) );
  INV_X1 U11144 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9109) );
  INV_X1 U11145 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13214) );
  INV_X1 U11146 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13147) );
  OAI21_X1 U11147 ( .B1(n9132), .B2(n13214), .A(n13147), .ZN(n8814) );
  AND2_X1 U11148 ( .A1(n8814), .A2(n9145), .ZN(n13504) );
  NAND2_X2 U11149 ( .A1(n13763), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U11150 ( .A1(n13504), .A2(n9183), .ZN(n8825) );
  INV_X1 U11151 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13681) );
  NAND2_X2 U11152 ( .A1(n12579), .A2(n13768), .ZN(n8904) );
  NAND2_X1 U11153 ( .A1(n9206), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11154 ( .A1(n9207), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U11155 ( .C1(n13681), .C2(n9451), .A(n8822), .B(n8821), .ZN(n8823)
         );
  INV_X1 U11156 ( .A(n8823), .ZN(n8824) );
  NAND2_X1 U11157 ( .A1(n8825), .A2(n8824), .ZN(n13512) );
  XNOR2_X1 U11158 ( .A(n13505), .B(n13483), .ZN(n13496) );
  INV_X1 U11159 ( .A(n13496), .ZN(n13499) );
  INV_X1 U11160 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8826) );
  OR2_X1 U11161 ( .A1(n8904), .A2(n8826), .ZN(n8832) );
  INV_X1 U11162 ( .A(n9453), .ZN(n8827) );
  NAND2_X1 U11163 ( .A1(n8827), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8831) );
  INV_X1 U11164 ( .A(n8869), .ZN(n8828) );
  NAND2_X1 U11165 ( .A1(n8828), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8830) );
  INV_X1 U11166 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14942) );
  INV_X1 U11167 ( .A(n9221), .ZN(n11216) );
  NAND2_X1 U11168 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8833) );
  NAND2_X1 U11169 ( .A1(n9221), .A2(n10663), .ZN(n8835) );
  NAND2_X1 U11170 ( .A1(n9592), .A2(SI_0_), .ZN(n8836) );
  XNOR2_X1 U11171 ( .A(n8836), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U11172 ( .A1(n8843), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n8841) );
  INV_X1 U11173 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U11174 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8837) );
  OAI21_X1 U11175 ( .B1(n8838), .B2(P2_IR_REG_30__SCAN_IN), .A(n8837), .ZN(
        n8839) );
  NAND2_X1 U11176 ( .A1(n8849), .A2(n8839), .ZN(n8840) );
  OAI21_X1 U11177 ( .B1(n8849), .B2(n8841), .A(n8840), .ZN(n8842) );
  NAND2_X1 U11178 ( .A1(n8842), .A2(n13768), .ZN(n8853) );
  AOI22_X1 U11179 ( .A1(n8843), .A2(P2_REG3_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n8848) );
  INV_X1 U11180 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11181 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_0__SCAN_IN), 
        .ZN(n8844) );
  OAI21_X1 U11182 ( .B1(n8845), .B2(P2_IR_REG_30__SCAN_IN), .A(n8844), .ZN(
        n8846) );
  NAND2_X1 U11183 ( .A1(n8849), .A2(n8846), .ZN(n8847) );
  OAI21_X1 U11184 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8851) );
  NAND2_X1 U11185 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  INV_X1 U11186 ( .A(n10715), .ZN(n13270) );
  NAND2_X1 U11187 ( .A1(n11276), .A2(n13270), .ZN(n11273) );
  INV_X1 U11188 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8855) );
  INV_X1 U11189 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11237) );
  INV_X1 U11190 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10462) );
  INV_X1 U11191 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8856) );
  OR2_X1 U11192 ( .A1(n9453), .A2(n8856), .ZN(n8857) );
  NAND4_X4 U11193 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n10668) );
  NAND2_X1 U11194 ( .A1(n8861), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8866) );
  INV_X1 U11195 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11196 ( .A1(n8863), .A2(n8862), .ZN(n8876) );
  NAND2_X1 U11197 ( .A1(n8876), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8864) );
  XNOR2_X1 U11198 ( .A(n8864), .B(P2_IR_REG_2__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U11199 ( .A1(n8899), .A2(n14958), .ZN(n8865) );
  OR2_X1 U11200 ( .A1(n10668), .A2(n6477), .ZN(n8867) );
  NAND2_X1 U11201 ( .A1(n8868), .A2(n8867), .ZN(n11224) );
  INV_X1 U11202 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10445) );
  OR2_X1 U11203 ( .A1(n9453), .A2(n10445), .ZN(n8873) );
  INV_X1 U11204 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10464) );
  OR2_X1 U11205 ( .A1(n8869), .A2(n10464), .ZN(n8872) );
  OR2_X1 U11206 ( .A1(n6499), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U11207 ( .A1(n9206), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8874) );
  INV_X1 U11208 ( .A(n8876), .ZN(n8878) );
  INV_X1 U11209 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11210 ( .A1(n8878), .A2(n8877), .ZN(n8890) );
  NAND2_X1 U11211 ( .A1(n8890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8880) );
  XNOR2_X1 U11212 ( .A(n8880), .B(n8879), .ZN(n13272) );
  OAI22_X1 U11213 ( .A1(n8898), .A2(n10342), .B1(n8875), .B2(n13272), .ZN(
        n8881) );
  NAND2_X1 U11214 ( .A1(n11224), .A2(n8883), .ZN(n8885) );
  OR2_X1 U11215 ( .A1(n13268), .A2(n11231), .ZN(n8884) );
  NAND2_X1 U11216 ( .A1(n8885), .A2(n8884), .ZN(n11260) );
  NAND2_X1 U11217 ( .A1(n9206), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8889) );
  INV_X1 U11218 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11266) );
  OR2_X1 U11219 ( .A1(n9453), .A2(n11266), .ZN(n8888) );
  XNOR2_X1 U11220 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n11269) );
  OR2_X1 U11221 ( .A1(n6499), .A2(n11269), .ZN(n8887) );
  INV_X1 U11222 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10466) );
  OR2_X1 U11223 ( .A1(n8869), .A2(n10466), .ZN(n8886) );
  NAND4_X2 U11224 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(n13267) );
  OAI21_X1 U11225 ( .B1(n8890), .B2(P2_IR_REG_3__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8891) );
  MUX2_X1 U11226 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8891), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8893) );
  NAND2_X1 U11227 ( .A1(n8893), .A2(n8892), .ZN(n13286) );
  NAND2_X1 U11228 ( .A1(n8861), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8894) );
  XNOR2_X1 U11229 ( .A(n13267), .B(n11268), .ZN(n11262) );
  INV_X1 U11230 ( .A(n11262), .ZN(n8896) );
  NAND2_X1 U11231 ( .A1(n10367), .A2(n9468), .ZN(n8902) );
  NAND2_X1 U11232 ( .A1(n8892), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8900) );
  XNOR2_X1 U11233 ( .A(n8900), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U11234 ( .A1(n9097), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9096), .B2(
        n10469), .ZN(n8901) );
  AOI21_X1 U11235 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8903) );
  NOR2_X1 U11236 ( .A1(n8903), .A2(n8915), .ZN(n11307) );
  NAND2_X1 U11237 ( .A1(n9183), .A2(n11307), .ZN(n8909) );
  INV_X1 U11238 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11302) );
  OR2_X1 U11239 ( .A1(n9453), .A2(n11302), .ZN(n8908) );
  INV_X1 U11240 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8905) );
  OR2_X1 U11241 ( .A1(n8904), .A2(n8905), .ZN(n8907) );
  INV_X1 U11242 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10468) );
  OR2_X1 U11243 ( .A1(n8869), .A2(n10468), .ZN(n8906) );
  NOR2_X1 U11244 ( .A1(n11306), .A2(n13266), .ZN(n8910) );
  OR2_X1 U11245 ( .A1(n8911), .A2(n8741), .ZN(n8912) );
  XNOR2_X1 U11246 ( .A(n8912), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U11247 ( .A1(n9097), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9096), .B2(
        n10488), .ZN(n8913) );
  NAND2_X1 U11248 ( .A1(n8828), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8920) );
  INV_X1 U11249 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11289) );
  OR2_X1 U11250 ( .A1(n9453), .A2(n11289), .ZN(n8919) );
  OAI21_X1 U11251 ( .B1(n8915), .B2(P2_REG3_REG_6__SCAN_IN), .A(n8928), .ZN(
        n11290) );
  OR2_X1 U11252 ( .A1(n6499), .A2(n11290), .ZN(n8918) );
  INV_X1 U11253 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8916) );
  OR2_X1 U11254 ( .A1(n8904), .A2(n8916), .ZN(n8917) );
  NAND4_X1 U11255 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n13265) );
  XNOR2_X1 U11256 ( .A(n11183), .B(n13265), .ZN(n11175) );
  NAND2_X1 U11257 ( .A1(n11183), .A2(n13265), .ZN(n8921) );
  NAND2_X1 U11258 ( .A1(n8922), .A2(n8921), .ZN(n11312) );
  OR2_X1 U11259 ( .A1(n10404), .A2(n9140), .ZN(n8926) );
  INV_X1 U11260 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U11261 ( .A1(n8911), .A2(n8923), .ZN(n8937) );
  NAND2_X1 U11262 ( .A1(n8937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8924) );
  XNOR2_X1 U11263 ( .A(n8924), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U11264 ( .A1(n9097), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9096), .B2(
        n10500), .ZN(n8925) );
  NAND2_X2 U11265 ( .A1(n8926), .A2(n8925), .ZN(n11332) );
  NAND2_X1 U11266 ( .A1(n8828), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8934) );
  INV_X1 U11267 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11323) );
  OR2_X1 U11268 ( .A1(n9453), .A2(n11323), .ZN(n8933) );
  AND2_X1 U11269 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  OR2_X1 U11270 ( .A1(n8929), .A2(n8943), .ZN(n11315) );
  OR2_X1 U11271 ( .A1(n6499), .A2(n11315), .ZN(n8932) );
  INV_X1 U11272 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8930) );
  OR2_X1 U11273 ( .A1(n8904), .A2(n8930), .ZN(n8931) );
  NAND4_X1 U11274 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(n13264) );
  INV_X1 U11275 ( .A(n13264), .ZN(n9325) );
  XNOR2_X1 U11276 ( .A(n11332), .B(n9325), .ZN(n11318) );
  NAND2_X1 U11277 ( .A1(n11312), .A2(n11318), .ZN(n8936) );
  NAND2_X1 U11278 ( .A1(n11332), .A2(n13264), .ZN(n8935) );
  OR2_X1 U11279 ( .A1(n10416), .A2(n9140), .ZN(n8942) );
  NAND2_X1 U11280 ( .A1(n8939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8938) );
  MUX2_X1 U11281 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8938), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8940) );
  NAND2_X1 U11282 ( .A1(n8940), .A2(n8955), .ZN(n10507) );
  INV_X1 U11283 ( .A(n10507), .ZN(n10528) );
  AOI22_X1 U11284 ( .A1(n9097), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9096), .B2(
        n10528), .ZN(n8941) );
  NAND2_X1 U11285 ( .A1(n9206), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8949) );
  INV_X1 U11286 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11392) );
  OR2_X1 U11287 ( .A1(n9453), .A2(n11392), .ZN(n8948) );
  OR2_X1 U11288 ( .A1(n8943), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11289 ( .A1(n8959), .A2(n8944), .ZN(n11391) );
  OR2_X1 U11290 ( .A1(n6499), .A2(n11391), .ZN(n8947) );
  INV_X1 U11291 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8945) );
  OR2_X1 U11292 ( .A1(n9451), .A2(n8945), .ZN(n8946) );
  NAND4_X1 U11293 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n8946), .ZN(n13263) );
  INV_X1 U11294 ( .A(n13263), .ZN(n11378) );
  NAND2_X1 U11295 ( .A1(n11396), .A2(n11378), .ZN(n9230) );
  OR2_X1 U11296 ( .A1(n11396), .A2(n11378), .ZN(n8950) );
  NAND2_X1 U11297 ( .A1(n9230), .A2(n8950), .ZN(n11387) );
  NAND2_X1 U11298 ( .A1(n11383), .A2(n11387), .ZN(n8952) );
  NAND2_X1 U11299 ( .A1(n11396), .A2(n13263), .ZN(n8951) );
  NAND2_X1 U11300 ( .A1(n8952), .A2(n8951), .ZN(n11481) );
  OR2_X1 U11301 ( .A1(n10442), .A2(n9140), .ZN(n8958) );
  NAND2_X1 U11302 ( .A1(n8955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8953) );
  MUX2_X1 U11303 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8953), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8954) );
  INV_X1 U11304 ( .A(n8954), .ZN(n8956) );
  NOR2_X1 U11305 ( .A1(n8955), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8968) );
  NOR2_X1 U11306 ( .A1(n8956), .A2(n8968), .ZN(n14978) );
  AOI22_X1 U11307 ( .A1(n9097), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9096), .B2(
        n14978), .ZN(n8957) );
  NAND2_X1 U11308 ( .A1(n9206), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8964) );
  INV_X1 U11309 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11490) );
  OR2_X1 U11310 ( .A1(n9453), .A2(n11490), .ZN(n8963) );
  NAND2_X1 U11311 ( .A1(n8959), .A2(n11379), .ZN(n8960) );
  NAND2_X1 U11312 ( .A1(n8972), .A2(n8960), .ZN(n11489) );
  OR2_X1 U11313 ( .A1(n6499), .A2(n11489), .ZN(n8962) );
  INV_X1 U11314 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10531) );
  OR2_X1 U11315 ( .A1(n9451), .A2(n10531), .ZN(n8961) );
  NAND4_X1 U11316 ( .A1(n8964), .A2(n8963), .A3(n8962), .A4(n8961), .ZN(n13262) );
  INV_X1 U11317 ( .A(n13262), .ZN(n11439) );
  NAND2_X1 U11318 ( .A1(n11701), .A2(n11439), .ZN(n9231) );
  OR2_X1 U11319 ( .A1(n11701), .A2(n11439), .ZN(n8965) );
  NAND2_X1 U11320 ( .A1(n11481), .A2(n11480), .ZN(n8967) );
  NAND2_X1 U11321 ( .A1(n11701), .A2(n13262), .ZN(n8966) );
  NAND2_X1 U11322 ( .A1(n10509), .A2(n9468), .ZN(n8971) );
  INV_X1 U11323 ( .A(n8968), .ZN(n8981) );
  NAND2_X1 U11324 ( .A1(n8981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8969) );
  XNOR2_X1 U11325 ( .A(n8969), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U11326 ( .A1(n9097), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9096), 
        .B2(n10554), .ZN(n8970) );
  NAND2_X1 U11327 ( .A1(n9206), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8977) );
  INV_X1 U11328 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11618) );
  OR2_X1 U11329 ( .A1(n9453), .A2(n11618), .ZN(n8976) );
  NAND2_X1 U11330 ( .A1(n8972), .A2(n11438), .ZN(n8973) );
  NAND2_X1 U11331 ( .A1(n8987), .A2(n8973), .ZN(n11617) );
  OR2_X1 U11332 ( .A1(n6499), .A2(n11617), .ZN(n8975) );
  INV_X1 U11333 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10527) );
  OR2_X1 U11334 ( .A1(n9451), .A2(n10527), .ZN(n8974) );
  NAND4_X1 U11335 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n13261) );
  NAND2_X1 U11336 ( .A1(n11620), .A2(n11788), .ZN(n9232) );
  OR2_X1 U11337 ( .A1(n11620), .A2(n11788), .ZN(n8978) );
  INV_X1 U11338 ( .A(n11613), .ZN(n8979) );
  NAND2_X1 U11339 ( .A1(n11620), .A2(n13261), .ZN(n8980) );
  NAND2_X1 U11340 ( .A1(n10517), .A2(n9468), .ZN(n8984) );
  OAI21_X1 U11341 ( .B1(n8981), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8982) );
  XNOR2_X1 U11342 ( .A(n8982), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U11343 ( .A1(n9097), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9096), 
        .B2(n13323), .ZN(n8983) );
  NAND2_X1 U11344 ( .A1(n9206), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8993) );
  INV_X1 U11345 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8985) );
  OR2_X1 U11346 ( .A1(n9453), .A2(n8985), .ZN(n8992) );
  AND2_X1 U11347 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  OR2_X1 U11348 ( .A1(n8988), .A2(n9002), .ZN(n11669) );
  OR2_X1 U11349 ( .A1(n6499), .A2(n11669), .ZN(n8991) );
  INV_X1 U11350 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8989) );
  OR2_X1 U11351 ( .A1(n9451), .A2(n8989), .ZN(n8990) );
  NAND4_X1 U11352 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n13260) );
  AND2_X1 U11353 ( .A1(n11902), .A2(n13260), .ZN(n8994) );
  OR2_X1 U11354 ( .A1(n11902), .A2(n13260), .ZN(n8995) );
  NAND2_X1 U11355 ( .A1(n10561), .A2(n9468), .ZN(n9001) );
  NOR2_X1 U11356 ( .A1(n8998), .A2(n8741), .ZN(n8996) );
  MUX2_X1 U11357 ( .A(n8741), .B(n8996), .S(P2_IR_REG_12__SCAN_IN), .Z(n8999)
         );
  NAND2_X1 U11358 ( .A1(n8998), .A2(n8997), .ZN(n9012) );
  INV_X1 U11359 ( .A(n9012), .ZN(n9028) );
  AOI22_X1 U11360 ( .A1(n9097), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9096), 
        .B2(n14994), .ZN(n9000) );
  NAND2_X1 U11361 ( .A1(n8828), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9010) );
  INV_X1 U11362 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13316) );
  OR2_X1 U11363 ( .A1(n9453), .A2(n13316), .ZN(n9009) );
  INV_X1 U11364 ( .A(n9002), .ZN(n9004) );
  INV_X1 U11365 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11366 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  NAND2_X1 U11367 ( .A1(n9018), .A2(n9005), .ZN(n14933) );
  OR2_X1 U11368 ( .A1(n6499), .A2(n14933), .ZN(n9008) );
  INV_X1 U11369 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9006) );
  OR2_X1 U11370 ( .A1(n8904), .A2(n9006), .ZN(n9007) );
  NAND4_X1 U11371 ( .A1(n9010), .A2(n9009), .A3(n9008), .A4(n9007), .ZN(n13259) );
  NOR2_X1 U11372 ( .A1(n14931), .A2(n13259), .ZN(n9011) );
  OAI22_X2 U11373 ( .A1(n11919), .A2(n9011), .B1(n14676), .B2(n11787), .ZN(
        n11914) );
  NAND2_X1 U11374 ( .A1(n10792), .A2(n9468), .ZN(n9015) );
  NAND2_X1 U11375 ( .A1(n9012), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9013) );
  XNOR2_X1 U11376 ( .A(n9013), .B(P2_IR_REG_13__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U11377 ( .A1(n9097), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9096), 
        .B2(n13343), .ZN(n9014) );
  NAND2_X1 U11378 ( .A1(n9206), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9024) );
  INV_X1 U11379 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11911) );
  OR2_X1 U11380 ( .A1(n9453), .A2(n11911), .ZN(n9023) );
  INV_X1 U11381 ( .A(n9016), .ZN(n9034) );
  INV_X1 U11382 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U11383 ( .A1(n9018), .A2(n9017), .ZN(n9019) );
  NAND2_X1 U11384 ( .A1(n9034), .A2(n9019), .ZN(n12101) );
  OR2_X1 U11385 ( .A1(n6499), .A2(n12101), .ZN(n9022) );
  INV_X1 U11386 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9020) );
  OR2_X1 U11387 ( .A1(n9451), .A2(n9020), .ZN(n9021) );
  NAND4_X1 U11388 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n13258) );
  AND2_X1 U11389 ( .A1(n12115), .A2(n13258), .ZN(n9026) );
  OR2_X1 U11390 ( .A1(n12115), .A2(n13258), .ZN(n9025) );
  NAND2_X1 U11391 ( .A1(n10890), .A2(n9468), .ZN(n9032) );
  INV_X1 U11392 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9027) );
  AND2_X1 U11393 ( .A1(n9028), .A2(n9027), .ZN(n9043) );
  INV_X1 U11394 ( .A(n9043), .ZN(n9029) );
  NAND2_X1 U11395 ( .A1(n9029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U11396 ( .A(n9030), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U11397 ( .A1(n9097), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9096), 
        .B2(n13349), .ZN(n9031) );
  NAND2_X1 U11398 ( .A1(n9207), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9040) );
  INV_X1 U11399 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11400 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  NAND2_X1 U11401 ( .A1(n9059), .A2(n9035), .ZN(n14652) );
  OR2_X1 U11402 ( .A1(n6499), .A2(n14652), .ZN(n9039) );
  INV_X1 U11403 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13346) );
  OR2_X1 U11404 ( .A1(n9451), .A2(n13346), .ZN(n9038) );
  INV_X1 U11405 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9036) );
  OR2_X1 U11406 ( .A1(n8904), .A2(n9036), .ZN(n9037) );
  NAND4_X1 U11407 ( .A1(n9040), .A2(n9039), .A3(n9038), .A4(n9037), .ZN(n13257) );
  INV_X1 U11408 ( .A(n13257), .ZN(n13247) );
  XNOR2_X1 U11409 ( .A(n14656), .B(n13247), .ZN(n14648) );
  INV_X1 U11410 ( .A(n14648), .ZN(n14660) );
  NAND2_X1 U11411 ( .A1(n14656), .A2(n13257), .ZN(n9041) );
  NAND2_X1 U11412 ( .A1(n11172), .A2(n9468), .ZN(n9046) );
  INV_X1 U11413 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11414 ( .A1(n9043), .A2(n9042), .ZN(n9053) );
  NAND2_X1 U11415 ( .A1(n9053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9044) );
  XNOR2_X1 U11416 ( .A(n9044), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U11417 ( .A1(n9097), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9096), 
        .B2(n15016), .ZN(n9045) );
  NAND2_X1 U11418 ( .A1(n9206), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9051) );
  INV_X1 U11419 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9047) );
  OR2_X1 U11420 ( .A1(n9453), .A2(n9047), .ZN(n9050) );
  INV_X1 U11421 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9058) );
  XNOR2_X1 U11422 ( .A(n9059), .B(n9058), .ZN(n13633) );
  OR2_X1 U11423 ( .A1(n6499), .A2(n13633), .ZN(n9049) );
  INV_X1 U11424 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15011) );
  OR2_X1 U11425 ( .A1(n9451), .A2(n15011), .ZN(n9048) );
  NAND4_X1 U11426 ( .A1(n9051), .A2(n9050), .A3(n9049), .A4(n9048), .ZN(n13613) );
  INV_X1 U11427 ( .A(n13613), .ZN(n14637) );
  XNOR2_X1 U11428 ( .A(n13721), .B(n14637), .ZN(n9518) );
  OR2_X1 U11429 ( .A1(n13721), .A2(n13613), .ZN(n9052) );
  NAND2_X1 U11430 ( .A1(n11256), .A2(n9468), .ZN(n9056) );
  NAND2_X1 U11431 ( .A1(n9068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9054) );
  XNOR2_X1 U11432 ( .A(n9054), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U11433 ( .A1(n9097), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9096), 
        .B2(n13368), .ZN(n9055) );
  NAND2_X1 U11434 ( .A1(n9207), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9066) );
  INV_X1 U11435 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9057) );
  OAI21_X1 U11436 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9060) );
  NAND2_X1 U11437 ( .A1(n9060), .A2(n9075), .ZN(n14647) );
  OR2_X1 U11438 ( .A1(n6499), .A2(n14647), .ZN(n9065) );
  INV_X1 U11439 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9061) );
  OR2_X1 U11440 ( .A1(n9451), .A2(n9061), .ZN(n9064) );
  INV_X1 U11441 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9062) );
  OR2_X1 U11442 ( .A1(n8904), .A2(n9062), .ZN(n9063) );
  NAND4_X1 U11443 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n13256) );
  INV_X1 U11444 ( .A(n13256), .ZN(n13246) );
  XNOR2_X1 U11445 ( .A(n14644), .B(n13246), .ZN(n13618) );
  NAND2_X1 U11446 ( .A1(n14644), .A2(n13256), .ZN(n9067) );
  NAND2_X1 U11447 ( .A1(n13617), .A2(n9067), .ZN(n13600) );
  NAND2_X1 U11448 ( .A1(n11355), .A2(n9468), .ZN(n9073) );
  OAI21_X1 U11449 ( .B1(n9068), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9070) );
  INV_X1 U11450 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U11451 ( .A1(n9070), .A2(n9069), .ZN(n9082) );
  OR2_X1 U11452 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  AND2_X1 U11453 ( .A1(n9082), .A2(n9071), .ZN(n15026) );
  AOI22_X1 U11454 ( .A1(n9097), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9096), 
        .B2(n15026), .ZN(n9072) );
  NAND2_X1 U11455 ( .A1(n9206), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9080) );
  INV_X1 U11456 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9074) );
  OR2_X1 U11457 ( .A1(n9453), .A2(n9074), .ZN(n9079) );
  INV_X1 U11458 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15024) );
  NAND2_X1 U11459 ( .A1(n9075), .A2(n15024), .ZN(n9076) );
  NAND2_X1 U11460 ( .A1(n9087), .A2(n9076), .ZN(n13603) );
  OR2_X1 U11461 ( .A1(n6499), .A2(n13603), .ZN(n9078) );
  INV_X1 U11462 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13371) );
  OR2_X1 U11463 ( .A1(n9451), .A2(n13371), .ZN(n9077) );
  NAND4_X1 U11464 ( .A1(n9080), .A2(n9079), .A3(n9078), .A4(n9077), .ZN(n13615) );
  INV_X1 U11465 ( .A(n13615), .ZN(n14636) );
  XNOR2_X1 U11466 ( .A(n13712), .B(n14636), .ZN(n13599) );
  NAND2_X1 U11467 ( .A1(n13712), .A2(n13615), .ZN(n9081) );
  NAND2_X1 U11468 ( .A1(n9082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  XNOR2_X1 U11469 ( .A(n9083), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U11470 ( .A1(n9096), .A2(n13365), .B1(n9097), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11471 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U11472 ( .A1(n9101), .A2(n9088), .ZN(n13583) );
  INV_X1 U11473 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15044) );
  OR2_X1 U11474 ( .A1(n9451), .A2(n15044), .ZN(n9089) );
  OAI21_X1 U11475 ( .B1(n13583), .B2(n6499), .A(n9089), .ZN(n9094) );
  INV_X1 U11476 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9092) );
  INV_X1 U11477 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9090) );
  OR2_X1 U11478 ( .A1(n9453), .A2(n9090), .ZN(n9091) );
  OAI21_X1 U11479 ( .B1(n8904), .B2(n9092), .A(n9091), .ZN(n9093) );
  INV_X1 U11480 ( .A(n13564), .ZN(n9242) );
  XNOR2_X1 U11481 ( .A(n13707), .B(n9242), .ZN(n13577) );
  INV_X1 U11482 ( .A(n13577), .ZN(n13589) );
  OR2_X1 U11483 ( .A1(n13707), .A2(n13564), .ZN(n9095) );
  NAND2_X1 U11484 ( .A1(n11745), .A2(n9468), .ZN(n9099) );
  AOI22_X1 U11485 ( .A1(n9097), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11210), 
        .B2(n9096), .ZN(n9098) );
  INV_X1 U11486 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9105) );
  INV_X1 U11487 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11488 ( .A1(n9101), .A2(n9100), .ZN(n9102) );
  NAND2_X1 U11489 ( .A1(n9110), .A2(n9102), .ZN(n13568) );
  OR2_X1 U11490 ( .A1(n13568), .A2(n6499), .ZN(n9104) );
  AOI22_X1 U11491 ( .A1(n9206), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n9207), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n9103) );
  OAI211_X1 U11492 ( .C1(n9451), .C2(n9105), .A(n9104), .B(n9103), .ZN(n13579)
         );
  NOR2_X1 U11493 ( .A1(n13702), .A2(n13579), .ZN(n9106) );
  INV_X1 U11494 ( .A(n13702), .ZN(n13571) );
  INV_X1 U11495 ( .A(n13579), .ZN(n9244) );
  OR2_X1 U11496 ( .A1(n11747), .A2(n9140), .ZN(n9108) );
  NAND2_X1 U11497 ( .A1(n9097), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U11498 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  AND2_X1 U11499 ( .A1(n9118), .A2(n9111), .ZN(n13552) );
  NAND2_X1 U11500 ( .A1(n13552), .A2(n9183), .ZN(n9114) );
  AOI22_X1 U11501 ( .A1(n9206), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n9207), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U11502 ( .A1(n8828), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9112) );
  OR2_X1 U11503 ( .A1(n12588), .A2(n9140), .ZN(n9116) );
  NAND2_X1 U11504 ( .A1(n9097), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9115) );
  INV_X1 U11505 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11506 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  NAND2_X1 U11507 ( .A1(n9132), .A2(n9119), .ZN(n13165) );
  OR2_X1 U11508 ( .A1(n13165), .A2(n6499), .ZN(n9124) );
  INV_X1 U11509 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13693) );
  NAND2_X1 U11510 ( .A1(n9206), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U11511 ( .A1(n9207), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9120) );
  OAI211_X1 U11512 ( .C1(n13693), .C2(n9451), .A(n9121), .B(n9120), .ZN(n9122)
         );
  INV_X1 U11513 ( .A(n9122), .ZN(n9123) );
  NAND2_X1 U11514 ( .A1(n9124), .A2(n9123), .ZN(n13558) );
  XNOR2_X1 U11515 ( .A(n13541), .B(n13558), .ZN(n13534) );
  INV_X1 U11516 ( .A(n13558), .ZN(n13514) );
  NAND2_X1 U11517 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U11518 ( .A1(n9129), .A2(n9128), .ZN(n12136) );
  NAND2_X1 U11519 ( .A1(n9097), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U11520 ( .A(n9132), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n13522) );
  NAND2_X1 U11521 ( .A1(n13522), .A2(n9183), .ZN(n9138) );
  INV_X1 U11522 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U11523 ( .A1(n9206), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U11524 ( .A1(n9207), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9133) );
  OAI211_X1 U11525 ( .C1(n9135), .C2(n9451), .A(n9134), .B(n9133), .ZN(n9136)
         );
  INV_X1 U11526 ( .A(n9136), .ZN(n9137) );
  XNOR2_X1 U11527 ( .A(n13748), .B(n13168), .ZN(n13511) );
  INV_X1 U11528 ( .A(n13511), .ZN(n13518) );
  NAND2_X1 U11529 ( .A1(n13748), .A2(n13168), .ZN(n9139) );
  NAND2_X1 U11530 ( .A1(n9097), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9141) );
  INV_X1 U11531 ( .A(n9145), .ZN(n9143) );
  NAND2_X1 U11532 ( .A1(n9143), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9159) );
  INV_X1 U11533 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11534 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  NAND2_X1 U11535 ( .A1(n9159), .A2(n9146), .ZN(n13196) );
  OR2_X1 U11536 ( .A1(n13196), .A2(n6499), .ZN(n9152) );
  INV_X1 U11537 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11538 ( .A1(n9206), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11539 ( .A1(n9207), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9147) );
  OAI211_X1 U11540 ( .C1(n9149), .C2(n9451), .A(n9148), .B(n9147), .ZN(n9150)
         );
  INV_X1 U11541 ( .A(n9150), .ZN(n9151) );
  INV_X1 U11542 ( .A(n13460), .ZN(n13255) );
  NAND2_X1 U11543 ( .A1(n13490), .A2(n13255), .ZN(n9153) );
  NAND2_X1 U11544 ( .A1(n13671), .A2(n13255), .ZN(n9154) );
  AND2_X2 U11545 ( .A1(n13475), .A2(n9154), .ZN(n13466) );
  NAND2_X1 U11546 ( .A1(n13779), .A2(n9468), .ZN(n9156) );
  NAND2_X1 U11547 ( .A1(n9097), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9155) );
  INV_X1 U11548 ( .A(n9159), .ZN(n9157) );
  NAND2_X1 U11549 ( .A1(n9157), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9171) );
  INV_X1 U11550 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U11551 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  NAND2_X1 U11552 ( .A1(n9171), .A2(n9160), .ZN(n13174) );
  OR2_X1 U11553 ( .A1(n13174), .A2(n6499), .ZN(n9166) );
  INV_X1 U11554 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11555 ( .A1(n9206), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11556 ( .A1(n9207), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9161) );
  OAI211_X1 U11557 ( .C1(n9163), .C2(n9451), .A(n9162), .B(n9161), .ZN(n9164)
         );
  INV_X1 U11558 ( .A(n9164), .ZN(n9165) );
  NAND2_X1 U11559 ( .A1(n9166), .A2(n9165), .ZN(n13481) );
  INV_X1 U11560 ( .A(n13458), .ZN(n13465) );
  OR2_X1 U11561 ( .A1(n13739), .A2(n13481), .ZN(n9167) );
  NAND2_X1 U11562 ( .A1(n13776), .A2(n9468), .ZN(n9169) );
  NAND2_X1 U11563 ( .A1(n9097), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9168) );
  INV_X1 U11564 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U11565 ( .A1(n9171), .A2(n9170), .ZN(n9172) );
  NAND2_X1 U11566 ( .A1(n13449), .A2(n9183), .ZN(n9178) );
  INV_X1 U11567 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U11568 ( .A1(n9206), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11569 ( .A1(n9207), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9173) );
  OAI211_X1 U11570 ( .C1(n9175), .C2(n9451), .A(n9174), .B(n9173), .ZN(n9176)
         );
  INV_X1 U11571 ( .A(n9176), .ZN(n9177) );
  OR2_X1 U11572 ( .A1(n13451), .A2(n13461), .ZN(n9179) );
  NAND2_X1 U11573 ( .A1(n13451), .A2(n13461), .ZN(n9180) );
  NAND2_X1 U11574 ( .A1(n9097), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9181) );
  NAND2_X2 U11575 ( .A1(n9182), .A2(n9181), .ZN(n13656) );
  XNOR2_X1 U11576 ( .A(n9196), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U11577 ( .A1(n13430), .A2(n9183), .ZN(n9189) );
  INV_X1 U11578 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U11579 ( .A1(n9206), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11580 ( .A1(n9207), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9184) );
  OAI211_X1 U11581 ( .C1(n9186), .C2(n9451), .A(n9185), .B(n9184), .ZN(n9187)
         );
  INV_X1 U11582 ( .A(n9187), .ZN(n9188) );
  NAND2_X1 U11583 ( .A1(n9189), .A2(n9188), .ZN(n13441) );
  NAND2_X1 U11584 ( .A1(n13656), .A2(n13441), .ZN(n9191) );
  NAND2_X1 U11585 ( .A1(n12425), .A2(n9468), .ZN(n9193) );
  NAND2_X1 U11586 ( .A1(n9097), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9192) );
  NAND2_X2 U11587 ( .A1(n9193), .A2(n9192), .ZN(n13733) );
  INV_X1 U11588 ( .A(n9196), .ZN(n9195) );
  AND2_X1 U11589 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9194) );
  NAND2_X1 U11590 ( .A1(n9195), .A2(n9194), .ZN(n13399) );
  INV_X1 U11591 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13135) );
  INV_X1 U11592 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12572) );
  OAI21_X1 U11593 ( .B1(n9196), .B2(n13135), .A(n12572), .ZN(n9197) );
  NAND2_X1 U11594 ( .A1(n13399), .A2(n9197), .ZN(n13420) );
  OR2_X1 U11595 ( .A1(n13420), .A2(n6499), .ZN(n9203) );
  INV_X1 U11596 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U11597 ( .A1(n9206), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U11598 ( .A1(n9207), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9198) );
  OAI211_X1 U11599 ( .C1(n9200), .C2(n9451), .A(n9199), .B(n9198), .ZN(n9201)
         );
  INV_X1 U11600 ( .A(n9201), .ZN(n9202) );
  NAND2_X1 U11601 ( .A1(n9203), .A2(n9202), .ZN(n13427) );
  NAND2_X1 U11602 ( .A1(n13733), .A2(n13427), .ZN(n9205) );
  NAND2_X1 U11603 ( .A1(n9205), .A2(n9204), .ZN(n13408) );
  OR2_X1 U11604 ( .A1(n13399), .A2(n6499), .ZN(n9213) );
  INV_X1 U11605 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9210) );
  NAND2_X1 U11606 ( .A1(n9206), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U11607 ( .A1(n9207), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9208) );
  OAI211_X1 U11608 ( .C1(n9210), .C2(n9451), .A(n9209), .B(n9208), .ZN(n9211)
         );
  INV_X1 U11609 ( .A(n9211), .ZN(n9212) );
  NAND2_X1 U11610 ( .A1(n9213), .A2(n9212), .ZN(n13254) );
  XNOR2_X1 U11611 ( .A(n13401), .B(n13254), .ZN(n9525) );
  INV_X1 U11612 ( .A(n9525), .ZN(n9214) );
  AND2_X2 U11613 ( .A1(n9216), .A2(n9215), .ZN(n9275) );
  XNOR2_X1 U11614 ( .A(n9275), .B(n9217), .ZN(n9218) );
  NAND2_X1 U11615 ( .A1(n8803), .A2(n11210), .ZN(n9220) );
  NAND2_X1 U11616 ( .A1(n9509), .A2(n11279), .ZN(n11278) );
  OR2_X1 U11617 ( .A1(n13269), .A2(n8834), .ZN(n9222) );
  INV_X1 U11618 ( .A(n6477), .ZN(n10641) );
  OR2_X1 U11619 ( .A1(n10668), .A2(n10641), .ZN(n9223) );
  NAND2_X1 U11620 ( .A1(n9224), .A2(n9223), .ZN(n11221) );
  NAND2_X1 U11621 ( .A1(n11221), .A2(n11225), .ZN(n9226) );
  OR2_X1 U11622 ( .A1(n6921), .A2(n13268), .ZN(n9225) );
  INV_X1 U11623 ( .A(n11268), .ZN(n15118) );
  OR2_X1 U11624 ( .A1(n13267), .A2(n15118), .ZN(n9227) );
  XNOR2_X1 U11625 ( .A(n13266), .B(n11306), .ZN(n11298) );
  INV_X1 U11626 ( .A(n13266), .ZN(n10703) );
  INV_X1 U11627 ( .A(n13265), .ZN(n10825) );
  NAND2_X1 U11628 ( .A1(n11183), .A2(n10825), .ZN(n9228) );
  AND2_X1 U11629 ( .A1(n11332), .A2(n9325), .ZN(n9229) );
  NAND2_X1 U11630 ( .A1(n11384), .A2(n9230), .ZN(n11483) );
  NAND2_X1 U11631 ( .A1(n11483), .A2(n11484), .ZN(n11482) );
  NAND2_X1 U11632 ( .A1(n11482), .A2(n9231), .ZN(n11609) );
  XNOR2_X1 U11633 ( .A(n11902), .B(n13260), .ZN(n11785) );
  INV_X1 U11634 ( .A(n13260), .ZN(n14922) );
  OR2_X1 U11635 ( .A1(n14931), .A2(n11787), .ZN(n9233) );
  NAND2_X1 U11636 ( .A1(n14931), .A2(n11787), .ZN(n9234) );
  INV_X1 U11637 ( .A(n13258), .ZN(n14919) );
  NAND2_X1 U11638 ( .A1(n12115), .A2(n14919), .ZN(n9507) );
  OR2_X1 U11639 ( .A1(n12115), .A2(n14919), .ZN(n9508) );
  NOR2_X1 U11640 ( .A1(n14656), .A2(n13247), .ZN(n9235) );
  NAND2_X1 U11641 ( .A1(n14656), .A2(n13247), .ZN(n9236) );
  AND2_X1 U11642 ( .A1(n13721), .A2(n14637), .ZN(n9237) );
  OR2_X1 U11643 ( .A1(n13721), .A2(n14637), .ZN(n9238) );
  NOR2_X1 U11644 ( .A1(n14644), .A2(n13246), .ZN(n9239) );
  INV_X1 U11645 ( .A(n14644), .ZN(n13625) );
  OR2_X1 U11646 ( .A1(n13712), .A2(n14636), .ZN(n9240) );
  NAND2_X1 U11647 ( .A1(n13707), .A2(n9242), .ZN(n9241) );
  OR2_X1 U11648 ( .A1(n13707), .A2(n9242), .ZN(n9243) );
  NOR2_X1 U11649 ( .A1(n13702), .A2(n9244), .ZN(n13530) );
  NAND2_X1 U11650 ( .A1(n13702), .A2(n9244), .ZN(n13531) );
  NAND2_X1 U11651 ( .A1(n13697), .A2(n13538), .ZN(n13532) );
  OR2_X1 U11652 ( .A1(n13697), .A2(n13538), .ZN(n9506) );
  NAND2_X1 U11653 ( .A1(n13755), .A2(n13558), .ZN(n9245) );
  NAND3_X1 U11654 ( .A1(n9246), .A2(n9506), .A3(n9245), .ZN(n9248) );
  NAND2_X1 U11655 ( .A1(n13541), .A2(n13514), .ZN(n9247) );
  NAND2_X1 U11656 ( .A1(n9248), .A2(n9247), .ZN(n13510) );
  NAND2_X1 U11657 ( .A1(n13510), .A2(n13511), .ZN(n9250) );
  NAND2_X1 U11658 ( .A1(n13748), .A2(n13536), .ZN(n9249) );
  OR2_X1 U11659 ( .A1(n13505), .A2(n13483), .ZN(n9251) );
  NAND2_X1 U11660 ( .A1(n13459), .A2(n13458), .ZN(n13457) );
  INV_X1 U11661 ( .A(n13481), .ZN(n13443) );
  NAND2_X1 U11662 ( .A1(n13739), .A2(n13443), .ZN(n9253) );
  NAND2_X1 U11663 ( .A1(n13457), .A2(n9253), .ZN(n13440) );
  OR2_X1 U11664 ( .A1(n13661), .A2(n13461), .ZN(n9505) );
  NAND2_X1 U11665 ( .A1(n13661), .A2(n13461), .ZN(n9504) );
  INV_X1 U11666 ( .A(n13441), .ZN(n13234) );
  AND2_X1 U11667 ( .A1(n13656), .A2(n13234), .ZN(n9254) );
  INV_X1 U11668 ( .A(n13427), .ZN(n13138) );
  NAND2_X1 U11669 ( .A1(n9217), .A2(n11210), .ZN(n9473) );
  NAND2_X1 U11670 ( .A1(n9529), .A2(n9512), .ZN(n9256) );
  INV_X1 U11671 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13650) );
  OR2_X1 U11672 ( .A1(n9451), .A2(n13650), .ZN(n9261) );
  INV_X1 U11673 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13393) );
  OR2_X1 U11674 ( .A1(n9453), .A2(n13393), .ZN(n9260) );
  INV_X1 U11675 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13730) );
  OR2_X1 U11676 ( .A1(n8904), .A2(n13730), .ZN(n9259) );
  AND3_X1 U11677 ( .A1(n9261), .A2(n9260), .A3(n9259), .ZN(n9472) );
  INV_X1 U11678 ( .A(n10677), .ZN(n9262) );
  INV_X1 U11679 ( .A(n13774), .ZN(n10474) );
  NAND2_X1 U11680 ( .A1(n10474), .A2(P2_B_REG_SCAN_IN), .ZN(n9264) );
  NAND2_X1 U11681 ( .A1(n13614), .A2(n9264), .ZN(n13386) );
  NOR2_X1 U11682 ( .A1(n9472), .A2(n13386), .ZN(n9265) );
  AOI21_X1 U11683 ( .B1(n13427), .B2(n13612), .A(n9265), .ZN(n9266) );
  NAND2_X1 U11684 ( .A1(n11275), .A2(n10641), .ZN(n11228) );
  INV_X1 U11685 ( .A(n11306), .ZN(n15127) );
  INV_X1 U11686 ( .A(n11183), .ZN(n11291) );
  OR2_X2 U11687 ( .A1(n11313), .A2(n11396), .ZN(n11488) );
  INV_X1 U11688 ( .A(n11620), .ZN(n15141) );
  INV_X1 U11689 ( .A(n11902), .ZN(n11899) );
  NAND2_X1 U11690 ( .A1(n13625), .A2(n13632), .ZN(n13621) );
  NAND2_X1 U11691 ( .A1(n13521), .A2(n13540), .ZN(n13520) );
  NAND2_X1 U11692 ( .A1(n9255), .A2(n13429), .ZN(n13417) );
  NOR2_X2 U11693 ( .A1(n13417), .A2(n13401), .ZN(n13392) );
  NAND2_X1 U11694 ( .A1(n13417), .A2(n13401), .ZN(n9270) );
  NAND3_X1 U11695 ( .A1(n9271), .A2(n6483), .A3(n9270), .ZN(n13404) );
  MUX2_X1 U11696 ( .A(n10715), .B(n9275), .S(n11276), .Z(n9278) );
  AND2_X1 U11697 ( .A1(n13270), .A2(n6502), .ZN(n9279) );
  OAI21_X1 U11698 ( .B1(n9217), .B2(n13379), .A(n9275), .ZN(n9277) );
  OAI21_X1 U11699 ( .B1(n9278), .B2(n9279), .A(n9277), .ZN(n9281) );
  INV_X1 U11700 ( .A(n11276), .ZN(n9510) );
  NAND2_X1 U11701 ( .A1(n9279), .A2(n9510), .ZN(n9280) );
  NAND2_X1 U11702 ( .A1(n9281), .A2(n9280), .ZN(n9289) );
  NAND2_X1 U11703 ( .A1(n13269), .A2(n6502), .ZN(n9283) );
  NAND2_X1 U11704 ( .A1(n10663), .A2(n9477), .ZN(n9282) );
  NAND2_X1 U11705 ( .A1(n9283), .A2(n9282), .ZN(n9288) );
  AOI22_X1 U11706 ( .A1(n13269), .A2(n9471), .B1(n10663), .B2(n6502), .ZN(
        n9284) );
  AOI21_X1 U11707 ( .B1(n9289), .B2(n9288), .A(n9284), .ZN(n9295) );
  AND2_X1 U11708 ( .A1(n6477), .A2(n6502), .ZN(n9285) );
  NAND2_X1 U11709 ( .A1(n10668), .A2(n6502), .ZN(n9287) );
  NAND2_X1 U11710 ( .A1(n6477), .A2(n9477), .ZN(n9286) );
  AOI22_X1 U11711 ( .A1(n13268), .A2(n9477), .B1(n11231), .B2(n6502), .ZN(
        n9297) );
  NAND2_X1 U11712 ( .A1(n13268), .A2(n6502), .ZN(n9291) );
  NAND2_X1 U11713 ( .A1(n11231), .A2(n9477), .ZN(n9290) );
  NAND2_X1 U11714 ( .A1(n9291), .A2(n9290), .ZN(n9296) );
  OAI21_X1 U11715 ( .B1(n9295), .B2(n9294), .A(n9293), .ZN(n9301) );
  INV_X1 U11716 ( .A(n9296), .ZN(n9299) );
  INV_X1 U11717 ( .A(n9297), .ZN(n9298) );
  NAND2_X1 U11718 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  NAND2_X1 U11719 ( .A1(n9301), .A2(n9300), .ZN(n9307) );
  NAND2_X1 U11720 ( .A1(n13267), .A2(n9477), .ZN(n9303) );
  NAND2_X1 U11721 ( .A1(n11268), .A2(n6502), .ZN(n9302) );
  NAND2_X1 U11722 ( .A1(n9303), .A2(n9302), .ZN(n9308) );
  NAND2_X1 U11723 ( .A1(n13267), .A2(n6502), .ZN(n9305) );
  NAND2_X1 U11724 ( .A1(n11268), .A2(n9477), .ZN(n9304) );
  NAND2_X1 U11725 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  INV_X1 U11726 ( .A(n9308), .ZN(n9309) );
  NAND2_X1 U11727 ( .A1(n11306), .A2(n9477), .ZN(n9311) );
  NAND2_X1 U11728 ( .A1(n13266), .A2(n6502), .ZN(n9310) );
  NAND2_X1 U11729 ( .A1(n9311), .A2(n9310), .ZN(n9313) );
  AOI22_X1 U11730 ( .A1(n11306), .A2(n6502), .B1(n13266), .B2(n9477), .ZN(
        n9312) );
  NOR2_X1 U11731 ( .A1(n9314), .A2(n9313), .ZN(n9315) );
  OR2_X1 U11732 ( .A1(n9316), .A2(n9315), .ZN(n9321) );
  NAND2_X1 U11733 ( .A1(n11183), .A2(n6502), .ZN(n9318) );
  NAND2_X1 U11734 ( .A1(n13265), .A2(n9477), .ZN(n9317) );
  NAND2_X1 U11735 ( .A1(n9318), .A2(n9317), .ZN(n9320) );
  AOI22_X1 U11736 ( .A1(n11183), .A2(n9471), .B1(n13265), .B2(n6502), .ZN(
        n9319) );
  NAND2_X1 U11737 ( .A1(n11332), .A2(n9471), .ZN(n9323) );
  NAND2_X1 U11738 ( .A1(n13264), .A2(n6502), .ZN(n9322) );
  NAND2_X1 U11739 ( .A1(n9323), .A2(n9322), .ZN(n9329) );
  NAND2_X1 U11740 ( .A1(n11332), .A2(n6502), .ZN(n9324) );
  OAI21_X1 U11741 ( .B1(n9325), .B2(n6502), .A(n9324), .ZN(n9326) );
  NAND2_X1 U11742 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  OAI21_X1 U11743 ( .B1(n9330), .B2(n9329), .A(n9328), .ZN(n9335) );
  NAND2_X1 U11744 ( .A1(n11396), .A2(n6502), .ZN(n9332) );
  NAND2_X1 U11745 ( .A1(n13263), .A2(n9477), .ZN(n9331) );
  NAND2_X1 U11746 ( .A1(n9332), .A2(n9331), .ZN(n9334) );
  AOI22_X1 U11747 ( .A1(n11396), .A2(n9471), .B1(n13263), .B2(n6502), .ZN(
        n9333) );
  INV_X1 U11748 ( .A(n9341), .ZN(n9339) );
  NAND2_X1 U11749 ( .A1(n11701), .A2(n9471), .ZN(n9337) );
  NAND2_X1 U11750 ( .A1(n13262), .A2(n6502), .ZN(n9336) );
  NAND2_X1 U11751 ( .A1(n9337), .A2(n9336), .ZN(n9340) );
  INV_X1 U11752 ( .A(n9340), .ZN(n9338) );
  NAND2_X1 U11753 ( .A1(n9339), .A2(n9338), .ZN(n9346) );
  NAND2_X1 U11754 ( .A1(n11701), .A2(n6502), .ZN(n9342) );
  OAI21_X1 U11755 ( .B1(n11439), .B2(n6502), .A(n9342), .ZN(n9343) );
  NAND2_X1 U11756 ( .A1(n9344), .A2(n9343), .ZN(n9345) );
  NAND2_X1 U11757 ( .A1(n11620), .A2(n6502), .ZN(n9348) );
  NAND2_X1 U11758 ( .A1(n13261), .A2(n9471), .ZN(n9347) );
  AOI22_X1 U11759 ( .A1(n11620), .A2(n9471), .B1(n13261), .B2(n6502), .ZN(
        n9349) );
  NAND2_X1 U11760 ( .A1(n11902), .A2(n9477), .ZN(n9351) );
  NAND2_X1 U11761 ( .A1(n13260), .A2(n6502), .ZN(n9350) );
  NAND2_X1 U11762 ( .A1(n9351), .A2(n9350), .ZN(n9356) );
  NAND2_X1 U11763 ( .A1(n9355), .A2(n9356), .ZN(n9354) );
  NAND2_X1 U11764 ( .A1(n11902), .A2(n6502), .ZN(n9352) );
  OAI21_X1 U11765 ( .B1(n14922), .B2(n6502), .A(n9352), .ZN(n9353) );
  NAND2_X1 U11766 ( .A1(n9354), .A2(n9353), .ZN(n9360) );
  INV_X1 U11767 ( .A(n9355), .ZN(n9358) );
  NAND2_X1 U11768 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  NAND2_X1 U11769 ( .A1(n9360), .A2(n9359), .ZN(n9365) );
  NAND2_X1 U11770 ( .A1(n14931), .A2(n6502), .ZN(n9362) );
  NAND2_X1 U11771 ( .A1(n13259), .A2(n9471), .ZN(n9361) );
  NAND2_X1 U11772 ( .A1(n9362), .A2(n9361), .ZN(n9364) );
  AOI22_X1 U11773 ( .A1(n14931), .A2(n9471), .B1(n13259), .B2(n6502), .ZN(
        n9363) );
  AOI21_X1 U11774 ( .B1(n9365), .B2(n9364), .A(n9363), .ZN(n9367) );
  NOR2_X1 U11775 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  OR2_X1 U11776 ( .A1(n9367), .A2(n9366), .ZN(n9375) );
  NAND2_X1 U11777 ( .A1(n12115), .A2(n9471), .ZN(n9369) );
  NAND2_X1 U11778 ( .A1(n13258), .A2(n6502), .ZN(n9368) );
  NAND2_X1 U11779 ( .A1(n9369), .A2(n9368), .ZN(n9374) );
  NAND2_X1 U11780 ( .A1(n9375), .A2(n9374), .ZN(n9372) );
  NAND2_X1 U11781 ( .A1(n12115), .A2(n6502), .ZN(n9370) );
  OAI21_X1 U11782 ( .B1(n14919), .B2(n6502), .A(n9370), .ZN(n9371) );
  NAND2_X1 U11783 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  NAND2_X1 U11784 ( .A1(n14656), .A2(n6502), .ZN(n9377) );
  NAND2_X1 U11785 ( .A1(n13257), .A2(n9471), .ZN(n9376) );
  NAND2_X1 U11786 ( .A1(n9377), .A2(n9376), .ZN(n9391) );
  AOI22_X1 U11787 ( .A1(n13712), .A2(n6502), .B1(n9471), .B2(n13615), .ZN(
        n9380) );
  NAND2_X1 U11788 ( .A1(n13712), .A2(n9471), .ZN(n9379) );
  NAND2_X1 U11789 ( .A1(n13615), .A2(n6502), .ZN(n9378) );
  NAND2_X1 U11790 ( .A1(n9379), .A2(n9378), .ZN(n9397) );
  NAND2_X1 U11791 ( .A1(n9380), .A2(n9397), .ZN(n9385) );
  AND2_X1 U11792 ( .A1(n13256), .A2(n9471), .ZN(n9381) );
  AOI21_X1 U11793 ( .B1(n14644), .B2(n6502), .A(n9381), .ZN(n9395) );
  NAND2_X1 U11794 ( .A1(n14644), .A2(n9471), .ZN(n9383) );
  NAND2_X1 U11795 ( .A1(n13256), .A2(n6502), .ZN(n9382) );
  NAND2_X1 U11796 ( .A1(n9383), .A2(n9382), .ZN(n9394) );
  NAND2_X1 U11797 ( .A1(n9395), .A2(n9394), .ZN(n9384) );
  AND2_X1 U11798 ( .A1(n9385), .A2(n9384), .ZN(n9400) );
  AND2_X1 U11799 ( .A1(n13613), .A2(n9471), .ZN(n9386) );
  AOI21_X1 U11800 ( .B1(n13721), .B2(n6502), .A(n9386), .ZN(n9393) );
  NAND2_X1 U11801 ( .A1(n13721), .A2(n9471), .ZN(n9388) );
  NAND2_X1 U11802 ( .A1(n13613), .A2(n6502), .ZN(n9387) );
  NAND2_X1 U11803 ( .A1(n9388), .A2(n9387), .ZN(n9392) );
  NAND2_X1 U11804 ( .A1(n9393), .A2(n9392), .ZN(n9389) );
  AOI22_X1 U11805 ( .A1(n14656), .A2(n9471), .B1(n13257), .B2(n6502), .ZN(
        n9390) );
  OAI22_X1 U11806 ( .A1(n9395), .A2(n9394), .B1(n9393), .B2(n9392), .ZN(n9399)
         );
  NOR2_X1 U11807 ( .A1(n13712), .A2(n13615), .ZN(n9396) );
  NOR2_X1 U11808 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  AOI21_X1 U11809 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9401) );
  NAND2_X1 U11810 ( .A1(n9402), .A2(n9401), .ZN(n9407) );
  NAND2_X1 U11811 ( .A1(n13707), .A2(n6502), .ZN(n9404) );
  NAND2_X1 U11812 ( .A1(n13564), .A2(n9471), .ZN(n9403) );
  NAND2_X1 U11813 ( .A1(n9404), .A2(n9403), .ZN(n9406) );
  AOI22_X1 U11814 ( .A1(n13707), .A2(n9471), .B1(n13564), .B2(n6502), .ZN(
        n9405) );
  NAND2_X1 U11815 ( .A1(n13702), .A2(n9471), .ZN(n9409) );
  NAND2_X1 U11816 ( .A1(n13579), .A2(n6502), .ZN(n9408) );
  NAND2_X1 U11817 ( .A1(n9409), .A2(n9408), .ZN(n9414) );
  AOI22_X1 U11818 ( .A1(n13702), .A2(n6502), .B1(n9471), .B2(n13579), .ZN(
        n9410) );
  NAND2_X1 U11819 ( .A1(n9412), .A2(n9411), .ZN(n9418) );
  INV_X1 U11820 ( .A(n9413), .ZN(n9416) );
  INV_X1 U11821 ( .A(n9414), .ZN(n9415) );
  NAND2_X1 U11822 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  NAND2_X1 U11823 ( .A1(n9418), .A2(n9417), .ZN(n9421) );
  OAI22_X1 U11824 ( .A1(n13554), .A2(n9471), .B1(n13538), .B2(n6502), .ZN(
        n9420) );
  INV_X1 U11825 ( .A(n13538), .ZN(n13565) );
  AOI22_X1 U11826 ( .A1(n13697), .A2(n9471), .B1(n13565), .B2(n6502), .ZN(
        n9419) );
  AOI22_X1 U11827 ( .A1(n13541), .A2(n9471), .B1(n13558), .B2(n6502), .ZN(
        n9424) );
  AOI22_X1 U11828 ( .A1(n13541), .A2(n6502), .B1(n9477), .B2(n13558), .ZN(
        n9422) );
  INV_X1 U11829 ( .A(n9422), .ZN(n9423) );
  OAI22_X1 U11830 ( .A1(n13521), .A2(n9477), .B1(n13536), .B2(n6502), .ZN(
        n9426) );
  AOI22_X1 U11831 ( .A1(n13748), .A2(n9471), .B1(n13168), .B2(n6502), .ZN(
        n9425) );
  AOI21_X1 U11832 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(n9428) );
  AOI22_X1 U11833 ( .A1(n13505), .A2(n9471), .B1(n13512), .B2(n6502), .ZN(
        n9430) );
  AOI22_X1 U11834 ( .A1(n13505), .A2(n6502), .B1(n9471), .B2(n13512), .ZN(
        n9432) );
  OAI22_X1 U11835 ( .A1(n13490), .A2(n9477), .B1(n13460), .B2(n6502), .ZN(
        n9433) );
  OAI22_X1 U11836 ( .A1(n13490), .A2(n6502), .B1(n13460), .B2(n9471), .ZN(
        n9434) );
  INV_X1 U11837 ( .A(n9437), .ZN(n9440) );
  AOI22_X1 U11838 ( .A1(n13739), .A2(n9471), .B1(n13481), .B2(n6502), .ZN(
        n9436) );
  INV_X1 U11839 ( .A(n9436), .ZN(n9439) );
  INV_X1 U11840 ( .A(n13739), .ZN(n13179) );
  OAI22_X1 U11841 ( .A1(n13179), .A2(n9477), .B1(n13443), .B2(n6502), .ZN(
        n9435) );
  OAI21_X1 U11842 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9443) );
  OAI22_X1 U11843 ( .A1(n13451), .A2(n9471), .B1(n13461), .B2(n6502), .ZN(
        n9444) );
  OAI22_X1 U11844 ( .A1(n13451), .A2(n6502), .B1(n13461), .B2(n9477), .ZN(
        n9442) );
  AOI22_X1 U11845 ( .A1(n13656), .A2(n9471), .B1(n13441), .B2(n6502), .ZN(
        n9461) );
  INV_X1 U11846 ( .A(n13656), .ZN(n13432) );
  OAI22_X1 U11847 ( .A1(n13432), .A2(n9471), .B1(n13234), .B2(n6502), .ZN(
        n9445) );
  AND2_X1 U11848 ( .A1(n13427), .A2(n9471), .ZN(n9446) );
  AOI21_X1 U11849 ( .B1(n13733), .B2(n6502), .A(n9446), .ZN(n9466) );
  NAND2_X1 U11850 ( .A1(n13733), .A2(n9477), .ZN(n9448) );
  NAND2_X1 U11851 ( .A1(n13427), .A2(n6502), .ZN(n9447) );
  NAND2_X1 U11852 ( .A1(n9448), .A2(n9447), .ZN(n9465) );
  NAND2_X1 U11853 ( .A1(n13762), .A2(n9468), .ZN(n9450) );
  NAND2_X1 U11854 ( .A1(n9097), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9449) );
  INV_X1 U11855 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13646) );
  NOR2_X1 U11856 ( .A1(n9451), .A2(n13646), .ZN(n9456) );
  INV_X1 U11857 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9452) );
  NOR2_X1 U11858 ( .A1(n9453), .A2(n9452), .ZN(n9455) );
  INV_X1 U11859 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13726) );
  NOR2_X1 U11860 ( .A1(n8904), .A2(n13726), .ZN(n9454) );
  OR3_X1 U11861 ( .A1(n9456), .A2(n9455), .A3(n9454), .ZN(n13388) );
  XNOR2_X1 U11862 ( .A(n13384), .B(n13388), .ZN(n9527) );
  AND2_X1 U11863 ( .A1(n13254), .A2(n6502), .ZN(n9457) );
  AOI21_X1 U11864 ( .B1(n13401), .B2(n9477), .A(n9457), .ZN(n9480) );
  NAND2_X1 U11865 ( .A1(n13401), .A2(n6502), .ZN(n9459) );
  NAND2_X1 U11866 ( .A1(n13254), .A2(n9477), .ZN(n9458) );
  NAND2_X1 U11867 ( .A1(n9459), .A2(n9458), .ZN(n9479) );
  NAND2_X1 U11868 ( .A1(n9480), .A2(n9479), .ZN(n9467) );
  OAI211_X1 U11869 ( .C1(n9466), .C2(n9465), .A(n9527), .B(n9467), .ZN(n9460)
         );
  AOI21_X1 U11870 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(n9463) );
  NAND2_X1 U11871 ( .A1(n9464), .A2(n9463), .ZN(n9488) );
  NAND4_X1 U11872 ( .A1(n9527), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n9486)
         );
  NAND2_X1 U11873 ( .A1(n12444), .A2(n9468), .ZN(n9470) );
  NAND2_X1 U11874 ( .A1(n9097), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9469) );
  OAI22_X1 U11875 ( .A1(n13731), .A2(n9471), .B1(n9472), .B2(n6502), .ZN(n9490) );
  INV_X1 U11876 ( .A(n9472), .ZN(n13253) );
  INV_X1 U11877 ( .A(n13388), .ZN(n9491) );
  OR2_X1 U11878 ( .A1(n9473), .A2(n9512), .ZN(n9475) );
  AND2_X1 U11879 ( .A1(n9529), .A2(n9531), .ZN(n9474) );
  AND2_X1 U11880 ( .A1(n9475), .A2(n9474), .ZN(n9476) );
  OAI21_X1 U11881 ( .B1(n9491), .B2(n9477), .A(n9476), .ZN(n9478) );
  AOI22_X1 U11882 ( .A1(n13396), .A2(n9471), .B1(n13253), .B2(n9478), .ZN(
        n9489) );
  OAI22_X1 U11883 ( .A1(n9490), .A2(n9489), .B1(n9480), .B2(n9479), .ZN(n9484)
         );
  MUX2_X1 U11884 ( .A(n13388), .B(n9471), .S(n13384), .Z(n9481) );
  OAI21_X1 U11885 ( .B1(n9491), .B2(n6502), .A(n9481), .ZN(n9483) );
  NAND2_X1 U11886 ( .A1(n9484), .A2(n9483), .ZN(n9485) );
  NAND2_X1 U11887 ( .A1(n9488), .A2(n9487), .ZN(n9496) );
  NAND2_X1 U11888 ( .A1(n9490), .A2(n9489), .ZN(n9495) );
  NOR2_X1 U11889 ( .A1(n9491), .A2(n6502), .ZN(n9493) );
  NOR2_X1 U11890 ( .A1(n13388), .A2(n9477), .ZN(n9492) );
  MUX2_X1 U11891 ( .A(n9493), .B(n9492), .S(n13384), .Z(n9494) );
  AOI21_X2 U11892 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9503) );
  INV_X1 U11893 ( .A(n9275), .ZN(n11206) );
  NAND2_X1 U11894 ( .A1(n9529), .A2(n13379), .ZN(n9497) );
  OAI211_X1 U11895 ( .C1(n9217), .C2(n11206), .A(n9531), .B(n9497), .ZN(n9498)
         );
  NAND2_X1 U11896 ( .A1(n9503), .A2(n9499), .ZN(n9500) );
  INV_X1 U11897 ( .A(n10682), .ZN(n10449) );
  AND2_X1 U11898 ( .A1(n10449), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9534) );
  NAND2_X1 U11899 ( .A1(n9500), .A2(n9534), .ZN(n9541) );
  INV_X1 U11900 ( .A(n9217), .ZN(n12137) );
  INV_X1 U11901 ( .A(n9529), .ZN(n11879) );
  MUX2_X1 U11902 ( .A(n12137), .B(n11879), .S(n9512), .Z(n9501) );
  NOR2_X1 U11903 ( .A1(n9501), .A2(n13379), .ZN(n9502) );
  NAND2_X1 U11904 ( .A1(n9503), .A2(n8803), .ZN(n9538) );
  XNOR2_X1 U11905 ( .A(n13396), .B(n13253), .ZN(n9528) );
  NAND2_X1 U11906 ( .A1(n9506), .A2(n13532), .ZN(n13548) );
  XNOR2_X1 U11907 ( .A(n14931), .B(n11787), .ZN(n11921) );
  NAND2_X1 U11908 ( .A1(n9508), .A2(n9507), .ZN(n11915) );
  NAND2_X1 U11909 ( .A1(n10715), .A2(n9510), .ZN(n9511) );
  NAND2_X1 U11910 ( .A1(n11273), .A2(n9511), .ZN(n15094) );
  AND4_X1 U11911 ( .A1(n9509), .A2(n9512), .A3(n11262), .A4(n15094), .ZN(n9514) );
  AND2_X1 U11912 ( .A1(n11225), .A2(n10637), .ZN(n9513) );
  NAND4_X1 U11913 ( .A1(n9514), .A2(n11175), .A3(n9513), .A4(n11298), .ZN(
        n9515) );
  NOR3_X1 U11914 ( .A1(n11387), .A2(n11318), .A3(n9515), .ZN(n9516) );
  NAND4_X1 U11915 ( .A1(n11785), .A2(n11484), .A3(n11613), .A4(n9516), .ZN(
        n9517) );
  OR4_X1 U11916 ( .A1(n14648), .A2(n11921), .A3(n11915), .A4(n9517), .ZN(n9519) );
  OR4_X1 U11917 ( .A1(n13599), .A2(n9519), .A3(n13618), .A4(n9518), .ZN(n9520)
         );
  NOR3_X1 U11918 ( .A1(n13548), .A2(n13577), .A3(n9520), .ZN(n9521) );
  XNOR2_X1 U11919 ( .A(n13702), .B(n13579), .ZN(n13572) );
  NAND4_X1 U11920 ( .A1(n13511), .A2(n9521), .A3(n13534), .A4(n13572), .ZN(
        n9522) );
  NOR3_X1 U11921 ( .A1(n13478), .A2(n13496), .A3(n9522), .ZN(n9523) );
  AND4_X1 U11922 ( .A1(n13433), .A2(n13452), .A3(n9523), .A4(n13458), .ZN(
        n9524) );
  AND2_X1 U11923 ( .A1(n9524), .A2(n13408), .ZN(n9526) );
  NAND4_X1 U11924 ( .A1(n9528), .A2(n9527), .A3(n9526), .A4(n9525), .ZN(n9530)
         );
  INV_X1 U11925 ( .A(n9534), .ZN(n12188) );
  NOR4_X1 U11926 ( .A1(n9530), .A2(n9529), .A3(n11210), .A4(n12188), .ZN(n9536) );
  INV_X1 U11927 ( .A(P2_B_REG_SCAN_IN), .ZN(n9533) );
  NOR4_X1 U11928 ( .A1(n15093), .A2(n13539), .A3(n13774), .A4(n9531), .ZN(
        n9532) );
  AOI211_X1 U11929 ( .C1(n9534), .C2(n12137), .A(n9533), .B(n9532), .ZN(n9535)
         );
  OAI21_X1 U11930 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(P2_U3328) );
  INV_X1 U11931 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12190) );
  INV_X1 U11932 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U11933 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12421), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11746), .ZN(n9940) );
  AOI22_X1 U11934 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11573), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7056), .ZN(n9923) );
  XNOR2_X1 U11935 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9888) );
  NAND2_X1 U11936 ( .A1(n9682), .A2(n9681), .ZN(n9545) );
  INV_X1 U11937 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U11938 ( .A1(n9543), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U11939 ( .A1(n9545), .A2(n9544), .ZN(n9703) );
  XNOR2_X1 U11940 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9701) );
  NAND2_X1 U11941 ( .A1(n9703), .A2(n9701), .ZN(n9548) );
  NAND2_X1 U11942 ( .A1(n9546), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U11943 ( .A1(n10342), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U11944 ( .A1(n10370), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9550) );
  NAND2_X1 U11945 ( .A1(n10403), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U11946 ( .A1(n9765), .A2(n9763), .ZN(n9555) );
  NAND2_X1 U11947 ( .A1(n10417), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9554) );
  XNOR2_X1 U11948 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9778) );
  NAND2_X1 U11949 ( .A1(n9779), .A2(n9778), .ZN(n9558) );
  NAND2_X1 U11950 ( .A1(n9556), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9557) );
  XNOR2_X1 U11951 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9794) );
  NAND2_X1 U11952 ( .A1(n9559), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9560) );
  XNOR2_X1 U11953 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9810) );
  XNOR2_X1 U11954 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9822) );
  NAND2_X1 U11955 ( .A1(n10795), .A2(n9564), .ZN(n9565) );
  XNOR2_X1 U11956 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9853) );
  INV_X1 U11957 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U11958 ( .A1(n9566), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9567) );
  XNOR2_X1 U11959 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9874) );
  AOI22_X1 U11960 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n11357), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7058), .ZN(n9909) );
  NAND2_X1 U11961 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n9573), .ZN(n9575) );
  NAND2_X1 U11962 ( .A1(n9960), .A2(n11744), .ZN(n9574) );
  INV_X1 U11963 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U11964 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11880), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12589), .ZN(n9972) );
  AOI22_X1 U11965 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12138), .B2(n7565), .ZN(n9988) );
  INV_X1 U11966 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U11967 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n12190), .B2(n12195), .ZN(n9610) );
  XNOR2_X1 U11968 ( .A(n12380), .B(n10004), .ZN(n12027) );
  NOR2_X1 U11969 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), 
        .ZN(n9578) );
  NOR2_X1 U11970 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n9579) );
  INV_X1 U11971 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9587) );
  AND2_X2 U11972 ( .A1(n10941), .A2(n10344), .ZN(n9704) );
  CLKBUF_X3 U11973 ( .A(n9704), .Z(n10076) );
  NAND2_X1 U11974 ( .A1(n12027), .A2(n10076), .ZN(n9594) );
  OR2_X1 U11975 ( .A1(n10033), .A2(n7569), .ZN(n9593) );
  NAND2_X1 U11976 ( .A1(n9596), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9597) );
  MUX2_X1 U11977 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9597), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9600) );
  INV_X1 U11978 ( .A(n13121), .ZN(n9602) );
  NAND2_X1 U11979 ( .A1(n10036), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9609) );
  INV_X1 U11980 ( .A(n12578), .ZN(n9605) );
  NAND2_X1 U11981 ( .A1(n9717), .A2(n9716), .ZN(n9719) );
  INV_X1 U11982 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U11983 ( .A1(n11835), .A2(n12012), .ZN(n9603) );
  INV_X1 U11984 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9932) );
  INV_X1 U11985 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12674) );
  AND2_X1 U11986 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9615), .ZN(n9604) );
  OR2_X1 U11987 ( .A1(n9604), .A2(n10010), .ZN(n12896) );
  NAND2_X1 U11988 ( .A1(n10063), .A2(n12896), .ZN(n9608) );
  NAND2_X1 U11989 ( .A1(n10098), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U11990 ( .A1(n10099), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9606) );
  XNOR2_X1 U11991 ( .A(n13019), .B(n12475), .ZN(n12892) );
  XNOR2_X1 U11992 ( .A(n9611), .B(n9610), .ZN(n11740) );
  NAND2_X1 U11993 ( .A1(n11740), .A2(n10076), .ZN(n9613) );
  OR2_X1 U11994 ( .A1(n6480), .A2(n8560), .ZN(n9612) );
  OR2_X1 U11995 ( .A1(n9994), .A2(n9614), .ZN(n9616) );
  NAND2_X1 U11996 ( .A1(n9616), .A2(n9615), .ZN(n12914) );
  NAND2_X1 U11997 ( .A1(n12914), .A2(n10063), .ZN(n9619) );
  AOI22_X1 U11998 ( .A1(n10036), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n10098), 
        .B2(P3_REG0_REG_23__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U11999 ( .A1(n10099), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9617) );
  NOR2_X1 U12000 ( .A1(n12603), .A2(n12659), .ZN(n12890) );
  NOR2_X1 U12001 ( .A1(n12892), .A2(n12890), .ZN(n10147) );
  NAND2_X1 U12002 ( .A1(n9623), .A2(n9927), .ZN(n9943) );
  INV_X1 U12003 ( .A(n9943), .ZN(n9624) );
  INV_X1 U12004 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9627) );
  INV_X2 U12005 ( .A(n10939), .ZN(n10294) );
  NAND2_X1 U12006 ( .A1(n13019), .A2(n12475), .ZN(n10148) );
  XOR2_X1 U12007 ( .A(n10294), .B(n10148), .Z(n10003) );
  INV_X1 U12008 ( .A(n9694), .ZN(n9895) );
  NAND2_X1 U12009 ( .A1(n10036), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12010 ( .A1(n9719), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9628) );
  AND2_X1 U12011 ( .A1(n9741), .A2(n9628), .ZN(n15194) );
  INV_X1 U12012 ( .A(n15194), .ZN(n11426) );
  NAND2_X1 U12013 ( .A1(n10063), .A2(n11426), .ZN(n9631) );
  NAND2_X1 U12014 ( .A1(n10098), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U12015 ( .A1(n10099), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9629) );
  NAND4_X1 U12016 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n12717) );
  XNOR2_X1 U12017 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9633) );
  XNOR2_X1 U12018 ( .A(n9634), .B(n9633), .ZN(n10386) );
  NAND2_X1 U12019 ( .A1(n10076), .A2(n10386), .ZN(n9642) );
  OR2_X1 U12020 ( .A1(n10033), .A2(n10387), .ZN(n9641) );
  INV_X1 U12021 ( .A(n9660), .ZN(n9636) );
  NOR2_X1 U12022 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9635) );
  NAND2_X1 U12023 ( .A1(n9636), .A2(n9635), .ZN(n9638) );
  NAND2_X1 U12024 ( .A1(n9638), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9637) );
  MUX2_X1 U12025 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9637), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n9639) );
  NAND2_X1 U12026 ( .A1(n9639), .A2(n9751), .ZN(n11095) );
  OR2_X1 U12027 ( .A1(n10941), .A2(n11095), .ZN(n9640) );
  AND2_X1 U12028 ( .A1(n12717), .A2(n11801), .ZN(n9736) );
  INV_X1 U12029 ( .A(n9736), .ZN(n10115) );
  XNOR2_X1 U12030 ( .A(n9644), .B(n7061), .ZN(n10385) );
  NAND2_X1 U12031 ( .A1(n9704), .A2(n10385), .ZN(n9647) );
  NAND2_X1 U12032 ( .A1(n6942), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9645) );
  XNOR2_X1 U12033 ( .A(n9645), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10962) );
  OR2_X1 U12034 ( .A1(n10941), .A2(n10962), .ZN(n9646) );
  OAI211_X1 U12035 ( .C1(n6480), .C2(SI_3_), .A(n9647), .B(n9646), .ZN(n10219)
         );
  NAND2_X1 U12036 ( .A1(n9693), .A2(n15203), .ZN(n9651) );
  NAND2_X1 U12037 ( .A1(n9694), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U12038 ( .A1(n9695), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U12039 ( .A1(n9696), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9648) );
  NAND4_X1 U12040 ( .A1(n9651), .A2(n9650), .A3(n9649), .A4(n9648), .ZN(n12721) );
  NAND2_X1 U12041 ( .A1(n10036), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9657) );
  AND2_X1 U12042 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9653) );
  OR2_X1 U12043 ( .A1(n9653), .A2(n9717), .ZN(n11154) );
  NAND2_X1 U12044 ( .A1(n10063), .A2(n11154), .ZN(n9656) );
  NAND2_X1 U12045 ( .A1(n10098), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U12046 ( .A1(n10099), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9654) );
  XNOR2_X1 U12047 ( .A(n9659), .B(n7064), .ZN(n10392) );
  NAND2_X1 U12048 ( .A1(n10076), .A2(n10392), .ZN(n9667) );
  OR2_X1 U12049 ( .A1(n10033), .A2(SI_4_), .ZN(n9666) );
  NAND2_X1 U12050 ( .A1(n9660), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9663) );
  INV_X1 U12051 ( .A(n9663), .ZN(n9661) );
  NAND2_X1 U12052 ( .A1(n9661), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9664) );
  INV_X1 U12053 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12054 ( .A1(n9663), .A2(n9662), .ZN(n9726) );
  OR2_X1 U12055 ( .A1(n10941), .A2(n10965), .ZN(n9665) );
  AND3_X2 U12056 ( .A1(n9667), .A2(n9666), .A3(n9665), .ZN(n11156) );
  NAND2_X1 U12057 ( .A1(n11248), .A2(n11156), .ZN(n10113) );
  INV_X1 U12058 ( .A(n11156), .ZN(n11166) );
  NAND2_X1 U12059 ( .A1(n12719), .A2(n11166), .ZN(n9731) );
  NAND2_X1 U12060 ( .A1(n10113), .A2(n9731), .ZN(n10221) );
  NAND2_X1 U12061 ( .A1(n9693), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U12062 ( .A1(n9694), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U12063 ( .A1(n9695), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U12064 ( .A1(n9696), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9668) );
  INV_X1 U12065 ( .A(n9681), .ZN(n9674) );
  NAND2_X1 U12066 ( .A1(n9672), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U12067 ( .A1(n9674), .A2(n9673), .ZN(n10393) );
  NAND2_X1 U12068 ( .A1(n9704), .A2(n10393), .ZN(n9676) );
  INV_X1 U12069 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10943) );
  OR2_X1 U12070 ( .A1(n10941), .A2(n10943), .ZN(n9675) );
  NAND2_X1 U12071 ( .A1(n10209), .A2(n10812), .ZN(n15322) );
  INV_X1 U12072 ( .A(n11445), .ZN(n9691) );
  NOR2_X1 U12073 ( .A1(n10209), .A2(n10812), .ZN(n10167) );
  NAND2_X1 U12074 ( .A1(n9696), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U12075 ( .A1(n9693), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U12076 ( .A1(n9695), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12077 ( .A1(n9694), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9677) );
  AND4_X2 U12078 ( .A1(n9680), .A2(n9679), .A3(n9678), .A4(n9677), .ZN(n10211)
         );
  XNOR2_X1 U12079 ( .A(n9682), .B(n9681), .ZN(n10398) );
  NAND2_X1 U12080 ( .A1(n9704), .A2(n10398), .ZN(n9688) );
  NAND2_X1 U12081 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9683) );
  MUX2_X1 U12082 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9683), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n9686) );
  INV_X1 U12083 ( .A(n9684), .ZN(n9685) );
  OR2_X1 U12084 ( .A1(n10941), .A2(n10959), .ZN(n9687) );
  NAND2_X1 U12085 ( .A1(n12723), .A2(n10212), .ZN(n10109) );
  NAND2_X1 U12086 ( .A1(n10109), .A2(n10579), .ZN(n10210) );
  NOR2_X1 U12087 ( .A1(n10167), .A2(n10181), .ZN(n9690) );
  INV_X1 U12088 ( .A(n10579), .ZN(n9689) );
  OAI33_X1 U12089 ( .A1(n9691), .A2(n10167), .A3(n15323), .B1(n10939), .B2(
        n9690), .B3(n9689), .ZN(n9692) );
  OAI21_X1 U12090 ( .B1(n11075), .B2(n15322), .A(n9692), .ZN(n9710) );
  NAND2_X1 U12091 ( .A1(n9693), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U12092 ( .A1(n9694), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U12093 ( .A1(n9695), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12094 ( .A1(n9696), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9697) );
  INV_X1 U12095 ( .A(n9701), .ZN(n9702) );
  XNOR2_X1 U12096 ( .A(n9703), .B(n9702), .ZN(n10390) );
  NAND2_X1 U12097 ( .A1(n9704), .A2(n10390), .ZN(n9708) );
  OR2_X1 U12098 ( .A1(n10058), .A2(SI_2_), .ZN(n9707) );
  NOR2_X1 U12099 ( .A1(n9684), .A2(n9589), .ZN(n9705) );
  OR2_X1 U12100 ( .A1(n10941), .A2(n10961), .ZN(n9706) );
  NAND2_X1 U12101 ( .A1(n11025), .A2(n10837), .ZN(n10110) );
  MUX2_X1 U12102 ( .A(n10579), .B(n10109), .S(n10294), .Z(n9709) );
  INV_X1 U12103 ( .A(n10110), .ZN(n9711) );
  OAI21_X1 U12104 ( .B1(n9715), .B2(n9711), .A(n10294), .ZN(n9712) );
  NAND2_X1 U12105 ( .A1(n12721), .A2(n10219), .ZN(n10111) );
  AOI21_X1 U12106 ( .B1(n10111), .B2(n9713), .A(n10294), .ZN(n9714) );
  NAND2_X1 U12107 ( .A1(n10036), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9723) );
  OR2_X1 U12108 ( .A1(n9717), .A2(n9716), .ZN(n9718) );
  NAND2_X1 U12109 ( .A1(n9719), .A2(n9718), .ZN(n11246) );
  NAND2_X1 U12110 ( .A1(n10063), .A2(n11246), .ZN(n9722) );
  NAND2_X1 U12111 ( .A1(n10098), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U12112 ( .A1(n9695), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9720) );
  NAND4_X1 U12113 ( .A1(n9723), .A2(n9722), .A3(n9721), .A4(n9720), .ZN(n12718) );
  XNOR2_X1 U12114 ( .A(n9725), .B(n6780), .ZN(n10397) );
  NAND2_X1 U12115 ( .A1(n10076), .A2(n10397), .ZN(n9730) );
  NAND2_X1 U12116 ( .A1(n9726), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9728) );
  XNOR2_X1 U12117 ( .A(n9728), .B(n9727), .ZN(n15240) );
  OR2_X1 U12118 ( .A1(n10941), .A2(n10966), .ZN(n9729) );
  XNOR2_X1 U12119 ( .A(n12718), .B(n11449), .ZN(n10168) );
  NAND2_X1 U12120 ( .A1(n11344), .A2(n9731), .ZN(n9732) );
  NOR2_X1 U12121 ( .A1(n12717), .A2(n11801), .ZN(n9737) );
  INV_X1 U12122 ( .A(n9737), .ZN(n10116) );
  INV_X1 U12123 ( .A(n12718), .ZN(n11803) );
  INV_X1 U12124 ( .A(n11449), .ZN(n11247) );
  NAND2_X1 U12125 ( .A1(n11803), .A2(n11247), .ZN(n10114) );
  OAI211_X1 U12126 ( .C1(n9734), .C2(n9732), .A(n10116), .B(n10114), .ZN(n9740) );
  INV_X1 U12127 ( .A(n10113), .ZN(n9733) );
  NOR3_X1 U12128 ( .A1(n9734), .A2(n9733), .A3(n10168), .ZN(n9735) );
  AOI211_X1 U12129 ( .C1(n12718), .C2(n11449), .A(n9736), .B(n9735), .ZN(n9738) );
  NOR2_X1 U12130 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  AND2_X1 U12131 ( .A1(n9741), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9742) );
  NOR2_X1 U12132 ( .A1(n9757), .A2(n9742), .ZN(n15168) );
  INV_X1 U12133 ( .A(n15168), .ZN(n9743) );
  NAND2_X1 U12134 ( .A1(n10063), .A2(n9743), .ZN(n9747) );
  NAND2_X1 U12135 ( .A1(n10036), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U12136 ( .A1(n10099), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U12137 ( .A1(n10098), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9744) );
  XNOR2_X1 U12138 ( .A(n9749), .B(n9748), .ZN(n10375) );
  NAND2_X1 U12139 ( .A1(n10076), .A2(n10375), .ZN(n9755) );
  OR2_X1 U12140 ( .A1(n10033), .A2(SI_7_), .ZN(n9754) );
  NAND2_X1 U12141 ( .A1(n9751), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9750) );
  MUX2_X1 U12142 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9750), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n9752) );
  NAND2_X1 U12143 ( .A1(n9752), .A2(n9780), .ZN(n11520) );
  OR2_X1 U12144 ( .A1(n10941), .A2(n11534), .ZN(n9753) );
  NAND2_X1 U12145 ( .A1(n11809), .A2(n15162), .ZN(n10118) );
  NAND2_X1 U12146 ( .A1(n11810), .A2(n11674), .ZN(n9770) );
  NAND2_X1 U12147 ( .A1(n10036), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9762) );
  NOR2_X1 U12148 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  OR2_X1 U12149 ( .A1(n9772), .A2(n9758), .ZN(n11646) );
  NAND2_X1 U12150 ( .A1(n10063), .A2(n11646), .ZN(n9761) );
  NAND2_X1 U12151 ( .A1(n10098), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12152 ( .A1(n10099), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9759) );
  INV_X1 U12153 ( .A(n9763), .ZN(n9764) );
  XNOR2_X1 U12154 ( .A(n9765), .B(n9764), .ZN(n10371) );
  NAND2_X1 U12155 ( .A1(n10076), .A2(n10371), .ZN(n9769) );
  NAND2_X1 U12156 ( .A1(n9780), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9767) );
  INV_X1 U12157 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9766) );
  OR2_X1 U12158 ( .A1(n10941), .A2(n15256), .ZN(n9768) );
  OAI211_X1 U12159 ( .C1(n10033), .C2(n10372), .A(n9769), .B(n9768), .ZN(
        n12618) );
  NAND2_X1 U12160 ( .A1(n11816), .A2(n12618), .ZN(n10119) );
  INV_X1 U12161 ( .A(n11816), .ZN(n12716) );
  INV_X1 U12162 ( .A(n12618), .ZN(n15351) );
  NAND2_X1 U12163 ( .A1(n12716), .A2(n15351), .ZN(n9786) );
  MUX2_X1 U12164 ( .A(n10118), .B(n9770), .S(n10294), .Z(n9771) );
  NAND2_X1 U12165 ( .A1(n10036), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9777) );
  OR2_X1 U12166 ( .A1(n9772), .A2(n8586), .ZN(n9773) );
  NAND2_X1 U12167 ( .A1(n9788), .A2(n9773), .ZN(n11820) );
  NAND2_X1 U12168 ( .A1(n10063), .A2(n11820), .ZN(n9776) );
  NAND2_X1 U12169 ( .A1(n10098), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12170 ( .A1(n10099), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9774) );
  NAND4_X1 U12171 ( .A1(n9777), .A2(n9776), .A3(n9775), .A4(n9774), .ZN(n12715) );
  XNOR2_X1 U12172 ( .A(n9779), .B(n9778), .ZN(n10347) );
  NAND2_X1 U12173 ( .A1(n10076), .A2(n10347), .ZN(n9785) );
  OR2_X1 U12174 ( .A1(n10033), .A2(SI_9_), .ZN(n9784) );
  OAI21_X1 U12175 ( .B1(n9780), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9782) );
  INV_X1 U12176 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9781) );
  XNOR2_X1 U12177 ( .A(n9782), .B(n9781), .ZN(n15284) );
  OR2_X1 U12178 ( .A1(n10941), .A2(n11544), .ZN(n9783) );
  NAND2_X1 U12179 ( .A1(n12715), .A2(n11799), .ZN(n10229) );
  OAI21_X1 U12180 ( .B1(n12715), .B2(n11799), .A(n10229), .ZN(n10228) );
  MUX2_X1 U12181 ( .A(n9786), .B(n10119), .S(n10294), .Z(n9787) );
  MUX2_X1 U12182 ( .A(n11799), .B(n12715), .S(n10294), .Z(n9802) );
  NAND2_X1 U12183 ( .A1(n10036), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U12184 ( .A1(n9788), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U12185 ( .A1(n9816), .A2(n9789), .ZN(n11937) );
  NAND2_X1 U12186 ( .A1(n10063), .A2(n11937), .ZN(n9792) );
  NAND2_X1 U12187 ( .A1(n10098), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U12188 ( .A1(n10099), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9790) );
  XNOR2_X1 U12189 ( .A(n9795), .B(n9794), .ZN(n10377) );
  NAND2_X1 U12190 ( .A1(n10076), .A2(n10377), .ZN(n9801) );
  OR2_X1 U12191 ( .A1(n10033), .A2(SI_10_), .ZN(n9800) );
  OR2_X1 U12192 ( .A1(n9620), .A2(n9589), .ZN(n9797) );
  MUX2_X1 U12193 ( .A(n9797), .B(P3_IR_REG_31__SCAN_IN), .S(n9796), .Z(n9798)
         );
  NAND2_X1 U12194 ( .A1(n9798), .A2(n10187), .ZN(n11830) );
  INV_X1 U12195 ( .A(n11830), .ZN(n11548) );
  OR2_X1 U12196 ( .A1(n10941), .A2(n11548), .ZN(n9799) );
  NAND2_X1 U12197 ( .A1(n12334), .A2(n11947), .ZN(n10122) );
  INV_X1 U12198 ( .A(n12334), .ZN(n12714) );
  NAND2_X1 U12199 ( .A1(n12714), .A2(n11936), .ZN(n10121) );
  NAND2_X1 U12200 ( .A1(n10122), .A2(n10121), .ZN(n11752) );
  AOI21_X1 U12201 ( .B1(n10229), .B2(n9802), .A(n11752), .ZN(n9804) );
  NOR2_X1 U12202 ( .A1(n12334), .A2(n10294), .ZN(n9803) );
  AOI22_X1 U12203 ( .A1(n9805), .A2(n9804), .B1(n9803), .B2(n11936), .ZN(n9832) );
  NAND2_X1 U12204 ( .A1(n10036), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9809) );
  XNOR2_X1 U12205 ( .A(n9816), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U12206 ( .A1(n10063), .A2(n12338), .ZN(n9808) );
  NAND2_X1 U12207 ( .A1(n10098), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12208 ( .A1(n10099), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9806) );
  XNOR2_X1 U12209 ( .A(n9811), .B(n9810), .ZN(n10379) );
  NAND2_X1 U12210 ( .A1(n10076), .A2(n10379), .ZN(n9815) );
  OR2_X1 U12211 ( .A1(n10033), .A2(SI_11_), .ZN(n9814) );
  NAND2_X1 U12212 ( .A1(n10187), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9812) );
  XNOR2_X1 U12213 ( .A(n9812), .B(n6851), .ZN(n12007) );
  INV_X1 U12214 ( .A(n12007), .ZN(n12015) );
  OR2_X1 U12215 ( .A1(n10941), .A2(n12015), .ZN(n9813) );
  NAND2_X1 U12216 ( .A1(n12352), .A2(n12331), .ZN(n10124) );
  INV_X1 U12217 ( .A(n12352), .ZN(n12713) );
  NAND2_X1 U12218 ( .A1(n12713), .A2(n14622), .ZN(n9833) );
  INV_X1 U12219 ( .A(n10122), .ZN(n9830) );
  NAND2_X1 U12220 ( .A1(n10036), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9821) );
  OAI21_X1 U12221 ( .B1(n9816), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12222 ( .A1(n9817), .A2(n9843), .ZN(n12354) );
  NAND2_X1 U12223 ( .A1(n10063), .A2(n12354), .ZN(n9820) );
  NAND2_X1 U12224 ( .A1(n10098), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U12225 ( .A1(n10099), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9818) );
  NAND4_X1 U12226 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n12712) );
  INV_X1 U12227 ( .A(n9822), .ZN(n9823) );
  XNOR2_X1 U12228 ( .A(n9824), .B(n9823), .ZN(n10400) );
  NAND2_X1 U12229 ( .A1(n10400), .A2(n10076), .ZN(n9829) );
  NAND2_X1 U12230 ( .A1(n6508), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9826) );
  INV_X1 U12231 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9825) );
  XNOR2_X1 U12232 ( .A(n9826), .B(n9825), .ZN(n12263) );
  OR2_X1 U12233 ( .A1(n10941), .A2(n12263), .ZN(n9828) );
  OR2_X1 U12234 ( .A1(n10033), .A2(n10401), .ZN(n9827) );
  NOR2_X1 U12235 ( .A1(n12712), .A2(n14617), .ZN(n9836) );
  AOI211_X1 U12236 ( .C1(n10172), .C2(n9830), .A(n6980), .B(n9836), .ZN(n9831)
         );
  OAI22_X1 U12237 ( .A1(n9832), .A2(n6978), .B1(n10939), .B2(n9831), .ZN(n9835) );
  NAND2_X1 U12238 ( .A1(n12712), .A2(n14617), .ZN(n10125) );
  AOI21_X1 U12239 ( .B1(n10125), .B2(n9833), .A(n10294), .ZN(n9834) );
  AOI21_X1 U12240 ( .B1(n9835), .B2(n10125), .A(n9834), .ZN(n9850) );
  INV_X1 U12241 ( .A(n9836), .ZN(n10126) );
  NOR2_X1 U12242 ( .A1(n10126), .A2(n10294), .ZN(n9849) );
  XNOR2_X1 U12243 ( .A(n9837), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U12244 ( .A1(n10441), .A2(n10076), .ZN(n9842) );
  OR2_X1 U12245 ( .A1(n6508), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12246 ( .A1(n9855), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9839) );
  XNOR2_X1 U12247 ( .A(n9839), .B(n9838), .ZN(n12732) );
  OAI22_X1 U12248 ( .A1(n10033), .A2(SI_13_), .B1(n12257), .B2(n10941), .ZN(
        n9840) );
  INV_X1 U12249 ( .A(n9840), .ZN(n9841) );
  NAND2_X1 U12250 ( .A1(n10036), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9848) );
  AND2_X1 U12251 ( .A1(n9843), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9844) );
  OR2_X1 U12252 ( .A1(n9844), .A2(n9865), .ZN(n12184) );
  NAND2_X1 U12253 ( .A1(n10063), .A2(n12184), .ZN(n9847) );
  NAND2_X1 U12254 ( .A1(n10098), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12255 ( .A1(n10099), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9845) );
  NAND4_X1 U12256 ( .A1(n9848), .A2(n9847), .A3(n9846), .A4(n9845), .ZN(n12711) );
  NOR2_X1 U12257 ( .A1(n12222), .A2(n12711), .ZN(n10127) );
  AND2_X1 U12258 ( .A1(n12222), .A2(n12711), .ZN(n9851) );
  NOR2_X1 U12259 ( .A1(n10127), .A2(n9851), .ZN(n12093) );
  OAI21_X1 U12260 ( .B1(n9850), .B2(n9849), .A(n12093), .ZN(n9872) );
  INV_X1 U12261 ( .A(n10127), .ZN(n9852) );
  INV_X1 U12262 ( .A(n9851), .ZN(n10128) );
  MUX2_X1 U12263 ( .A(n9852), .B(n10128), .S(n10294), .Z(n9871) );
  XNOR2_X1 U12264 ( .A(n9854), .B(n9853), .ZN(n10508) );
  NAND2_X1 U12265 ( .A1(n10508), .A2(n10076), .ZN(n9863) );
  NOR2_X1 U12266 ( .A1(n9855), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U12267 ( .A1(n9858), .A2(n9589), .ZN(n9856) );
  MUX2_X1 U12268 ( .A(n9589), .B(n9856), .S(P3_IR_REG_14__SCAN_IN), .Z(n9860)
         );
  NAND2_X1 U12269 ( .A1(n9858), .A2(n9857), .ZN(n9891) );
  INV_X1 U12270 ( .A(n9891), .ZN(n9859) );
  NOR2_X1 U12271 ( .A1(n9860), .A2(n9859), .ZN(n12735) );
  OAI22_X1 U12272 ( .A1(n10033), .A2(SI_14_), .B1(n12735), .B2(n10941), .ZN(
        n9861) );
  INV_X1 U12273 ( .A(n9861), .ZN(n9862) );
  NAND2_X1 U12274 ( .A1(n10036), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9870) );
  OR2_X1 U12275 ( .A1(n9865), .A2(n9864), .ZN(n9866) );
  NAND2_X1 U12276 ( .A1(n9881), .A2(n9866), .ZN(n12284) );
  NAND2_X1 U12277 ( .A1(n10063), .A2(n12284), .ZN(n9869) );
  NAND2_X1 U12278 ( .A1(n10098), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12279 ( .A1(n10099), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9867) );
  NAND4_X1 U12280 ( .A1(n9870), .A2(n9869), .A3(n9868), .A4(n9867), .ZN(n12710) );
  OR2_X1 U12281 ( .A1(n12330), .A2(n12710), .ZN(n10130) );
  NAND2_X1 U12282 ( .A1(n12330), .A2(n12710), .ZN(n9873) );
  NAND2_X1 U12283 ( .A1(n10130), .A2(n9873), .ZN(n12143) );
  INV_X1 U12284 ( .A(n9873), .ZN(n10131) );
  MUX2_X1 U12285 ( .A(n6995), .B(n10131), .S(n10294), .Z(n9887) );
  INV_X1 U12286 ( .A(n9874), .ZN(n9875) );
  XNOR2_X1 U12287 ( .A(n9876), .B(n9875), .ZN(n10521) );
  NAND2_X1 U12288 ( .A1(n10521), .A2(n10076), .ZN(n9880) );
  NAND2_X1 U12289 ( .A1(n9891), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9877) );
  XNOR2_X1 U12290 ( .A(n9877), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12785) );
  OAI22_X1 U12291 ( .A1(n10033), .A2(n10522), .B1(n10941), .B2(n12798), .ZN(
        n9878) );
  INV_X1 U12292 ( .A(n9878), .ZN(n9879) );
  NAND2_X1 U12293 ( .A1(n9880), .A2(n9879), .ZN(n12370) );
  NAND2_X1 U12294 ( .A1(n10036), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U12295 ( .A1(n9881), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12296 ( .A1(n9896), .A2(n9882), .ZN(n12374) );
  NAND2_X1 U12297 ( .A1(n10063), .A2(n12374), .ZN(n9885) );
  NAND2_X1 U12298 ( .A1(n10098), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U12299 ( .A1(n10099), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9883) );
  OR2_X1 U12300 ( .A1(n12370), .A2(n12408), .ZN(n9903) );
  NAND2_X1 U12301 ( .A1(n12370), .A2(n12408), .ZN(n10132) );
  INV_X1 U12302 ( .A(n9888), .ZN(n9889) );
  XNOR2_X1 U12303 ( .A(n9890), .B(n9889), .ZN(n10545) );
  NAND2_X1 U12304 ( .A1(n9911), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9893) );
  INV_X1 U12305 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9892) );
  XNOR2_X1 U12306 ( .A(n9893), .B(n9892), .ZN(n12801) );
  OAI22_X1 U12307 ( .A1(n10033), .A2(n10546), .B1(n10941), .B2(n12801), .ZN(
        n9894) );
  AOI21_X1 U12308 ( .B1(n10545), .B2(n10076), .A(n9894), .ZN(n12404) );
  NAND2_X1 U12309 ( .A1(n10036), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9902) );
  INV_X1 U12310 ( .A(n9915), .ZN(n9898) );
  NAND2_X1 U12311 ( .A1(n9896), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U12312 ( .A1(n9898), .A2(n9897), .ZN(n12405) );
  NAND2_X1 U12313 ( .A1(n10063), .A2(n12405), .ZN(n9901) );
  NAND2_X1 U12314 ( .A1(n10099), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U12315 ( .A1(n10098), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9899) );
  NAND4_X1 U12316 ( .A1(n9902), .A2(n9901), .A3(n9900), .A4(n9899), .ZN(n12708) );
  AND2_X1 U12317 ( .A1(n12404), .A2(n12708), .ZN(n9907) );
  INV_X1 U12318 ( .A(n9903), .ZN(n9904) );
  OAI21_X1 U12319 ( .B1(n9907), .B2(n9904), .A(n10294), .ZN(n9905) );
  INV_X1 U12320 ( .A(n12404), .ZN(n13054) );
  AOI21_X1 U12321 ( .B1(n10134), .B2(n10132), .A(n10294), .ZN(n9908) );
  INV_X1 U12322 ( .A(n9907), .ZN(n10133) );
  XOR2_X1 U12323 ( .A(n9910), .B(n9909), .Z(n10796) );
  OAI21_X1 U12324 ( .B1(n9911), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9912) );
  XNOR2_X1 U12325 ( .A(n9912), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14583) );
  OAI22_X1 U12326 ( .A1(n6480), .A2(n10797), .B1(n10941), .B2(n12803), .ZN(
        n9913) );
  NAND2_X1 U12327 ( .A1(n10036), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U12328 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  OR2_X1 U12329 ( .A1(n9933), .A2(n9916), .ZN(n12995) );
  NAND2_X1 U12330 ( .A1(n10063), .A2(n12995), .ZN(n9919) );
  NAND2_X1 U12331 ( .A1(n10098), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U12332 ( .A1(n10099), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9917) );
  NAND4_X1 U12333 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), .ZN(n12707) );
  NAND2_X1 U12334 ( .A1(n13105), .A2(n12707), .ZN(n9955) );
  INV_X1 U12335 ( .A(n13105), .ZN(n12650) );
  NAND2_X1 U12336 ( .A1(n12650), .A2(n12978), .ZN(n10135) );
  NAND2_X1 U12337 ( .A1(n9955), .A2(n10135), .ZN(n12988) );
  INV_X1 U12338 ( .A(n12988), .ZN(n12993) );
  INV_X1 U12339 ( .A(n10135), .ZN(n9921) );
  AOI22_X1 U12340 ( .A1(n9922), .A2(n12993), .B1(n9921), .B2(n10294), .ZN(
        n9939) );
  INV_X1 U12341 ( .A(n9923), .ZN(n9924) );
  XNOR2_X1 U12342 ( .A(n9925), .B(n9924), .ZN(n10831) );
  NAND2_X1 U12343 ( .A1(n10831), .A2(n10076), .ZN(n9931) );
  NAND2_X1 U12344 ( .A1(n9926), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9928) );
  XNOR2_X1 U12345 ( .A(n9928), .B(n9927), .ZN(n12818) );
  OAI22_X1 U12346 ( .A1(n6480), .A2(n10832), .B1(n10941), .B2(n12818), .ZN(
        n9929) );
  INV_X1 U12347 ( .A(n9929), .ZN(n9930) );
  NAND2_X1 U12348 ( .A1(n9931), .A2(n9930), .ZN(n12683) );
  NAND2_X1 U12349 ( .A1(n10036), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9938) );
  OR2_X1 U12350 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  NAND2_X1 U12351 ( .A1(n9949), .A2(n9934), .ZN(n12982) );
  NAND2_X1 U12352 ( .A1(n10063), .A2(n12982), .ZN(n9937) );
  NAND2_X1 U12353 ( .A1(n10098), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U12354 ( .A1(n10099), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9935) );
  NAND2_X1 U12355 ( .A1(n12683), .A2(n12991), .ZN(n9957) );
  NAND2_X1 U12356 ( .A1(n10136), .A2(n9957), .ZN(n10243) );
  NOR2_X1 U12357 ( .A1(n9939), .A2(n10243), .ZN(n9971) );
  INV_X1 U12358 ( .A(n9957), .ZN(n9956) );
  INV_X1 U12359 ( .A(n9940), .ZN(n9941) );
  XNOR2_X1 U12360 ( .A(n9942), .B(n9941), .ZN(n11030) );
  NAND2_X1 U12361 ( .A1(n11030), .A2(n10076), .ZN(n9948) );
  NAND2_X1 U12362 ( .A1(n9943), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9945) );
  XNOR2_X2 U12363 ( .A(n9945), .B(n9944), .ZN(n12822) );
  OAI22_X1 U12364 ( .A1(n10033), .A2(n11032), .B1(n12822), .B2(n10941), .ZN(
        n9946) );
  INV_X1 U12365 ( .A(n9946), .ZN(n9947) );
  NAND2_X1 U12366 ( .A1(n9949), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12367 ( .A1(n9963), .A2(n9950), .ZN(n12969) );
  NAND2_X1 U12368 ( .A1(n10063), .A2(n12969), .ZN(n9954) );
  NAND2_X1 U12369 ( .A1(n10036), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U12370 ( .A1(n10099), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12371 ( .A1(n10098), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9951) );
  OR2_X1 U12372 ( .A1(n13095), .A2(n12979), .ZN(n10138) );
  OAI211_X1 U12373 ( .C1(n9956), .C2(n9955), .A(n10138), .B(n10136), .ZN(n9959) );
  NAND2_X1 U12374 ( .A1(n13095), .A2(n12979), .ZN(n10139) );
  NAND2_X1 U12375 ( .A1(n10139), .A2(n9957), .ZN(n9958) );
  MUX2_X1 U12376 ( .A(n9959), .B(n9958), .S(n10294), .Z(n9970) );
  XNOR2_X1 U12377 ( .A(n9960), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U12378 ( .A1(n11335), .A2(n10076), .ZN(n9962) );
  OR2_X1 U12379 ( .A1(n6480), .A2(n11336), .ZN(n9961) );
  AND2_X1 U12380 ( .A1(n9963), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9964) );
  OR2_X1 U12381 ( .A1(n9964), .A2(n9978), .ZN(n12945) );
  NAND2_X1 U12382 ( .A1(n12945), .A2(n10063), .ZN(n9968) );
  NAND2_X1 U12383 ( .A1(n10098), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U12384 ( .A1(n10036), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U12385 ( .A1(n10099), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9965) );
  NAND4_X1 U12386 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n12961) );
  NAND2_X1 U12387 ( .A1(n13092), .A2(n12961), .ZN(n10140) );
  NAND2_X1 U12388 ( .A1(n12950), .A2(n12934), .ZN(n9985) );
  MUX2_X1 U12389 ( .A(n10139), .B(n10138), .S(n10294), .Z(n9969) );
  OAI211_X1 U12390 ( .C1(n9971), .C2(n9970), .A(n10176), .B(n9969), .ZN(n9987)
         );
  INV_X1 U12391 ( .A(n9972), .ZN(n9973) );
  XNOR2_X1 U12392 ( .A(n9974), .B(n9973), .ZN(n11400) );
  NAND2_X1 U12393 ( .A1(n11400), .A2(n10076), .ZN(n9976) );
  OR2_X1 U12394 ( .A1(n10033), .A2(n11402), .ZN(n9975) );
  NOR2_X1 U12395 ( .A1(n9978), .A2(n9977), .ZN(n9979) );
  OR2_X1 U12396 ( .A1(n9992), .A2(n9979), .ZN(n12937) );
  NAND2_X1 U12397 ( .A1(n12937), .A2(n10063), .ZN(n9984) );
  NAND2_X1 U12398 ( .A1(n10036), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12399 ( .A1(n10099), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9980) );
  AND2_X1 U12400 ( .A1(n9981), .A2(n9980), .ZN(n9983) );
  NAND2_X1 U12401 ( .A1(n10098), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12402 ( .A1(n12625), .A2(n12944), .ZN(n10141) );
  MUX2_X1 U12403 ( .A(n10140), .B(n9985), .S(n10294), .Z(n9986) );
  NAND3_X1 U12404 ( .A1(n9987), .A2(n12936), .A3(n9986), .ZN(n9999) );
  XNOR2_X1 U12405 ( .A(n9989), .B(n9988), .ZN(n11444) );
  NAND2_X1 U12406 ( .A1(n11444), .A2(n10076), .ZN(n9991) );
  OR2_X1 U12407 ( .A1(n6480), .A2(n7184), .ZN(n9990) );
  NOR2_X1 U12408 ( .A1(n9992), .A2(n12674), .ZN(n9993) );
  OR2_X1 U12409 ( .A1(n9994), .A2(n9993), .ZN(n12924) );
  NAND2_X1 U12410 ( .A1(n12924), .A2(n10063), .ZN(n9997) );
  AOI22_X1 U12411 ( .A1(n10036), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n10098), 
        .B2(P3_REG0_REG_22__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U12412 ( .A1(n10099), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U12413 ( .A1(n12675), .A2(n12933), .ZN(n10144) );
  MUX2_X1 U12414 ( .A(n10141), .B(n10142), .S(n10294), .Z(n9998) );
  NAND3_X1 U12415 ( .A1(n9999), .A2(n12923), .A3(n9998), .ZN(n10001) );
  XNOR2_X1 U12416 ( .A(n12603), .B(n12659), .ZN(n12907) );
  INV_X1 U12417 ( .A(n12907), .ZN(n12902) );
  MUX2_X1 U12418 ( .A(n10145), .B(n10144), .S(n10294), .Z(n10000) );
  INV_X1 U12419 ( .A(n12603), .ZN(n13080) );
  NOR3_X1 U12420 ( .A1(n13080), .A2(n10294), .A3(n12704), .ZN(n10002) );
  NAND2_X1 U12421 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n10005), .ZN(n10006) );
  INV_X1 U12422 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13782) );
  INV_X1 U12423 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U12424 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13782), .B2(n14526), .ZN(n10007) );
  XNOR2_X1 U12425 ( .A(n10020), .B(n10007), .ZN(n12166) );
  NAND2_X1 U12426 ( .A1(n12166), .A2(n10076), .ZN(n10009) );
  OR2_X1 U12427 ( .A1(n10033), .A2(n12169), .ZN(n10008) );
  NAND2_X1 U12428 ( .A1(n10036), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n10015) );
  INV_X1 U12429 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12641) );
  NAND2_X1 U12430 ( .A1(n10010), .A2(n12641), .ZN(n10023) );
  OR2_X1 U12431 ( .A1(n10010), .A2(n12641), .ZN(n10011) );
  NAND2_X1 U12432 ( .A1(n10023), .A2(n10011), .ZN(n12881) );
  NAND2_X1 U12433 ( .A1(n10063), .A2(n12881), .ZN(n10014) );
  NAND2_X1 U12434 ( .A1(n10098), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U12435 ( .A1(n10099), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n10012) );
  NAND3_X1 U12436 ( .A1(n12479), .A2(n12865), .A3(n10294), .ZN(n10017) );
  INV_X1 U12437 ( .A(n12865), .ZN(n12703) );
  NAND3_X1 U12438 ( .A1(n13075), .A2(n10939), .A3(n12703), .ZN(n10016) );
  NAND2_X1 U12439 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13782), .ZN(n10019) );
  AOI22_X1 U12440 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13777), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14519), .ZN(n10029) );
  XNOR2_X1 U12441 ( .A(n10030), .B(n10029), .ZN(n12252) );
  NAND2_X1 U12442 ( .A1(n12252), .A2(n10076), .ZN(n10022) );
  OR2_X1 U12443 ( .A1(n6480), .A2(n8689), .ZN(n10021) );
  NAND2_X1 U12444 ( .A1(n10036), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n10028) );
  NAND2_X1 U12445 ( .A1(n10023), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U12446 ( .A1(n10037), .A2(n10024), .ZN(n12869) );
  NAND2_X1 U12447 ( .A1(n10063), .A2(n12869), .ZN(n10027) );
  NAND2_X1 U12448 ( .A1(n10098), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U12449 ( .A1(n10099), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n10025) );
  NAND4_X1 U12450 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n12702) );
  NOR2_X1 U12451 ( .A1(n13071), .A2(n12702), .ZN(n10150) );
  INV_X1 U12452 ( .A(n13071), .ZN(n10251) );
  NOR2_X1 U12453 ( .A1(n10251), .A2(n10252), .ZN(n10151) );
  NOR2_X1 U12454 ( .A1(n10150), .A2(n10151), .ZN(n12868) );
  MUX2_X1 U12455 ( .A(n10151), .B(n10150), .S(n10294), .Z(n10043) );
  NAND2_X1 U12456 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  AOI22_X1 U12457 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13775), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14518), .ZN(n10032) );
  XNOR2_X1 U12458 ( .A(n10045), .B(n10032), .ZN(n12446) );
  NAND2_X1 U12459 ( .A1(n12446), .A2(n10076), .ZN(n10035) );
  NAND2_X1 U12460 ( .A1(n10036), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n10042) );
  AND2_X1 U12461 ( .A1(n10037), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12462 ( .A1(n10063), .A2(n12858), .ZN(n10041) );
  NAND2_X1 U12463 ( .A1(n10099), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U12464 ( .A1(n10098), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U12465 ( .A1(n12857), .A2(n12866), .ZN(n10153) );
  OAI21_X1 U12466 ( .B1(n12857), .B2(n12866), .A(n10153), .ZN(n10152) );
  AOI211_X1 U12467 ( .C1(n10044), .C2(n12868), .A(n10043), .B(n10152), .ZN(
        n10069) );
  NOR3_X1 U12468 ( .A1(n12857), .A2(n10939), .A3(n12866), .ZN(n10068) );
  NOR2_X1 U12469 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n14518), .ZN(n10046) );
  INV_X1 U12470 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10054) );
  NAND2_X1 U12471 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n10054), .ZN(n10048) );
  INV_X1 U12472 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12426) );
  INV_X1 U12473 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13767) );
  INV_X1 U12474 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14515) );
  AOI22_X1 U12475 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13767), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14515), .ZN(n10072) );
  XNOR2_X1 U12476 ( .A(n10075), .B(n10072), .ZN(n13120) );
  NAND2_X1 U12477 ( .A1(n13120), .A2(n10076), .ZN(n10050) );
  OR2_X1 U12478 ( .A1(n6480), .A2(n13124), .ZN(n10049) );
  NAND2_X1 U12479 ( .A1(n10050), .A2(n10049), .ZN(n10300) );
  NAND2_X1 U12480 ( .A1(n10063), .A2(n14604), .ZN(n10103) );
  NAND2_X1 U12481 ( .A1(n10036), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U12482 ( .A1(n10099), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U12483 ( .A1(n10098), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U12484 ( .A1(n10300), .A2(n12837), .ZN(n10157) );
  AOI22_X1 U12485 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n10054), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n12426), .ZN(n10055) );
  INV_X1 U12486 ( .A(n10055), .ZN(n10056) );
  XNOR2_X1 U12487 ( .A(n10057), .B(n10056), .ZN(n13126) );
  NAND2_X1 U12488 ( .A1(n13126), .A2(n10076), .ZN(n10060) );
  OR2_X1 U12489 ( .A1(n10033), .A2(n13128), .ZN(n10059) );
  NAND2_X1 U12490 ( .A1(n10036), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U12491 ( .A1(n10061), .A2(n8562), .ZN(n10062) );
  NAND2_X1 U12492 ( .A1(n10063), .A2(n12844), .ZN(n10066) );
  NAND2_X1 U12493 ( .A1(n10099), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10065) );
  NAND2_X1 U12494 ( .A1(n10098), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10064) );
  NAND4_X1 U12495 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n12700) );
  OAI211_X1 U12496 ( .C1(n10069), .C2(n10068), .A(n10266), .B(n12842), .ZN(
        n10085) );
  INV_X1 U12497 ( .A(n12700), .ZN(n12596) );
  NOR2_X1 U12498 ( .A1(n13003), .A2(n12596), .ZN(n10070) );
  NAND2_X1 U12499 ( .A1(n13003), .A2(n12596), .ZN(n10154) );
  OAI21_X1 U12500 ( .B1(n10070), .B2(n10153), .A(n10154), .ZN(n10071) );
  MUX2_X1 U12501 ( .A(n10071), .B(n10070), .S(n10294), .Z(n10082) );
  INV_X1 U12502 ( .A(n10072), .ZN(n10074) );
  NAND2_X1 U12503 ( .A1(n14515), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10073) );
  INV_X1 U12504 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U12505 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n10093), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n12445), .ZN(n10091) );
  NAND2_X1 U12506 ( .A1(n12575), .A2(n10076), .ZN(n10078) );
  OR2_X1 U12507 ( .A1(n6480), .A2(n12576), .ZN(n10077) );
  NAND2_X1 U12508 ( .A1(n10098), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U12509 ( .A1(n10036), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U12510 ( .A1(n10099), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U12511 ( .A1(n14615), .A2(n11285), .ZN(n10159) );
  NAND2_X1 U12512 ( .A1(n10087), .A2(n10159), .ZN(n10179) );
  AOI21_X1 U12513 ( .B1(n10266), .B2(n10082), .A(n10179), .ZN(n10084) );
  MUX2_X1 U12514 ( .A(n10157), .B(n10155), .S(n10294), .Z(n10083) );
  INV_X1 U12515 ( .A(n10088), .ZN(n10086) );
  NAND2_X1 U12516 ( .A1(n10086), .A2(n10159), .ZN(n10090) );
  INV_X1 U12517 ( .A(n10087), .ZN(n10162) );
  NOR2_X1 U12518 ( .A1(n10088), .A2(n10162), .ZN(n10089) );
  MUX2_X1 U12519 ( .A(n10090), .B(n10089), .S(n10939), .Z(n10105) );
  INV_X1 U12520 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10544) );
  INV_X1 U12521 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U12522 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n10544), .B2(n10094), .ZN(n10095) );
  NOR2_X1 U12523 ( .A1(n6480), .A2(n13119), .ZN(n10097) );
  AOI21_X1 U12524 ( .B1(n13113), .B2(n10076), .A(n10097), .ZN(n14610) );
  NAND2_X1 U12525 ( .A1(n10098), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U12526 ( .A1(n10036), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U12527 ( .A1(n10099), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10100) );
  NAND4_X1 U12528 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n14603) );
  INV_X1 U12529 ( .A(n14603), .ZN(n10104) );
  NAND2_X1 U12530 ( .A1(n11338), .A2(n12822), .ZN(n10296) );
  INV_X1 U12531 ( .A(n15322), .ZN(n10166) );
  NAND2_X1 U12532 ( .A1(n10166), .A2(n10109), .ZN(n10582) );
  NAND2_X1 U12533 ( .A1(n10582), .A2(n10579), .ZN(n15301) );
  NAND2_X1 U12534 ( .A1(n15301), .A2(n15300), .ZN(n15299) );
  NAND2_X1 U12535 ( .A1(n15299), .A2(n10110), .ZN(n11020) );
  NAND2_X1 U12536 ( .A1(n11020), .A2(n11024), .ZN(n11019) );
  NAND2_X1 U12537 ( .A1(n11019), .A2(n10112), .ZN(n11078) );
  INV_X1 U12538 ( .A(n10221), .ZN(n11080) );
  NAND2_X1 U12539 ( .A1(n11078), .A2(n11080), .ZN(n11077) );
  NAND2_X1 U12540 ( .A1(n10117), .A2(n10116), .ZN(n11404) );
  NAND2_X1 U12541 ( .A1(n11404), .A2(n11808), .ZN(n11403) );
  NAND2_X1 U12542 ( .A1(n11403), .A2(n10118), .ZN(n11638) );
  INV_X1 U12543 ( .A(n11799), .ZN(n15358) );
  NAND2_X1 U12544 ( .A1(n12715), .A2(n15358), .ZN(n10120) );
  INV_X1 U12545 ( .A(n12715), .ZN(n11939) );
  NAND2_X1 U12546 ( .A1(n11753), .A2(n10121), .ZN(n10123) );
  NAND2_X1 U12547 ( .A1(n10123), .A2(n10122), .ZN(n11951) );
  NAND2_X1 U12548 ( .A1(n12362), .A2(n12361), .ZN(n12360) );
  NAND2_X1 U12549 ( .A1(n12360), .A2(n10134), .ZN(n12994) );
  NAND2_X1 U12550 ( .A1(n12994), .A2(n12993), .ZN(n12992) );
  NAND2_X1 U12551 ( .A1(n12992), .A2(n10135), .ZN(n12981) );
  NAND2_X1 U12552 ( .A1(n10137), .A2(n10136), .ZN(n12968) );
  NAND2_X1 U12553 ( .A1(n10138), .A2(n10139), .ZN(n12967) );
  NAND2_X1 U12554 ( .A1(n10143), .A2(n10142), .ZN(n12922) );
  NAND2_X1 U12555 ( .A1(n12922), .A2(n10144), .ZN(n10146) );
  NAND2_X1 U12556 ( .A1(n10146), .A2(n10145), .ZN(n12903) );
  NAND2_X1 U12557 ( .A1(n12903), .A2(n12902), .ZN(n12905) );
  NAND2_X1 U12558 ( .A1(n12905), .A2(n10147), .ZN(n12894) );
  INV_X1 U12559 ( .A(n12876), .ZN(n10149) );
  NAND2_X1 U12560 ( .A1(n12851), .A2(n10153), .ZN(n12843) );
  NAND2_X1 U12561 ( .A1(n12843), .A2(n12842), .ZN(n12841) );
  INV_X1 U12562 ( .A(n14615), .ZN(n10158) );
  OAI211_X1 U12563 ( .C1(n10158), .C2(n14603), .A(n10164), .B(n10157), .ZN(
        n10160) );
  INV_X1 U12564 ( .A(n11338), .ZN(n10180) );
  AND2_X1 U12565 ( .A1(n11075), .A2(n10180), .ZN(n10258) );
  NOR2_X1 U12566 ( .A1(n6584), .A2(n15323), .ZN(n10165) );
  NAND4_X1 U12567 ( .A1(n10165), .A2(n11080), .A3(n15300), .A4(n10228), .ZN(
        n10170) );
  NOR2_X1 U12568 ( .A1(n10167), .A2(n10166), .ZN(n10815) );
  NAND4_X1 U12569 ( .A1(n10815), .A2(n11808), .A3(n11642), .A4(n11024), .ZN(
        n10169) );
  NOR4_X1 U12570 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n11752), .ZN(
        n10171) );
  AND4_X1 U12571 ( .A1(n12093), .A2(n10172), .A3(n11991), .A4(n10171), .ZN(
        n10173) );
  NAND4_X1 U12572 ( .A1(n12361), .A2(n12296), .A3(n6895), .A4(n10173), .ZN(
        n10174) );
  NOR4_X1 U12573 ( .A1(n12967), .A2(n10243), .A3(n12988), .A4(n10174), .ZN(
        n10175) );
  NAND4_X1 U12574 ( .A1(n12936), .A2(n10176), .A3(n12923), .A4(n10175), .ZN(
        n10177) );
  NOR4_X1 U12575 ( .A1(n12892), .A2(n12876), .A3(n12907), .A4(n10177), .ZN(
        n10178) );
  XNOR2_X1 U12576 ( .A(n6509), .B(n12822), .ZN(n10182) );
  AOI21_X1 U12577 ( .B1(n10184), .B2(n10258), .A(n10183), .ZN(n10185) );
  INV_X1 U12578 ( .A(n10187), .ZN(n10189) );
  NAND2_X1 U12579 ( .A1(n6637), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U12580 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10190), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n10191) );
  AND2_X1 U12581 ( .A1(n10191), .A2(n10198), .ZN(n10204) );
  AND2_X1 U12582 ( .A1(n10204), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10936) );
  INV_X1 U12583 ( .A(n12254), .ZN(n10203) );
  INV_X1 U12584 ( .A(n10195), .ZN(n10200) );
  NAND2_X1 U12585 ( .A1(n10200), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10196) );
  MUX2_X1 U12586 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10196), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n10197) );
  NAND2_X1 U12587 ( .A1(n10192), .A2(n10197), .ZN(n12167) );
  NAND2_X1 U12588 ( .A1(n10198), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U12589 ( .A1(n12167), .A2(n12028), .ZN(n10202) );
  NAND2_X1 U12590 ( .A1(n10203), .A2(n10202), .ZN(n10565) );
  INV_X1 U12591 ( .A(n10204), .ZN(n10938) );
  INV_X1 U12592 ( .A(n10296), .ZN(n10596) );
  AND2_X1 U12593 ( .A1(n10939), .A2(n10596), .ZN(n10808) );
  NAND2_X1 U12594 ( .A1(n10937), .A2(n10808), .ZN(n10569) );
  INV_X1 U12595 ( .A(n10205), .ZN(n10907) );
  NOR3_X1 U12596 ( .A1(n10569), .A2(n10907), .A3(n6501), .ZN(n10208) );
  INV_X1 U12597 ( .A(n10936), .ZN(n11741) );
  OAI21_X1 U12598 ( .B1(n11445), .B2(n11741), .A(P3_B_REG_SCAN_IN), .ZN(n10207) );
  OR2_X1 U12599 ( .A1(n10209), .A2(n11089), .ZN(n15316) );
  NAND2_X1 U12600 ( .A1(n10210), .A2(n15316), .ZN(n10213) );
  NAND2_X1 U12601 ( .A1(n10211), .A2(n10212), .ZN(n10580) );
  NAND2_X1 U12602 ( .A1(n10213), .A2(n10580), .ZN(n15298) );
  NAND2_X1 U12603 ( .A1(n15298), .A2(n10214), .ZN(n10216) );
  NAND2_X1 U12604 ( .A1(n11025), .A2(n15309), .ZN(n10215) );
  NAND2_X1 U12605 ( .A1(n10216), .A2(n10215), .ZN(n11023) );
  INV_X1 U12606 ( .A(n11023), .ZN(n10218) );
  NAND2_X1 U12607 ( .A1(n10218), .A2(n10217), .ZN(n11021) );
  NAND2_X1 U12608 ( .A1(n12721), .A2(n9652), .ZN(n10220) );
  NAND2_X1 U12609 ( .A1(n11021), .A2(n10220), .ZN(n11079) );
  OR2_X1 U12610 ( .A1(n11248), .A2(n11166), .ZN(n10222) );
  NAND2_X1 U12611 ( .A1(n11803), .A2(n11449), .ZN(n10223) );
  INV_X1 U12612 ( .A(n11801), .ZN(n15185) );
  NAND2_X1 U12613 ( .A1(n12717), .A2(n15185), .ZN(n10224) );
  NAND2_X1 U12614 ( .A1(n11419), .A2(n10224), .ZN(n11407) );
  INV_X1 U12615 ( .A(n11808), .ZN(n11406) );
  OR2_X1 U12616 ( .A1(n11809), .A2(n11674), .ZN(n10225) );
  NAND2_X1 U12617 ( .A1(n11816), .A2(n15351), .ZN(n10227) );
  INV_X1 U12618 ( .A(n10228), .ZN(n11730) );
  NAND2_X1 U12619 ( .A1(n11731), .A2(n11730), .ZN(n11729) );
  NAND2_X1 U12620 ( .A1(n11729), .A2(n10229), .ZN(n11750) );
  NAND2_X1 U12621 ( .A1(n11750), .A2(n11752), .ZN(n11749) );
  OR2_X1 U12622 ( .A1(n12334), .A2(n11936), .ZN(n10230) );
  NAND2_X1 U12623 ( .A1(n11749), .A2(n10230), .ZN(n11952) );
  NAND2_X1 U12624 ( .A1(n12352), .A2(n14622), .ZN(n10231) );
  NAND2_X1 U12625 ( .A1(n11952), .A2(n10231), .ZN(n10233) );
  OR2_X1 U12626 ( .A1(n12352), .A2(n14622), .ZN(n10232) );
  NAND2_X1 U12627 ( .A1(n11988), .A2(n6981), .ZN(n10236) );
  INV_X1 U12628 ( .A(n14617), .ZN(n10234) );
  NAND2_X1 U12629 ( .A1(n10234), .A2(n12712), .ZN(n10235) );
  INV_X1 U12630 ( .A(n12711), .ZN(n12179) );
  INV_X1 U12631 ( .A(n12710), .ZN(n12283) );
  OR2_X1 U12632 ( .A1(n12330), .A2(n12283), .ZN(n10237) );
  NAND2_X1 U12633 ( .A1(n12139), .A2(n10237), .ZN(n12293) );
  OR2_X1 U12634 ( .A1(n12370), .A2(n12709), .ZN(n10238) );
  NAND2_X1 U12635 ( .A1(n12293), .A2(n10238), .ZN(n10240) );
  NAND2_X1 U12636 ( .A1(n12370), .A2(n12709), .ZN(n10239) );
  NAND2_X1 U12637 ( .A1(n10240), .A2(n10239), .ZN(n12357) );
  INV_X1 U12638 ( .A(n12361), .ZN(n10241) );
  OR2_X1 U12639 ( .A1(n12404), .A2(n12990), .ZN(n10242) );
  INV_X1 U12640 ( .A(n12976), .ZN(n10244) );
  OR2_X1 U12641 ( .A1(n12683), .A2(n12964), .ZN(n10245) );
  NAND2_X1 U12642 ( .A1(n13095), .A2(n12706), .ZN(n10246) );
  NAND2_X1 U12643 ( .A1(n12960), .A2(n10246), .ZN(n12942) );
  NAND2_X1 U12644 ( .A1(n12950), .A2(n12961), .ZN(n10247) );
  OR2_X1 U12645 ( .A1(n12625), .A2(n12705), .ZN(n10248) );
  NAND2_X1 U12646 ( .A1(n12675), .A2(n12909), .ZN(n10249) );
  INV_X1 U12647 ( .A(n13019), .ZN(n12898) );
  NAND2_X1 U12648 ( .A1(n12886), .A2(n7497), .ZN(n12877) );
  NOR2_X1 U12649 ( .A1(n12857), .A2(n12701), .ZN(n12836) );
  NOR2_X1 U12650 ( .A1(n12835), .A2(n10255), .ZN(n10257) );
  XNOR2_X1 U12651 ( .A(n10257), .B(n10256), .ZN(n10264) );
  INV_X1 U12652 ( .A(n10258), .ZN(n10259) );
  NAND2_X1 U12653 ( .A1(n11445), .A2(n10576), .ZN(n10308) );
  NAND2_X1 U12654 ( .A1(n10941), .A2(n10973), .ZN(n10260) );
  INV_X1 U12655 ( .A(P3_B_REG_SCAN_IN), .ZN(n10261) );
  NOR2_X1 U12656 ( .A1(n6501), .A2(n10261), .ZN(n10262) );
  OR2_X1 U12657 ( .A1(n15303), .A2(n10262), .ZN(n14601) );
  NAND3_X1 U12658 ( .A1(n10973), .A2(n10941), .A3(n10939), .ZN(n15302) );
  OAI22_X1 U12659 ( .A1(n11285), .A2(n14601), .B1(n12596), .B2(n15302), .ZN(
        n10263) );
  XOR2_X1 U12660 ( .A(n10266), .B(n10265), .Z(n12581) );
  AND2_X1 U12661 ( .A1(n10181), .A2(n11338), .ZN(n10292) );
  INV_X1 U12662 ( .A(n10292), .ZN(n10267) );
  XNOR2_X1 U12663 ( .A(n11445), .B(n10267), .ZN(n10269) );
  NAND2_X1 U12664 ( .A1(n10181), .A2(n12822), .ZN(n10268) );
  NAND2_X1 U12665 ( .A1(n10269), .A2(n10268), .ZN(n10588) );
  AND2_X1 U12666 ( .A1(n15357), .A2(n10596), .ZN(n10270) );
  NAND2_X1 U12667 ( .A1(n10588), .A2(n10270), .ZN(n10273) );
  NOR2_X1 U12668 ( .A1(n11338), .A2(n10576), .ZN(n10271) );
  AND2_X1 U12669 ( .A1(n11445), .A2(n10271), .ZN(n10295) );
  INV_X1 U12670 ( .A(n10295), .ZN(n10272) );
  OR2_X1 U12671 ( .A1(n15327), .A2(n11445), .ZN(n15359) );
  NAND2_X1 U12672 ( .A1(n12587), .A2(n6546), .ZN(n10313) );
  XNOR2_X1 U12673 ( .A(n12028), .B(P3_B_REG_SCAN_IN), .ZN(n10274) );
  INV_X1 U12674 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U12675 ( .A1(n10355), .A2(n10275), .ZN(n10277) );
  NAND2_X1 U12676 ( .A1(n12254), .A2(n12167), .ZN(n10276) );
  NAND2_X1 U12677 ( .A1(n10277), .A2(n10276), .ZN(n10801) );
  INV_X1 U12678 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U12679 ( .A1(n12254), .A2(n12028), .ZN(n10279) );
  NOR2_X1 U12680 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n10284) );
  NOR4_X1 U12681 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10283) );
  NOR4_X1 U12682 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n10282) );
  NOR4_X1 U12683 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10281) );
  NAND4_X1 U12684 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n10290) );
  NOR4_X1 U12685 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n10288) );
  NOR4_X1 U12686 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n10287) );
  NOR4_X1 U12687 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n10286) );
  NOR4_X1 U12688 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n10285) );
  NAND4_X1 U12689 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10289) );
  OAI21_X1 U12690 ( .B1(n10290), .B2(n10289), .A(n10355), .ZN(n10309) );
  AND2_X1 U12691 ( .A1(n10937), .A2(n10309), .ZN(n10291) );
  OAI211_X1 U12692 ( .C1(n10292), .C2(n11445), .A(n10308), .B(n10296), .ZN(
        n10293) );
  NAND2_X1 U12693 ( .A1(n10294), .A2(n10293), .ZN(n10298) );
  OR2_X1 U12694 ( .A1(n10939), .A2(n10295), .ZN(n10802) );
  NAND2_X1 U12695 ( .A1(n10939), .A2(n10296), .ZN(n10803) );
  NAND2_X1 U12696 ( .A1(n10802), .A2(n10803), .ZN(n10297) );
  AOI22_X1 U12697 ( .A1(n10801), .A2(n10298), .B1(n10574), .B2(n10297), .ZN(
        n10299) );
  NAND2_X1 U12698 ( .A1(n10313), .A2(n15374), .ZN(n10305) );
  INV_X1 U12699 ( .A(n10300), .ZN(n12583) );
  INV_X1 U12700 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10302) );
  NOR2_X1 U12701 ( .A1(n15374), .A2(n10302), .ZN(n10303) );
  NAND2_X1 U12702 ( .A1(n10305), .A2(n10304), .ZN(P3_U3488) );
  INV_X1 U12703 ( .A(n10306), .ZN(n10307) );
  NAND2_X1 U12704 ( .A1(n10307), .A2(n10309), .ZN(n10599) );
  NOR2_X1 U12705 ( .A1(n7354), .A2(n10308), .ZN(n10589) );
  NOR2_X1 U12706 ( .A1(n10589), .A2(n10808), .ZN(n10311) );
  INV_X1 U12707 ( .A(n10588), .ZN(n10310) );
  NAND3_X1 U12708 ( .A1(n10801), .A2(n10574), .A3(n10309), .ZN(n10598) );
  OAI22_X1 U12709 ( .A1(n10599), .A2(n10311), .B1(n10310), .B2(n10598), .ZN(
        n10312) );
  NAND2_X1 U12710 ( .A1(n10313), .A2(n15365), .ZN(n10317) );
  INV_X1 U12711 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U12712 ( .A1(n10314), .A2(n7477), .ZN(n10316) );
  NAND2_X1 U12713 ( .A1(n10317), .A2(n10316), .ZN(P3_U3456) );
  NAND2_X1 U12714 ( .A1(n10865), .A2(n10858), .ZN(n10318) );
  NAND2_X1 U12715 ( .A1(n10850), .A2(n10335), .ZN(n10860) );
  INV_X2 U12716 ( .A(n14393), .ZN(n14377) );
  NOR2_X2 U12717 ( .A1(n10325), .A2(n10846), .ZN(n14397) );
  NOR2_X1 U12718 ( .A1(n10887), .A2(n11743), .ZN(n10324) );
  OAI22_X1 U12719 ( .A1(n10327), .A2(n14386), .B1(n10326), .B2(n10325), .ZN(
        n10328) );
  AOI21_X1 U12720 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14377), .A(n10328), 
        .ZN(n10329) );
  OAI21_X1 U12721 ( .B1(n6799), .B2(n14394), .A(n10329), .ZN(n10330) );
  AOI21_X1 U12722 ( .B1(n10331), .B2(n14397), .A(n10330), .ZN(n10332) );
  INV_X1 U12723 ( .A(n10333), .ZN(n10334) );
  INV_X1 U12724 ( .A(n10336), .ZN(n10337) );
  OR2_X1 U12725 ( .A1(n10683), .A2(n10337), .ZN(n12419) );
  INV_X2 U12726 ( .A(n12419), .ZN(P2_U3947) );
  AND2_X1 U12727 ( .A1(n9592), .A2(P2_U3088), .ZN(n12187) );
  INV_X2 U12728 ( .A(n12187), .ZN(n13781) );
  AND2_X1 U12729 ( .A1(n10344), .A2(P2_U3088), .ZN(n13770) );
  AOI22_X1 U12730 ( .A1(n13770), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n14958), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10338) );
  OAI21_X1 U12731 ( .B1(n10349), .B2(n13781), .A(n10338), .ZN(P2_U3325) );
  INV_X1 U12732 ( .A(n14090), .ZN(n10339) );
  NAND2_X1 U12733 ( .A1(n10344), .A2(P1_U3086), .ZN(n14521) );
  INV_X1 U12734 ( .A(n14521), .ZN(n12191) );
  INV_X1 U12735 ( .A(n12191), .ZN(n14525) );
  OAI222_X1 U12736 ( .A1(P1_U3086), .A2(n10339), .B1(n14525), .B2(n12424), 
        .C1(n7503), .C2(n14527), .ZN(P1_U3354) );
  INV_X1 U12737 ( .A(n14120), .ZN(n10340) );
  OAI222_X1 U12738 ( .A1(n14527), .A2(n6723), .B1(n14525), .B2(n10341), .C1(
        n10340), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X2 U12739 ( .A(n13770), .ZN(n13783) );
  OAI222_X1 U12740 ( .A1(n13783), .A2(n10342), .B1(n13781), .B2(n10341), .C1(
        n13272), .C2(P2_U3088), .ZN(P2_U3324) );
  OAI222_X1 U12741 ( .A1(n13783), .A2(n10343), .B1(n13781), .B2(n10351), .C1(
        n13286), .C2(P2_U3088), .ZN(P2_U3323) );
  NAND2_X1 U12742 ( .A1(n10344), .A2(P3_U3151), .ZN(n13130) );
  OAI222_X1 U12743 ( .A1(n13130), .A2(n10347), .B1(n13125), .B2(n10346), .C1(
        n15284), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U12744 ( .A(n14113), .ZN(n10348) );
  OAI222_X1 U12745 ( .A1(n14527), .A2(n10350), .B1(n14521), .B2(n10349), .C1(
        n10348), .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U12746 ( .A1(n14527), .A2(n6711), .B1(n14521), .B2(n10351), .C1(
        n14774), .C2(P1_U3086), .ZN(P1_U3351) );
  NAND2_X1 U12747 ( .A1(n10354), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10352) );
  OAI21_X1 U12748 ( .B1(n10801), .B2(n10354), .A(n10352), .ZN(P3_U3377) );
  NAND2_X1 U12749 ( .A1(n10354), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10353) );
  OAI21_X1 U12750 ( .B1(n10574), .B2(n10354), .A(n10353), .ZN(P3_U3376) );
  INV_X1 U12751 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U12752 ( .A1(n10419), .A2(n10356), .ZN(P3_U3258) );
  INV_X1 U12753 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10357) );
  NOR2_X1 U12754 ( .A1(n10419), .A2(n10357), .ZN(P3_U3248) );
  INV_X1 U12755 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10358) );
  NOR2_X1 U12756 ( .A1(n10419), .A2(n10358), .ZN(P3_U3247) );
  INV_X1 U12757 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10359) );
  NOR2_X1 U12758 ( .A1(n10419), .A2(n10359), .ZN(P3_U3250) );
  INV_X1 U12759 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10360) );
  NOR2_X1 U12760 ( .A1(n10419), .A2(n10360), .ZN(P3_U3261) );
  INV_X1 U12761 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10361) );
  NOR2_X1 U12762 ( .A1(n10419), .A2(n10361), .ZN(P3_U3249) );
  INV_X1 U12763 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10362) );
  NOR2_X1 U12764 ( .A1(n10419), .A2(n10362), .ZN(P3_U3246) );
  INV_X1 U12765 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10363) );
  NOR2_X1 U12766 ( .A1(n10419), .A2(n10363), .ZN(P3_U3259) );
  INV_X1 U12767 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10364) );
  NOR2_X1 U12768 ( .A1(n10419), .A2(n10364), .ZN(P3_U3253) );
  INV_X1 U12769 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10365) );
  NOR2_X1 U12770 ( .A1(n10419), .A2(n10365), .ZN(P3_U3251) );
  INV_X1 U12771 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10366) );
  NOR2_X1 U12772 ( .A1(n10419), .A2(n10366), .ZN(P3_U3260) );
  INV_X1 U12773 ( .A(n10629), .ZN(n10777) );
  INV_X1 U12774 ( .A(n10367), .ZN(n10369) );
  INV_X1 U12775 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10368) );
  OAI222_X1 U12776 ( .A1(P1_U3086), .A2(n10777), .B1(n14521), .B2(n10369), 
        .C1(n10368), .C2(n14527), .ZN(P1_U3350) );
  INV_X1 U12777 ( .A(n10469), .ZN(n13300) );
  OAI222_X1 U12778 ( .A1(n13783), .A2(n10370), .B1(n13781), .B2(n10369), .C1(
        n13300), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U12779 ( .A(n13130), .ZN(n13112) );
  INV_X1 U12780 ( .A(n10371), .ZN(n10373) );
  OAI222_X1 U12781 ( .A1(n13123), .A2(n10373), .B1(n13125), .B2(n10372), .C1(
        n15256), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12782 ( .A(SI_7_), .ZN(n10374) );
  OAI222_X1 U12783 ( .A1(n13123), .A2(n10375), .B1(n13125), .B2(n10374), .C1(
        n11520), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12784 ( .A(SI_10_), .ZN(n10376) );
  OAI222_X1 U12785 ( .A1(n13123), .A2(n10377), .B1(n13125), .B2(n10376), .C1(
        n11830), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U12786 ( .A1(n13123), .A2(n10379), .B1(n12007), .B2(P3_U3151), 
        .C1(n13125), .C2(n10378), .ZN(P3_U3284) );
  INV_X1 U12787 ( .A(n10650), .ZN(n10645) );
  OAI222_X1 U12788 ( .A1(n14527), .A2(n10380), .B1(n14521), .B2(n10382), .C1(
        n10645), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12789 ( .A(n10488), .ZN(n10381) );
  OAI222_X1 U12790 ( .A1(n13783), .A2(n10383), .B1(n13781), .B2(n10382), .C1(
        n10381), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12791 ( .A(n10962), .ZN(n15206) );
  INV_X1 U12792 ( .A(SI_3_), .ZN(n10384) );
  OAI222_X1 U12793 ( .A1(n15206), .A2(P3_U3151), .B1(n13123), .B2(n10385), 
        .C1(n10384), .C2(n13125), .ZN(P3_U3292) );
  INV_X1 U12794 ( .A(n10386), .ZN(n10388) );
  OAI222_X1 U12795 ( .A1(n11095), .A2(P3_U3151), .B1(n13123), .B2(n10388), 
        .C1(n10387), .C2(n13125), .ZN(P3_U3289) );
  INV_X1 U12796 ( .A(n10961), .ZN(n11001) );
  OAI222_X1 U12797 ( .A1(n11001), .A2(P3_U3151), .B1(n13123), .B2(n10390), 
        .C1(n10389), .C2(n13125), .ZN(P3_U3293) );
  INV_X1 U12798 ( .A(n10965), .ZN(n15223) );
  INV_X1 U12799 ( .A(SI_4_), .ZN(n10391) );
  OAI222_X1 U12800 ( .A1(n15223), .A2(P3_U3151), .B1(n13123), .B2(n10392), 
        .C1(n10391), .C2(n13125), .ZN(P3_U3291) );
  INV_X1 U12801 ( .A(n10393), .ZN(n10395) );
  OAI222_X1 U12802 ( .A1(n10943), .A2(P3_U3151), .B1(n13123), .B2(n10395), 
        .C1(n10394), .C2(n13125), .ZN(P3_U3295) );
  OAI222_X1 U12803 ( .A1(n15240), .A2(P3_U3151), .B1(n13123), .B2(n10397), 
        .C1(n10396), .C2(n13125), .ZN(P3_U3290) );
  INV_X1 U12804 ( .A(n10398), .ZN(n10399) );
  INV_X1 U12805 ( .A(n10400), .ZN(n10402) );
  OAI222_X1 U12806 ( .A1(n13123), .A2(n10402), .B1(n12263), .B2(P3_U3151), 
        .C1(n10401), .C2(n13125), .ZN(P3_U3283) );
  INV_X1 U12807 ( .A(n10652), .ZN(n10743) );
  OAI222_X1 U12808 ( .A1(n14527), .A2(n10403), .B1(n14525), .B2(n10404), .C1(
        n10743), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12809 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10405) );
  INV_X1 U12810 ( .A(n10500), .ZN(n10456) );
  OAI222_X1 U12811 ( .A1(n13783), .A2(n10405), .B1(n13781), .B2(n10404), .C1(
        n10456), .C2(P2_U3088), .ZN(P2_U3320) );
  AND2_X2 U12812 ( .A1(n10407), .A2(n10406), .ZN(n14844) );
  INV_X1 U12813 ( .A(n10408), .ZN(n10409) );
  OAI22_X1 U12814 ( .A1(n14844), .A2(P1_D_REG_0__SCAN_IN), .B1(n10413), .B2(
        n10409), .ZN(n10410) );
  INV_X1 U12815 ( .A(n10410), .ZN(P1_U3445) );
  INV_X1 U12816 ( .A(n10411), .ZN(n10412) );
  OAI22_X1 U12817 ( .A1(n14844), .A2(P1_D_REG_1__SCAN_IN), .B1(n10413), .B2(
        n10412), .ZN(n10414) );
  INV_X1 U12818 ( .A(n10414), .ZN(P1_U3446) );
  INV_X1 U12819 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10415) );
  OAI222_X1 U12820 ( .A1(n13783), .A2(n10415), .B1(n13781), .B2(n10416), .C1(
        n10507), .C2(P2_U3088), .ZN(P2_U3319) );
  OAI222_X1 U12821 ( .A1(n14527), .A2(n10417), .B1(n14525), .B2(n10416), .C1(
        n10748), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U12822 ( .A(n14527), .ZN(n14509) );
  AOI22_X1 U12823 ( .A1(n14138), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14509), .ZN(n10418) );
  OAI21_X1 U12824 ( .B1(n10442), .B2(n14521), .A(n10418), .ZN(P1_U3346) );
  CLKBUF_X1 U12825 ( .A(n10419), .Z(n10439) );
  INV_X1 U12826 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10420) );
  NOR2_X1 U12827 ( .A1(n10439), .A2(n10420), .ZN(P3_U3255) );
  INV_X1 U12828 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10421) );
  NOR2_X1 U12829 ( .A1(n10439), .A2(n10421), .ZN(P3_U3262) );
  INV_X1 U12830 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10422) );
  NOR2_X1 U12831 ( .A1(n10439), .A2(n10422), .ZN(P3_U3237) );
  INV_X1 U12832 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10423) );
  NOR2_X1 U12833 ( .A1(n10439), .A2(n10423), .ZN(P3_U3254) );
  INV_X1 U12834 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10424) );
  NOR2_X1 U12835 ( .A1(n10439), .A2(n10424), .ZN(P3_U3263) );
  INV_X1 U12836 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10425) );
  NOR2_X1 U12837 ( .A1(n10439), .A2(n10425), .ZN(P3_U3252) );
  INV_X1 U12838 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10426) );
  NOR2_X1 U12839 ( .A1(n10439), .A2(n10426), .ZN(P3_U3257) );
  INV_X1 U12840 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10427) );
  NOR2_X1 U12841 ( .A1(n10439), .A2(n10427), .ZN(P3_U3256) );
  INV_X1 U12842 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10428) );
  NOR2_X1 U12843 ( .A1(n10439), .A2(n10428), .ZN(P3_U3245) );
  INV_X1 U12844 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10429) );
  NOR2_X1 U12845 ( .A1(n10439), .A2(n10429), .ZN(P3_U3244) );
  INV_X1 U12846 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10430) );
  NOR2_X1 U12847 ( .A1(n10439), .A2(n10430), .ZN(P3_U3243) );
  INV_X1 U12848 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10431) );
  NOR2_X1 U12849 ( .A1(n10439), .A2(n10431), .ZN(P3_U3242) );
  INV_X1 U12850 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10432) );
  NOR2_X1 U12851 ( .A1(n10439), .A2(n10432), .ZN(P3_U3241) );
  INV_X1 U12852 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10433) );
  NOR2_X1 U12853 ( .A1(n10439), .A2(n10433), .ZN(P3_U3240) );
  INV_X1 U12854 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10434) );
  NOR2_X1 U12855 ( .A1(n10439), .A2(n10434), .ZN(P3_U3239) );
  INV_X1 U12856 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10435) );
  NOR2_X1 U12857 ( .A1(n10439), .A2(n10435), .ZN(P3_U3238) );
  INV_X1 U12858 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10436) );
  NOR2_X1 U12859 ( .A1(n10439), .A2(n10436), .ZN(P3_U3236) );
  INV_X1 U12860 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10437) );
  NOR2_X1 U12861 ( .A1(n10439), .A2(n10437), .ZN(P3_U3235) );
  INV_X1 U12862 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10438) );
  NOR2_X1 U12863 ( .A1(n10439), .A2(n10438), .ZN(P3_U3234) );
  OAI222_X1 U12864 ( .A1(n12732), .A2(P3_U3151), .B1(n13123), .B2(n10441), 
        .C1(n10440), .C2(n13125), .ZN(P3_U3282) );
  INV_X1 U12865 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10443) );
  INV_X1 U12866 ( .A(n14978), .ZN(n10532) );
  OAI222_X1 U12867 ( .A1(n13783), .A2(n10443), .B1(n13781), .B2(n10442), .C1(
        n10532), .C2(P2_U3088), .ZN(P2_U3318) );
  INV_X1 U12868 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10444) );
  MUX2_X1 U12869 ( .A(n10444), .B(P2_REG2_REG_1__SCAN_IN), .S(n14944), .Z(
        n14951) );
  NAND2_X1 U12870 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n14950) );
  NOR2_X1 U12871 ( .A1(n14951), .A2(n14950), .ZN(n14949) );
  AOI21_X1 U12872 ( .B1(n14944), .B2(P2_REG2_REG_1__SCAN_IN), .A(n14949), .ZN(
        n14963) );
  MUX2_X1 U12873 ( .A(n8856), .B(P2_REG2_REG_2__SCAN_IN), .S(n14958), .Z(
        n14962) );
  OR2_X1 U12874 ( .A1(n14963), .A2(n14962), .ZN(n14965) );
  NAND2_X1 U12875 ( .A1(n14958), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13279) );
  MUX2_X1 U12876 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10445), .S(n13272), .Z(
        n13278) );
  NOR2_X1 U12877 ( .A1(n13272), .A2(n10445), .ZN(n13293) );
  MUX2_X1 U12878 ( .A(n11266), .B(P2_REG2_REG_4__SCAN_IN), .S(n13286), .Z(
        n13292) );
  INV_X1 U12879 ( .A(n13286), .ZN(n10446) );
  NAND2_X1 U12880 ( .A1(n10446), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13308) );
  MUX2_X1 U12881 ( .A(n11302), .B(P2_REG2_REG_5__SCAN_IN), .S(n10469), .Z(
        n13307) );
  AOI21_X1 U12882 ( .B1(n13309), .B2(n13308), .A(n13307), .ZN(n13306) );
  NOR2_X1 U12883 ( .A1(n13300), .A2(n11302), .ZN(n10483) );
  MUX2_X1 U12884 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11289), .S(n10488), .Z(
        n10482) );
  OAI21_X1 U12885 ( .B1(n13306), .B2(n10483), .A(n10482), .ZN(n10481) );
  NAND2_X1 U12886 ( .A1(n10488), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U12887 ( .A(n11323), .B(P2_REG2_REG_7__SCAN_IN), .S(n10500), .Z(
        n10447) );
  AOI21_X1 U12888 ( .B1(n10481), .B2(n10448), .A(n10447), .ZN(n10494) );
  NAND3_X1 U12889 ( .A1(n10481), .A2(n10448), .A3(n10447), .ZN(n10453) );
  OAI21_X1 U12890 ( .B1(n10677), .B2(n10449), .A(n8875), .ZN(n10452) );
  INV_X1 U12891 ( .A(n10683), .ZN(n10450) );
  NAND2_X1 U12892 ( .A1(n10450), .A2(n10682), .ZN(n10451) );
  NAND2_X1 U12893 ( .A1(n10452), .A2(n10451), .ZN(n10455) );
  NOR2_X1 U12894 ( .A1(n9258), .A2(P2_U3088), .ZN(n13769) );
  AND2_X1 U12895 ( .A1(n10455), .A2(n13769), .ZN(n10473) );
  AND2_X1 U12896 ( .A1(n10473), .A2(n10474), .ZN(n15033) );
  NAND2_X1 U12897 ( .A1(n10453), .A2(n15033), .ZN(n10480) );
  NAND2_X1 U12898 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11069) );
  INV_X1 U12899 ( .A(n11069), .ZN(n10458) );
  AND2_X1 U12900 ( .A1(n9258), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10454) );
  NOR2_X1 U12901 ( .A1(n15048), .A2(n10456), .ZN(n10457) );
  AOI211_X1 U12902 ( .C1(n15051), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10458), .B(
        n10457), .ZN(n10479) );
  INV_X1 U12903 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10459) );
  MUX2_X1 U12904 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10459), .S(n10500), .Z(
        n10477) );
  INV_X1 U12905 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10460) );
  XNOR2_X1 U12906 ( .A(n14944), .B(n10460), .ZN(n14941) );
  AND2_X1 U12907 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14940) );
  NAND2_X1 U12908 ( .A1(n14941), .A2(n14940), .ZN(n14939) );
  NAND2_X1 U12909 ( .A1(n14944), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U12910 ( .A1(n14939), .A2(n10461), .ZN(n14956) );
  XNOR2_X1 U12911 ( .A(n14958), .B(n10462), .ZN(n14957) );
  NAND2_X1 U12912 ( .A1(n14956), .A2(n14957), .ZN(n14955) );
  NAND2_X1 U12913 ( .A1(n14958), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U12914 ( .A1(n14955), .A2(n10463), .ZN(n13276) );
  XNOR2_X1 U12915 ( .A(n13272), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n13277) );
  NAND2_X1 U12916 ( .A1(n13276), .A2(n13277), .ZN(n13275) );
  OR2_X1 U12917 ( .A1(n13272), .A2(n10464), .ZN(n10465) );
  NAND2_X1 U12918 ( .A1(n13275), .A2(n10465), .ZN(n13290) );
  XNOR2_X1 U12919 ( .A(n13286), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n13291) );
  NAND2_X1 U12920 ( .A1(n13290), .A2(n13291), .ZN(n13289) );
  OR2_X1 U12921 ( .A1(n13286), .A2(n10466), .ZN(n10467) );
  NAND2_X1 U12922 ( .A1(n13289), .A2(n10467), .ZN(n13304) );
  XNOR2_X1 U12923 ( .A(n10469), .B(n10468), .ZN(n13305) );
  NAND2_X1 U12924 ( .A1(n13304), .A2(n13305), .ZN(n13303) );
  NAND2_X1 U12925 ( .A1(n10469), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U12926 ( .A1(n13303), .A2(n10470), .ZN(n10490) );
  INV_X1 U12927 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10471) );
  MUX2_X1 U12928 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10471), .S(n10488), .Z(
        n10491) );
  NAND2_X1 U12929 ( .A1(n10490), .A2(n10491), .ZN(n10489) );
  NAND2_X1 U12930 ( .A1(n10488), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U12931 ( .A1(n10489), .A2(n10472), .ZN(n10476) );
  INV_X1 U12932 ( .A(n10473), .ZN(n10475) );
  NAND2_X1 U12933 ( .A1(n10476), .A2(n10477), .ZN(n10502) );
  OAI211_X1 U12934 ( .C1(n10477), .C2(n10476), .A(n15021), .B(n10502), .ZN(
        n10478) );
  OAI211_X1 U12935 ( .C1(n10494), .C2(n10480), .A(n10479), .B(n10478), .ZN(
        P2_U3221) );
  NAND2_X1 U12936 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10880) );
  OAI21_X1 U12937 ( .B1(n15039), .B2(n8513), .A(n10880), .ZN(n10487) );
  INV_X1 U12938 ( .A(n10481), .ZN(n10485) );
  NOR3_X1 U12939 ( .A1(n13306), .A2(n10483), .A3(n10482), .ZN(n10484) );
  NOR3_X1 U12940 ( .A1(n15053), .A2(n10485), .A3(n10484), .ZN(n10486) );
  AOI211_X1 U12941 ( .C1(n15027), .C2(n10488), .A(n10487), .B(n10486), .ZN(
        n10493) );
  OAI211_X1 U12942 ( .C1(n10491), .C2(n10490), .A(n15021), .B(n10489), .ZN(
        n10492) );
  NAND2_X1 U12943 ( .A1(n10493), .A2(n10492), .ZN(P2_U3220) );
  NAND2_X1 U12944 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11194) );
  AOI21_X1 U12945 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10500), .A(n10494), .ZN(
        n10496) );
  MUX2_X1 U12946 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11392), .S(n10507), .Z(
        n10495) );
  NOR2_X1 U12947 ( .A1(n10496), .A2(n10495), .ZN(n10524) );
  AOI211_X1 U12948 ( .C1(n10496), .C2(n10495), .A(n15053), .B(n10524), .ZN(
        n10497) );
  INV_X1 U12949 ( .A(n10497), .ZN(n10498) );
  OAI211_X1 U12950 ( .C1(n14548), .C2(n15039), .A(n11194), .B(n10498), .ZN(
        n10499) );
  INV_X1 U12951 ( .A(n10499), .ZN(n10506) );
  MUX2_X1 U12952 ( .A(n8945), .B(P2_REG1_REG_8__SCAN_IN), .S(n10507), .Z(
        n10504) );
  NAND2_X1 U12953 ( .A1(n10500), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U12954 ( .A1(n10502), .A2(n10501), .ZN(n10503) );
  NAND2_X1 U12955 ( .A1(n10503), .A2(n10504), .ZN(n10530) );
  OAI211_X1 U12956 ( .C1(n10504), .C2(n10503), .A(n15021), .B(n10530), .ZN(
        n10505) );
  OAI211_X1 U12957 ( .C1(n15048), .C2(n10507), .A(n10506), .B(n10505), .ZN(
        P2_U3222) );
  INV_X1 U12958 ( .A(n12735), .ZN(n12756) );
  OAI222_X1 U12959 ( .A1(n13123), .A2(n10508), .B1(n13125), .B2(n7197), .C1(
        n12756), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12960 ( .A(n10509), .ZN(n10515) );
  AOI22_X1 U12961 ( .A1(n10785), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14509), .ZN(n10510) );
  OAI21_X1 U12962 ( .B1(n10515), .B2(n14521), .A(n10510), .ZN(P1_U3345) );
  OR2_X1 U12963 ( .A1(n10861), .A2(n10511), .ZN(n10513) );
  NAND2_X1 U12964 ( .A1(n10513), .A2(n10512), .ZN(n10604) );
  AND2_X1 U12965 ( .A1(n10860), .A2(n12193), .ZN(n10603) );
  INV_X1 U12966 ( .A(n10603), .ZN(n10514) );
  AND2_X1 U12967 ( .A1(n10604), .A2(n10514), .ZN(n14757) );
  NOR2_X1 U12968 ( .A1(n14757), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12969 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10516) );
  INV_X1 U12970 ( .A(n10554), .ZN(n10539) );
  OAI222_X1 U12971 ( .A1(n13783), .A2(n10516), .B1(n13781), .B2(n10515), .C1(
        P2_U3088), .C2(n10539), .ZN(P2_U3317) );
  INV_X1 U12972 ( .A(n10517), .ZN(n10519) );
  INV_X1 U12973 ( .A(n11126), .ZN(n11138) );
  OAI222_X1 U12974 ( .A1(n14527), .A2(n10518), .B1(n14525), .B2(n10519), .C1(
        P1_U3086), .C2(n11138), .ZN(P1_U3344) );
  INV_X1 U12975 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10520) );
  INV_X1 U12976 ( .A(n13323), .ZN(n13315) );
  OAI222_X1 U12977 ( .A1(n13783), .A2(n10520), .B1(n13781), .B2(n10519), .C1(
        P2_U3088), .C2(n13315), .ZN(P2_U3316) );
  INV_X1 U12978 ( .A(n10521), .ZN(n10523) );
  OAI222_X1 U12979 ( .A1(n13130), .A2(n10523), .B1(n13125), .B2(n10522), .C1(
        n12798), .C2(P3_U3151), .ZN(P3_U3280) );
  AOI21_X1 U12980 ( .B1(n10528), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10524), .ZN(
        n14971) );
  MUX2_X1 U12981 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11490), .S(n14978), .Z(
        n14970) );
  NAND2_X1 U12982 ( .A1(n14971), .A2(n14970), .ZN(n14969) );
  OAI21_X1 U12983 ( .B1(n14978), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14969), .ZN(
        n10526) );
  MUX2_X1 U12984 ( .A(n11618), .B(P2_REG2_REG_10__SCAN_IN), .S(n10554), .Z(
        n10525) );
  NOR2_X1 U12985 ( .A1(n10526), .A2(n10525), .ZN(n10548) );
  AOI211_X1 U12986 ( .C1(n10526), .C2(n10525), .A(n15053), .B(n10548), .ZN(
        n10542) );
  MUX2_X1 U12987 ( .A(n10527), .B(P2_REG1_REG_10__SCAN_IN), .S(n10554), .Z(
        n10536) );
  NAND2_X1 U12988 ( .A1(n10528), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U12989 ( .A1(n10530), .A2(n10529), .ZN(n14974) );
  MUX2_X1 U12990 ( .A(n10531), .B(P2_REG1_REG_9__SCAN_IN), .S(n14978), .Z(
        n14973) );
  OR2_X1 U12991 ( .A1(n14974), .A2(n14973), .ZN(n14976) );
  NAND2_X1 U12992 ( .A1(n10532), .A2(n10531), .ZN(n10533) );
  NAND2_X1 U12993 ( .A1(n14976), .A2(n10533), .ZN(n10535) );
  OR2_X1 U12994 ( .A1(n10535), .A2(n10536), .ZN(n10556) );
  INV_X1 U12995 ( .A(n10556), .ZN(n10534) );
  AOI211_X1 U12996 ( .C1(n10536), .C2(n10535), .A(n15042), .B(n10534), .ZN(
        n10541) );
  NOR2_X1 U12997 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11438), .ZN(n10537) );
  AOI21_X1 U12998 ( .B1(n15051), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10537), 
        .ZN(n10538) );
  OAI21_X1 U12999 ( .B1(n10539), .B2(n15048), .A(n10538), .ZN(n10540) );
  OR3_X1 U13000 ( .A1(n10542), .A2(n10541), .A3(n10540), .ZN(P2_U3224) );
  NAND2_X1 U13001 ( .A1(n14179), .A2(n14102), .ZN(n10543) );
  OAI21_X1 U13002 ( .B1(P1_U4016), .B2(n10544), .A(n10543), .ZN(P1_U3591) );
  INV_X1 U13003 ( .A(n10545), .ZN(n10547) );
  OAI222_X1 U13004 ( .A1(n13123), .A2(n10547), .B1(n13125), .B2(n10546), .C1(
        n12801), .C2(P3_U3151), .ZN(P3_U3279) );
  AOI21_X1 U13005 ( .B1(n10554), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10548), 
        .ZN(n10550) );
  MUX2_X1 U13006 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n8985), .S(n13323), .Z(
        n10549) );
  NAND2_X1 U13007 ( .A1(n10550), .A2(n10549), .ZN(n14989) );
  OAI21_X1 U13008 ( .B1(n10550), .B2(n10549), .A(n14989), .ZN(n10553) );
  AND2_X1 U13009 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11671) );
  AOI21_X1 U13010 ( .B1(n15051), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n11671), 
        .ZN(n10551) );
  OAI21_X1 U13011 ( .B1(n13315), .B2(n15048), .A(n10551), .ZN(n10552) );
  AOI21_X1 U13012 ( .B1(n10553), .B2(n15033), .A(n10552), .ZN(n10560) );
  NAND2_X1 U13013 ( .A1(n10554), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U13014 ( .A1(n10556), .A2(n10555), .ZN(n10558) );
  MUX2_X1 U13015 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8989), .S(n13323), .Z(
        n10557) );
  NAND2_X1 U13016 ( .A1(n10558), .A2(n10557), .ZN(n13325) );
  OAI211_X1 U13017 ( .C1(n10558), .C2(n10557), .A(n13325), .B(n15021), .ZN(
        n10559) );
  NAND2_X1 U13018 ( .A1(n10560), .A2(n10559), .ZN(P2_U3225) );
  INV_X1 U13019 ( .A(n14788), .ZN(n11132) );
  INV_X1 U13020 ( .A(n10561), .ZN(n10562) );
  OAI222_X1 U13021 ( .A1(P1_U3086), .A2(n11132), .B1(n14525), .B2(n10562), 
        .C1(n9561), .C2(n14527), .ZN(P1_U3343) );
  INV_X1 U13022 ( .A(n14994), .ZN(n13317) );
  OAI222_X1 U13023 ( .A1(n13783), .A2(n10563), .B1(n13781), .B2(n10562), .C1(
        n13317), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U13024 ( .A1(n13168), .A2(P2_U3947), .ZN(n10564) );
  OAI21_X1 U13025 ( .B1(P2_U3947), .B2(n7565), .A(n10564), .ZN(P2_U3553) );
  NAND2_X1 U13026 ( .A1(n10599), .A2(n10588), .ZN(n10568) );
  NAND2_X1 U13027 ( .A1(n10565), .A2(n10803), .ZN(n10566) );
  AOI21_X1 U13028 ( .B1(n10598), .B2(n10589), .A(n10566), .ZN(n10567) );
  NAND2_X1 U13029 ( .A1(n10568), .A2(n10567), .ZN(n10572) );
  INV_X1 U13030 ( .A(n10569), .ZN(n10570) );
  AND2_X1 U13031 ( .A1(n10598), .A2(n10570), .ZN(n10571) );
  AOI21_X1 U13032 ( .B1(n10572), .B2(P3_STATE_REG_SCAN_IN), .A(n10571), .ZN(
        n11155) );
  AND2_X1 U13033 ( .A1(n11155), .A2(n10573), .ZN(n10841) );
  INV_X1 U13034 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13035 ( .A1(n10181), .A2(n10576), .ZN(n10577) );
  NAND2_X1 U13036 ( .A1(n10577), .A2(n11338), .ZN(n10578) );
  NAND2_X1 U13037 ( .A1(n15316), .A2(n11800), .ZN(n10583) );
  NAND3_X1 U13038 ( .A1(n12723), .A2(n11800), .A3(n15326), .ZN(n10581) );
  INV_X1 U13039 ( .A(n10584), .ZN(n10587) );
  NAND3_X1 U13040 ( .A1(n15323), .A2(n15322), .A3(n12485), .ZN(n10586) );
  OAI21_X1 U13041 ( .B1(n10587), .B2(n15316), .A(n10586), .ZN(n10593) );
  NAND2_X1 U13042 ( .A1(n10588), .A2(n15357), .ZN(n10591) );
  INV_X1 U13043 ( .A(n10589), .ZN(n10590) );
  OAI22_X1 U13044 ( .A1(n10599), .A2(n10591), .B1(n10590), .B2(n10598), .ZN(
        n10592) );
  OAI21_X1 U13045 ( .B1(n10840), .B2(n10593), .A(n15180), .ZN(n10602) );
  OR2_X1 U13046 ( .A1(n10209), .A2(n15302), .ZN(n10595) );
  OR2_X1 U13047 ( .A1(n11025), .A2(n15303), .ZN(n10594) );
  NAND2_X1 U13048 ( .A1(n10595), .A2(n10594), .ZN(n15319) );
  NAND2_X1 U13049 ( .A1(n10937), .A2(n10596), .ZN(n10597) );
  INV_X1 U13050 ( .A(n15189), .ZN(n15178) );
  NAND2_X1 U13051 ( .A1(n10599), .A2(n15327), .ZN(n10600) );
  AOI22_X1 U13052 ( .A1(n15319), .A2(n15178), .B1(n15186), .B2(n15326), .ZN(
        n10601) );
  OAI211_X1 U13053 ( .C1(n10841), .C2(n11007), .A(n10602), .B(n10601), .ZN(
        P3_U3162) );
  INV_X1 U13054 ( .A(n14516), .ZN(n14749) );
  NAND2_X1 U13055 ( .A1(n14101), .A2(n14749), .ZN(n10605) );
  NOR2_X2 U13056 ( .A1(n14760), .A2(n10605), .ZN(n14771) );
  INV_X1 U13057 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10606) );
  MUX2_X1 U13058 ( .A(n10606), .B(P1_REG2_REG_4__SCAN_IN), .S(n14774), .Z(
        n10614) );
  INV_X1 U13059 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10607) );
  MUX2_X1 U13060 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10607), .S(n14120), .Z(
        n14122) );
  INV_X1 U13061 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10608) );
  XNOR2_X1 U13062 ( .A(n14113), .B(n10608), .ZN(n14109) );
  AND2_X1 U13063 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10609) );
  NAND2_X1 U13064 ( .A1(n14090), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10610) );
  OAI211_X1 U13065 ( .C1(n14090), .C2(P1_REG2_REG_1__SCAN_IN), .A(n10609), .B(
        n10610), .ZN(n14091) );
  NAND2_X1 U13066 ( .A1(n14091), .A2(n10610), .ZN(n14107) );
  NAND2_X1 U13067 ( .A1(n14109), .A2(n14107), .ZN(n10612) );
  NAND2_X1 U13068 ( .A1(n14113), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13069 ( .A1(n10612), .A2(n10611), .ZN(n14121) );
  NAND2_X1 U13070 ( .A1(n14122), .A2(n14121), .ZN(n14767) );
  NAND2_X1 U13071 ( .A1(n14120), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U13072 ( .A1(n14767), .A2(n14766), .ZN(n10613) );
  NAND2_X1 U13073 ( .A1(n10614), .A2(n10613), .ZN(n14770) );
  INV_X1 U13074 ( .A(n14770), .ZN(n10769) );
  NOR2_X1 U13075 ( .A1(n14774), .A2(n10606), .ZN(n10768) );
  INV_X1 U13076 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11464) );
  MUX2_X1 U13077 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11464), .S(n10629), .Z(
        n10767) );
  OAI21_X1 U13078 ( .B1(n10769), .B2(n10768), .A(n10767), .ZN(n10766) );
  NAND2_X1 U13079 ( .A1(n10629), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10617) );
  INV_X1 U13080 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10615) );
  MUX2_X1 U13081 ( .A(n10615), .B(P1_REG2_REG_6__SCAN_IN), .S(n10650), .Z(
        n10616) );
  AOI21_X1 U13082 ( .B1(n10766), .B2(n10617), .A(n10616), .ZN(n10739) );
  AND3_X1 U13083 ( .A1(n10766), .A2(n10617), .A3(n10616), .ZN(n10618) );
  NOR3_X1 U13084 ( .A1(n14807), .A2(n10739), .A3(n10618), .ZN(n10633) );
  INV_X1 U13085 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10619) );
  MUX2_X1 U13086 ( .A(n10619), .B(P1_REG1_REG_6__SCAN_IN), .S(n10650), .Z(
        n10631) );
  INV_X1 U13087 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11636) );
  MUX2_X1 U13088 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n11636), .S(n14120), .Z(
        n14118) );
  INV_X1 U13089 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10620) );
  XNOR2_X1 U13090 ( .A(n14090), .B(n10620), .ZN(n14089) );
  AND2_X1 U13091 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14088) );
  NAND2_X1 U13092 ( .A1(n14089), .A2(n14088), .ZN(n14087) );
  NAND2_X1 U13093 ( .A1(n14090), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U13094 ( .A1(n14087), .A2(n10621), .ZN(n14105) );
  INV_X1 U13095 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10622) );
  XNOR2_X1 U13096 ( .A(n14113), .B(n10622), .ZN(n14106) );
  NAND2_X1 U13097 ( .A1(n14105), .A2(n14106), .ZN(n14104) );
  NAND2_X1 U13098 ( .A1(n14113), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10623) );
  NAND2_X1 U13099 ( .A1(n14104), .A2(n10623), .ZN(n14117) );
  NAND2_X1 U13100 ( .A1(n14120), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U13101 ( .A1(n14761), .A2(n14762), .ZN(n10626) );
  INV_X1 U13102 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10624) );
  MUX2_X1 U13103 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10624), .S(n14774), .Z(
        n14763) );
  INV_X1 U13104 ( .A(n14763), .ZN(n10625) );
  NAND2_X1 U13105 ( .A1(n10626), .A2(n10625), .ZN(n14765) );
  INV_X1 U13106 ( .A(n14765), .ZN(n10627) );
  XOR2_X1 U13107 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10629), .Z(n10765) );
  NAND2_X1 U13108 ( .A1(n10764), .A2(n10765), .ZN(n10763) );
  OAI21_X1 U13109 ( .B1(n10629), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10763), .ZN(
        n10630) );
  NOR2_X1 U13110 ( .A1(n10630), .A2(n10631), .ZN(n10649) );
  AOI211_X1 U13111 ( .C1(n10631), .C2(n10630), .A(n10649), .B(n14168), .ZN(
        n10632) );
  NOR2_X1 U13112 ( .A1(n10633), .A2(n10632), .ZN(n10636) );
  NAND2_X1 U13113 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11852) );
  INV_X1 U13114 ( .A(n11852), .ZN(n10634) );
  AOI21_X1 U13115 ( .B1(n14757), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10634), .ZN(
        n10635) );
  OAI211_X1 U13116 ( .C1(n10645), .C2(n14775), .A(n10636), .B(n10635), .ZN(
        P1_U3249) );
  XNOR2_X1 U13117 ( .A(n10638), .B(n10637), .ZN(n11243) );
  AOI21_X1 U13118 ( .B1(n9219), .B2(n15123), .A(n11243), .ZN(n10643) );
  AOI22_X1 U13119 ( .A1(n13612), .A2(n13269), .B1(n13268), .B2(n13614), .ZN(
        n10732) );
  OAI21_X1 U13120 ( .B1(n10640), .B2(n13593), .A(n10732), .ZN(n11236) );
  OAI211_X1 U13121 ( .C1(n11275), .C2(n10641), .A(n11228), .B(n6483), .ZN(
        n11238) );
  OAI21_X1 U13122 ( .B1(n10641), .B2(n15140), .A(n11238), .ZN(n10642) );
  NOR3_X1 U13123 ( .A1(n10643), .A2(n11236), .A3(n10642), .ZN(n15107) );
  NAND2_X1 U13124 ( .A1(n15154), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10644) );
  OAI21_X1 U13125 ( .B1(n15107), .B2(n15154), .A(n10644), .ZN(P2_U3501) );
  NOR2_X1 U13126 ( .A1(n10645), .A2(n10615), .ZN(n10738) );
  INV_X1 U13127 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11502) );
  MUX2_X1 U13128 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11502), .S(n10652), .Z(
        n10737) );
  OAI21_X1 U13129 ( .B1(n10739), .B2(n10738), .A(n10737), .ZN(n10736) );
  NAND2_X1 U13130 ( .A1(n10652), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10647) );
  INV_X1 U13131 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10747) );
  MUX2_X1 U13132 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10747), .S(n10748), .Z(
        n10646) );
  AOI21_X1 U13133 ( .B1(n10736), .B2(n10647), .A(n10646), .ZN(n14137) );
  NAND3_X1 U13134 ( .A1(n10736), .A2(n10647), .A3(n10646), .ZN(n10648) );
  NAND2_X1 U13135 ( .A1(n14771), .A2(n10648), .ZN(n10661) );
  INV_X1 U13136 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10651) );
  MUX2_X1 U13137 ( .A(n10651), .B(P1_REG1_REG_7__SCAN_IN), .S(n10652), .Z(
        n10734) );
  NOR2_X1 U13138 ( .A1(n10735), .A2(n10734), .ZN(n10733) );
  INV_X1 U13139 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10653) );
  MUX2_X1 U13140 ( .A(n10653), .B(P1_REG1_REG_8__SCAN_IN), .S(n10748), .Z(
        n10654) );
  NAND2_X1 U13141 ( .A1(n10655), .A2(n10654), .ZN(n10752) );
  OAI21_X1 U13142 ( .B1(n10655), .B2(n10654), .A(n10752), .ZN(n10656) );
  INV_X1 U13143 ( .A(n14168), .ZN(n14801) );
  NAND2_X1 U13144 ( .A1(n10656), .A2(n14801), .ZN(n10660) );
  NAND2_X1 U13145 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12073) );
  INV_X1 U13146 ( .A(n12073), .ZN(n10658) );
  NOR2_X1 U13147 ( .A1(n14775), .A2(n10748), .ZN(n10657) );
  AOI211_X1 U13148 ( .C1(n14757), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10658), .B(
        n10657), .ZN(n10659) );
  OAI211_X1 U13149 ( .C1(n14137), .C2(n10661), .A(n10660), .B(n10659), .ZN(
        P1_U3251) );
  NAND2_X2 U13150 ( .A1(n10662), .A2(n11206), .ZN(n10879) );
  OAI21_X1 U13151 ( .B1(n12547), .B2(n11276), .A(n10709), .ZN(n10719) );
  NAND2_X1 U13152 ( .A1(n10719), .A2(n10720), .ZN(n10718) );
  NAND2_X1 U13153 ( .A1(n10718), .A2(n10667), .ZN(n10726) );
  XNOR2_X1 U13154 ( .A(n6477), .B(n10879), .ZN(n10670) );
  NOR2_X1 U13155 ( .A1(n10673), .A2(n10672), .ZN(n10727) );
  NAND2_X1 U13156 ( .A1(n10726), .A2(n10727), .ZN(n10725) );
  INV_X1 U13157 ( .A(n10673), .ZN(n10674) );
  XOR2_X1 U13158 ( .A(n10694), .B(n10695), .Z(n10697) );
  XNOR2_X1 U13159 ( .A(n10698), .B(n10697), .ZN(n10693) );
  NAND3_X1 U13160 ( .A1(n10675), .A2(n11203), .A3(n11202), .ZN(n10681) );
  INV_X1 U13161 ( .A(n10681), .ZN(n10676) );
  NAND2_X1 U13162 ( .A1(n10676), .A2(n15090), .ZN(n10686) );
  NAND2_X1 U13163 ( .A1(n15140), .A2(n10677), .ZN(n10678) );
  INV_X1 U13164 ( .A(n13267), .ZN(n10826) );
  INV_X1 U13165 ( .A(n13614), .ZN(n13537) );
  OAI22_X1 U13166 ( .A1(n6671), .A2(n13539), .B1(n10826), .B2(n13537), .ZN(
        n11222) );
  INV_X1 U13167 ( .A(n10686), .ZN(n10680) );
  AND2_X1 U13168 ( .A1(n10680), .A2(n10679), .ZN(n13249) );
  NAND2_X1 U13169 ( .A1(n10681), .A2(n10687), .ZN(n10685) );
  AND3_X1 U13170 ( .A1(n11201), .A2(n10683), .A3(n10682), .ZN(n10684) );
  NAND2_X1 U13171 ( .A1(n10685), .A2(n10684), .ZN(n10712) );
  NOR2_X1 U13172 ( .A1(n14934), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10691) );
  OR2_X1 U13173 ( .A1(n11208), .A2(n8803), .ZN(n11229) );
  OR2_X1 U13174 ( .A1(n10686), .A2(n11229), .ZN(n10689) );
  INV_X1 U13175 ( .A(n10687), .ZN(n10688) );
  INV_X1 U13176 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13271) );
  OAI22_X1 U13177 ( .A1(n13252), .A2(n6921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13271), .ZN(n10690) );
  AOI211_X1 U13178 ( .C1(n11222), .C2(n13249), .A(n10691), .B(n10690), .ZN(
        n10692) );
  OAI21_X1 U13179 ( .B1(n10693), .B2(n14926), .A(n10692), .ZN(P2_U3190) );
  INV_X1 U13180 ( .A(n10694), .ZN(n10696) );
  XNOR2_X1 U13181 ( .A(n11268), .B(n12547), .ZN(n10700) );
  NAND2_X1 U13182 ( .A1(n13267), .A2(n12562), .ZN(n10699) );
  NAND2_X1 U13183 ( .A1(n10700), .A2(n10699), .ZN(n10819) );
  OAI21_X1 U13184 ( .B1(n10700), .B2(n10699), .A(n10819), .ZN(n10701) );
  AOI21_X1 U13185 ( .B1(n10702), .B2(n10701), .A(n6469), .ZN(n10708) );
  INV_X1 U13186 ( .A(n13268), .ZN(n10704) );
  OAI22_X1 U13187 ( .A1(n10704), .A2(n13539), .B1(n10703), .B2(n13537), .ZN(
        n11264) );
  NOR2_X1 U13188 ( .A1(n14934), .A2(n11269), .ZN(n10706) );
  NAND2_X1 U13189 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n13285) );
  OAI21_X1 U13190 ( .B1(n13252), .B2(n15118), .A(n13285), .ZN(n10705) );
  AOI211_X1 U13191 ( .C1(n11264), .C2(n13249), .A(n10706), .B(n10705), .ZN(
        n10707) );
  OAI21_X1 U13192 ( .B1(n10708), .B2(n14926), .A(n10707), .ZN(P2_U3202) );
  NAND2_X1 U13193 ( .A1(n13249), .A2(n13614), .ZN(n14920) );
  INV_X1 U13194 ( .A(n10709), .ZN(n10711) );
  NOR3_X1 U13195 ( .A1(n10715), .A2(n11276), .A3(n6483), .ZN(n10710) );
  OAI21_X1 U13196 ( .B1(n10711), .B2(n10710), .A(n13243), .ZN(n10714) );
  OR2_X1 U13197 ( .A1(n10712), .A2(P2_U3088), .ZN(n10729) );
  AOI22_X1 U13198 ( .A1(n14930), .A2(n11276), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n10729), .ZN(n10713) );
  OAI211_X1 U13199 ( .C1(n11216), .C2(n14920), .A(n10714), .B(n10713), .ZN(
        P2_U3204) );
  NAND2_X1 U13200 ( .A1(n10668), .A2(n13614), .ZN(n10717) );
  OR2_X1 U13201 ( .A1(n10715), .A2(n13539), .ZN(n10716) );
  NAND2_X1 U13202 ( .A1(n10717), .A2(n10716), .ZN(n11280) );
  INV_X1 U13203 ( .A(n11280), .ZN(n10724) );
  INV_X1 U13204 ( .A(n13249), .ZN(n11070) );
  OAI21_X1 U13205 ( .B1(n10720), .B2(n10719), .A(n10718), .ZN(n10721) );
  NAND2_X1 U13206 ( .A1(n10721), .A2(n13243), .ZN(n10723) );
  AOI22_X1 U13207 ( .A1(n14930), .A2(n10663), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n10729), .ZN(n10722) );
  OAI211_X1 U13208 ( .C1(n10724), .C2(n11070), .A(n10723), .B(n10722), .ZN(
        P2_U3194) );
  OAI21_X1 U13209 ( .B1(n10727), .B2(n10726), .A(n10725), .ZN(n10728) );
  NAND2_X1 U13210 ( .A1(n10728), .A2(n13243), .ZN(n10731) );
  AOI22_X1 U13211 ( .A1(n14930), .A2(n6477), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n10729), .ZN(n10730) );
  OAI211_X1 U13212 ( .C1(n10732), .C2(n11070), .A(n10731), .B(n10730), .ZN(
        P2_U3209) );
  AOI211_X1 U13213 ( .C1(n10735), .C2(n10734), .A(n14168), .B(n10733), .ZN(
        n10746) );
  INV_X1 U13214 ( .A(n10736), .ZN(n10741) );
  NOR3_X1 U13215 ( .A1(n10739), .A2(n10738), .A3(n10737), .ZN(n10740) );
  NOR3_X1 U13216 ( .A1(n14807), .A2(n10741), .A3(n10740), .ZN(n10745) );
  NAND2_X1 U13217 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U13218 ( .A1(n14757), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10742) );
  OAI211_X1 U13219 ( .C1(n14775), .C2(n10743), .A(n12081), .B(n10742), .ZN(
        n10744) );
  OR3_X1 U13220 ( .A1(n10746), .A2(n10745), .A3(n10744), .ZN(P1_U3250) );
  NOR2_X1 U13221 ( .A1(n10748), .A2(n10747), .ZN(n14132) );
  INV_X1 U13222 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10749) );
  MUX2_X1 U13223 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10749), .S(n14138), .Z(
        n10750) );
  OAI21_X1 U13224 ( .B1(n14137), .B2(n14132), .A(n10750), .ZN(n14135) );
  NAND2_X1 U13225 ( .A1(n14138), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10782) );
  INV_X1 U13226 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10751) );
  MUX2_X1 U13227 ( .A(n10751), .B(P1_REG2_REG_10__SCAN_IN), .S(n10785), .Z(
        n10781) );
  AOI21_X1 U13228 ( .B1(n14135), .B2(n10782), .A(n10781), .ZN(n10784) );
  AOI21_X1 U13229 ( .B1(n10785), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10784), 
        .ZN(n11135) );
  INV_X1 U13230 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11137) );
  MUX2_X1 U13231 ( .A(n11137), .B(P1_REG2_REG_11__SCAN_IN), .S(n11126), .Z(
        n11134) );
  XNOR2_X1 U13232 ( .A(n11135), .B(n11134), .ZN(n10762) );
  OAI21_X1 U13233 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10753), .A(n10752), .ZN(
        n14128) );
  MUX2_X1 U13234 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14914), .S(n14138), .Z(
        n14129) );
  NAND2_X1 U13235 ( .A1(n14128), .A2(n14129), .ZN(n14127) );
  OAI21_X1 U13236 ( .B1(n14138), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14127), .ZN(
        n10779) );
  INV_X1 U13237 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10754) );
  MUX2_X1 U13238 ( .A(n10754), .B(P1_REG1_REG_10__SCAN_IN), .S(n10785), .Z(
        n10780) );
  NOR2_X1 U13239 ( .A1(n10779), .A2(n10780), .ZN(n10778) );
  INV_X1 U13240 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10755) );
  MUX2_X1 U13241 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10755), .S(n11126), .Z(
        n10756) );
  NAND2_X1 U13242 ( .A1(n10757), .A2(n10756), .ZN(n11125) );
  OAI21_X1 U13243 ( .B1(n10757), .B2(n10756), .A(n11125), .ZN(n10758) );
  NAND2_X1 U13244 ( .A1(n10758), .A2(n14801), .ZN(n10761) );
  AND2_X1 U13245 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12313) );
  NOR2_X1 U13246 ( .A1(n14775), .A2(n11138), .ZN(n10759) );
  AOI211_X1 U13247 ( .C1(n14757), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n12313), 
        .B(n10759), .ZN(n10760) );
  OAI211_X1 U13248 ( .C1(n14807), .C2(n10762), .A(n10761), .B(n10760), .ZN(
        P1_U3254) );
  OAI21_X1 U13249 ( .B1(n10765), .B2(n10764), .A(n10763), .ZN(n10773) );
  INV_X1 U13250 ( .A(n10766), .ZN(n10771) );
  NOR3_X1 U13251 ( .A1(n10769), .A2(n10768), .A3(n10767), .ZN(n10770) );
  NOR3_X1 U13252 ( .A1(n14807), .A2(n10771), .A3(n10770), .ZN(n10772) );
  AOI21_X1 U13253 ( .B1(n14801), .B2(n10773), .A(n10772), .ZN(n10776) );
  NAND2_X1 U13254 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11602) );
  INV_X1 U13255 ( .A(n11602), .ZN(n10774) );
  AOI21_X1 U13256 ( .B1(n14757), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10774), .ZN(
        n10775) );
  OAI211_X1 U13257 ( .C1(n10777), .C2(n14775), .A(n10776), .B(n10775), .ZN(
        P1_U3248) );
  AOI211_X1 U13258 ( .C1(n10780), .C2(n10779), .A(n14168), .B(n10778), .ZN(
        n10791) );
  AND3_X1 U13259 ( .A1(n14135), .A2(n10782), .A3(n10781), .ZN(n10783) );
  NOR3_X1 U13260 ( .A1(n10784), .A2(n10783), .A3(n14807), .ZN(n10790) );
  INV_X1 U13261 ( .A(n10785), .ZN(n10788) );
  NOR2_X1 U13262 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10786), .ZN(n12207) );
  AOI21_X1 U13263 ( .B1(n14757), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n12207), 
        .ZN(n10787) );
  OAI21_X1 U13264 ( .B1(n14775), .B2(n10788), .A(n10787), .ZN(n10789) );
  OR3_X1 U13265 ( .A1(n10791), .A2(n10790), .A3(n10789), .ZN(P1_U3253) );
  INV_X1 U13266 ( .A(n10792), .ZN(n10794) );
  INV_X1 U13267 ( .A(n13343), .ZN(n13318) );
  OAI222_X1 U13268 ( .A1(n13783), .A2(n6774), .B1(n13781), .B2(n10794), .C1(
        n13318), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13269 ( .A(n11775), .ZN(n10793) );
  OAI222_X1 U13270 ( .A1(n14527), .A2(n10795), .B1(n14525), .B2(n10794), .C1(
        n10793), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13271 ( .A(n10796), .ZN(n10798) );
  OAI222_X1 U13272 ( .A1(n13123), .A2(n10798), .B1(n13125), .B2(n10797), .C1(
        n12803), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13273 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10957) );
  AND2_X2 U13274 ( .A1(n10799), .A2(n15311), .ZN(n15331) );
  INV_X1 U13275 ( .A(n10802), .ZN(n10800) );
  NAND2_X1 U13276 ( .A1(n10801), .A2(n10800), .ZN(n10805) );
  NAND2_X1 U13277 ( .A1(n10574), .A2(n10802), .ZN(n10804) );
  AND3_X1 U13278 ( .A1(n10805), .A2(n10804), .A3(n10803), .ZN(n10806) );
  INV_X1 U13279 ( .A(n10808), .ZN(n10809) );
  NAND2_X1 U13280 ( .A1(n10809), .A2(n15357), .ZN(n10810) );
  OAI22_X1 U13281 ( .A1(n10815), .A2(n10810), .B1(n10211), .B2(n15303), .ZN(
        n11091) );
  NAND2_X1 U13282 ( .A1(n11091), .A2(n15334), .ZN(n10814) );
  NAND2_X1 U13283 ( .A1(n15325), .A2(n15327), .ZN(n10811) );
  INV_X1 U13284 ( .A(n12997), .ZN(n14607) );
  AOI22_X1 U13285 ( .A1(n14607), .A2(n10812), .B1(n15331), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10813) );
  OAI211_X1 U13286 ( .C1(n10957), .C2(n15334), .A(n10814), .B(n10813), .ZN(
        P3_U3233) );
  INV_X1 U13287 ( .A(n10815), .ZN(n10817) );
  INV_X1 U13288 ( .A(n15186), .ZN(n15170) );
  NOR2_X2 U13289 ( .A1(n15189), .A2(n15303), .ZN(n12692) );
  INV_X1 U13290 ( .A(n12692), .ZN(n11817) );
  OAI22_X1 U13291 ( .A1(n15170), .A2(n11089), .B1(n11817), .B2(n10211), .ZN(
        n10816) );
  AOI21_X1 U13292 ( .B1(n10817), .B2(n15180), .A(n10816), .ZN(n10818) );
  OAI21_X1 U13293 ( .B1(n10841), .B2(n11365), .A(n10818), .ZN(P3_U3172) );
  XNOR2_X1 U13294 ( .A(n11306), .B(n12547), .ZN(n10822) );
  NAND2_X1 U13295 ( .A1(n13266), .A2(n12562), .ZN(n10821) );
  NAND2_X1 U13296 ( .A1(n10822), .A2(n10821), .ZN(n10876) );
  OAI21_X1 U13297 ( .B1(n10822), .B2(n10821), .A(n10876), .ZN(n10823) );
  AOI21_X1 U13298 ( .B1(n10824), .B2(n10823), .A(n10878), .ZN(n10830) );
  OAI22_X1 U13299 ( .A1(n10826), .A2(n13539), .B1(n10825), .B2(n13537), .ZN(
        n11300) );
  NAND2_X1 U13300 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n13299) );
  INV_X1 U13301 ( .A(n14934), .ZN(n13235) );
  NAND2_X1 U13302 ( .A1(n13235), .A2(n11307), .ZN(n10827) );
  OAI211_X1 U13303 ( .C1(n15127), .C2(n13252), .A(n13299), .B(n10827), .ZN(
        n10828) );
  AOI21_X1 U13304 ( .B1(n11300), .B2(n13249), .A(n10828), .ZN(n10829) );
  OAI21_X1 U13305 ( .B1(n10830), .B2(n14926), .A(n10829), .ZN(P2_U3199) );
  INV_X1 U13306 ( .A(n10831), .ZN(n10833) );
  OAI222_X1 U13307 ( .A1(n13123), .A2(n10833), .B1(n13125), .B2(n10832), .C1(
        n12818), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13308 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10834) );
  OAI22_X1 U13309 ( .A1(n13110), .A2(n11089), .B1(n15365), .B2(n10834), .ZN(
        n10835) );
  AOI21_X1 U13310 ( .B1(n11091), .B2(n15365), .A(n10835), .ZN(n10836) );
  INV_X1 U13311 ( .A(n10836), .ZN(P3_U3390) );
  XNOR2_X1 U13312 ( .A(n10837), .B(n10585), .ZN(n11157) );
  XNOR2_X1 U13313 ( .A(n11157), .B(n11025), .ZN(n11159) );
  INV_X1 U13314 ( .A(n10838), .ZN(n10839) );
  XOR2_X1 U13315 ( .A(n11159), .B(n11160), .Z(n10845) );
  NAND2_X1 U13316 ( .A1(n15178), .A2(n12963), .ZN(n12694) );
  INV_X1 U13317 ( .A(n12694), .ZN(n12619) );
  INV_X1 U13318 ( .A(n12721), .ZN(n15304) );
  OAI22_X1 U13319 ( .A1(n15170), .A2(n15309), .B1(n11817), .B2(n15304), .ZN(
        n10843) );
  NOR2_X1 U13320 ( .A1(n10841), .A2(n10984), .ZN(n10842) );
  AOI211_X1 U13321 ( .C1(n12619), .C2(n12723), .A(n10843), .B(n10842), .ZN(
        n10844) );
  OAI21_X1 U13322 ( .B1(n10845), .B2(n15172), .A(n10844), .ZN(P3_U3177) );
  AND2_X4 U13323 ( .A1(n10848), .A2(n10850), .ZN(n13935) );
  AND2_X4 U13324 ( .A1(n10846), .A2(n13935), .ZN(n13932) );
  INV_X1 U13325 ( .A(n10850), .ZN(n10847) );
  OR2_X2 U13326 ( .A1(n10848), .A2(n10847), .ZN(n13855) );
  OAI22_X1 U13327 ( .A1(n11860), .A2(n13855), .B1(n14752), .B2(n10850), .ZN(
        n10849) );
  AOI21_X1 U13328 ( .B1(n13932), .B2(n8099), .A(n10849), .ZN(n10855) );
  NAND2_X1 U13329 ( .A1(n8099), .A2(n11847), .ZN(n10854) );
  INV_X1 U13330 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10851) );
  OAI22_X1 U13331 ( .A1(n11860), .A2(n13838), .B1(n10851), .B2(n10850), .ZN(
        n10852) );
  INV_X1 U13332 ( .A(n10852), .ZN(n10853) );
  NAND2_X1 U13333 ( .A1(n10854), .A2(n10853), .ZN(n10892) );
  NOR2_X1 U13334 ( .A1(n10855), .A2(n10892), .ZN(n10856) );
  OR2_X1 U13335 ( .A1(n10893), .A2(n10856), .ZN(n14099) );
  NAND3_X1 U13336 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n10870) );
  OR2_X1 U13337 ( .A1(n10870), .A2(n10860), .ZN(n10868) );
  INV_X1 U13338 ( .A(n10868), .ZN(n10863) );
  AND2_X1 U13339 ( .A1(n14875), .A2(n10861), .ZN(n10862) );
  OR2_X1 U13340 ( .A1(n10865), .A2(n10864), .ZN(n10866) );
  INV_X1 U13341 ( .A(n14049), .ZN(n14691) );
  INV_X2 U13342 ( .A(n14351), .ZN(n14362) );
  NAND2_X1 U13343 ( .A1(n14691), .A2(n14362), .ZN(n14030) );
  INV_X1 U13344 ( .A(n14030), .ZN(n14055) );
  AOI22_X1 U13345 ( .A1(n14099), .A2(n14689), .B1(n14055), .B2(n7088), .ZN(
        n10875) );
  NAND2_X1 U13346 ( .A1(n10868), .A2(n14386), .ZN(n12148) );
  NAND2_X1 U13347 ( .A1(n10870), .A2(n10869), .ZN(n10872) );
  NAND2_X1 U13348 ( .A1(n10872), .A2(n10871), .ZN(n11599) );
  OR2_X1 U13349 ( .A1(n11599), .A2(P1_U3086), .ZN(n11120) );
  AOI22_X1 U13350 ( .A1(n14687), .A2(n10873), .B1(n11120), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U13351 ( .A1(n10875), .A2(n10874), .ZN(P1_U3232) );
  INV_X1 U13352 ( .A(n10876), .ZN(n10877) );
  XNOR2_X1 U13353 ( .A(n12518), .B(n11183), .ZN(n11065) );
  NAND2_X1 U13354 ( .A1(n13265), .A2(n12562), .ZN(n11064) );
  XNOR2_X1 U13355 ( .A(n11065), .B(n11064), .ZN(n11067) );
  XNOR2_X1 U13356 ( .A(n11068), .B(n11067), .ZN(n10884) );
  OAI21_X1 U13357 ( .B1(n14934), .B2(n11290), .A(n10880), .ZN(n10882) );
  AOI22_X1 U13358 ( .A1(n13612), .A2(n13266), .B1(n13264), .B2(n13614), .ZN(
        n11179) );
  NOR2_X1 U13359 ( .A1(n11179), .A2(n11070), .ZN(n10881) );
  AOI211_X1 U13360 ( .C1(n11183), .C2(n14930), .A(n10882), .B(n10881), .ZN(
        n10883) );
  OAI21_X1 U13361 ( .B1(n10884), .B2(n14926), .A(n10883), .ZN(P2_U3211) );
  INV_X1 U13362 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10889) );
  AND2_X1 U13363 ( .A1(n7088), .A2(n14362), .ZN(n10885) );
  AOI21_X1 U13364 ( .B1(n11865), .B2(n14384), .A(n10885), .ZN(n11862) );
  NAND2_X1 U13365 ( .A1(n11865), .A2(n14904), .ZN(n10886) );
  OAI211_X1 U13366 ( .C1(n10887), .C2(n11860), .A(n11862), .B(n10886), .ZN(
        n14485) );
  NAND2_X1 U13367 ( .A1(n14485), .A2(n14504), .ZN(n10888) );
  OAI21_X1 U13368 ( .B1(n14504), .B2(n10889), .A(n10888), .ZN(P1_U3459) );
  INV_X1 U13369 ( .A(n10890), .ZN(n11034) );
  AOI22_X1 U13370 ( .A1(n14151), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n14509), .ZN(n10891) );
  OAI21_X1 U13371 ( .B1(n11034), .B2(n14521), .A(n10891), .ZN(P1_U3341) );
  INV_X1 U13372 ( .A(n14687), .ZN(n14059) );
  INV_X1 U13373 ( .A(n10892), .ZN(n10894) );
  AOI21_X1 U13374 ( .B1(n10894), .B2(n12151), .A(n10893), .ZN(n11115) );
  INV_X2 U13375 ( .A(n7488), .ZN(n12151) );
  XNOR2_X1 U13376 ( .A(n10895), .B(n12151), .ZN(n10898) );
  XNOR2_X1 U13377 ( .A(n10898), .B(n10897), .ZN(n11114) );
  OAI22_X1 U13378 ( .A1(n11115), .A2(n11114), .B1(n10898), .B2(n10897), .ZN(
        n11584) );
  OAI22_X1 U13379 ( .A1(n11117), .A2(n13855), .B1(n14845), .B2(n13838), .ZN(
        n10899) );
  XNOR2_X1 U13380 ( .A(n10899), .B(n12151), .ZN(n11580) );
  NOR2_X1 U13381 ( .A1(n14845), .A2(n13855), .ZN(n10900) );
  AOI21_X1 U13382 ( .B1(n13932), .B2(n14086), .A(n10900), .ZN(n11581) );
  XNOR2_X1 U13383 ( .A(n11580), .B(n11581), .ZN(n11583) );
  XNOR2_X1 U13384 ( .A(n10901), .B(n11583), .ZN(n10902) );
  NAND2_X1 U13385 ( .A1(n10902), .A2(n14689), .ZN(n10906) );
  NAND2_X1 U13386 ( .A1(n7088), .A2(n14364), .ZN(n10904) );
  NAND2_X1 U13387 ( .A1(n14085), .A2(n14362), .ZN(n10903) );
  NAND2_X1 U13388 ( .A1(n10904), .A2(n10903), .ZN(n11563) );
  AOI22_X1 U13389 ( .A1(n14691), .A2(n11563), .B1(n11120), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10905) );
  OAI211_X1 U13390 ( .C1(n14845), .C2(n14059), .A(n10906), .B(n10905), .ZN(
        P1_U3237) );
  MUX2_X1 U13391 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12823), .Z(n11533) );
  XNOR2_X1 U13392 ( .A(n11533), .B(n11534), .ZN(n11531) );
  INV_X1 U13393 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10909) );
  INV_X1 U13394 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10908) );
  MUX2_X1 U13395 ( .A(n10909), .B(n10908), .S(n12823), .Z(n10910) );
  INV_X1 U13396 ( .A(n10959), .ZN(n11015) );
  INV_X1 U13397 ( .A(n10910), .ZN(n10911) );
  NAND2_X1 U13398 ( .A1(n10911), .A2(n10959), .ZN(n10912) );
  NAND2_X1 U13399 ( .A1(n10994), .A2(n10912), .ZN(n11004) );
  INV_X1 U13400 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10913) );
  MUX2_X1 U13401 ( .A(n10957), .B(n10913), .S(n12823), .Z(n11361) );
  NAND2_X1 U13402 ( .A1(n11361), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11003) );
  OR2_X1 U13403 ( .A1(n11004), .A2(n11003), .ZN(n10993) );
  NAND2_X1 U13404 ( .A1(n10993), .A2(n10994), .ZN(n10917) );
  INV_X1 U13405 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10960) );
  INV_X1 U13406 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10945) );
  MUX2_X1 U13407 ( .A(n10960), .B(n10945), .S(n12823), .Z(n10914) );
  NAND2_X1 U13408 ( .A1(n10914), .A2(n10961), .ZN(n15199) );
  INV_X1 U13409 ( .A(n10914), .ZN(n10915) );
  NAND2_X1 U13410 ( .A1(n10915), .A2(n11001), .ZN(n10916) );
  AND2_X1 U13411 ( .A1(n15199), .A2(n10916), .ZN(n10995) );
  NAND2_X1 U13412 ( .A1(n10917), .A2(n10995), .ZN(n15200) );
  NAND2_X1 U13413 ( .A1(n15200), .A2(n15199), .ZN(n10923) );
  INV_X1 U13414 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10919) );
  INV_X1 U13415 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10918) );
  MUX2_X1 U13416 ( .A(n10919), .B(n10918), .S(n12823), .Z(n10920) );
  NAND2_X1 U13417 ( .A1(n10920), .A2(n10962), .ZN(n10924) );
  INV_X1 U13418 ( .A(n10920), .ZN(n10921) );
  NAND2_X1 U13419 ( .A1(n10921), .A2(n15206), .ZN(n10922) );
  AND2_X1 U13420 ( .A1(n10924), .A2(n10922), .ZN(n15197) );
  NAND2_X1 U13421 ( .A1(n10923), .A2(n15197), .ZN(n15202) );
  NAND2_X1 U13422 ( .A1(n15202), .A2(n10924), .ZN(n15219) );
  MUX2_X1 U13423 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12823), .Z(n10925) );
  XNOR2_X1 U13424 ( .A(n10925), .B(n10965), .ZN(n15218) );
  NAND2_X1 U13425 ( .A1(n15219), .A2(n15218), .ZN(n15217) );
  INV_X1 U13426 ( .A(n10925), .ZN(n10926) );
  NAND2_X1 U13427 ( .A1(n10926), .A2(n10965), .ZN(n10927) );
  NAND2_X1 U13428 ( .A1(n15217), .A2(n10927), .ZN(n15239) );
  MUX2_X1 U13429 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12823), .Z(n10928) );
  NAND2_X1 U13430 ( .A1(n10928), .A2(n15240), .ZN(n15237) );
  NAND2_X1 U13431 ( .A1(n15239), .A2(n15237), .ZN(n10930) );
  INV_X1 U13432 ( .A(n10928), .ZN(n10929) );
  NAND2_X1 U13433 ( .A1(n10929), .A2(n10966), .ZN(n15236) );
  NAND2_X1 U13434 ( .A1(n10930), .A2(n15236), .ZN(n11094) );
  MUX2_X1 U13435 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12823), .Z(n10931) );
  INV_X1 U13436 ( .A(n11095), .ZN(n10932) );
  XNOR2_X1 U13437 ( .A(n10931), .B(n10932), .ZN(n11093) );
  NAND2_X1 U13438 ( .A1(n11094), .A2(n11093), .ZN(n10935) );
  INV_X1 U13439 ( .A(n10931), .ZN(n10933) );
  NAND2_X1 U13440 ( .A1(n10933), .A2(n10932), .ZN(n10934) );
  NAND2_X1 U13441 ( .A1(n10935), .A2(n10934), .ZN(n11532) );
  XOR2_X1 U13442 ( .A(n11531), .B(n11532), .Z(n10980) );
  NAND2_X1 U13443 ( .A1(P3_U3897), .A2(n6501), .ZN(n15241) );
  OR2_X1 U13444 ( .A1(n10937), .A2(n10936), .ZN(n10955) );
  NAND2_X1 U13445 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  AND2_X1 U13446 ( .A1(n10941), .A2(n10940), .ZN(n10953) );
  NAND2_X1 U13447 ( .A1(n10955), .A2(n10953), .ZN(n10974) );
  NOR2_X2 U13448 ( .A1(n10974), .A2(n10907), .ZN(n15287) );
  NAND2_X1 U13449 ( .A1(n11095), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10951) );
  INV_X1 U13450 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10942) );
  MUX2_X1 U13451 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10942), .S(n11095), .Z(
        n11104) );
  INV_X1 U13452 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U13453 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10943), .ZN(n11364) );
  NOR2_X1 U13454 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11364), .ZN(n10944) );
  NAND2_X1 U13455 ( .A1(n11006), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11005) );
  OAI21_X1 U13456 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n11364), .A(n11005), .ZN(
        n10982) );
  AOI22_X1 U13457 ( .A1(n15209), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n15206), 
        .B2(n10946), .ZN(n15228) );
  MUX2_X1 U13458 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10948), .S(n10965), .Z(
        n15227) );
  INV_X1 U13459 ( .A(n15226), .ZN(n10947) );
  OAI21_X1 U13460 ( .B1(n10965), .B2(n10948), .A(n10947), .ZN(n10949) );
  NAND2_X1 U13461 ( .A1(n15240), .A2(n10949), .ZN(n10950) );
  XNOR2_X1 U13462 ( .A(n10949), .B(n10966), .ZN(n15247) );
  NAND2_X1 U13463 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15247), .ZN(n15246) );
  NAND2_X1 U13464 ( .A1(n10950), .A2(n15246), .ZN(n11105) );
  NAND2_X1 U13465 ( .A1(n11104), .A2(n11105), .ZN(n11103) );
  NAND2_X1 U13466 ( .A1(n10951), .A2(n11103), .ZN(n11519) );
  XNOR2_X1 U13467 ( .A(n11519), .B(n11534), .ZN(n10952) );
  NAND2_X1 U13468 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10952), .ZN(n11521) );
  OAI21_X1 U13469 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10952), .A(n11521), .ZN(
        n10978) );
  MUX2_X1 U13470 ( .A(n12720), .B(n10974), .S(n6501), .Z(n15285) );
  INV_X1 U13471 ( .A(n10953), .ZN(n10954) );
  AOI22_X1 U13472 ( .A1(n15245), .A2(P3_ADDR_REG_7__SCAN_IN), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(P3_U3151), .ZN(n10956) );
  OAI21_X1 U13473 ( .B1(n15285), .B2(n11520), .A(n10956), .ZN(n10977) );
  INV_X1 U13474 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15235) );
  NOR2_X1 U13475 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10957), .ZN(n11358) );
  NAND2_X1 U13476 ( .A1(n9684), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10958) );
  OAI21_X1 U13477 ( .B1(n10959), .B2(n11358), .A(n10958), .ZN(n11010) );
  NOR2_X1 U13478 ( .A1(n11010), .A2(n10909), .ZN(n11009) );
  INV_X1 U13479 ( .A(n10963), .ZN(n10964) );
  NOR2_X1 U13480 ( .A1(n15196), .A2(n10919), .ZN(n15195) );
  INV_X1 U13481 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11084) );
  XNOR2_X1 U13482 ( .A(n10965), .B(n11084), .ZN(n15216) );
  NOR2_X1 U13483 ( .A1(n15235), .A2(n15234), .ZN(n15233) );
  NAND2_X1 U13484 ( .A1(n11095), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10970) );
  OR2_X1 U13485 ( .A1(n11095), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13486 ( .A1(n10970), .A2(n10968), .ZN(n11099) );
  INV_X1 U13487 ( .A(n11099), .ZN(n10969) );
  INV_X1 U13488 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10971) );
  AOI21_X1 U13489 ( .B1(n10972), .B2(n10971), .A(n11509), .ZN(n10975) );
  NOR2_X1 U13490 ( .A1(n10975), .A2(n15291), .ZN(n10976) );
  AOI211_X1 U13491 ( .C1(n15287), .C2(n10978), .A(n10977), .B(n10976), .ZN(
        n10979) );
  OAI21_X1 U13492 ( .B1(n10980), .B2(n15241), .A(n10979), .ZN(P3_U3189) );
  OAI21_X1 U13493 ( .B1(n10983), .B2(n10982), .A(n10981), .ZN(n10992) );
  OAI22_X1 U13494 ( .A1(n15296), .A2(n10985), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10984), .ZN(n10991) );
  AOI21_X1 U13495 ( .B1(n10988), .B2(n10987), .A(n10986), .ZN(n10989) );
  NOR2_X1 U13496 ( .A1(n15291), .A2(n10989), .ZN(n10990) );
  AOI211_X1 U13497 ( .C1(n15287), .C2(n10992), .A(n10991), .B(n10990), .ZN(
        n11000) );
  INV_X1 U13498 ( .A(n10993), .ZN(n11002) );
  INV_X1 U13499 ( .A(n10994), .ZN(n10996) );
  NOR3_X1 U13500 ( .A1(n11002), .A2(n10996), .A3(n10995), .ZN(n10998) );
  INV_X1 U13501 ( .A(n15200), .ZN(n10997) );
  OAI21_X1 U13502 ( .B1(n10998), .B2(n10997), .A(n15280), .ZN(n10999) );
  OAI211_X1 U13503 ( .C1(n15285), .C2(n11001), .A(n11000), .B(n10999), .ZN(
        P3_U3184) );
  AOI21_X1 U13504 ( .B1(n11004), .B2(n11003), .A(n11002), .ZN(n11018) );
  OAI21_X1 U13505 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n11006), .A(n11005), .ZN(
        n11014) );
  OAI22_X1 U13506 ( .A1(n15296), .A2(n11008), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11007), .ZN(n11013) );
  AOI21_X1 U13507 ( .B1(n10909), .B2(n11010), .A(n11009), .ZN(n11011) );
  NOR2_X1 U13508 ( .A1(n15291), .A2(n11011), .ZN(n11012) );
  AOI211_X1 U13509 ( .C1(n15287), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        n11017) );
  INV_X1 U13510 ( .A(n15285), .ZN(n14584) );
  NAND2_X1 U13511 ( .A1(n14584), .A2(n11015), .ZN(n11016) );
  OAI211_X1 U13512 ( .C1(n11018), .C2(n15241), .A(n11017), .B(n11016), .ZN(
        P3_U3183) );
  OAI21_X1 U13513 ( .B1(n11020), .B2(n11024), .A(n11019), .ZN(n11578) );
  INV_X1 U13514 ( .A(n11021), .ZN(n11022) );
  AOI211_X1 U13515 ( .C1(n11024), .C2(n11023), .A(n15308), .B(n11022), .ZN(
        n11026) );
  OAI22_X1 U13516 ( .A1(n11248), .A2(n15303), .B1(n11025), .B2(n15302), .ZN(
        n15177) );
  OR2_X1 U13517 ( .A1(n11026), .A2(n15177), .ZN(n11575) );
  AOI21_X1 U13518 ( .B1(n15339), .B2(n11578), .A(n11575), .ZN(n11048) );
  INV_X1 U13519 ( .A(n9652), .ZN(n15169) );
  INV_X1 U13520 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11027) );
  OAI22_X1 U13521 ( .A1(n13110), .A2(n15169), .B1(n15365), .B2(n11027), .ZN(
        n11028) );
  INV_X1 U13522 ( .A(n11028), .ZN(n11029) );
  OAI21_X1 U13523 ( .B1(n11048), .B2(n15363), .A(n11029), .ZN(P3_U3399) );
  INV_X1 U13524 ( .A(n11030), .ZN(n11031) );
  OAI222_X1 U13525 ( .A1(P3_U3151), .A2(n12822), .B1(n13125), .B2(n11032), 
        .C1(n13123), .C2(n11031), .ZN(P3_U3276) );
  INV_X1 U13526 ( .A(n13349), .ZN(n15005) );
  INV_X1 U13527 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11033) );
  OAI222_X1 U13528 ( .A1(P2_U3088), .A2(n15005), .B1(n13781), .B2(n11034), 
        .C1(n11033), .C2(n13783), .ZN(P2_U3313) );
  INV_X1 U13529 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n11045) );
  OAI21_X1 U13530 ( .B1(n11039), .B2(n11036), .A(n11035), .ZN(n11706) );
  NOR2_X1 U13531 ( .A1(n11704), .A2(n11860), .ZN(n11037) );
  NOR2_X1 U13532 ( .A1(n11568), .A2(n11037), .ZN(n11707) );
  INV_X1 U13533 ( .A(n11707), .ZN(n11038) );
  OAI22_X1 U13534 ( .A1(n11038), .A2(n10323), .B1(n11704), .B2(n14875), .ZN(
        n11043) );
  INV_X1 U13535 ( .A(n8099), .ZN(n11116) );
  INV_X1 U13536 ( .A(n14384), .ZN(n14348) );
  XNOR2_X1 U13537 ( .A(n11707), .B(n7088), .ZN(n11041) );
  INV_X1 U13538 ( .A(n11039), .ZN(n11040) );
  MUX2_X1 U13539 ( .A(n11041), .B(n11040), .S(n8099), .Z(n11042) );
  OAI222_X1 U13540 ( .A1(n14353), .A2(n11116), .B1(n14351), .B2(n11117), .C1(
        n14348), .C2(n11042), .ZN(n11712) );
  AOI211_X1 U13541 ( .C1(n14904), .C2(n11706), .A(n11043), .B(n11712), .ZN(
        n11220) );
  OR2_X1 U13542 ( .A1(n11220), .A2(n14905), .ZN(n11044) );
  OAI21_X1 U13543 ( .B1(n14504), .B2(n11045), .A(n11044), .ZN(P1_U3462) );
  OAI22_X1 U13544 ( .A1(n13062), .A2(n15169), .B1(n15374), .B2(n10918), .ZN(
        n11046) );
  INV_X1 U13545 ( .A(n11046), .ZN(n11047) );
  OAI21_X1 U13546 ( .B1(n11048), .B2(n15371), .A(n11047), .ZN(P3_U3462) );
  INV_X1 U13547 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11063) );
  OAI21_X1 U13548 ( .B1(n11051), .B2(n11050), .A(n6474), .ZN(n11052) );
  NAND2_X1 U13549 ( .A1(n11052), .A2(n14879), .ZN(n11058) );
  XNOR2_X1 U13550 ( .A(n11054), .B(n11053), .ZN(n11055) );
  NAND2_X1 U13551 ( .A1(n11055), .A2(n14384), .ZN(n11057) );
  AOI22_X1 U13552 ( .A1(n14084), .A2(n14362), .B1(n14364), .B2(n14086), .ZN(
        n11056) );
  NAND3_X1 U13553 ( .A1(n11058), .A2(n11057), .A3(n11056), .ZN(n12412) );
  INV_X1 U13554 ( .A(n12412), .ZN(n11061) );
  AND2_X1 U13555 ( .A1(n11567), .A2(n13916), .ZN(n11059) );
  NOR2_X1 U13556 ( .A1(n11682), .A2(n11059), .ZN(n12413) );
  AOI22_X1 U13557 ( .A1(n12413), .A2(n14883), .B1(n14882), .B2(n13916), .ZN(
        n11060) );
  NAND2_X1 U13558 ( .A1(n11061), .A2(n11060), .ZN(n11634) );
  NAND2_X1 U13559 ( .A1(n11634), .A2(n14504), .ZN(n11062) );
  OAI21_X1 U13560 ( .B1(n14504), .B2(n11063), .A(n11062), .ZN(P1_U3468) );
  INV_X1 U13561 ( .A(n11064), .ZN(n11066) );
  XNOR2_X1 U13562 ( .A(n11332), .B(n12518), .ZN(n11186) );
  NAND2_X1 U13563 ( .A1(n13264), .A2(n12562), .ZN(n11187) );
  XOR2_X1 U13564 ( .A(n11186), .B(n11187), .Z(n11188) );
  XNOR2_X1 U13565 ( .A(n11189), .B(n11188), .ZN(n11074) );
  OAI21_X1 U13566 ( .B1(n14934), .B2(n11315), .A(n11069), .ZN(n11072) );
  AOI22_X1 U13567 ( .A1(n13614), .A2(n13263), .B1(n13265), .B2(n13612), .ZN(
        n11320) );
  NOR2_X1 U13568 ( .A1(n11320), .A2(n11070), .ZN(n11071) );
  AOI211_X1 U13569 ( .C1(n11332), .C2(n14930), .A(n11072), .B(n11071), .ZN(
        n11073) );
  OAI21_X1 U13570 ( .B1(n11074), .B2(n14926), .A(n11073), .ZN(P2_U3185) );
  NAND2_X1 U13571 ( .A1(n11075), .A2(n15311), .ZN(n15312) );
  NAND2_X1 U13572 ( .A1(n12912), .A2(n15312), .ZN(n11076) );
  INV_X1 U13573 ( .A(n12999), .ZN(n11088) );
  OAI21_X1 U13574 ( .B1(n11078), .B2(n11080), .A(n11077), .ZN(n11148) );
  INV_X1 U13575 ( .A(n11148), .ZN(n11087) );
  INV_X1 U13576 ( .A(n11079), .ZN(n11081) );
  AOI21_X1 U13577 ( .B1(n11081), .B2(n11080), .A(n15308), .ZN(n11083) );
  OAI22_X1 U13578 ( .A1(n11803), .A2(n15303), .B1(n15304), .B2(n15302), .ZN(
        n11168) );
  AOI21_X1 U13579 ( .B1(n11083), .B2(n11082), .A(n11168), .ZN(n11146) );
  MUX2_X1 U13580 ( .A(n11084), .B(n11146), .S(n15334), .Z(n11086) );
  AOI22_X1 U13581 ( .A1(n14607), .A2(n11156), .B1(n15331), .B2(n11154), .ZN(
        n11085) );
  OAI211_X1 U13582 ( .C1(n11088), .C2(n11087), .A(n11086), .B(n11085), .ZN(
        P3_U3229) );
  OAI22_X1 U13583 ( .A1(n13062), .A2(n11089), .B1(n15374), .B2(n10913), .ZN(
        n11090) );
  AOI21_X1 U13584 ( .B1(n11091), .B2(n15374), .A(n11090), .ZN(n11092) );
  INV_X1 U13585 ( .A(n11092), .ZN(P3_U3459) );
  XNOR2_X1 U13586 ( .A(n11094), .B(n11093), .ZN(n11112) );
  NOR2_X1 U13587 ( .A1(n15285), .A2(n11095), .ZN(n11111) );
  INV_X1 U13588 ( .A(n11096), .ZN(n11100) );
  INV_X1 U13589 ( .A(n11097), .ZN(n11098) );
  AOI21_X1 U13590 ( .B1(n11100), .B2(n11099), .A(n11098), .ZN(n11101) );
  INV_X1 U13591 ( .A(n11101), .ZN(n11102) );
  NAND2_X1 U13592 ( .A1(n14593), .A2(n11102), .ZN(n11109) );
  AND2_X1 U13593 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n15184) );
  AOI21_X1 U13594 ( .B1(n15245), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n15184), .ZN(
        n11108) );
  OAI21_X1 U13595 ( .B1(n11105), .B2(n11104), .A(n11103), .ZN(n11106) );
  NAND2_X1 U13596 ( .A1(n15287), .A2(n11106), .ZN(n11107) );
  NAND3_X1 U13597 ( .A1(n11109), .A2(n11108), .A3(n11107), .ZN(n11110) );
  AOI211_X1 U13598 ( .C1(n11112), .C2(n15280), .A(n11111), .B(n11110), .ZN(
        n11113) );
  INV_X1 U13599 ( .A(n11113), .ZN(P3_U3188) );
  XOR2_X1 U13600 ( .A(n11115), .B(n11114), .Z(n11122) );
  NOR2_X1 U13601 ( .A1(n14059), .A2(n11704), .ZN(n11119) );
  NAND2_X1 U13602 ( .A1(n14691), .A2(n14364), .ZN(n14057) );
  OAI22_X1 U13603 ( .A1(n11117), .A2(n14030), .B1(n14057), .B2(n11116), .ZN(
        n11118) );
  AOI211_X1 U13604 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n11120), .A(n11119), .B(
        n11118), .ZN(n11121) );
  OAI21_X1 U13605 ( .B1(n11122), .B2(n14065), .A(n11121), .ZN(P1_U3222) );
  INV_X1 U13606 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n14018) );
  NOR2_X1 U13607 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14018), .ZN(n11123) );
  AOI21_X1 U13608 ( .B1(n14757), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11123), 
        .ZN(n11124) );
  INV_X1 U13609 ( .A(n11124), .ZN(n11131) );
  INV_X1 U13610 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14561) );
  AOI22_X1 U13611 ( .A1(n14788), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14561), 
        .B2(n11132), .ZN(n14786) );
  OAI21_X1 U13612 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n14788), .A(n14784), 
        .ZN(n11129) );
  INV_X1 U13613 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11127) );
  MUX2_X1 U13614 ( .A(n11127), .B(P1_REG1_REG_13__SCAN_IN), .S(n11775), .Z(
        n11128) );
  NOR2_X1 U13615 ( .A1(n11129), .A2(n11128), .ZN(n11774) );
  AOI211_X1 U13616 ( .C1(n11129), .C2(n11128), .A(n11774), .B(n14168), .ZN(
        n11130) );
  AOI211_X1 U13617 ( .C1(n14804), .C2(n11775), .A(n11131), .B(n11130), .ZN(
        n11145) );
  NOR2_X1 U13618 ( .A1(n14788), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11139) );
  INV_X1 U13619 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U13620 ( .A1(n14788), .A2(n11133), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n11132), .ZN(n14783) );
  OR2_X1 U13621 ( .A1(n11135), .A2(n11134), .ZN(n11136) );
  OAI21_X1 U13622 ( .B1(n11138), .B2(n11137), .A(n11136), .ZN(n14782) );
  NOR2_X1 U13623 ( .A1(n14783), .A2(n14782), .ZN(n14781) );
  NOR2_X1 U13624 ( .A1(n11139), .A2(n14781), .ZN(n11143) );
  INV_X1 U13625 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11140) );
  MUX2_X1 U13626 ( .A(n11140), .B(P1_REG2_REG_13__SCAN_IN), .S(n11775), .Z(
        n11141) );
  INV_X1 U13627 ( .A(n11141), .ZN(n11142) );
  NAND2_X1 U13628 ( .A1(n11142), .A2(n11143), .ZN(n11759) );
  OAI211_X1 U13629 ( .C1(n11143), .C2(n11142), .A(n14771), .B(n11759), .ZN(
        n11144) );
  NAND2_X1 U13630 ( .A1(n11145), .A2(n11144), .ZN(P1_U3256) );
  INV_X1 U13631 ( .A(n11146), .ZN(n11147) );
  AOI21_X1 U13632 ( .B1(n15339), .B2(n11148), .A(n11147), .ZN(n11153) );
  INV_X1 U13633 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11149) );
  OAI22_X1 U13634 ( .A1(n13110), .A2(n11166), .B1(n15365), .B2(n11149), .ZN(
        n11150) );
  INV_X1 U13635 ( .A(n11150), .ZN(n11151) );
  OAI21_X1 U13636 ( .B1(n11153), .B2(n15363), .A(n11151), .ZN(P3_U3402) );
  INV_X1 U13637 ( .A(n13062), .ZN(n13044) );
  AOI22_X1 U13638 ( .A1(n13044), .A2(n11156), .B1(n15371), .B2(
        P3_REG1_REG_4__SCAN_IN), .ZN(n11152) );
  OAI21_X1 U13639 ( .B1(n11153), .B2(n15371), .A(n11152), .ZN(P3_U3463) );
  INV_X1 U13640 ( .A(n11154), .ZN(n11171) );
  XNOR2_X1 U13641 ( .A(n11156), .B(n10585), .ZN(n11244) );
  XNOR2_X1 U13642 ( .A(n12719), .B(n11244), .ZN(n11164) );
  INV_X1 U13643 ( .A(n11157), .ZN(n11158) );
  XNOR2_X1 U13644 ( .A(n10219), .B(n10585), .ZN(n11161) );
  XNOR2_X1 U13645 ( .A(n11161), .B(n12721), .ZN(n15174) );
  OAI21_X1 U13646 ( .B1(n11164), .B2(n11163), .A(n11245), .ZN(n11165) );
  NAND2_X1 U13647 ( .A1(n11165), .A2(n15180), .ZN(n11170) );
  OAI22_X1 U13648 ( .A1(n15170), .A2(n11166), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15220), .ZN(n11167) );
  AOI21_X1 U13649 ( .B1(n15178), .B2(n11168), .A(n11167), .ZN(n11169) );
  OAI211_X1 U13650 ( .C1(n11171), .C2(n15193), .A(n11170), .B(n11169), .ZN(
        P3_U3170) );
  INV_X1 U13651 ( .A(n11172), .ZN(n11199) );
  AOI22_X1 U13652 ( .A1(n14803), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n14509), .ZN(n11173) );
  OAI21_X1 U13653 ( .B1(n11199), .B2(n14521), .A(n11173), .ZN(P1_U3340) );
  XNOR2_X1 U13654 ( .A(n11174), .B(n11175), .ZN(n11286) );
  INV_X1 U13655 ( .A(n11304), .ZN(n11177) );
  INV_X1 U13656 ( .A(n11314), .ZN(n11176) );
  AOI211_X1 U13657 ( .C1(n11183), .C2(n11177), .A(n12562), .B(n11176), .ZN(
        n11293) );
  XNOR2_X1 U13658 ( .A(n11178), .B(n6837), .ZN(n11180) );
  OAI21_X1 U13659 ( .B1(n11180), .B2(n13593), .A(n11179), .ZN(n11287) );
  AOI211_X1 U13660 ( .C1(n15137), .C2(n11286), .A(n11293), .B(n11287), .ZN(
        n11185) );
  OAI22_X1 U13661 ( .A1(n13754), .A2(n11291), .B1(n15147), .B2(n8916), .ZN(
        n11181) );
  INV_X1 U13662 ( .A(n11181), .ZN(n11182) );
  OAI21_X1 U13663 ( .B1(n11185), .B2(n15145), .A(n11182), .ZN(P2_U3448) );
  AOI22_X1 U13664 ( .A1(n13688), .A2(n11183), .B1(n15154), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11184) );
  OAI21_X1 U13665 ( .B1(n11185), .B2(n15154), .A(n11184), .ZN(P2_U3505) );
  XNOR2_X1 U13666 ( .A(n11396), .B(n12547), .ZN(n11191) );
  NAND2_X1 U13667 ( .A1(n13263), .A2(n12562), .ZN(n11190) );
  NOR2_X1 U13668 ( .A1(n11191), .A2(n11190), .ZN(n11372) );
  NAND2_X1 U13669 ( .A1(n11191), .A2(n11190), .ZN(n11373) );
  INV_X1 U13670 ( .A(n11373), .ZN(n11192) );
  NOR2_X1 U13671 ( .A1(n11372), .A2(n11192), .ZN(n11193) );
  XNOR2_X1 U13672 ( .A(n11374), .B(n11193), .ZN(n11198) );
  NAND2_X1 U13673 ( .A1(n13249), .A2(n13612), .ZN(n14921) );
  INV_X1 U13674 ( .A(n14921), .ZN(n13220) );
  INV_X1 U13675 ( .A(n14920), .ZN(n13219) );
  AOI22_X1 U13676 ( .A1(n13220), .A2(n13264), .B1(n13219), .B2(n13262), .ZN(
        n11195) );
  OAI211_X1 U13677 ( .C1(n11391), .C2(n14934), .A(n11195), .B(n11194), .ZN(
        n11196) );
  AOI21_X1 U13678 ( .B1(n11396), .B2(n14930), .A(n11196), .ZN(n11197) );
  OAI21_X1 U13679 ( .B1(n11198), .B2(n14926), .A(n11197), .ZN(P2_U3193) );
  INV_X1 U13680 ( .A(n15016), .ZN(n13350) );
  OAI222_X1 U13681 ( .A1(n13783), .A2(n11200), .B1(n13781), .B2(n11199), .C1(
        n13350), .C2(P2_U3088), .ZN(P2_U3312) );
  AND2_X1 U13682 ( .A1(n11201), .A2(n15089), .ZN(n11204) );
  NAND4_X1 U13683 ( .A1(n11204), .A2(n15090), .A3(n11203), .A4(n11202), .ZN(
        n11205) );
  OR2_X1 U13684 ( .A1(n11206), .A2(n13379), .ZN(n11226) );
  INV_X1 U13685 ( .A(n11226), .ZN(n11207) );
  NAND2_X1 U13686 ( .A1(n7490), .A2(n11207), .ZN(n13495) );
  INV_X1 U13687 ( .A(n11208), .ZN(n11209) );
  AND2_X1 U13688 ( .A1(n11276), .A2(n11209), .ZN(n15096) );
  OAI21_X1 U13689 ( .B1(n14668), .B2(n8803), .A(n13525), .ZN(n11214) );
  INV_X1 U13690 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11212) );
  INV_X1 U13691 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11211) );
  OAI22_X1 U13692 ( .A1(n7490), .A2(n11212), .B1(n11211), .B2(n13419), .ZN(
        n11213) );
  AOI21_X1 U13693 ( .B1(n15096), .B2(n11214), .A(n11213), .ZN(n11218) );
  INV_X1 U13694 ( .A(n9219), .ZN(n15106) );
  NOR2_X1 U13695 ( .A1(n15106), .A2(n9268), .ZN(n11215) );
  OAI22_X1 U13696 ( .A1(n11216), .A2(n13537), .B1(n11215), .B2(n15094), .ZN(
        n15095) );
  NAND2_X1 U13697 ( .A1(n15095), .A2(n7490), .ZN(n11217) );
  OAI211_X1 U13698 ( .C1(n13495), .C2(n15094), .A(n11218), .B(n11217), .ZN(
        P2_U3265) );
  NAND2_X1 U13699 ( .A1(n14917), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11219) );
  OAI21_X1 U13700 ( .B1(n11220), .B2(n14917), .A(n11219), .ZN(P1_U3529) );
  XNOR2_X1 U13701 ( .A(n11221), .B(n11225), .ZN(n11223) );
  AOI21_X1 U13702 ( .B1(n11223), .B2(n9268), .A(n11222), .ZN(n15110) );
  XNOR2_X1 U13703 ( .A(n11224), .B(n11225), .ZN(n15108) );
  INV_X1 U13704 ( .A(n15108), .ZN(n11234) );
  AND2_X1 U13705 ( .A1(n9219), .A2(n11226), .ZN(n11227) );
  OAI211_X1 U13706 ( .C1(n6922), .C2(n6921), .A(n6483), .B(n11267), .ZN(n15109) );
  OAI22_X1 U13707 ( .A1(n7490), .A2(n10445), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n13419), .ZN(n11230) );
  AOI21_X1 U13708 ( .B1(n14655), .B2(n11231), .A(n11230), .ZN(n11232) );
  OAI21_X1 U13709 ( .B1(n15109), .B2(n13525), .A(n11232), .ZN(n11233) );
  AOI21_X1 U13710 ( .B1(n11234), .B2(n14665), .A(n11233), .ZN(n11235) );
  OAI21_X1 U13711 ( .B1(n14668), .B2(n15110), .A(n11235), .ZN(P2_U3262) );
  NAND2_X1 U13712 ( .A1(n11236), .A2(n7490), .ZN(n11242) );
  OAI22_X1 U13713 ( .A1(n7490), .A2(n8856), .B1(n11237), .B2(n13419), .ZN(
        n11240) );
  NOR2_X1 U13714 ( .A1(n11238), .A2(n13525), .ZN(n11239) );
  AOI211_X1 U13715 ( .C1(n14655), .C2(n6477), .A(n11240), .B(n11239), .ZN(
        n11241) );
  OAI211_X1 U13716 ( .C1(n13641), .C2(n11243), .A(n11242), .B(n11241), .ZN(
        P2_U3263) );
  XNOR2_X1 U13717 ( .A(n11449), .B(n12485), .ZN(n11802) );
  XNOR2_X1 U13718 ( .A(n11803), .B(n11802), .ZN(n11805) );
  XNOR2_X1 U13719 ( .A(n11806), .B(n11805), .ZN(n11254) );
  INV_X1 U13720 ( .A(n11246), .ZN(n11448) );
  AOI22_X1 U13721 ( .A1(n15186), .A2(n11247), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11252) );
  OR2_X1 U13722 ( .A1(n11248), .A2(n15302), .ZN(n11250) );
  INV_X1 U13723 ( .A(n15303), .ZN(n12962) );
  NAND2_X1 U13724 ( .A1(n12717), .A2(n12962), .ZN(n11249) );
  NAND2_X1 U13725 ( .A1(n11250), .A2(n11249), .ZN(n11345) );
  NAND2_X1 U13726 ( .A1(n11345), .A2(n15178), .ZN(n11251) );
  OAI211_X1 U13727 ( .C1(n15193), .C2(n11448), .A(n11252), .B(n11251), .ZN(
        n11253) );
  AOI21_X1 U13728 ( .B1(n11254), .B2(n15180), .A(n11253), .ZN(n11255) );
  INV_X1 U13729 ( .A(n11255), .ZN(P3_U3167) );
  INV_X1 U13730 ( .A(n13368), .ZN(n13361) );
  INV_X1 U13731 ( .A(n11256), .ZN(n11258) );
  OAI222_X1 U13732 ( .A1(P2_U3088), .A2(n13361), .B1(n13781), .B2(n11258), 
        .C1(n11257), .C2(n13783), .ZN(P2_U3311) );
  OAI222_X1 U13733 ( .A1(n14527), .A2(n11259), .B1(n14525), .B2(n11258), .C1(
        n11772), .C2(P1_U3086), .ZN(P1_U3339) );
  XNOR2_X1 U13734 ( .A(n11261), .B(n11262), .ZN(n15114) );
  XNOR2_X1 U13735 ( .A(n11263), .B(n11262), .ZN(n11265) );
  AOI21_X1 U13736 ( .B1(n11265), .B2(n9268), .A(n11264), .ZN(n15117) );
  MUX2_X1 U13737 ( .A(n11266), .B(n15117), .S(n7490), .Z(n11272) );
  AOI211_X1 U13738 ( .C1(n11268), .C2(n11267), .A(n12562), .B(n11303), .ZN(
        n15115) );
  OAI22_X1 U13739 ( .A1(n13636), .A2(n15118), .B1(n13419), .B2(n11269), .ZN(
        n11270) );
  AOI21_X1 U13740 ( .B1(n15115), .B2(n14664), .A(n11270), .ZN(n11271) );
  OAI211_X1 U13741 ( .C1(n13641), .C2(n15114), .A(n11272), .B(n11271), .ZN(
        P2_U3261) );
  INV_X1 U13742 ( .A(n11273), .ZN(n11274) );
  AOI21_X1 U13743 ( .B1(n11274), .B2(n9509), .A(n6643), .ZN(n15102) );
  AOI211_X1 U13744 ( .C1(n11276), .C2(n10663), .A(n12562), .B(n11275), .ZN(
        n15099) );
  OAI22_X1 U13745 ( .A1(n13636), .A2(n8834), .B1(n14942), .B2(n13419), .ZN(
        n11277) );
  AOI21_X1 U13746 ( .B1(n15099), .B2(n14664), .A(n11277), .ZN(n11283) );
  OAI21_X1 U13747 ( .B1(n11279), .B2(n9509), .A(n11278), .ZN(n11281) );
  AOI21_X1 U13748 ( .B1(n11281), .B2(n9268), .A(n11280), .ZN(n15098) );
  MUX2_X1 U13749 ( .A(n15098), .B(n10444), .S(n14668), .Z(n11282) );
  OAI211_X1 U13750 ( .C1(n15102), .C2(n13641), .A(n11283), .B(n11282), .ZN(
        P2_U3264) );
  NAND2_X1 U13751 ( .A1(n12720), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11284) );
  OAI21_X1 U13752 ( .B1(n11285), .B2(n12720), .A(n11284), .ZN(P3_U3521) );
  INV_X1 U13753 ( .A(n11286), .ZN(n11296) );
  INV_X1 U13754 ( .A(n11287), .ZN(n11288) );
  MUX2_X1 U13755 ( .A(n11289), .B(n11288), .S(n7490), .Z(n11295) );
  OAI22_X1 U13756 ( .A1(n11291), .A2(n13636), .B1(n13419), .B2(n11290), .ZN(
        n11292) );
  AOI21_X1 U13757 ( .B1(n11293), .B2(n14664), .A(n11292), .ZN(n11294) );
  OAI211_X1 U13758 ( .C1(n11296), .C2(n13641), .A(n11295), .B(n11294), .ZN(
        P2_U3259) );
  XNOR2_X1 U13759 ( .A(n11297), .B(n11298), .ZN(n15122) );
  XNOR2_X1 U13760 ( .A(n11299), .B(n11298), .ZN(n11301) );
  AOI21_X1 U13761 ( .B1(n11301), .B2(n9268), .A(n11300), .ZN(n15126) );
  MUX2_X1 U13762 ( .A(n11302), .B(n15126), .S(n7490), .Z(n11311) );
  INV_X1 U13763 ( .A(n11303), .ZN(n11305) );
  AOI211_X1 U13764 ( .C1(n11306), .C2(n11305), .A(n12562), .B(n11304), .ZN(
        n15124) );
  INV_X1 U13765 ( .A(n11307), .ZN(n11308) );
  OAI22_X1 U13766 ( .A1(n15127), .A2(n13636), .B1(n13419), .B2(n11308), .ZN(
        n11309) );
  AOI21_X1 U13767 ( .B1(n15124), .B2(n14664), .A(n11309), .ZN(n11310) );
  OAI211_X1 U13768 ( .C1(n13641), .C2(n15122), .A(n11311), .B(n11310), .ZN(
        P2_U3260) );
  XOR2_X1 U13769 ( .A(n11312), .B(n11318), .Z(n11329) );
  INV_X1 U13770 ( .A(n11329), .ZN(n11326) );
  INV_X1 U13771 ( .A(n11313), .ZN(n11393) );
  AOI211_X1 U13772 ( .C1(n11332), .C2(n11314), .A(n12562), .B(n11393), .ZN(
        n11328) );
  INV_X1 U13773 ( .A(n11332), .ZN(n11316) );
  OAI22_X1 U13774 ( .A1(n11316), .A2(n13636), .B1(n13419), .B2(n11315), .ZN(
        n11317) );
  AOI21_X1 U13775 ( .B1(n11328), .B2(n14664), .A(n11317), .ZN(n11325) );
  XNOR2_X1 U13776 ( .A(n11319), .B(n11318), .ZN(n11321) );
  OAI21_X1 U13777 ( .B1(n11321), .B2(n13593), .A(n11320), .ZN(n11327) );
  INV_X1 U13778 ( .A(n11327), .ZN(n11322) );
  MUX2_X1 U13779 ( .A(n11323), .B(n11322), .S(n7490), .Z(n11324) );
  OAI211_X1 U13780 ( .C1(n11326), .C2(n13641), .A(n11325), .B(n11324), .ZN(
        P2_U3258) );
  AOI211_X1 U13781 ( .C1(n15137), .C2(n11329), .A(n11328), .B(n11327), .ZN(
        n11334) );
  AOI22_X1 U13782 ( .A1(n11332), .A2(n13688), .B1(n15154), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11330) );
  OAI21_X1 U13783 ( .B1(n11334), .B2(n15154), .A(n11330), .ZN(P2_U3506) );
  NOR2_X1 U13784 ( .A1(n15147), .A2(n8930), .ZN(n11331) );
  AOI21_X1 U13785 ( .B1(n11332), .B2(n13749), .A(n11331), .ZN(n11333) );
  OAI21_X1 U13786 ( .B1(n11334), .B2(n15145), .A(n11333), .ZN(P2_U3451) );
  INV_X1 U13787 ( .A(n11335), .ZN(n11337) );
  OAI222_X1 U13788 ( .A1(n11338), .A2(P3_U3151), .B1(n13123), .B2(n11337), 
        .C1(n11336), .C2(n13125), .ZN(P3_U3275) );
  OAI21_X1 U13789 ( .B1(n11340), .B2(n11344), .A(n11339), .ZN(n11453) );
  INV_X1 U13790 ( .A(n11341), .ZN(n11342) );
  AOI21_X1 U13791 ( .B1(n11344), .B2(n11343), .A(n11342), .ZN(n11347) );
  INV_X1 U13792 ( .A(n11345), .ZN(n11346) );
  OAI21_X1 U13793 ( .B1(n11347), .B2(n15308), .A(n11346), .ZN(n11450) );
  AOI21_X1 U13794 ( .B1(n15339), .B2(n11453), .A(n11450), .ZN(n11354) );
  INV_X1 U13795 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11348) );
  OAI22_X1 U13796 ( .A1(n13110), .A2(n11449), .B1(n15365), .B2(n11348), .ZN(
        n11349) );
  INV_X1 U13797 ( .A(n11349), .ZN(n11350) );
  OAI21_X1 U13798 ( .B1(n11354), .B2(n15363), .A(n11350), .ZN(P3_U3405) );
  INV_X1 U13799 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11351) );
  OAI22_X1 U13800 ( .A1(n13062), .A2(n11449), .B1(n15374), .B2(n11351), .ZN(
        n11352) );
  INV_X1 U13801 ( .A(n11352), .ZN(n11353) );
  OAI21_X1 U13802 ( .B1(n11354), .B2(n15371), .A(n11353), .ZN(P3_U3464) );
  INV_X1 U13803 ( .A(n11355), .ZN(n11356) );
  INV_X1 U13804 ( .A(n12239), .ZN(n12244) );
  OAI222_X1 U13805 ( .A1(n14527), .A2(n7058), .B1(n14525), .B2(n11356), .C1(
        n12244), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13806 ( .A(n15026), .ZN(n13363) );
  OAI222_X1 U13807 ( .A1(n13783), .A2(n11357), .B1(n13781), .B2(n11356), .C1(
        n13363), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13808 ( .A(n11358), .ZN(n11371) );
  INV_X1 U13809 ( .A(n11361), .ZN(n11359) );
  NAND2_X1 U13810 ( .A1(n15280), .A2(n11359), .ZN(n11363) );
  INV_X1 U13811 ( .A(n15287), .ZN(n15257) );
  NAND3_X1 U13812 ( .A1(n15291), .A2(n15241), .A3(n15257), .ZN(n11360) );
  AOI21_X1 U13813 ( .B1(n11361), .B2(n11360), .A(n14584), .ZN(n11362) );
  MUX2_X1 U13814 ( .A(n11363), .B(n11362), .S(P3_IR_REG_0__SCAN_IN), .Z(n11370) );
  INV_X1 U13815 ( .A(n11364), .ZN(n11368) );
  OAI22_X1 U13816 ( .A1(n15296), .A2(n11366), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11365), .ZN(n11367) );
  AOI21_X1 U13817 ( .B1(n15287), .B2(n11368), .A(n11367), .ZN(n11369) );
  OAI211_X1 U13818 ( .C1(n15291), .C2(n11371), .A(n11370), .B(n11369), .ZN(
        P3_U3182) );
  XNOR2_X1 U13819 ( .A(n11701), .B(n12518), .ZN(n11429) );
  NAND2_X1 U13820 ( .A1(n13262), .A2(n12562), .ZN(n11430) );
  XNOR2_X1 U13821 ( .A(n11429), .B(n11430), .ZN(n11375) );
  NAND2_X1 U13822 ( .A1(n11376), .A2(n11375), .ZN(n11433) );
  OAI21_X1 U13823 ( .B1(n11376), .B2(n11375), .A(n11433), .ZN(n11377) );
  NAND2_X1 U13824 ( .A1(n11377), .A2(n13243), .ZN(n11382) );
  OAI22_X1 U13825 ( .A1(n11378), .A2(n13539), .B1(n11788), .B2(n13537), .ZN(
        n11485) );
  OAI22_X1 U13826 ( .A1(n14934), .A2(n11489), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11379), .ZN(n11380) );
  AOI21_X1 U13827 ( .B1(n11485), .B2(n13249), .A(n11380), .ZN(n11381) );
  OAI211_X1 U13828 ( .C1(n6932), .C2(n13252), .A(n11382), .B(n11381), .ZN(
        P2_U3203) );
  XOR2_X1 U13829 ( .A(n11383), .B(n11387), .Z(n15134) );
  INV_X1 U13830 ( .A(n15134), .ZN(n11399) );
  INV_X1 U13831 ( .A(n11384), .ZN(n11385) );
  AOI21_X1 U13832 ( .B1(n11387), .B2(n11386), .A(n11385), .ZN(n11390) );
  NAND2_X1 U13833 ( .A1(n15134), .A2(n15106), .ZN(n11389) );
  AOI22_X1 U13834 ( .A1(n13612), .A2(n13264), .B1(n13262), .B2(n13614), .ZN(
        n11388) );
  OAI211_X1 U13835 ( .C1(n13593), .C2(n11390), .A(n11389), .B(n11388), .ZN(
        n15132) );
  NAND2_X1 U13836 ( .A1(n15132), .A2(n7490), .ZN(n11398) );
  OAI22_X1 U13837 ( .A1(n7490), .A2(n11392), .B1(n11391), .B2(n13419), .ZN(
        n11395) );
  INV_X1 U13838 ( .A(n11396), .ZN(n15131) );
  OAI211_X1 U13839 ( .C1(n11393), .C2(n15131), .A(n6483), .B(n11488), .ZN(
        n15130) );
  NOR2_X1 U13840 ( .A1(n15130), .A2(n13525), .ZN(n11394) );
  AOI211_X1 U13841 ( .C1(n14655), .C2(n11396), .A(n11395), .B(n11394), .ZN(
        n11397) );
  OAI211_X1 U13842 ( .C1(n11399), .C2(n13495), .A(n11398), .B(n11397), .ZN(
        P2_U3257) );
  INV_X1 U13843 ( .A(n11400), .ZN(n11401) );
  OAI222_X1 U13844 ( .A1(P3_U3151), .A2(n10181), .B1(n13125), .B2(n11402), 
        .C1(n13123), .C2(n11401), .ZN(P3_U3274) );
  OAI21_X1 U13845 ( .B1(n11404), .B2(n11808), .A(n11403), .ZN(n11678) );
  OAI211_X1 U13846 ( .C1(n11407), .C2(n11406), .A(n11405), .B(n15317), .ZN(
        n11410) );
  OR2_X1 U13847 ( .A1(n11816), .A2(n15303), .ZN(n11409) );
  NAND2_X1 U13848 ( .A1(n12717), .A2(n12963), .ZN(n11408) );
  AND2_X1 U13849 ( .A1(n11409), .A2(n11408), .ZN(n15165) );
  NAND2_X1 U13850 ( .A1(n11410), .A2(n15165), .ZN(n11675) );
  AOI21_X1 U13851 ( .B1(n15339), .B2(n11678), .A(n11675), .ZN(n11417) );
  INV_X1 U13852 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11411) );
  OAI22_X1 U13853 ( .A1(n13110), .A2(n11674), .B1(n15365), .B2(n11411), .ZN(
        n11412) );
  INV_X1 U13854 ( .A(n11412), .ZN(n11413) );
  OAI21_X1 U13855 ( .B1(n11417), .B2(n15363), .A(n11413), .ZN(P3_U3411) );
  INV_X1 U13856 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11414) );
  OAI22_X1 U13857 ( .A1(n13062), .A2(n11674), .B1(n15374), .B2(n11414), .ZN(
        n11415) );
  INV_X1 U13858 ( .A(n11415), .ZN(n11416) );
  OAI21_X1 U13859 ( .B1(n11417), .B2(n15371), .A(n11416), .ZN(P3_U3466) );
  XNOR2_X1 U13860 ( .A(n11418), .B(n6584), .ZN(n15345) );
  NOR2_X1 U13861 ( .A1(n13001), .A2(n15312), .ZN(n15332) );
  INV_X1 U13862 ( .A(n15332), .ZN(n11739) );
  OAI211_X1 U13863 ( .C1(n11420), .C2(n6584), .A(n11419), .B(n15317), .ZN(
        n11421) );
  AOI22_X1 U13864 ( .A1(n11810), .A2(n12962), .B1(n12963), .B2(n12718), .ZN(
        n15190) );
  OAI211_X1 U13865 ( .C1(n12912), .C2(n15345), .A(n11421), .B(n15190), .ZN(
        n15347) );
  INV_X1 U13866 ( .A(n15347), .ZN(n11423) );
  INV_X1 U13867 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11422) );
  MUX2_X1 U13868 ( .A(n11423), .B(n11422), .S(n13001), .Z(n11428) );
  NAND2_X1 U13869 ( .A1(n15185), .A2(n15325), .ZN(n15346) );
  NOR3_X1 U13870 ( .A1(n15346), .A2(n15311), .A3(n11424), .ZN(n11425) );
  AOI21_X1 U13871 ( .B1(n15331), .B2(n11426), .A(n11425), .ZN(n11427) );
  OAI211_X1 U13872 ( .C1(n15345), .C2(n11739), .A(n11428), .B(n11427), .ZN(
        P3_U3227) );
  INV_X1 U13873 ( .A(n11429), .ZN(n11431) );
  XNOR2_X1 U13874 ( .A(n11620), .B(n12547), .ZN(n11435) );
  NAND2_X1 U13875 ( .A1(n13261), .A2(n12562), .ZN(n11434) );
  NOR2_X1 U13876 ( .A1(n11435), .A2(n11434), .ZN(n11662) );
  AOI21_X1 U13877 ( .B1(n11435), .B2(n11434), .A(n11662), .ZN(n11436) );
  OAI211_X1 U13878 ( .C1(n11437), .C2(n11436), .A(n11664), .B(n13243), .ZN(
        n11443) );
  OAI22_X1 U13879 ( .A1(n14934), .A2(n11617), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11438), .ZN(n11441) );
  OAI22_X1 U13880 ( .A1(n11439), .A2(n14921), .B1(n14920), .B2(n14922), .ZN(
        n11440) );
  AOI211_X1 U13881 ( .C1(n11620), .C2(n14930), .A(n11441), .B(n11440), .ZN(
        n11442) );
  NAND2_X1 U13882 ( .A1(n11443), .A2(n11442), .ZN(P2_U3189) );
  INV_X1 U13883 ( .A(n11444), .ZN(n11447) );
  OAI22_X1 U13884 ( .A1(n11445), .A2(P3_U3151), .B1(SI_22_), .B2(n13125), .ZN(
        n11446) );
  AOI21_X1 U13885 ( .B1(n11447), .B2(n13112), .A(n11446), .ZN(P3_U3273) );
  OAI22_X1 U13886 ( .A1(n12997), .A2(n11449), .B1(n11448), .B2(n12946), .ZN(
        n11452) );
  MUX2_X1 U13887 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n11450), .S(n15334), .Z(
        n11451) );
  AOI211_X1 U13888 ( .C1(n12999), .C2(n11453), .A(n11452), .B(n11451), .ZN(
        n11454) );
  INV_X1 U13889 ( .A(n11454), .ZN(P3_U3228) );
  XOR2_X1 U13890 ( .A(n11459), .B(n11455), .Z(n14861) );
  INV_X1 U13891 ( .A(n11456), .ZN(n11457) );
  AOI21_X1 U13892 ( .B1(n11459), .B2(n11458), .A(n11457), .ZN(n11462) );
  OR2_X1 U13893 ( .A1(n11591), .A2(n14353), .ZN(n11461) );
  NAND2_X1 U13894 ( .A1(n14082), .A2(n14362), .ZN(n11460) );
  AND2_X1 U13895 ( .A1(n11461), .A2(n11460), .ZN(n11603) );
  OAI21_X1 U13896 ( .B1(n11462), .B2(n14348), .A(n11603), .ZN(n14856) );
  INV_X1 U13897 ( .A(n14856), .ZN(n11463) );
  MUX2_X1 U13898 ( .A(n11464), .B(n11463), .S(n14393), .Z(n11468) );
  XNOR2_X1 U13899 ( .A(n11681), .B(n11596), .ZN(n14858) );
  INV_X1 U13900 ( .A(n11605), .ZN(n11465) );
  OAI22_X1 U13901 ( .A1(n14394), .A2(n11596), .B1(n14386), .B2(n11465), .ZN(
        n11466) );
  AOI21_X1 U13902 ( .B1(n14858), .B2(n14397), .A(n11466), .ZN(n11467) );
  OAI211_X1 U13903 ( .C1(n14861), .C2(n14400), .A(n11468), .B(n11467), .ZN(
        P1_U3288) );
  XNOR2_X1 U13904 ( .A(n11469), .B(n11470), .ZN(n14868) );
  XNOR2_X1 U13905 ( .A(n11471), .B(n11470), .ZN(n11472) );
  AOI222_X1 U13906 ( .A1(n14384), .A2(n11472), .B1(n14083), .B2(n14364), .C1(
        n14081), .C2(n14362), .ZN(n14867) );
  MUX2_X1 U13907 ( .A(n10615), .B(n14867), .S(n14393), .Z(n11479) );
  NAND2_X1 U13908 ( .A1(n11473), .A2(n14864), .ZN(n11474) );
  AND2_X1 U13909 ( .A1(n11503), .A2(n11474), .ZN(n14865) );
  INV_X1 U13910 ( .A(n11856), .ZN(n11475) );
  OAI22_X1 U13911 ( .A1(n14394), .A2(n11476), .B1(n11475), .B2(n14386), .ZN(
        n11477) );
  AOI21_X1 U13912 ( .B1(n14865), .B2(n14397), .A(n11477), .ZN(n11478) );
  OAI211_X1 U13913 ( .C1(n14400), .C2(n14868), .A(n11479), .B(n11478), .ZN(
        P1_U3287) );
  XNOR2_X1 U13914 ( .A(n11481), .B(n11480), .ZN(n11694) );
  OAI21_X1 U13915 ( .B1(n11484), .B2(n11483), .A(n11482), .ZN(n11486) );
  AOI21_X1 U13916 ( .B1(n11486), .B2(n9268), .A(n11485), .ZN(n11487) );
  OAI21_X1 U13917 ( .B1(n11694), .B2(n9219), .A(n11487), .ZN(n11695) );
  NAND2_X1 U13918 ( .A1(n11695), .A2(n7490), .ZN(n11494) );
  AOI211_X1 U13919 ( .C1(n11701), .C2(n11488), .A(n12562), .B(n11615), .ZN(
        n11696) );
  NOR2_X1 U13920 ( .A1(n6932), .A2(n13636), .ZN(n11492) );
  OAI22_X1 U13921 ( .A1(n7490), .A2(n11490), .B1(n11489), .B2(n13419), .ZN(
        n11491) );
  AOI211_X1 U13922 ( .C1(n11696), .C2(n14664), .A(n11492), .B(n11491), .ZN(
        n11493) );
  OAI211_X1 U13923 ( .C1(n11694), .C2(n13495), .A(n11494), .B(n11493), .ZN(
        P2_U3256) );
  XOR2_X1 U13924 ( .A(n11495), .B(n11497), .Z(n14871) );
  XOR2_X1 U13925 ( .A(n11497), .B(n11496), .Z(n11501) );
  NAND2_X1 U13926 ( .A1(n14082), .A2(n14364), .ZN(n11499) );
  NAND2_X1 U13927 ( .A1(n14080), .A2(n14362), .ZN(n11498) );
  AND2_X1 U13928 ( .A1(n11499), .A2(n11498), .ZN(n12083) );
  INV_X1 U13929 ( .A(n12083), .ZN(n11500) );
  AOI21_X1 U13930 ( .B1(n11501), .B2(n14384), .A(n11500), .ZN(n14874) );
  MUX2_X1 U13931 ( .A(n14874), .B(n11502), .S(n14377), .Z(n11508) );
  AND2_X1 U13932 ( .A1(n11503), .A2(n12089), .ZN(n11504) );
  NOR2_X1 U13933 ( .A1(n11657), .A2(n11504), .ZN(n14872) );
  INV_X1 U13934 ( .A(n12089), .ZN(n14876) );
  INV_X1 U13935 ( .A(n11505), .ZN(n12080) );
  OAI22_X1 U13936 ( .A1(n14394), .A2(n14876), .B1(n14386), .B2(n12080), .ZN(
        n11506) );
  AOI21_X1 U13937 ( .B1(n14872), .B2(n14397), .A(n11506), .ZN(n11507) );
  OAI211_X1 U13938 ( .C1(n14400), .C2(n14871), .A(n11508), .B(n11507), .ZN(
        P1_U3286) );
  NOR2_X1 U13939 ( .A1(n11534), .A2(n6597), .ZN(n11510) );
  NAND2_X1 U13940 ( .A1(n15256), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11512) );
  OR2_X1 U13941 ( .A1(n15256), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11511) );
  NAND2_X1 U13942 ( .A1(n11512), .A2(n11511), .ZN(n15259) );
  NOR2_X1 U13943 ( .A1(n11544), .A2(n11513), .ZN(n11515) );
  INV_X1 U13944 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15270) );
  NAND2_X1 U13945 ( .A1(n11830), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11823) );
  OAI21_X1 U13946 ( .B1(n11830), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11823), 
        .ZN(n11517) );
  INV_X1 U13947 ( .A(n11824), .ZN(n11516) );
  AOI21_X1 U13948 ( .B1(n11518), .B2(n11517), .A(n11516), .ZN(n11557) );
  NAND2_X1 U13949 ( .A1(n15256), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11523) );
  MUX2_X1 U13950 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n15369), .S(n15256), .Z(
        n15255) );
  NAND2_X1 U13951 ( .A1(n11520), .A2(n11519), .ZN(n11522) );
  NAND2_X1 U13952 ( .A1(n11522), .A2(n11521), .ZN(n15254) );
  NAND2_X1 U13953 ( .A1(n15284), .A2(n11524), .ZN(n11525) );
  NAND2_X1 U13954 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15283), .ZN(n15282) );
  NAND2_X1 U13955 ( .A1(n11525), .A2(n15282), .ZN(n11527) );
  INV_X1 U13956 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11546) );
  MUX2_X1 U13957 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11546), .S(n11830), .Z(
        n11526) );
  NAND2_X1 U13958 ( .A1(n11526), .A2(n11527), .ZN(n11831) );
  OAI21_X1 U13959 ( .B1(n11527), .B2(n11526), .A(n11831), .ZN(n11530) );
  NAND2_X1 U13960 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11944)
         );
  NAND2_X1 U13961 ( .A1(n15245), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11528) );
  OAI211_X1 U13962 ( .C1(n15285), .C2(n11830), .A(n11944), .B(n11528), .ZN(
        n11529) );
  AOI21_X1 U13963 ( .B1(n11530), .B2(n15287), .A(n11529), .ZN(n11556) );
  NAND2_X1 U13964 ( .A1(n11532), .A2(n11531), .ZN(n11537) );
  INV_X1 U13965 ( .A(n11533), .ZN(n11535) );
  NAND2_X1 U13966 ( .A1(n11535), .A2(n11534), .ZN(n11536) );
  NAND2_X1 U13967 ( .A1(n11537), .A2(n11536), .ZN(n15253) );
  MUX2_X1 U13968 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12823), .Z(n11538) );
  INV_X1 U13969 ( .A(n15256), .ZN(n11539) );
  XNOR2_X1 U13970 ( .A(n11538), .B(n11539), .ZN(n15252) );
  NAND2_X1 U13971 ( .A1(n15253), .A2(n15252), .ZN(n11542) );
  INV_X1 U13972 ( .A(n11538), .ZN(n11540) );
  NAND2_X1 U13973 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  NAND2_X1 U13974 ( .A1(n11542), .A2(n11541), .ZN(n15278) );
  MUX2_X1 U13975 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12823), .Z(n11543) );
  NAND2_X1 U13976 ( .A1(n11543), .A2(n15284), .ZN(n15272) );
  INV_X1 U13977 ( .A(n11543), .ZN(n11545) );
  AND2_X1 U13978 ( .A1(n11545), .A2(n11544), .ZN(n15274) );
  INV_X1 U13979 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11547) );
  MUX2_X1 U13980 ( .A(n11547), .B(n11546), .S(n12823), .Z(n11549) );
  NAND2_X1 U13981 ( .A1(n11549), .A2(n11548), .ZN(n11826) );
  INV_X1 U13982 ( .A(n11549), .ZN(n11550) );
  NAND2_X1 U13983 ( .A1(n11550), .A2(n11830), .ZN(n11551) );
  AND2_X1 U13984 ( .A1(n11826), .A2(n11551), .ZN(n11552) );
  OAI21_X1 U13985 ( .B1(n15276), .B2(n15274), .A(n11552), .ZN(n11827) );
  INV_X1 U13986 ( .A(n11827), .ZN(n11554) );
  NOR3_X1 U13987 ( .A1(n15276), .A2(n15274), .A3(n11552), .ZN(n11553) );
  OAI21_X1 U13988 ( .B1(n11554), .B2(n11553), .A(n15280), .ZN(n11555) );
  OAI211_X1 U13989 ( .C1(n11557), .C2(n15291), .A(n11556), .B(n11555), .ZN(
        P3_U3192) );
  XNOR2_X1 U13990 ( .A(n11559), .B(n11558), .ZN(n11566) );
  OAI21_X1 U13991 ( .B1(n11562), .B2(n11561), .A(n11560), .ZN(n11564) );
  AOI21_X1 U13992 ( .B1(n11564), .B2(n14879), .A(n11563), .ZN(n11565) );
  OAI21_X1 U13993 ( .B1(n14348), .B2(n11566), .A(n11565), .ZN(n14847) );
  NAND2_X1 U13994 ( .A1(n14847), .A2(n14393), .ZN(n11572) );
  INV_X1 U13995 ( .A(n14397), .ZN(n14319) );
  OAI21_X1 U13996 ( .B1(n11568), .B2(n14845), .A(n11567), .ZN(n14846) );
  INV_X1 U13997 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11569) );
  OAI22_X1 U13998 ( .A1(n14319), .A2(n14846), .B1(n11569), .B2(n14386), .ZN(
        n11570) );
  AOI21_X1 U13999 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n14377), .A(n11570), .ZN(
        n11571) );
  OAI211_X1 U14000 ( .C1(n14845), .C2(n14394), .A(n11572), .B(n11571), .ZN(
        P1_U3291) );
  INV_X1 U14001 ( .A(n13365), .ZN(n15047) );
  OAI222_X1 U14002 ( .A1(n13783), .A2(n11573), .B1(n13781), .B2(n11574), .C1(
        n15047), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U14003 ( .A(n14162), .ZN(n14156) );
  OAI222_X1 U14004 ( .A1(n14527), .A2(n7056), .B1(n14525), .B2(n11574), .C1(
        n14156), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI22_X1 U14005 ( .A1(n12997), .A2(n15169), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n12946), .ZN(n11577) );
  MUX2_X1 U14006 ( .A(n11575), .B(P3_REG2_REG_3__SCAN_IN), .S(n13001), .Z(
        n11576) );
  AOI211_X1 U14007 ( .C1(n12999), .C2(n11578), .A(n11577), .B(n11576), .ZN(
        n11579) );
  INV_X1 U14008 ( .A(n11579), .ZN(P3_U3230) );
  INV_X1 U14009 ( .A(n11580), .ZN(n11582) );
  AOI22_X1 U14010 ( .A1(n13932), .A2(n14085), .B1(n13933), .B2(n13916), .ZN(
        n11586) );
  AOI22_X1 U14011 ( .A1(n14085), .A2(n11847), .B1(n13935), .B2(n13916), .ZN(
        n11585) );
  XNOR2_X1 U14012 ( .A(n11585), .B(n12151), .ZN(n11587) );
  XOR2_X1 U14013 ( .A(n11586), .B(n11587), .Z(n13914) );
  NOR2_X1 U14014 ( .A1(n14850), .A2(n13855), .ZN(n11589) );
  AOI21_X1 U14015 ( .B1(n14084), .B2(n13932), .A(n11589), .ZN(n11593) );
  OAI22_X1 U14016 ( .A1(n11591), .A2(n13855), .B1(n14850), .B2(n13838), .ZN(
        n11592) );
  XOR2_X1 U14017 ( .A(n12151), .B(n11592), .Z(n11627) );
  NOR2_X1 U14018 ( .A1(n11626), .A2(n11627), .ZN(n11625) );
  AND2_X1 U14019 ( .A1(n11594), .A2(n11590), .ZN(n11595) );
  NOR2_X2 U14020 ( .A1(n11625), .A2(n11595), .ZN(n11844) );
  OAI22_X1 U14021 ( .A1(n11854), .A2(n13855), .B1(n11596), .B2(n13838), .ZN(
        n11597) );
  XOR2_X1 U14022 ( .A(n12151), .B(n11597), .Z(n11843) );
  AOI22_X1 U14023 ( .A1(n13932), .A2(n14083), .B1(n13933), .B2(n11600), .ZN(
        n11845) );
  XNOR2_X1 U14024 ( .A(n11843), .B(n11845), .ZN(n11598) );
  XNOR2_X1 U14025 ( .A(n11844), .B(n11598), .ZN(n11607) );
  AND2_X1 U14026 ( .A1(n11600), .A2(n14882), .ZN(n14857) );
  NAND2_X1 U14027 ( .A1(n12148), .A2(n14857), .ZN(n11601) );
  OAI211_X1 U14028 ( .C1(n11603), .C2(n14049), .A(n11602), .B(n11601), .ZN(
        n11604) );
  AOI21_X1 U14029 ( .B1(n11605), .B2(n14063), .A(n11604), .ZN(n11606) );
  OAI21_X1 U14030 ( .B1(n11607), .B2(n14065), .A(n11606), .ZN(P1_U3227) );
  OAI21_X1 U14031 ( .B1(n11613), .B2(n11609), .A(n11608), .ZN(n11610) );
  NAND2_X1 U14032 ( .A1(n11610), .A2(n9268), .ZN(n11612) );
  AOI22_X1 U14033 ( .A1(n13612), .A2(n13262), .B1(n13260), .B2(n13614), .ZN(
        n11611) );
  NAND2_X1 U14034 ( .A1(n11612), .A2(n11611), .ZN(n15143) );
  INV_X1 U14035 ( .A(n15143), .ZN(n11624) );
  XNOR2_X1 U14036 ( .A(n11614), .B(n11613), .ZN(n15138) );
  OAI21_X1 U14037 ( .B1(n11615), .B2(n15141), .A(n6483), .ZN(n11616) );
  OR2_X1 U14038 ( .A1(n11792), .A2(n11616), .ZN(n15139) );
  OAI22_X1 U14039 ( .A1(n7490), .A2(n11618), .B1(n11617), .B2(n13419), .ZN(
        n11619) );
  AOI21_X1 U14040 ( .B1(n11620), .B2(n14655), .A(n11619), .ZN(n11621) );
  OAI21_X1 U14041 ( .B1(n15139), .B2(n13525), .A(n11621), .ZN(n11622) );
  AOI21_X1 U14042 ( .B1(n15138), .B2(n14665), .A(n11622), .ZN(n11623) );
  OAI21_X1 U14043 ( .B1(n11624), .B2(n14668), .A(n11623), .ZN(P2_U3255) );
  AOI211_X1 U14044 ( .C1(n11627), .C2(n11626), .A(n14065), .B(n11625), .ZN(
        n11633) );
  NAND2_X1 U14045 ( .A1(n14055), .A2(n14083), .ZN(n11628) );
  NAND2_X1 U14046 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14779) );
  OAI211_X1 U14047 ( .C1(n11629), .C2(n14057), .A(n11628), .B(n14779), .ZN(
        n11632) );
  OAI22_X1 U14048 ( .A1(n14059), .A2(n14850), .B1(n11630), .B2(n14696), .ZN(
        n11631) );
  OR3_X1 U14049 ( .A1(n11633), .A2(n11632), .A3(n11631), .ZN(P1_U3230) );
  NAND2_X1 U14050 ( .A1(n11634), .A2(n14916), .ZN(n11635) );
  OAI21_X1 U14051 ( .B1(n14916), .B2(n11636), .A(n11635), .ZN(P1_U3531) );
  OAI21_X1 U14052 ( .B1(n11638), .B2(n11642), .A(n11637), .ZN(n15354) );
  INV_X1 U14053 ( .A(n15354), .ZN(n11650) );
  INV_X1 U14054 ( .A(n11639), .ZN(n11640) );
  AOI21_X1 U14055 ( .B1(n11642), .B2(n11641), .A(n11640), .ZN(n11645) );
  INV_X1 U14056 ( .A(n12912), .ZN(n15324) );
  OAI22_X1 U14057 ( .A1(n11939), .A2(n15303), .B1(n11809), .B2(n15302), .ZN(
        n11643) );
  AOI21_X1 U14058 ( .B1(n15354), .B2(n15324), .A(n11643), .ZN(n11644) );
  OAI21_X1 U14059 ( .B1(n11645), .B2(n15308), .A(n11644), .ZN(n15352) );
  NAND2_X1 U14060 ( .A1(n15352), .A2(n15334), .ZN(n11649) );
  INV_X1 U14061 ( .A(n11646), .ZN(n12620) );
  OAI22_X1 U14062 ( .A1(n12997), .A2(n15351), .B1(n12620), .B2(n12946), .ZN(
        n11647) );
  AOI21_X1 U14063 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13001), .A(n11647), .ZN(
        n11648) );
  OAI211_X1 U14064 ( .C1(n11650), .C2(n11739), .A(n11649), .B(n11648), .ZN(
        P3_U3225) );
  XNOR2_X1 U14065 ( .A(n11651), .B(n11652), .ZN(n14887) );
  XNOR2_X1 U14066 ( .A(n11654), .B(n11653), .ZN(n11656) );
  AOI22_X1 U14067 ( .A1(n14362), .A2(n14079), .B1(n14081), .B2(n14364), .ZN(
        n12074) );
  INV_X1 U14068 ( .A(n12074), .ZN(n11655) );
  AOI21_X1 U14069 ( .B1(n11656), .B2(n14384), .A(n11655), .ZN(n14886) );
  MUX2_X1 U14070 ( .A(n14886), .B(n10747), .S(n14377), .Z(n11661) );
  XNOR2_X1 U14071 ( .A(n11657), .B(n14881), .ZN(n14884) );
  INV_X1 U14072 ( .A(n12076), .ZN(n11658) );
  OAI22_X1 U14073 ( .A1(n12079), .A2(n14394), .B1(n11658), .B2(n14386), .ZN(
        n11659) );
  AOI21_X1 U14074 ( .B1(n14884), .B2(n14397), .A(n11659), .ZN(n11660) );
  OAI211_X1 U14075 ( .C1(n14400), .C2(n14887), .A(n11661), .B(n11660), .ZN(
        P1_U3285) );
  INV_X1 U14076 ( .A(n11662), .ZN(n11663) );
  NAND2_X1 U14077 ( .A1(n11664), .A2(n11663), .ZN(n11668) );
  XNOR2_X1 U14078 ( .A(n11902), .B(n12547), .ZN(n11666) );
  NAND2_X1 U14079 ( .A1(n13260), .A2(n12562), .ZN(n11665) );
  NOR2_X1 U14080 ( .A1(n11666), .A2(n11665), .ZN(n12104) );
  AOI21_X1 U14081 ( .B1(n11666), .B2(n11665), .A(n12104), .ZN(n11667) );
  OAI211_X1 U14082 ( .C1(n11668), .C2(n11667), .A(n12106), .B(n13243), .ZN(
        n11673) );
  INV_X1 U14083 ( .A(n11669), .ZN(n11794) );
  OAI22_X1 U14084 ( .A1(n11788), .A2(n14921), .B1(n14920), .B2(n11787), .ZN(
        n11670) );
  AOI211_X1 U14085 ( .C1(n11794), .C2(n13235), .A(n11671), .B(n11670), .ZN(
        n11672) );
  OAI211_X1 U14086 ( .C1(n11899), .C2(n13252), .A(n11673), .B(n11672), .ZN(
        P2_U3208) );
  OAI22_X1 U14087 ( .A1(n12997), .A2(n11674), .B1(n15168), .B2(n12946), .ZN(
        n11677) );
  MUX2_X1 U14088 ( .A(n11675), .B(P3_REG2_REG_7__SCAN_IN), .S(n13001), .Z(
        n11676) );
  AOI211_X1 U14089 ( .C1(n12999), .C2(n11678), .A(n11677), .B(n11676), .ZN(
        n11679) );
  INV_X1 U14090 ( .A(n11679), .ZN(P3_U3226) );
  XOR2_X1 U14091 ( .A(n6496), .B(n11686), .Z(n14854) );
  OAI21_X1 U14092 ( .B1(n11682), .B2(n14850), .A(n11681), .ZN(n14851) );
  INV_X1 U14093 ( .A(n14386), .ZN(n14369) );
  AOI22_X1 U14094 ( .A1(n14322), .A2(n11684), .B1(n11683), .B2(n14369), .ZN(
        n11685) );
  OAI21_X1 U14095 ( .B1(n14319), .B2(n14851), .A(n11685), .ZN(n11692) );
  XNOR2_X1 U14096 ( .A(n11687), .B(n11686), .ZN(n11688) );
  NAND2_X1 U14097 ( .A1(n11688), .A2(n14384), .ZN(n11690) );
  AOI22_X1 U14098 ( .A1(n14362), .A2(n14083), .B1(n14085), .B2(n14364), .ZN(
        n11689) );
  NAND2_X1 U14099 ( .A1(n11690), .A2(n11689), .ZN(n14852) );
  MUX2_X1 U14100 ( .A(n14852), .B(P1_REG2_REG_4__SCAN_IN), .S(n14377), .Z(
        n11691) );
  AOI211_X1 U14101 ( .C1(n14325), .C2(n14854), .A(n11692), .B(n11691), .ZN(
        n11693) );
  INV_X1 U14102 ( .A(n11693), .ZN(P1_U3289) );
  INV_X1 U14103 ( .A(n11694), .ZN(n11697) );
  INV_X1 U14104 ( .A(n15123), .ZN(n15135) );
  AOI211_X1 U14105 ( .C1(n11697), .C2(n15135), .A(n11696), .B(n11695), .ZN(
        n11703) );
  INV_X1 U14106 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11698) );
  NOR2_X1 U14107 ( .A1(n15147), .A2(n11698), .ZN(n11699) );
  AOI21_X1 U14108 ( .B1(n11701), .B2(n13749), .A(n11699), .ZN(n11700) );
  OAI21_X1 U14109 ( .B1(n11703), .B2(n15145), .A(n11700), .ZN(P2_U3457) );
  AOI22_X1 U14110 ( .A1(n11701), .A2(n13688), .B1(n15154), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11702) );
  OAI21_X1 U14111 ( .B1(n11703), .B2(n15154), .A(n11702), .ZN(P2_U3508) );
  INV_X1 U14112 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11710) );
  INV_X1 U14113 ( .A(n11704), .ZN(n11705) );
  AOI22_X1 U14114 ( .A1(n14325), .A2(n11706), .B1(n14322), .B2(n11705), .ZN(
        n11709) );
  AOI22_X1 U14115 ( .A1(n14397), .A2(n11707), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14369), .ZN(n11708) );
  OAI211_X1 U14116 ( .C1(n11710), .C2(n14393), .A(n11709), .B(n11708), .ZN(
        n11711) );
  AOI21_X1 U14117 ( .B1(n11712), .B2(n14393), .A(n11711), .ZN(n11713) );
  INV_X1 U14118 ( .A(n11713), .ZN(P1_U3292) );
  XNOR2_X1 U14119 ( .A(n6494), .B(n11715), .ZN(n14891) );
  INV_X1 U14120 ( .A(n14891), .ZN(n11727) );
  XNOR2_X1 U14121 ( .A(n11716), .B(n11717), .ZN(n11718) );
  NAND2_X1 U14122 ( .A1(n11718), .A2(n14384), .ZN(n11720) );
  AOI22_X1 U14123 ( .A1(n14362), .A2(n14078), .B1(n14080), .B2(n14364), .ZN(
        n11719) );
  NAND2_X1 U14124 ( .A1(n11720), .A2(n11719), .ZN(n14896) );
  NAND2_X1 U14125 ( .A1(n11721), .A2(n12153), .ZN(n11722) );
  NAND2_X1 U14126 ( .A1(n11868), .A2(n11722), .ZN(n14893) );
  AOI22_X1 U14127 ( .A1(n14377), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n12163), 
        .B2(n14369), .ZN(n11724) );
  NAND2_X1 U14128 ( .A1(n12153), .A2(n14322), .ZN(n11723) );
  OAI211_X1 U14129 ( .C1(n14893), .C2(n14319), .A(n11724), .B(n11723), .ZN(
        n11725) );
  AOI21_X1 U14130 ( .B1(n14896), .B2(n14393), .A(n11725), .ZN(n11726) );
  OAI21_X1 U14131 ( .B1(n14400), .B2(n11727), .A(n11726), .ZN(P1_U3284) );
  XNOR2_X1 U14132 ( .A(n11728), .B(n11730), .ZN(n15360) );
  OAI211_X1 U14133 ( .C1(n11731), .C2(n11730), .A(n11729), .B(n15317), .ZN(
        n11734) );
  OAI22_X1 U14134 ( .A1(n12334), .A2(n15303), .B1(n11816), .B2(n15302), .ZN(
        n11732) );
  INV_X1 U14135 ( .A(n11732), .ZN(n11733) );
  OAI211_X1 U14136 ( .C1(n12912), .C2(n15360), .A(n11734), .B(n11733), .ZN(
        n15362) );
  NAND2_X1 U14137 ( .A1(n15362), .A2(n15334), .ZN(n11738) );
  INV_X1 U14138 ( .A(n11820), .ZN(n11735) );
  OAI22_X1 U14139 ( .A1(n12997), .A2(n15358), .B1(n11735), .B2(n12946), .ZN(
        n11736) );
  AOI21_X1 U14140 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n13001), .A(n11736), .ZN(
        n11737) );
  OAI211_X1 U14141 ( .C1(n15360), .C2(n11739), .A(n11738), .B(n11737), .ZN(
        P3_U3224) );
  NAND2_X1 U14142 ( .A1(n11740), .A2(n13112), .ZN(n11742) );
  OAI211_X1 U14143 ( .C1(n8560), .C2(n13125), .A(n11742), .B(n11741), .ZN(
        P3_U3272) );
  OAI222_X1 U14144 ( .A1(n14527), .A2(n11744), .B1(n14525), .B2(n11747), .C1(
        n11743), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U14145 ( .A(n11745), .ZN(n12420) );
  OAI222_X1 U14146 ( .A1(n14527), .A2(n11746), .B1(n14521), .B2(n12420), .C1(
        P1_U3086), .C2(n14172), .ZN(P1_U3336) );
  OAI222_X1 U14147 ( .A1(n13783), .A2(n11748), .B1(P2_U3088), .B2(n8803), .C1(
        n13781), .C2(n11747), .ZN(P2_U3307) );
  OAI211_X1 U14148 ( .C1(n11752), .C2(n11750), .A(n11749), .B(n15317), .ZN(
        n11751) );
  AOI22_X1 U14149 ( .A1(n12713), .A2(n12962), .B1(n12963), .B2(n12715), .ZN(
        n11945) );
  NAND2_X1 U14150 ( .A1(n11751), .A2(n11945), .ZN(n11930) );
  INV_X1 U14151 ( .A(n11930), .ZN(n11757) );
  XOR2_X1 U14152 ( .A(n11753), .B(n11752), .Z(n11931) );
  AOI22_X1 U14153 ( .A1(n13001), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15331), 
        .B2(n11937), .ZN(n11754) );
  OAI21_X1 U14154 ( .B1(n11936), .B2(n12997), .A(n11754), .ZN(n11755) );
  AOI21_X1 U14155 ( .B1(n11931), .B2(n12999), .A(n11755), .ZN(n11756) );
  OAI21_X1 U14156 ( .B1(n11757), .B2(n13001), .A(n11756), .ZN(P3_U3223) );
  INV_X1 U14157 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11758) );
  NAND2_X1 U14158 ( .A1(n14151), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11761) );
  MUX2_X1 U14159 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11758), .S(n14151), .Z(
        n14144) );
  NAND2_X1 U14160 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11775), .ZN(n11760) );
  NAND2_X1 U14161 ( .A1(n11760), .A2(n11759), .ZN(n14145) );
  NAND2_X1 U14162 ( .A1(n14144), .A2(n14145), .ZN(n14143) );
  NAND2_X1 U14163 ( .A1(n11761), .A2(n14143), .ZN(n11762) );
  INV_X1 U14164 ( .A(n11762), .ZN(n11764) );
  INV_X1 U14165 ( .A(n14803), .ZN(n11763) );
  XNOR2_X1 U14166 ( .A(n11762), .B(n14803), .ZN(n14797) );
  NOR2_X1 U14167 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14797), .ZN(n14796) );
  AOI21_X1 U14168 ( .B1(n11764), .B2(n11763), .A(n14796), .ZN(n11768) );
  INV_X1 U14169 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11766) );
  NOR2_X1 U14170 ( .A1(n11772), .A2(n11766), .ZN(n11765) );
  AOI21_X1 U14171 ( .B1(n11766), .B2(n11772), .A(n11765), .ZN(n11767) );
  NAND2_X1 U14172 ( .A1(n11767), .A2(n11768), .ZN(n11963) );
  OAI211_X1 U14173 ( .C1(n11768), .C2(n11767), .A(n14771), .B(n11963), .ZN(
        n11771) );
  NAND2_X1 U14174 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13980)
         );
  INV_X1 U14175 ( .A(n13980), .ZN(n11769) );
  AOI21_X1 U14176 ( .B1(n14757), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11769), 
        .ZN(n11770) );
  OAI211_X1 U14177 ( .C1(n14775), .C2(n11772), .A(n11771), .B(n11770), .ZN(
        n11782) );
  OR2_X1 U14178 ( .A1(n14151), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11776) );
  INV_X1 U14179 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11773) );
  MUX2_X1 U14180 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11773), .S(n14151), .Z(
        n14149) );
  NAND2_X1 U14181 ( .A1(n14149), .A2(n14148), .ZN(n14147) );
  NAND2_X1 U14182 ( .A1(n11776), .A2(n14147), .ZN(n11777) );
  INV_X1 U14183 ( .A(n11777), .ZN(n11778) );
  XNOR2_X1 U14184 ( .A(n11777), .B(n14803), .ZN(n14800) );
  INV_X1 U14185 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U14186 ( .A1(n14800), .A2(n14799), .ZN(n14798) );
  OAI21_X1 U14187 ( .B1(n11778), .B2(n14803), .A(n14798), .ZN(n11780) );
  XNOR2_X1 U14188 ( .A(n11965), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11779) );
  NOR2_X1 U14189 ( .A1(n11779), .A2(n11780), .ZN(n11960) );
  AOI211_X1 U14190 ( .C1(n11780), .C2(n11779), .A(n11960), .B(n14168), .ZN(
        n11781) );
  OR2_X1 U14191 ( .A1(n11782), .A2(n11781), .ZN(P1_U3259) );
  XOR2_X1 U14192 ( .A(n11783), .B(n11785), .Z(n11894) );
  OAI21_X1 U14193 ( .B1(n11786), .B2(n11785), .A(n11784), .ZN(n11790) );
  OAI22_X1 U14194 ( .A1(n11788), .A2(n13539), .B1(n11787), .B2(n13537), .ZN(
        n11789) );
  AOI21_X1 U14195 ( .B1(n11790), .B2(n9268), .A(n11789), .ZN(n11791) );
  OAI21_X1 U14196 ( .B1(n11894), .B2(n9219), .A(n11791), .ZN(n11895) );
  NAND2_X1 U14197 ( .A1(n11895), .A2(n7490), .ZN(n11798) );
  INV_X1 U14198 ( .A(n11792), .ZN(n11793) );
  AOI211_X1 U14199 ( .C1(n11902), .C2(n11793), .A(n12562), .B(n6633), .ZN(
        n11896) );
  INV_X1 U14200 ( .A(n13419), .ZN(n14654) );
  AOI22_X1 U14201 ( .A1(n14668), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n14654), 
        .B2(n11794), .ZN(n11795) );
  OAI21_X1 U14202 ( .B1(n11899), .B2(n13636), .A(n11795), .ZN(n11796) );
  AOI21_X1 U14203 ( .B1(n11896), .B2(n14664), .A(n11796), .ZN(n11797) );
  OAI211_X1 U14204 ( .C1(n11894), .C2(n13495), .A(n11798), .B(n11797), .ZN(
        P2_U3254) );
  XNOR2_X1 U14205 ( .A(n11799), .B(n12485), .ZN(n11938) );
  XNOR2_X1 U14206 ( .A(n11938), .B(n11939), .ZN(n11815) );
  XNOR2_X1 U14207 ( .A(n12618), .B(n12485), .ZN(n11813) );
  XNOR2_X1 U14208 ( .A(n11801), .B(n12485), .ZN(n11807) );
  INV_X1 U14209 ( .A(n11802), .ZN(n11804) );
  XOR2_X1 U14210 ( .A(n12717), .B(n11807), .Z(n15182) );
  XNOR2_X1 U14211 ( .A(n11808), .B(n12485), .ZN(n15158) );
  INV_X1 U14212 ( .A(n15158), .ZN(n11811) );
  XNOR2_X1 U14213 ( .A(n12716), .B(n11813), .ZN(n12615) );
  AOI21_X1 U14214 ( .B1(n11815), .B2(n11814), .A(n11941), .ZN(n11822) );
  OAI22_X1 U14215 ( .A1(n11817), .A2(n12334), .B1(n11816), .B2(n12694), .ZN(
        n11819) );
  OAI22_X1 U14216 ( .A1(n15170), .A2(n15358), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8586), .ZN(n11818) );
  AOI211_X1 U14217 ( .C1(n12696), .C2(n11820), .A(n11819), .B(n11818), .ZN(
        n11821) );
  OAI21_X1 U14218 ( .B1(n11822), .B2(n15172), .A(n11821), .ZN(P3_U3171) );
  INV_X1 U14219 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11955) );
  AOI21_X1 U14220 ( .B1(n11955), .B2(n11825), .A(n12001), .ZN(n11842) );
  NAND2_X1 U14221 ( .A1(n11827), .A2(n11826), .ZN(n11829) );
  MUX2_X1 U14222 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12823), .Z(n12014) );
  XNOR2_X1 U14223 ( .A(n12014), .B(n12015), .ZN(n11828) );
  NAND2_X1 U14224 ( .A1(n11829), .A2(n11828), .ZN(n12019) );
  OAI21_X1 U14225 ( .B1(n11829), .B2(n11828), .A(n12019), .ZN(n11840) );
  NAND2_X1 U14226 ( .A1(n11830), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U14227 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11833), .ZN(n12008) );
  OAI21_X1 U14228 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11833), .A(n12008), 
        .ZN(n11834) );
  NAND2_X1 U14229 ( .A1(n11834), .A2(n15287), .ZN(n11838) );
  NOR2_X1 U14230 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11835), .ZN(n11836) );
  AOI21_X1 U14231 ( .B1(n15245), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11836), 
        .ZN(n11837) );
  OAI211_X1 U14232 ( .C1(n15285), .C2(n12007), .A(n11838), .B(n11837), .ZN(
        n11839) );
  AOI21_X1 U14233 ( .B1(n15280), .B2(n11840), .A(n11839), .ZN(n11841) );
  OAI21_X1 U14234 ( .B1(n11842), .B2(n15291), .A(n11841), .ZN(P3_U3193) );
  INV_X1 U14235 ( .A(n11845), .ZN(n11846) );
  AOI22_X1 U14236 ( .A1(n13932), .A2(n14082), .B1(n14864), .B2(n13933), .ZN(
        n12054) );
  NAND2_X1 U14237 ( .A1(n14864), .A2(n13935), .ZN(n11849) );
  NAND2_X1 U14238 ( .A1(n14082), .A2(n13933), .ZN(n11848) );
  NAND2_X1 U14239 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  XNOR2_X1 U14240 ( .A(n11850), .B(n12151), .ZN(n12052) );
  XOR2_X1 U14241 ( .A(n12054), .B(n12052), .Z(n12055) );
  XNOR2_X1 U14242 ( .A(n12056), .B(n12055), .ZN(n11859) );
  OR2_X1 U14243 ( .A1(n14030), .A2(n11851), .ZN(n11853) );
  OAI211_X1 U14244 ( .C1(n11854), .C2(n14057), .A(n11853), .B(n11852), .ZN(
        n11855) );
  INV_X1 U14245 ( .A(n11855), .ZN(n11858) );
  AOI22_X1 U14246 ( .A1(n11856), .A2(n14063), .B1(n14687), .B2(n14864), .ZN(
        n11857) );
  OAI211_X1 U14247 ( .C1(n11859), .C2(n14065), .A(n11858), .B(n11857), .ZN(
        P1_U3239) );
  AOI21_X1 U14248 ( .B1(n14319), .B2(n14394), .A(n11860), .ZN(n11864) );
  AOI22_X1 U14249 ( .A1(n14377), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14369), .ZN(n11861) );
  OAI21_X1 U14250 ( .B1(n14377), .B2(n11862), .A(n11861), .ZN(n11863) );
  AOI211_X1 U14251 ( .C1(n14325), .C2(n11865), .A(n11864), .B(n11863), .ZN(
        n11866) );
  INV_X1 U14252 ( .A(n11866), .ZN(P1_U3293) );
  XOR2_X1 U14253 ( .A(n11867), .B(n11870), .Z(n14898) );
  AOI211_X1 U14254 ( .C1(n12200), .C2(n11868), .A(n10323), .B(n11887), .ZN(
        n11869) );
  AOI21_X1 U14255 ( .B1(n14362), .B2(n14077), .A(n11869), .ZN(n14900) );
  AOI21_X1 U14256 ( .B1(n11871), .B2(n11870), .A(n14348), .ZN(n11873) );
  AOI22_X1 U14257 ( .A1(n11873), .A2(n11872), .B1(n14364), .B2(n14079), .ZN(
        n14901) );
  OAI21_X1 U14258 ( .B1(n11874), .B2(n14900), .A(n14901), .ZN(n11877) );
  AOI22_X1 U14259 ( .A1(n14377), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n12211), 
        .B2(n14369), .ZN(n11875) );
  OAI21_X1 U14260 ( .B1(n6815), .B2(n14394), .A(n11875), .ZN(n11876) );
  AOI21_X1 U14261 ( .B1(n11877), .B2(n14393), .A(n11876), .ZN(n11878) );
  OAI21_X1 U14262 ( .B1(n14898), .B2(n14400), .A(n11878), .ZN(P1_U3283) );
  OAI222_X1 U14263 ( .A1(n13783), .A2(n11880), .B1(P2_U3088), .B2(n11879), 
        .C1(n13781), .C2(n12588), .ZN(P2_U3306) );
  XNOR2_X1 U14264 ( .A(n11881), .B(n11886), .ZN(n11882) );
  NAND2_X1 U14265 ( .A1(n11882), .A2(n14384), .ZN(n11884) );
  AOI22_X1 U14266 ( .A1(n14362), .A2(n14076), .B1(n14078), .B2(n14364), .ZN(
        n11883) );
  NAND2_X1 U14267 ( .A1(n11884), .A2(n11883), .ZN(n14720) );
  INV_X1 U14268 ( .A(n14720), .ZN(n11893) );
  XNOR2_X1 U14269 ( .A(n11885), .B(n11886), .ZN(n14715) );
  NOR2_X1 U14270 ( .A1(n11887), .A2(n14716), .ZN(n11888) );
  OR2_X1 U14271 ( .A1(n11974), .A2(n11888), .ZN(n14717) );
  AOI22_X1 U14272 ( .A1(n14377), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12314), 
        .B2(n14369), .ZN(n11890) );
  NAND2_X1 U14273 ( .A1(n12319), .A2(n14322), .ZN(n11889) );
  OAI211_X1 U14274 ( .C1(n14717), .C2(n14319), .A(n11890), .B(n11889), .ZN(
        n11891) );
  AOI21_X1 U14275 ( .B1(n14715), .B2(n14325), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14276 ( .B1(n11893), .B2(n14377), .A(n11892), .ZN(P1_U3282) );
  INV_X1 U14277 ( .A(n11894), .ZN(n11897) );
  AOI211_X1 U14278 ( .C1(n15135), .C2(n11897), .A(n11896), .B(n11895), .ZN(
        n11904) );
  INV_X1 U14279 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11898) );
  OAI22_X1 U14280 ( .A1(n11899), .A2(n13754), .B1(n15147), .B2(n11898), .ZN(
        n11900) );
  INV_X1 U14281 ( .A(n11900), .ZN(n11901) );
  OAI21_X1 U14282 ( .B1(n11904), .B2(n15145), .A(n11901), .ZN(P2_U3463) );
  AOI22_X1 U14283 ( .A1(n11902), .A2(n13688), .B1(n15154), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11903) );
  OAI21_X1 U14284 ( .B1(n11904), .B2(n15154), .A(n11903), .ZN(P2_U3510) );
  XNOR2_X1 U14285 ( .A(n11905), .B(n11915), .ZN(n11909) );
  NAND2_X1 U14286 ( .A1(n13259), .A2(n13612), .ZN(n11907) );
  NAND2_X1 U14287 ( .A1(n13257), .A2(n13614), .ZN(n11906) );
  NAND2_X1 U14288 ( .A1(n11907), .A2(n11906), .ZN(n12099) );
  INV_X1 U14289 ( .A(n12099), .ZN(n11908) );
  OAI21_X1 U14290 ( .B1(n11909), .B2(n13593), .A(n11908), .ZN(n12044) );
  INV_X1 U14291 ( .A(n12044), .ZN(n11918) );
  AOI211_X1 U14292 ( .C1(n12115), .C2(n11925), .A(n12562), .B(n6632), .ZN(
        n12045) );
  INV_X1 U14293 ( .A(n12115), .ZN(n11910) );
  NOR2_X1 U14294 ( .A1(n11910), .A2(n13636), .ZN(n11913) );
  OAI22_X1 U14295 ( .A1(n7490), .A2(n11911), .B1(n12101), .B2(n13419), .ZN(
        n11912) );
  AOI211_X1 U14296 ( .C1(n12045), .C2(n14664), .A(n11913), .B(n11912), .ZN(
        n11917) );
  XOR2_X1 U14297 ( .A(n11915), .B(n11914), .Z(n12046) );
  NAND2_X1 U14298 ( .A1(n12046), .A2(n14665), .ZN(n11916) );
  OAI211_X1 U14299 ( .C1(n11918), .C2(n14668), .A(n11917), .B(n11916), .ZN(
        P2_U3252) );
  XOR2_X1 U14300 ( .A(n11919), .B(n11921), .Z(n14674) );
  XOR2_X1 U14301 ( .A(n11921), .B(n11920), .Z(n11923) );
  OAI22_X1 U14302 ( .A1(n14922), .A2(n13539), .B1(n14919), .B2(n13537), .ZN(
        n11922) );
  AOI21_X1 U14303 ( .B1(n11923), .B2(n9268), .A(n11922), .ZN(n11924) );
  OAI21_X1 U14304 ( .B1(n14674), .B2(n9219), .A(n11924), .ZN(n14677) );
  NAND2_X1 U14305 ( .A1(n14677), .A2(n7490), .ZN(n11929) );
  OAI22_X1 U14306 ( .A1(n7490), .A2(n13316), .B1(n14933), .B2(n13419), .ZN(
        n11927) );
  OAI211_X1 U14307 ( .C1(n14676), .C2(n6633), .A(n6483), .B(n11925), .ZN(
        n14675) );
  NOR2_X1 U14308 ( .A1(n14675), .A2(n13525), .ZN(n11926) );
  AOI211_X1 U14309 ( .C1(n14655), .C2(n14931), .A(n11927), .B(n11926), .ZN(
        n11928) );
  OAI211_X1 U14310 ( .C1(n14674), .C2(n13495), .A(n11929), .B(n11928), .ZN(
        P2_U3253) );
  AOI21_X1 U14311 ( .B1(n11931), .B2(n15339), .A(n11930), .ZN(n11933) );
  MUX2_X1 U14312 ( .A(n11546), .B(n11933), .S(n15374), .Z(n11932) );
  OAI21_X1 U14313 ( .B1(n13062), .B2(n11936), .A(n11932), .ZN(P3_U3469) );
  INV_X1 U14314 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11934) );
  MUX2_X1 U14315 ( .A(n11934), .B(n11933), .S(n15365), .Z(n11935) );
  OAI21_X1 U14316 ( .B1(n13110), .B2(n11936), .A(n11935), .ZN(P3_U3420) );
  INV_X1 U14317 ( .A(n11937), .ZN(n11950) );
  XNOR2_X1 U14318 ( .A(n11947), .B(n12485), .ZN(n12170) );
  XNOR2_X1 U14319 ( .A(n12714), .B(n12170), .ZN(n11942) );
  OAI211_X1 U14320 ( .C1(n11943), .C2(n11942), .A(n12172), .B(n15180), .ZN(
        n11949) );
  OAI21_X1 U14321 ( .B1(n11945), .B2(n15189), .A(n11944), .ZN(n11946) );
  AOI21_X1 U14322 ( .B1(n11947), .B2(n15186), .A(n11946), .ZN(n11948) );
  OAI211_X1 U14323 ( .C1(n11950), .C2(n15193), .A(n11949), .B(n11948), .ZN(
        P3_U3157) );
  XNOR2_X1 U14324 ( .A(n11951), .B(n6978), .ZN(n14624) );
  INV_X1 U14325 ( .A(n12712), .ZN(n12175) );
  XNOR2_X1 U14326 ( .A(n11952), .B(n6978), .ZN(n11953) );
  OAI222_X1 U14327 ( .A1(n15303), .A2(n12175), .B1(n15302), .B2(n12334), .C1(
        n11953), .C2(n15308), .ZN(n14626) );
  NAND2_X1 U14328 ( .A1(n14626), .A2(n15334), .ZN(n11958) );
  INV_X1 U14329 ( .A(n12338), .ZN(n11954) );
  OAI22_X1 U14330 ( .A1(n15334), .A2(n11955), .B1(n11954), .B2(n12946), .ZN(
        n11956) );
  AOI21_X1 U14331 ( .B1(n12331), .B2(n14607), .A(n11956), .ZN(n11957) );
  OAI211_X1 U14332 ( .C1(n11088), .C2(n14624), .A(n11958), .B(n11957), .ZN(
        P3_U3222) );
  NAND2_X1 U14333 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13991)
         );
  NAND2_X1 U14334 ( .A1(n14757), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n11959) );
  OAI211_X1 U14335 ( .C1(n14775), .C2(n12244), .A(n13991), .B(n11959), .ZN(
        n11973) );
  XNOR2_X1 U14336 ( .A(n12239), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11961) );
  NOR2_X1 U14337 ( .A1(n11961), .A2(n11962), .ZN(n12238) );
  AOI211_X1 U14338 ( .C1(n11962), .C2(n11961), .A(n12238), .B(n14168), .ZN(
        n11972) );
  INV_X1 U14339 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12245) );
  INV_X1 U14340 ( .A(n11963), .ZN(n11964) );
  AOI21_X1 U14341 ( .B1(n11965), .B2(P1_REG2_REG_16__SCAN_IN), .A(n11964), 
        .ZN(n11967) );
  NOR2_X1 U14342 ( .A1(n12244), .A2(n12245), .ZN(n11966) );
  AOI211_X1 U14343 ( .C1(n12245), .C2(n12244), .A(n11967), .B(n11966), .ZN(
        n12242) );
  INV_X1 U14344 ( .A(n11967), .ZN(n11969) );
  NOR2_X1 U14345 ( .A1(n12244), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11968) );
  AOI211_X1 U14346 ( .C1(n12244), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11969), 
        .B(n11968), .ZN(n11970) );
  NOR3_X1 U14347 ( .A1(n14807), .A2(n12242), .A3(n11970), .ZN(n11971) );
  OR3_X1 U14348 ( .A1(n11973), .A2(n11972), .A3(n11971), .ZN(P1_U3260) );
  OR2_X1 U14349 ( .A1(n11974), .A2(n14556), .ZN(n11975) );
  NAND2_X1 U14350 ( .A1(n12037), .A2(n11975), .ZN(n14557) );
  XNOR2_X1 U14351 ( .A(n11976), .B(n11977), .ZN(n11983) );
  XNOR2_X1 U14352 ( .A(n11979), .B(n11978), .ZN(n11981) );
  OAI22_X1 U14353 ( .A1(n13794), .A2(n14351), .B1(n12395), .B2(n14353), .ZN(
        n11980) );
  AOI21_X1 U14354 ( .B1(n11981), .B2(n14384), .A(n11980), .ZN(n11982) );
  OAI21_X1 U14355 ( .B1(n14860), .B2(n11983), .A(n11982), .ZN(n14558) );
  NAND2_X1 U14356 ( .A1(n14558), .A2(n14393), .ZN(n11987) );
  OAI22_X1 U14357 ( .A1(n14393), .A2(n11133), .B1(n11984), .B2(n14386), .ZN(
        n11985) );
  AOI21_X1 U14358 ( .B1(n12387), .B2(n14322), .A(n11985), .ZN(n11986) );
  OAI211_X1 U14359 ( .C1(n14319), .C2(n14557), .A(n11987), .B(n11986), .ZN(
        P1_U3281) );
  XNOR2_X1 U14360 ( .A(n11988), .B(n6981), .ZN(n11989) );
  OAI222_X1 U14361 ( .A1(n15302), .A2(n12352), .B1(n15303), .B2(n12179), .C1(
        n11989), .C2(n15308), .ZN(n14618) );
  INV_X1 U14362 ( .A(n14618), .ZN(n11996) );
  OAI21_X1 U14363 ( .B1(n11992), .B2(n11991), .A(n11990), .ZN(n14620) );
  AOI22_X1 U14364 ( .A1(n13001), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15331), 
        .B2(n12354), .ZN(n11993) );
  OAI21_X1 U14365 ( .B1(n14617), .B2(n12997), .A(n11993), .ZN(n11994) );
  AOI21_X1 U14366 ( .B1(n14620), .B2(n12999), .A(n11994), .ZN(n11995) );
  OAI21_X1 U14367 ( .B1(n11996), .B2(n13001), .A(n11995), .ZN(P3_U3221) );
  INV_X1 U14368 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11997) );
  OR2_X1 U14369 ( .A1(n12263), .A2(n11997), .ZN(n11999) );
  NAND2_X1 U14370 ( .A1(n12263), .A2(n11997), .ZN(n11998) );
  AND2_X1 U14371 ( .A1(n11999), .A2(n11998), .ZN(n12004) );
  INV_X1 U14372 ( .A(n12256), .ZN(n12002) );
  AOI21_X1 U14373 ( .B1(n12004), .B2(n12003), .A(n12002), .ZN(n12026) );
  NOR2_X1 U14374 ( .A1(n12263), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12005) );
  AOI21_X1 U14375 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12263), .A(n12005), 
        .ZN(n12011) );
  NAND2_X1 U14376 ( .A1(n12007), .A2(n12006), .ZN(n12009) );
  NAND2_X1 U14377 ( .A1(n12009), .A2(n12008), .ZN(n12010) );
  NAND2_X1 U14378 ( .A1(n12010), .A2(n12011), .ZN(n12260) );
  OAI21_X1 U14379 ( .B1(n12011), .B2(n12010), .A(n12260), .ZN(n12024) );
  NOR2_X1 U14380 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12012), .ZN(n12349) );
  AOI21_X1 U14381 ( .B1(n15245), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12349), 
        .ZN(n12013) );
  OAI21_X1 U14382 ( .B1(n15285), .B2(n12263), .A(n12013), .ZN(n12023) );
  INV_X1 U14383 ( .A(n12014), .ZN(n12016) );
  NAND2_X1 U14384 ( .A1(n12016), .A2(n12015), .ZN(n12018) );
  MUX2_X1 U14385 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12823), .Z(n12264) );
  XOR2_X1 U14386 ( .A(n12263), .B(n12264), .Z(n12017) );
  NAND3_X1 U14387 ( .A1(n12019), .A2(n12018), .A3(n12017), .ZN(n12267) );
  INV_X1 U14388 ( .A(n12267), .ZN(n12021) );
  AOI21_X1 U14389 ( .B1(n12019), .B2(n12018), .A(n12017), .ZN(n12020) );
  NOR3_X1 U14390 ( .A1(n12021), .A2(n12020), .A3(n15241), .ZN(n12022) );
  AOI211_X1 U14391 ( .C1(n15287), .C2(n12024), .A(n12023), .B(n12022), .ZN(
        n12025) );
  OAI21_X1 U14392 ( .B1(n12026), .B2(n15291), .A(n12025), .ZN(P3_U3194) );
  INV_X1 U14393 ( .A(n12027), .ZN(n12029) );
  OAI222_X1 U14394 ( .A1(n13123), .A2(n12029), .B1(n13125), .B2(n7569), .C1(
        n12028), .C2(P3_U3151), .ZN(P3_U3271) );
  XNOR2_X1 U14395 ( .A(n12030), .B(n12036), .ZN(n12031) );
  NAND2_X1 U14396 ( .A1(n12031), .A2(n14384), .ZN(n12034) );
  NAND2_X1 U14397 ( .A1(n14074), .A2(n14362), .ZN(n12033) );
  NAND2_X1 U14398 ( .A1(n14076), .A2(n14364), .ZN(n12032) );
  AND2_X1 U14399 ( .A1(n12033), .A2(n12032), .ZN(n14019) );
  NAND2_X1 U14400 ( .A1(n12034), .A2(n14019), .ZN(n14714) );
  INV_X1 U14401 ( .A(n14714), .ZN(n12043) );
  XNOR2_X1 U14402 ( .A(n12035), .B(n12036), .ZN(n14709) );
  NAND2_X1 U14403 ( .A1(n12037), .A2(n14710), .ZN(n12038) );
  NAND2_X1 U14404 ( .A1(n12121), .A2(n12038), .ZN(n14711) );
  AOI22_X1 U14405 ( .A1(n14377), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n14021), 
        .B2(n14369), .ZN(n12040) );
  NAND2_X1 U14406 ( .A1(n14710), .A2(n14322), .ZN(n12039) );
  OAI211_X1 U14407 ( .C1(n14711), .C2(n14319), .A(n12040), .B(n12039), .ZN(
        n12041) );
  AOI21_X1 U14408 ( .B1(n14709), .B2(n14325), .A(n12041), .ZN(n12042) );
  OAI21_X1 U14409 ( .B1(n12043), .B2(n14377), .A(n12042), .ZN(P1_U3280) );
  AOI211_X1 U14410 ( .C1(n12046), .C2(n15137), .A(n12045), .B(n12044), .ZN(
        n12051) );
  AOI22_X1 U14411 ( .A1(n12115), .A2(n13688), .B1(n15154), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12047) );
  OAI21_X1 U14412 ( .B1(n12051), .B2(n15154), .A(n12047), .ZN(P2_U3512) );
  INV_X1 U14413 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12048) );
  NOR2_X1 U14414 ( .A1(n15147), .A2(n12048), .ZN(n12049) );
  AOI21_X1 U14415 ( .B1(n12115), .B2(n13749), .A(n12049), .ZN(n12050) );
  OAI21_X1 U14416 ( .B1(n12051), .B2(n15145), .A(n12050), .ZN(P2_U3469) );
  INV_X1 U14417 ( .A(n12052), .ZN(n12053) );
  NAND2_X1 U14418 ( .A1(n12089), .A2(n13935), .ZN(n12058) );
  NAND2_X1 U14419 ( .A1(n14081), .A2(n13933), .ZN(n12057) );
  NAND2_X1 U14420 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  XNOR2_X1 U14421 ( .A(n12059), .B(n12151), .ZN(n12062) );
  AOI22_X1 U14422 ( .A1(n12089), .A2(n13933), .B1(n13932), .B2(n14081), .ZN(
        n12060) );
  XNOR2_X1 U14423 ( .A(n12062), .B(n12060), .ZN(n12084) );
  INV_X1 U14424 ( .A(n12060), .ZN(n12061) );
  NAND2_X1 U14425 ( .A1(n14881), .A2(n13935), .ZN(n12064) );
  NAND2_X1 U14426 ( .A1(n14080), .A2(n13933), .ZN(n12063) );
  NAND2_X1 U14427 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  XNOR2_X1 U14428 ( .A(n12065), .B(n12151), .ZN(n12069) );
  NAND2_X1 U14429 ( .A1(n14881), .A2(n13933), .ZN(n12067) );
  NAND2_X1 U14430 ( .A1(n13932), .A2(n14080), .ZN(n12066) );
  NAND2_X1 U14431 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  NOR2_X1 U14432 ( .A1(n12069), .A2(n12068), .ZN(n12154) );
  AOI21_X1 U14433 ( .B1(n12069), .B2(n12068), .A(n12154), .ZN(n12070) );
  NAND2_X1 U14434 ( .A1(n12071), .A2(n12070), .ZN(n12156) );
  OAI21_X1 U14435 ( .B1(n12071), .B2(n12070), .A(n12156), .ZN(n12072) );
  NAND2_X1 U14436 ( .A1(n12072), .A2(n14689), .ZN(n12078) );
  OAI21_X1 U14437 ( .B1(n12074), .B2(n14049), .A(n12073), .ZN(n12075) );
  AOI21_X1 U14438 ( .B1(n12076), .B2(n14063), .A(n12075), .ZN(n12077) );
  OAI211_X1 U14439 ( .C1(n12079), .C2(n14059), .A(n12078), .B(n12077), .ZN(
        P1_U3221) );
  OR2_X1 U14440 ( .A1(n14696), .A2(n12080), .ZN(n12082) );
  OAI211_X1 U14441 ( .C1(n12083), .C2(n14049), .A(n12082), .B(n12081), .ZN(
        n12088) );
  XNOR2_X1 U14442 ( .A(n12085), .B(n12084), .ZN(n12086) );
  NOR2_X1 U14443 ( .A1(n12086), .A2(n14065), .ZN(n12087) );
  AOI211_X1 U14444 ( .C1(n14687), .C2(n12089), .A(n12088), .B(n12087), .ZN(
        n12090) );
  INV_X1 U14445 ( .A(n12090), .ZN(P1_U3213) );
  XOR2_X1 U14446 ( .A(n12093), .B(n12091), .Z(n12092) );
  AOI22_X1 U14447 ( .A1(n12963), .A2(n12712), .B1(n12710), .B2(n12962), .ZN(
        n12181) );
  OAI21_X1 U14448 ( .B1(n12092), .B2(n15308), .A(n12181), .ZN(n12215) );
  INV_X1 U14449 ( .A(n12215), .ZN(n12098) );
  XNOR2_X1 U14450 ( .A(n12094), .B(n12093), .ZN(n12216) );
  AOI22_X1 U14451 ( .A1(n13001), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15331), 
        .B2(n12184), .ZN(n12095) );
  OAI21_X1 U14452 ( .B1(n12222), .B2(n12997), .A(n12095), .ZN(n12096) );
  AOI21_X1 U14453 ( .B1(n12216), .B2(n12999), .A(n12096), .ZN(n12097) );
  OAI21_X1 U14454 ( .B1(n12098), .B2(n13001), .A(n12097), .ZN(P3_U3220) );
  NAND2_X1 U14455 ( .A1(n12099), .A2(n13249), .ZN(n12100) );
  NAND2_X1 U14456 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n13321)
         );
  OAI211_X1 U14457 ( .C1(n14934), .C2(n12101), .A(n12100), .B(n13321), .ZN(
        n12114) );
  XNOR2_X1 U14458 ( .A(n12115), .B(n12518), .ZN(n12103) );
  AND2_X1 U14459 ( .A1(n13258), .A2(n12562), .ZN(n12102) );
  NAND2_X1 U14460 ( .A1(n12103), .A2(n12102), .ZN(n12128) );
  OAI21_X1 U14461 ( .B1(n12103), .B2(n12102), .A(n12128), .ZN(n12112) );
  INV_X1 U14462 ( .A(n12104), .ZN(n12105) );
  NAND2_X1 U14463 ( .A1(n13259), .A2(n12562), .ZN(n12107) );
  XNOR2_X1 U14464 ( .A(n14931), .B(n12518), .ZN(n12109) );
  XOR2_X1 U14465 ( .A(n12107), .B(n12109), .Z(n14924) );
  INV_X1 U14466 ( .A(n12107), .ZN(n12108) );
  NAND2_X1 U14467 ( .A1(n14923), .A2(n12110), .ZN(n12111) );
  AOI211_X1 U14468 ( .C1(n12112), .C2(n12111), .A(n14926), .B(n12130), .ZN(
        n12113) );
  AOI211_X1 U14469 ( .C1(n12115), .C2(n14930), .A(n12114), .B(n12113), .ZN(
        n12116) );
  INV_X1 U14470 ( .A(n12116), .ZN(P2_U3206) );
  XNOR2_X1 U14471 ( .A(n12117), .B(n12120), .ZN(n12118) );
  OAI22_X1 U14472 ( .A1(n13794), .A2(n14353), .B1(n13977), .B2(n14351), .ZN(
        n14692) );
  AOI21_X1 U14473 ( .B1(n12118), .B2(n14384), .A(n14692), .ZN(n14705) );
  XNOR2_X1 U14474 ( .A(n12119), .B(n12120), .ZN(n14708) );
  INV_X1 U14475 ( .A(n12121), .ZN(n12122) );
  OAI21_X1 U14476 ( .B1(n14703), .B2(n12122), .A(n12232), .ZN(n14704) );
  AOI22_X1 U14477 ( .A1(n14377), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n12123), 
        .B2(n14369), .ZN(n12125) );
  NAND2_X1 U14478 ( .A1(n14688), .A2(n14322), .ZN(n12124) );
  OAI211_X1 U14479 ( .C1(n14704), .C2(n14319), .A(n12125), .B(n12124), .ZN(
        n12126) );
  AOI21_X1 U14480 ( .B1(n14708), .B2(n14325), .A(n12126), .ZN(n12127) );
  OAI21_X1 U14481 ( .B1(n14705), .B2(n14377), .A(n12127), .ZN(P1_U3279) );
  INV_X1 U14482 ( .A(n12128), .ZN(n12129) );
  NAND2_X1 U14483 ( .A1(n13257), .A2(n12562), .ZN(n12501) );
  XNOR2_X1 U14484 ( .A(n12500), .B(n12501), .ZN(n12131) );
  OAI21_X1 U14485 ( .B1(n6627), .B2(n12131), .A(n12504), .ZN(n12132) );
  NAND2_X1 U14486 ( .A1(n12132), .A2(n13243), .ZN(n12135) );
  OAI22_X1 U14487 ( .A1(n14637), .A2(n13537), .B1(n14919), .B2(n13539), .ZN(
        n14650) );
  NAND2_X1 U14488 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n15004)
         );
  OAI21_X1 U14489 ( .B1(n14934), .B2(n14652), .A(n15004), .ZN(n12133) );
  AOI21_X1 U14490 ( .B1(n14650), .B2(n13249), .A(n12133), .ZN(n12134) );
  OAI211_X1 U14491 ( .C1(n6678), .C2(n13252), .A(n12135), .B(n12134), .ZN(
        P2_U3187) );
  OAI222_X1 U14492 ( .A1(n13783), .A2(n12138), .B1(P2_U3088), .B2(n12137), 
        .C1(n13781), .C2(n12136), .ZN(P2_U3305) );
  OAI211_X1 U14493 ( .C1(n6628), .C2(n12143), .A(n12139), .B(n15317), .ZN(
        n12142) );
  OR2_X1 U14494 ( .A1(n12408), .A2(n15303), .ZN(n12141) );
  NAND2_X1 U14495 ( .A1(n12711), .A2(n12963), .ZN(n12140) );
  AND2_X1 U14496 ( .A1(n12141), .A2(n12140), .ZN(n12285) );
  XNOR2_X1 U14497 ( .A(n12144), .B(n12143), .ZN(n12322) );
  AOI22_X1 U14498 ( .A1(n13001), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15331), 
        .B2(n12284), .ZN(n12145) );
  OAI21_X1 U14499 ( .B1(n12330), .B2(n12997), .A(n12145), .ZN(n12146) );
  AOI21_X1 U14500 ( .B1(n12322), .B2(n12999), .A(n12146), .ZN(n12147) );
  OAI21_X1 U14501 ( .B1(n12324), .B2(n13001), .A(n12147), .ZN(P3_U3219) );
  INV_X1 U14502 ( .A(n12148), .ZN(n12214) );
  NAND2_X1 U14503 ( .A1(n12153), .A2(n14882), .ZN(n14892) );
  NAND2_X1 U14504 ( .A1(n12153), .A2(n13935), .ZN(n12150) );
  NAND2_X1 U14505 ( .A1(n14079), .A2(n13933), .ZN(n12149) );
  NAND2_X1 U14506 ( .A1(n12150), .A2(n12149), .ZN(n12152) );
  XNOR2_X1 U14507 ( .A(n12152), .B(n12151), .ZN(n12196) );
  AOI22_X1 U14508 ( .A1(n12153), .A2(n13933), .B1(n13932), .B2(n14079), .ZN(
        n12197) );
  XNOR2_X1 U14509 ( .A(n12196), .B(n12197), .ZN(n12158) );
  INV_X1 U14510 ( .A(n12154), .ZN(n12155) );
  NAND2_X1 U14511 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  NAND2_X1 U14512 ( .A1(n12157), .A2(n12158), .ZN(n12204) );
  OAI21_X1 U14513 ( .B1(n12158), .B2(n12157), .A(n12204), .ZN(n12159) );
  NAND2_X1 U14514 ( .A1(n12159), .A2(n14689), .ZN(n12165) );
  AND2_X1 U14515 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14131) );
  AOI21_X1 U14516 ( .B1(n14055), .B2(n14078), .A(n14131), .ZN(n12160) );
  OAI21_X1 U14517 ( .B1(n12161), .B2(n14057), .A(n12160), .ZN(n12162) );
  AOI21_X1 U14518 ( .B1(n12163), .B2(n14063), .A(n12162), .ZN(n12164) );
  OAI211_X1 U14519 ( .C1(n12214), .C2(n14892), .A(n12165), .B(n12164), .ZN(
        P1_U3231) );
  INV_X1 U14520 ( .A(n12166), .ZN(n12168) );
  OAI222_X1 U14521 ( .A1(n13125), .A2(n12169), .B1(n13123), .B2(n12168), .C1(
        P3_U3151), .C2(n12167), .ZN(P3_U3270) );
  OR2_X1 U14522 ( .A1(n12170), .A2(n12334), .ZN(n12171) );
  XNOR2_X1 U14523 ( .A(n14617), .B(n11800), .ZN(n12176) );
  NAND2_X1 U14524 ( .A1(n12176), .A2(n12175), .ZN(n12343) );
  XNOR2_X1 U14525 ( .A(n12331), .B(n11800), .ZN(n12341) );
  NOR2_X1 U14526 ( .A1(n12173), .A2(n12352), .ZN(n12177) );
  NOR2_X1 U14527 ( .A1(n12176), .A2(n12175), .ZN(n12344) );
  AOI21_X1 U14528 ( .B1(n12177), .B2(n12343), .A(n12344), .ZN(n12178) );
  XNOR2_X1 U14529 ( .A(n12222), .B(n12485), .ZN(n12280) );
  XNOR2_X1 U14530 ( .A(n12280), .B(n12179), .ZN(n12180) );
  XNOR2_X1 U14531 ( .A(n12279), .B(n12180), .ZN(n12186) );
  OAI22_X1 U14532 ( .A1(n12181), .A2(n15189), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12270), .ZN(n12183) );
  NOR2_X1 U14533 ( .A1(n12222), .A2(n15170), .ZN(n12182) );
  AOI211_X1 U14534 ( .C1(n12184), .C2(n12696), .A(n12183), .B(n12182), .ZN(
        n12185) );
  OAI21_X1 U14535 ( .B1(n12186), .B2(n15172), .A(n12185), .ZN(P3_U3174) );
  NAND2_X1 U14536 ( .A1(n12192), .A2(n12187), .ZN(n12189) );
  OAI211_X1 U14537 ( .C1(n12190), .C2(n13783), .A(n12189), .B(n12188), .ZN(
        P2_U3304) );
  NAND2_X1 U14538 ( .A1(n12192), .A2(n12191), .ZN(n12194) );
  OAI211_X1 U14539 ( .C1(n12195), .C2(n14527), .A(n12194), .B(n12193), .ZN(
        P1_U3332) );
  NAND2_X1 U14540 ( .A1(n12200), .A2(n14882), .ZN(n14899) );
  INV_X1 U14541 ( .A(n12196), .ZN(n12198) );
  NAND2_X1 U14542 ( .A1(n12198), .A2(n12197), .ZN(n12202) );
  AND2_X1 U14543 ( .A1(n12204), .A2(n12202), .ZN(n12206) );
  NOR2_X1 U14544 ( .A1(n13854), .A2(n12317), .ZN(n12199) );
  AOI21_X1 U14545 ( .B1(n12200), .B2(n13933), .A(n12199), .ZN(n12304) );
  AOI22_X1 U14546 ( .A1(n12200), .A2(n13935), .B1(n13933), .B2(n14078), .ZN(
        n12201) );
  XNOR2_X1 U14547 ( .A(n12201), .B(n12151), .ZN(n12303) );
  XOR2_X1 U14548 ( .A(n12304), .B(n12303), .Z(n12205) );
  OAI211_X1 U14549 ( .C1(n12206), .C2(n12205), .A(n14689), .B(n12308), .ZN(
        n12213) );
  AOI21_X1 U14550 ( .B1(n14055), .B2(n14077), .A(n12207), .ZN(n12208) );
  OAI21_X1 U14551 ( .B1(n12209), .B2(n14057), .A(n12208), .ZN(n12210) );
  AOI21_X1 U14552 ( .B1(n12211), .B2(n14063), .A(n12210), .ZN(n12212) );
  OAI211_X1 U14553 ( .C1(n12214), .C2(n14899), .A(n12213), .B(n12212), .ZN(
        P1_U3217) );
  INV_X1 U14554 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12217) );
  AOI21_X1 U14555 ( .B1(n12216), .B2(n15339), .A(n12215), .ZN(n12219) );
  MUX2_X1 U14556 ( .A(n12217), .B(n12219), .S(n15374), .Z(n12218) );
  OAI21_X1 U14557 ( .B1(n13062), .B2(n12222), .A(n12218), .ZN(P3_U3472) );
  INV_X1 U14558 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12220) );
  MUX2_X1 U14559 ( .A(n12220), .B(n12219), .S(n15365), .Z(n12221) );
  OAI21_X1 U14560 ( .B1(n13110), .B2(n12222), .A(n12221), .ZN(P3_U3429) );
  XNOR2_X1 U14561 ( .A(n12224), .B(n12223), .ZN(n12225) );
  NAND2_X1 U14562 ( .A1(n12225), .A2(n14384), .ZN(n12227) );
  AOI22_X1 U14563 ( .A1(n14362), .A2(n14365), .B1(n14074), .B2(n14364), .ZN(
        n12226) );
  NAND2_X1 U14564 ( .A1(n12229), .A2(n12228), .ZN(n12230) );
  NAND2_X1 U14565 ( .A1(n12231), .A2(n12230), .ZN(n14700) );
  AND2_X1 U14566 ( .A1(n13812), .A2(n12232), .ZN(n12233) );
  OR2_X1 U14567 ( .A1(n12233), .A2(n14389), .ZN(n14698) );
  AOI22_X1 U14568 ( .A1(n14377), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14062), 
        .B2(n14369), .ZN(n12235) );
  NAND2_X1 U14569 ( .A1(n13812), .A2(n14322), .ZN(n12234) );
  OAI211_X1 U14570 ( .C1(n14698), .C2(n14319), .A(n12235), .B(n12234), .ZN(
        n12236) );
  AOI21_X1 U14571 ( .B1(n14700), .B2(n14325), .A(n12236), .ZN(n12237) );
  OAI21_X1 U14572 ( .B1(n14702), .B2(n14377), .A(n12237), .ZN(P1_U3278) );
  XNOR2_X1 U14573 ( .A(n14157), .B(n14156), .ZN(n12241) );
  INV_X1 U14574 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n12240) );
  NOR2_X1 U14575 ( .A1(n12240), .A2(n12241), .ZN(n14159) );
  AOI211_X1 U14576 ( .C1(n12241), .C2(n12240), .A(n14159), .B(n14168), .ZN(
        n12251) );
  INV_X1 U14577 ( .A(n12242), .ZN(n12243) );
  OAI21_X1 U14578 ( .B1(n12245), .B2(n12244), .A(n12243), .ZN(n14161) );
  XNOR2_X1 U14579 ( .A(n14161), .B(n14156), .ZN(n12246) );
  NAND2_X1 U14580 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n12246), .ZN(n14164) );
  OAI211_X1 U14581 ( .C1(n12246), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14771), 
        .B(n14164), .ZN(n12249) );
  NAND2_X1 U14582 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14040)
         );
  INV_X1 U14583 ( .A(n14040), .ZN(n12247) );
  AOI21_X1 U14584 ( .B1(n14757), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n12247), 
        .ZN(n12248) );
  OAI211_X1 U14585 ( .C1(n14775), .C2(n14156), .A(n12249), .B(n12248), .ZN(
        n12250) );
  OR2_X1 U14586 ( .A1(n12251), .A2(n12250), .ZN(P1_U3261) );
  INV_X1 U14587 ( .A(n12252), .ZN(n12253) );
  OAI222_X1 U14588 ( .A1(n12254), .A2(P3_U3151), .B1(n13123), .B2(n12253), 
        .C1(n8689), .C2(n13125), .ZN(P3_U3269) );
  INV_X1 U14589 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U14590 ( .A1(n12263), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12255) );
  AOI21_X1 U14591 ( .B1(n12259), .B2(n12258), .A(n12725), .ZN(n12277) );
  INV_X1 U14592 ( .A(n12263), .ZN(n12261) );
  INV_X1 U14593 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14621) );
  XNOR2_X1 U14594 ( .A(n12731), .B(n12257), .ZN(n12262) );
  NAND2_X1 U14595 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12262), .ZN(n12733) );
  OAI21_X1 U14596 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12262), .A(n12733), 
        .ZN(n12275) );
  NAND2_X1 U14597 ( .A1(n12264), .A2(n12263), .ZN(n12266) );
  MUX2_X1 U14598 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12823), .Z(n12739) );
  XNOR2_X1 U14599 ( .A(n12739), .B(n12257), .ZN(n12265) );
  NAND3_X1 U14600 ( .A1(n12267), .A2(n12266), .A3(n12265), .ZN(n12745) );
  INV_X1 U14601 ( .A(n12745), .ZN(n12269) );
  AOI21_X1 U14602 ( .B1(n12267), .B2(n12266), .A(n12265), .ZN(n12268) );
  OAI21_X1 U14603 ( .B1(n12269), .B2(n12268), .A(n15280), .ZN(n12273) );
  NOR2_X1 U14604 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12270), .ZN(n12271) );
  AOI21_X1 U14605 ( .B1(n15245), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12271), 
        .ZN(n12272) );
  OAI211_X1 U14606 ( .C1(n15285), .C2(n12732), .A(n12273), .B(n12272), .ZN(
        n12274) );
  AOI21_X1 U14607 ( .B1(n15287), .B2(n12275), .A(n12274), .ZN(n12276) );
  OAI21_X1 U14608 ( .B1(n12277), .B2(n15291), .A(n12276), .ZN(P3_U3195) );
  NAND2_X1 U14609 ( .A1(n12280), .A2(n12711), .ZN(n12281) );
  XNOR2_X1 U14610 ( .A(n12330), .B(n12485), .ZN(n12368) );
  XNOR2_X1 U14611 ( .A(n12368), .B(n12283), .ZN(n12366) );
  XNOR2_X1 U14612 ( .A(n12367), .B(n12366), .ZN(n12292) );
  INV_X1 U14613 ( .A(n12330), .ZN(n12290) );
  INV_X1 U14614 ( .A(n12284), .ZN(n12288) );
  INV_X1 U14615 ( .A(n12285), .ZN(n12286) );
  NAND2_X1 U14616 ( .A1(n12286), .A2(n15178), .ZN(n12287) );
  NAND2_X1 U14617 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12738)
         );
  OAI211_X1 U14618 ( .C1(n15193), .C2(n12288), .A(n12287), .B(n12738), .ZN(
        n12289) );
  AOI21_X1 U14619 ( .B1(n12290), .B2(n15186), .A(n12289), .ZN(n12291) );
  OAI21_X1 U14620 ( .B1(n12292), .B2(n15172), .A(n12291), .ZN(P3_U3155) );
  XOR2_X1 U14621 ( .A(n12293), .B(n12296), .Z(n12294) );
  AOI22_X1 U14622 ( .A1(n12963), .A2(n12710), .B1(n12708), .B2(n12962), .ZN(
        n12371) );
  OAI21_X1 U14623 ( .B1(n12294), .B2(n15308), .A(n12371), .ZN(n13058) );
  INV_X1 U14624 ( .A(n13058), .ZN(n12301) );
  OAI21_X1 U14625 ( .B1(n12297), .B2(n12296), .A(n12295), .ZN(n13059) );
  INV_X1 U14626 ( .A(n12370), .ZN(n13111) );
  AOI22_X1 U14627 ( .A1(n13001), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15331), 
        .B2(n12374), .ZN(n12298) );
  OAI21_X1 U14628 ( .B1(n13111), .B2(n12997), .A(n12298), .ZN(n12299) );
  AOI21_X1 U14629 ( .B1(n13059), .B2(n12999), .A(n12299), .ZN(n12300) );
  OAI21_X1 U14630 ( .B1(n12301), .B2(n13001), .A(n12300), .ZN(P3_U3218) );
  AOI22_X1 U14631 ( .A1(n12319), .A2(n13935), .B1(n13933), .B2(n14077), .ZN(
        n12302) );
  XNOR2_X1 U14632 ( .A(n12302), .B(n12151), .ZN(n12384) );
  AOI22_X1 U14633 ( .A1(n12319), .A2(n13933), .B1(n13932), .B2(n14077), .ZN(
        n12383) );
  XNOR2_X1 U14634 ( .A(n12384), .B(n12383), .ZN(n12312) );
  INV_X1 U14635 ( .A(n12303), .ZN(n12306) );
  INV_X1 U14636 ( .A(n12304), .ZN(n12305) );
  INV_X1 U14637 ( .A(n12391), .ZN(n12310) );
  AOI21_X1 U14638 ( .B1(n12312), .B2(n12311), .A(n12310), .ZN(n12321) );
  AOI21_X1 U14639 ( .B1(n14055), .B2(n14076), .A(n12313), .ZN(n12316) );
  NAND2_X1 U14640 ( .A1(n14063), .A2(n12314), .ZN(n12315) );
  OAI211_X1 U14641 ( .C1(n12317), .C2(n14057), .A(n12316), .B(n12315), .ZN(
        n12318) );
  AOI21_X1 U14642 ( .B1(n12319), .B2(n14687), .A(n12318), .ZN(n12320) );
  OAI21_X1 U14643 ( .B1(n12321), .B2(n14065), .A(n12320), .ZN(P1_U3236) );
  INV_X1 U14644 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14645 ( .A1(n12322), .A2(n15339), .ZN(n12323) );
  AND2_X1 U14646 ( .A1(n12324), .A2(n12323), .ZN(n12327) );
  MUX2_X1 U14647 ( .A(n12325), .B(n12327), .S(n15374), .Z(n12326) );
  OAI21_X1 U14648 ( .B1(n13062), .B2(n12330), .A(n12326), .ZN(P3_U3473) );
  INV_X1 U14649 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12328) );
  MUX2_X1 U14650 ( .A(n12328), .B(n12327), .S(n15365), .Z(n12329) );
  OAI21_X1 U14651 ( .B1(n13110), .B2(n12330), .A(n12329), .ZN(P3_U3432) );
  AOI22_X1 U14652 ( .A1(n12692), .A2(n12712), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12333) );
  NAND2_X1 U14653 ( .A1(n15186), .A2(n12331), .ZN(n12332) );
  OAI211_X1 U14654 ( .C1(n12334), .C2(n12694), .A(n12333), .B(n12332), .ZN(
        n12337) );
  XNOR2_X1 U14655 ( .A(n12342), .B(n12341), .ZN(n12335) );
  NOR2_X1 U14656 ( .A1(n12335), .A2(n12352), .ZN(n12340) );
  AOI211_X1 U14657 ( .C1(n12352), .C2(n12335), .A(n15172), .B(n12340), .ZN(
        n12336) );
  AOI211_X1 U14658 ( .C1(n12338), .C2(n12696), .A(n12337), .B(n12336), .ZN(
        n12339) );
  INV_X1 U14659 ( .A(n12339), .ZN(P3_U3176) );
  AOI21_X1 U14660 ( .B1(n12342), .B2(n12341), .A(n12340), .ZN(n12347) );
  INV_X1 U14661 ( .A(n12343), .ZN(n12345) );
  NOR2_X1 U14662 ( .A1(n12344), .A2(n12345), .ZN(n12346) );
  OAI22_X1 U14663 ( .A1(n12347), .A2(n12346), .B1(n12345), .B2(n12279), .ZN(
        n12348) );
  NAND2_X1 U14664 ( .A1(n12348), .A2(n15180), .ZN(n12356) );
  NAND2_X1 U14665 ( .A1(n12692), .A2(n12711), .ZN(n12351) );
  INV_X1 U14666 ( .A(n12349), .ZN(n12350) );
  OAI211_X1 U14667 ( .C1(n12352), .C2(n12694), .A(n12351), .B(n12350), .ZN(
        n12353) );
  AOI21_X1 U14668 ( .B1(n12696), .B2(n12354), .A(n12353), .ZN(n12355) );
  OAI211_X1 U14669 ( .C1(n14617), .C2(n15170), .A(n12356), .B(n12355), .ZN(
        P3_U3164) );
  XNOR2_X1 U14670 ( .A(n12358), .B(n12361), .ZN(n12359) );
  AOI222_X1 U14671 ( .A1(n15317), .A2(n12359), .B1(n12707), .B2(n12962), .C1(
        n12709), .C2(n12963), .ZN(n13057) );
  OAI21_X1 U14672 ( .B1(n12362), .B2(n12361), .A(n12360), .ZN(n13055) );
  AOI22_X1 U14673 ( .A1(n13001), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15331), 
        .B2(n12405), .ZN(n12363) );
  OAI21_X1 U14674 ( .B1(n12404), .B2(n12997), .A(n12363), .ZN(n12364) );
  AOI21_X1 U14675 ( .B1(n13055), .B2(n12999), .A(n12364), .ZN(n12365) );
  OAI21_X1 U14676 ( .B1(n13057), .B2(n13001), .A(n12365), .ZN(P3_U3217) );
  NAND2_X1 U14677 ( .A1(n12368), .A2(n12710), .ZN(n12369) );
  XNOR2_X1 U14678 ( .A(n12370), .B(n12485), .ZN(n12402) );
  XNOR2_X1 U14679 ( .A(n12402), .B(n12709), .ZN(n12400) );
  XNOR2_X1 U14680 ( .A(n12401), .B(n12400), .ZN(n12376) );
  OAI22_X1 U14681 ( .A1(n12371), .A2(n15189), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12765), .ZN(n12373) );
  NOR2_X1 U14682 ( .A1(n13111), .A2(n15170), .ZN(n12372) );
  AOI211_X1 U14683 ( .C1(n12374), .C2(n12696), .A(n12373), .B(n12372), .ZN(
        n12375) );
  OAI21_X1 U14684 ( .B1(n12376), .B2(n15172), .A(n12375), .ZN(P3_U3181) );
  OAI222_X1 U14685 ( .A1(P2_U3088), .A2(n12378), .B1(n13781), .B2(n12381), 
        .C1(n12377), .C2(n13783), .ZN(P2_U3303) );
  INV_X1 U14686 ( .A(n12379), .ZN(n12382) );
  OAI222_X1 U14687 ( .A1(n12382), .A2(P1_U3086), .B1(n14525), .B2(n12381), 
        .C1(n12380), .C2(n14527), .ZN(P1_U3331) );
  NAND2_X1 U14688 ( .A1(n12384), .A2(n12383), .ZN(n12389) );
  AND2_X1 U14689 ( .A1(n12391), .A2(n12389), .ZN(n12393) );
  NOR2_X1 U14690 ( .A1(n13854), .A2(n12385), .ZN(n12386) );
  AOI21_X1 U14691 ( .B1(n12387), .B2(n13933), .A(n12386), .ZN(n13789) );
  AOI22_X1 U14692 ( .A1(n12387), .A2(n13935), .B1(n13933), .B2(n14076), .ZN(
        n12388) );
  XNOR2_X1 U14693 ( .A(n12388), .B(n12151), .ZN(n13788) );
  XOR2_X1 U14694 ( .A(n13789), .B(n13788), .Z(n12392) );
  NAND2_X1 U14695 ( .A1(n12391), .A2(n12390), .ZN(n13793) );
  OAI211_X1 U14696 ( .C1(n12393), .C2(n12392), .A(n14689), .B(n13793), .ZN(
        n12399) );
  NAND2_X1 U14697 ( .A1(n14055), .A2(n14075), .ZN(n12394) );
  NAND2_X1 U14698 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14793)
         );
  OAI211_X1 U14699 ( .C1(n12395), .C2(n14057), .A(n12394), .B(n14793), .ZN(
        n12396) );
  AOI21_X1 U14700 ( .B1(n12397), .B2(n14063), .A(n12396), .ZN(n12398) );
  OAI211_X1 U14701 ( .C1(n14556), .C2(n14059), .A(n12399), .B(n12398), .ZN(
        P1_U3224) );
  INV_X1 U14702 ( .A(n12402), .ZN(n12403) );
  XNOR2_X1 U14703 ( .A(n12404), .B(n12485), .ZN(n12453) );
  XNOR2_X1 U14704 ( .A(n12453), .B(n12990), .ZN(n12451) );
  XNOR2_X1 U14705 ( .A(n12452), .B(n12451), .ZN(n12411) );
  NAND2_X1 U14706 ( .A1(n12696), .A2(n12405), .ZN(n12407) );
  AOI22_X1 U14707 ( .A1(n12692), .A2(n12707), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12406) );
  OAI211_X1 U14708 ( .C1(n12408), .C2(n12694), .A(n12407), .B(n12406), .ZN(
        n12409) );
  AOI21_X1 U14709 ( .B1(n13054), .B2(n15186), .A(n12409), .ZN(n12410) );
  OAI21_X1 U14710 ( .B1(n12411), .B2(n15172), .A(n12410), .ZN(P3_U3166) );
  MUX2_X1 U14711 ( .A(n12412), .B(P1_REG2_REG_3__SCAN_IN), .S(n14377), .Z(
        n12418) );
  NAND2_X1 U14712 ( .A1(n12413), .A2(n14397), .ZN(n12416) );
  OR2_X1 U14713 ( .A1(n14394), .A2(n12414), .ZN(n12415) );
  OAI211_X1 U14714 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14386), .A(n12416), .B(
        n12415), .ZN(n12417) );
  OR2_X1 U14715 ( .A1(n12418), .A2(n12417), .ZN(P1_U3290) );
  AND2_X1 U14716 ( .A1(n15039), .A2(n12419), .ZN(P2_U3087) );
  OAI222_X1 U14717 ( .A1(n13783), .A2(n12421), .B1(n13781), .B2(n12420), .C1(
        n13379), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U14718 ( .A1(n12720), .A2(P3_DATAO_REG_0__SCAN_IN), .ZN(n12422) );
  OAI21_X1 U14719 ( .B1(n10209), .B2(n12720), .A(n12422), .ZN(P3_U3491) );
  AOI22_X1 U14720 ( .A1(n13770), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n14944), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n12423) );
  OAI21_X1 U14721 ( .B1(n12424), .B2(n13781), .A(n12423), .ZN(P2_U3326) );
  INV_X1 U14722 ( .A(n12425), .ZN(n13772) );
  OAI222_X1 U14723 ( .A1(n14527), .A2(n12426), .B1(n14525), .B2(n13772), .C1(
        P1_U3086), .C2(n7828), .ZN(P1_U3327) );
  XNOR2_X1 U14724 ( .A(n12427), .B(n12439), .ZN(n12431) );
  NAND2_X1 U14725 ( .A1(n14068), .A2(n14362), .ZN(n12429) );
  NAND2_X1 U14726 ( .A1(n12429), .A2(n12428), .ZN(n12430) );
  INV_X1 U14727 ( .A(n14188), .ZN(n12434) );
  INV_X1 U14728 ( .A(n12432), .ZN(n12433) );
  AOI21_X1 U14729 ( .B1(n14409), .B2(n12434), .A(n12433), .ZN(n14410) );
  AOI22_X1 U14730 ( .A1(n13942), .A2(n14369), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n14377), .ZN(n12435) );
  OAI21_X1 U14731 ( .B1(n12436), .B2(n14394), .A(n12435), .ZN(n12437) );
  AOI21_X1 U14732 ( .B1(n14410), .B2(n14397), .A(n12437), .ZN(n12442) );
  NAND2_X1 U14733 ( .A1(n12440), .A2(n12439), .ZN(n14408) );
  NAND3_X1 U14734 ( .A1(n6495), .A2(n14325), .A3(n14408), .ZN(n12441) );
  OAI211_X1 U14735 ( .C1(n14412), .C2(n14377), .A(n12442), .B(n12441), .ZN(
        P1_U3265) );
  INV_X1 U14736 ( .A(n12444), .ZN(n12580) );
  INV_X1 U14737 ( .A(n12446), .ZN(n12448) );
  OAI222_X1 U14738 ( .A1(n12823), .A2(P3_U3151), .B1(n13123), .B2(n12448), 
        .C1(n12447), .C2(n13125), .ZN(P3_U3268) );
  XNOR2_X1 U14739 ( .A(n12700), .B(n11800), .ZN(n12449) );
  XNOR2_X1 U14740 ( .A(n13003), .B(n12449), .ZN(n12494) );
  INV_X1 U14741 ( .A(n12494), .ZN(n12450) );
  NAND2_X1 U14742 ( .A1(n12450), .A2(n15180), .ZN(n12499) );
  NAND2_X1 U14743 ( .A1(n12452), .A2(n12451), .ZN(n12455) );
  NAND2_X1 U14744 ( .A1(n12453), .A2(n12708), .ZN(n12454) );
  NAND2_X1 U14745 ( .A1(n12455), .A2(n12454), .ZN(n12645) );
  XNOR2_X1 U14746 ( .A(n13105), .B(n12485), .ZN(n12456) );
  XNOR2_X1 U14747 ( .A(n12456), .B(n12978), .ZN(n12646) );
  NAND2_X1 U14748 ( .A1(n12645), .A2(n12646), .ZN(n12458) );
  NAND2_X1 U14749 ( .A1(n12456), .A2(n12707), .ZN(n12457) );
  XNOR2_X1 U14750 ( .A(n12683), .B(n12485), .ZN(n12459) );
  XNOR2_X1 U14751 ( .A(n12459), .B(n12964), .ZN(n12680) );
  INV_X1 U14752 ( .A(n12459), .ZN(n12460) );
  NAND2_X1 U14753 ( .A1(n12460), .A2(n12964), .ZN(n12461) );
  XNOR2_X1 U14754 ( .A(n13095), .B(n12485), .ZN(n12462) );
  XNOR2_X1 U14755 ( .A(n12462), .B(n12706), .ZN(n12606) );
  INV_X1 U14756 ( .A(n12462), .ZN(n12463) );
  XNOR2_X1 U14757 ( .A(n13092), .B(n12485), .ZN(n12464) );
  XNOR2_X1 U14758 ( .A(n12464), .B(n12934), .ZN(n12666) );
  INV_X1 U14759 ( .A(n12464), .ZN(n12465) );
  NOR2_X1 U14760 ( .A1(n12465), .A2(n12934), .ZN(n12466) );
  XNOR2_X1 U14761 ( .A(n12625), .B(n11800), .ZN(n12467) );
  NOR2_X1 U14762 ( .A1(n12467), .A2(n12705), .ZN(n12468) );
  AOI21_X1 U14763 ( .B1(n12467), .B2(n12705), .A(n12468), .ZN(n12628) );
  INV_X1 U14764 ( .A(n12468), .ZN(n12469) );
  NAND2_X1 U14765 ( .A1(n12626), .A2(n12469), .ZN(n12471) );
  XNOR2_X1 U14766 ( .A(n12675), .B(n12485), .ZN(n12470) );
  XNOR2_X1 U14767 ( .A(n12603), .B(n12485), .ZN(n12472) );
  XNOR2_X1 U14768 ( .A(n13019), .B(n12485), .ZN(n12474) );
  NAND2_X1 U14769 ( .A1(n12474), .A2(n12475), .ZN(n12635) );
  INV_X1 U14770 ( .A(n12474), .ZN(n12476) );
  INV_X1 U14771 ( .A(n12475), .ZN(n12908) );
  NAND2_X1 U14772 ( .A1(n12476), .A2(n12908), .ZN(n12477) );
  NAND2_X1 U14773 ( .A1(n12634), .A2(n12635), .ZN(n12483) );
  XNOR2_X1 U14774 ( .A(n12479), .B(n12485), .ZN(n12480) );
  NAND2_X1 U14775 ( .A1(n12480), .A2(n12865), .ZN(n12484) );
  INV_X1 U14776 ( .A(n12480), .ZN(n12481) );
  NAND2_X1 U14777 ( .A1(n12481), .A2(n12703), .ZN(n12482) );
  AND2_X1 U14778 ( .A1(n12484), .A2(n12482), .ZN(n12636) );
  NAND2_X1 U14779 ( .A1(n12638), .A2(n12484), .ZN(n12689) );
  XNOR2_X1 U14780 ( .A(n13071), .B(n12485), .ZN(n12486) );
  NOR2_X1 U14781 ( .A1(n12486), .A2(n12702), .ZN(n12487) );
  AOI21_X1 U14782 ( .B1(n12486), .B2(n12702), .A(n12487), .ZN(n12690) );
  NAND2_X1 U14783 ( .A1(n12689), .A2(n12690), .ZN(n12688) );
  INV_X1 U14784 ( .A(n12487), .ZN(n12488) );
  NAND2_X1 U14785 ( .A1(n12688), .A2(n12488), .ZN(n12590) );
  XNOR2_X1 U14786 ( .A(n12857), .B(n11800), .ZN(n12493) );
  NOR2_X1 U14787 ( .A1(n12493), .A2(n12701), .ZN(n12489) );
  AOI21_X1 U14788 ( .B1(n12493), .B2(n12701), .A(n12489), .ZN(n12591) );
  NAND2_X1 U14789 ( .A1(n12590), .A2(n12591), .ZN(n12595) );
  INV_X1 U14790 ( .A(n12489), .ZN(n12490) );
  NAND2_X1 U14791 ( .A1(n12696), .A2(n12844), .ZN(n12492) );
  INV_X1 U14792 ( .A(n12837), .ZN(n12699) );
  AOI22_X1 U14793 ( .A1(n12699), .A2(n12692), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12491) );
  OAI211_X1 U14794 ( .C1(n12866), .C2(n12694), .A(n12492), .B(n12491), .ZN(
        n12496) );
  NOR4_X1 U14795 ( .A1(n12494), .A2(n12493), .A3(n12701), .A4(n15172), .ZN(
        n12495) );
  AOI211_X1 U14796 ( .C1(n15186), .C2(n13003), .A(n12496), .B(n12495), .ZN(
        n12497) );
  OAI211_X1 U14797 ( .C1(n12499), .C2(n12595), .A(n12498), .B(n12497), .ZN(
        P3_U3160) );
  INV_X1 U14798 ( .A(n12500), .ZN(n12502) );
  NAND2_X1 U14799 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  XNOR2_X1 U14800 ( .A(n13721), .B(n12518), .ZN(n12506) );
  NOR2_X1 U14801 ( .A1(n14637), .A2(n6483), .ZN(n13244) );
  NAND2_X1 U14802 ( .A1(n13245), .A2(n13244), .ZN(n13241) );
  INV_X1 U14803 ( .A(n12505), .ZN(n12507) );
  NAND2_X1 U14804 ( .A1(n12507), .A2(n12506), .ZN(n12508) );
  NAND2_X1 U14805 ( .A1(n13256), .A2(n12562), .ZN(n12511) );
  XNOR2_X1 U14806 ( .A(n14644), .B(n12518), .ZN(n12510) );
  XOR2_X1 U14807 ( .A(n12511), .B(n12510), .Z(n14640) );
  INV_X1 U14808 ( .A(n12510), .ZN(n12512) );
  NAND2_X1 U14809 ( .A1(n12512), .A2(n12511), .ZN(n13182) );
  XNOR2_X1 U14810 ( .A(n13712), .B(n12518), .ZN(n12514) );
  NAND2_X1 U14811 ( .A1(n13615), .A2(n12562), .ZN(n12515) );
  XNOR2_X1 U14812 ( .A(n12514), .B(n12515), .ZN(n13183) );
  INV_X1 U14813 ( .A(n12514), .ZN(n12516) );
  NAND2_X1 U14814 ( .A1(n12516), .A2(n12515), .ZN(n12517) );
  INV_X1 U14815 ( .A(n13222), .ZN(n12522) );
  XNOR2_X1 U14816 ( .A(n12518), .B(n13707), .ZN(n12520) );
  AND2_X1 U14817 ( .A1(n13564), .A2(n12562), .ZN(n12519) );
  NAND2_X1 U14818 ( .A1(n12520), .A2(n12519), .ZN(n12523) );
  OAI21_X1 U14819 ( .B1(n12520), .B2(n12519), .A(n12523), .ZN(n13226) );
  NAND2_X1 U14820 ( .A1(n13579), .A2(n12562), .ZN(n12525) );
  XNOR2_X1 U14821 ( .A(n13702), .B(n12518), .ZN(n12524) );
  XOR2_X1 U14822 ( .A(n12525), .B(n12524), .Z(n13156) );
  INV_X1 U14823 ( .A(n12524), .ZN(n12526) );
  NAND2_X1 U14824 ( .A1(n12526), .A2(n12525), .ZN(n13204) );
  NAND2_X1 U14825 ( .A1(n13153), .A2(n13204), .ZN(n12527) );
  XNOR2_X1 U14826 ( .A(n13554), .B(n12518), .ZN(n12530) );
  NOR2_X1 U14827 ( .A1(n13538), .A2(n6483), .ZN(n12528) );
  XNOR2_X1 U14828 ( .A(n12530), .B(n12528), .ZN(n13203) );
  INV_X1 U14829 ( .A(n12528), .ZN(n12529) );
  NAND2_X1 U14830 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  XNOR2_X1 U14831 ( .A(n13541), .B(n12518), .ZN(n12535) );
  NAND2_X1 U14832 ( .A1(n13558), .A2(n12562), .ZN(n12533) );
  XOR2_X1 U14833 ( .A(n12535), .B(n12533), .Z(n13162) );
  INV_X1 U14834 ( .A(n13162), .ZN(n12532) );
  INV_X1 U14835 ( .A(n12533), .ZN(n12534) );
  NAND2_X1 U14836 ( .A1(n12535), .A2(n12534), .ZN(n12536) );
  NAND2_X1 U14837 ( .A1(n13163), .A2(n12536), .ZN(n12537) );
  XNOR2_X1 U14838 ( .A(n13521), .B(n12518), .ZN(n12538) );
  XNOR2_X1 U14839 ( .A(n12537), .B(n12538), .ZN(n13213) );
  NOR2_X1 U14840 ( .A1(n13536), .A2(n6483), .ZN(n13212) );
  NAND2_X1 U14841 ( .A1(n13213), .A2(n13212), .ZN(n13211) );
  INV_X1 U14842 ( .A(n12538), .ZN(n12539) );
  NAND2_X1 U14843 ( .A1(n12537), .A2(n12539), .ZN(n12540) );
  XNOR2_X1 U14844 ( .A(n13505), .B(n12547), .ZN(n12542) );
  XNOR2_X1 U14845 ( .A(n12541), .B(n12542), .ZN(n13142) );
  NAND2_X1 U14846 ( .A1(n13512), .A2(n12562), .ZN(n13145) );
  INV_X1 U14847 ( .A(n12542), .ZN(n12543) );
  NOR2_X1 U14848 ( .A1(n13460), .A2(n6483), .ZN(n12545) );
  XNOR2_X1 U14849 ( .A(n13490), .B(n12547), .ZN(n12544) );
  NAND2_X1 U14850 ( .A1(n12544), .A2(n12545), .ZN(n12546) );
  OAI21_X1 U14851 ( .B1(n12545), .B2(n12544), .A(n12546), .ZN(n13193) );
  NAND2_X1 U14852 ( .A1(n13194), .A2(n12546), .ZN(n13171) );
  XNOR2_X1 U14853 ( .A(n13739), .B(n12547), .ZN(n12550) );
  NAND2_X1 U14854 ( .A1(n13481), .A2(n12562), .ZN(n12549) );
  NOR2_X1 U14855 ( .A1(n12550), .A2(n12549), .ZN(n12551) );
  AOI21_X1 U14856 ( .B1(n12550), .B2(n12549), .A(n12551), .ZN(n13173) );
  INV_X1 U14857 ( .A(n12551), .ZN(n12552) );
  XNOR2_X1 U14858 ( .A(n13661), .B(n12518), .ZN(n12554) );
  NOR2_X1 U14859 ( .A1(n13461), .A2(n6483), .ZN(n12555) );
  XNOR2_X1 U14860 ( .A(n12554), .B(n12555), .ZN(n13233) );
  INV_X1 U14861 ( .A(n13233), .ZN(n12553) );
  INV_X1 U14862 ( .A(n12554), .ZN(n12557) );
  INV_X1 U14863 ( .A(n12555), .ZN(n12556) );
  NAND2_X1 U14864 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  XNOR2_X1 U14865 ( .A(n13656), .B(n12518), .ZN(n12560) );
  AND2_X1 U14866 ( .A1(n13441), .A2(n12562), .ZN(n12559) );
  NAND2_X1 U14867 ( .A1(n12560), .A2(n12559), .ZN(n12561) );
  OAI21_X1 U14868 ( .B1(n12560), .B2(n12559), .A(n12561), .ZN(n13132) );
  NAND2_X1 U14869 ( .A1(n13427), .A2(n12562), .ZN(n12563) );
  XNOR2_X1 U14870 ( .A(n12563), .B(n12518), .ZN(n12566) );
  NOR3_X1 U14871 ( .A1(n9255), .A2(n12566), .A3(n14930), .ZN(n12564) );
  AOI21_X1 U14872 ( .B1(n9255), .B2(n12566), .A(n12564), .ZN(n12569) );
  NAND3_X1 U14873 ( .A1(n13733), .A2(n13252), .A3(n12566), .ZN(n12565) );
  OAI21_X1 U14874 ( .B1(n13733), .B2(n12566), .A(n12565), .ZN(n12567) );
  OAI21_X1 U14875 ( .B1(n9255), .B2(n13252), .A(n14926), .ZN(n12568) );
  NAND2_X1 U14876 ( .A1(n13441), .A2(n13612), .ZN(n12571) );
  NAND2_X1 U14877 ( .A1(n13254), .A2(n13614), .ZN(n12570) );
  NAND2_X1 U14878 ( .A1(n12571), .A2(n12570), .ZN(n13412) );
  OAI22_X1 U14879 ( .A1(n13420), .A2(n14934), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12572), .ZN(n12573) );
  AOI21_X1 U14880 ( .B1(n13412), .B2(n13249), .A(n12573), .ZN(n12574) );
  INV_X1 U14881 ( .A(n12575), .ZN(n12577) );
  OAI222_X1 U14882 ( .A1(n12578), .A2(P3_U3151), .B1(n13123), .B2(n12577), 
        .C1(n12576), .C2(n13125), .ZN(P3_U3265) );
  OAI222_X1 U14883 ( .A1(n13781), .A2(n12580), .B1(P2_U3088), .B2(n12579), 
        .C1(n10093), .C2(n13783), .ZN(P2_U3297) );
  INV_X1 U14884 ( .A(n12581), .ZN(n12585) );
  AOI22_X1 U14885 ( .A1(n13001), .A2(P3_REG2_REG_29__SCAN_IN), .B1(n14604), 
        .B2(n15331), .ZN(n12582) );
  OAI21_X1 U14886 ( .B1(n12583), .B2(n12997), .A(n12582), .ZN(n12584) );
  AOI21_X1 U14887 ( .B1(n12585), .B2(n12999), .A(n12584), .ZN(n12586) );
  OAI21_X1 U14888 ( .B1(n12587), .B2(n13001), .A(n12586), .ZN(P3_U3204) );
  OAI222_X1 U14889 ( .A1(n14527), .A2(n12589), .B1(n14521), .B2(n12588), .C1(
        n8092), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U14890 ( .A(n12590), .ZN(n12593) );
  INV_X1 U14891 ( .A(n12591), .ZN(n12592) );
  NAND2_X1 U14892 ( .A1(n12593), .A2(n12592), .ZN(n12594) );
  OAI22_X1 U14893 ( .A1(n10252), .A2(n15302), .B1(n12596), .B2(n15303), .ZN(
        n12854) );
  AOI22_X1 U14894 ( .A1(n12854), .A2(n15178), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12597) );
  INV_X1 U14895 ( .A(n12598), .ZN(n12656) );
  AOI21_X1 U14896 ( .B1(n12704), .B2(n12599), .A(n12656), .ZN(n12605) );
  NAND2_X1 U14897 ( .A1(n12696), .A2(n12914), .ZN(n12601) );
  AOI22_X1 U14898 ( .A1(n12908), .A2(n12692), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12600) );
  OAI211_X1 U14899 ( .C1(n12933), .C2(n12694), .A(n12601), .B(n12600), .ZN(
        n12602) );
  AOI21_X1 U14900 ( .B1(n12603), .B2(n15186), .A(n12602), .ZN(n12604) );
  OAI21_X1 U14901 ( .B1(n12605), .B2(n15172), .A(n12604), .ZN(P3_U3156) );
  XNOR2_X1 U14902 ( .A(n12607), .B(n12606), .ZN(n12613) );
  NAND2_X1 U14903 ( .A1(n12696), .A2(n12969), .ZN(n12610) );
  NOR2_X1 U14904 ( .A1(n12608), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12820) );
  AOI21_X1 U14905 ( .B1(n12692), .B2(n12961), .A(n12820), .ZN(n12609) );
  OAI211_X1 U14906 ( .C1(n12991), .C2(n12694), .A(n12610), .B(n12609), .ZN(
        n12611) );
  AOI21_X1 U14907 ( .B1(n13095), .B2(n15186), .A(n12611), .ZN(n12612) );
  OAI21_X1 U14908 ( .B1(n12613), .B2(n15172), .A(n12612), .ZN(P3_U3159) );
  OAI211_X1 U14909 ( .C1(n12616), .C2(n12615), .A(n12614), .B(n15180), .ZN(
        n12624) );
  NAND2_X1 U14910 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15266) );
  INV_X1 U14911 ( .A(n15266), .ZN(n12617) );
  AOI21_X1 U14912 ( .B1(n15186), .B2(n12618), .A(n12617), .ZN(n12623) );
  AOI22_X1 U14913 ( .A1(n11810), .A2(n12619), .B1(n12692), .B2(n12715), .ZN(
        n12622) );
  OR2_X1 U14914 ( .A1(n15193), .A2(n12620), .ZN(n12621) );
  NAND4_X1 U14915 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        P3_U3161) );
  INV_X1 U14916 ( .A(n12625), .ZN(n13088) );
  OAI21_X1 U14917 ( .B1(n12628), .B2(n12627), .A(n12626), .ZN(n12629) );
  NAND2_X1 U14918 ( .A1(n12629), .A2(n15180), .ZN(n12633) );
  AOI22_X1 U14919 ( .A1(n12909), .A2(n12692), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12630) );
  OAI21_X1 U14920 ( .B1(n12934), .B2(n12694), .A(n12630), .ZN(n12631) );
  AOI21_X1 U14921 ( .B1(n12937), .B2(n12696), .A(n12631), .ZN(n12632) );
  OAI211_X1 U14922 ( .C1(n13088), .C2(n15170), .A(n12633), .B(n12632), .ZN(
        P3_U3163) );
  INV_X1 U14923 ( .A(n12634), .ZN(n12657) );
  INV_X1 U14924 ( .A(n12635), .ZN(n12637) );
  NOR3_X1 U14925 ( .A1(n12657), .A2(n12637), .A3(n12636), .ZN(n12640) );
  INV_X1 U14926 ( .A(n12638), .ZN(n12639) );
  OAI21_X1 U14927 ( .B1(n12640), .B2(n12639), .A(n15180), .ZN(n12644) );
  AOI22_X1 U14928 ( .A1(n12908), .A2(n12963), .B1(n12962), .B2(n12702), .ZN(
        n12878) );
  OAI22_X1 U14929 ( .A1(n12878), .A2(n15189), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12641), .ZN(n12642) );
  AOI21_X1 U14930 ( .B1(n12881), .B2(n12696), .A(n12642), .ZN(n12643) );
  OAI211_X1 U14931 ( .C1(n13075), .C2(n15170), .A(n12644), .B(n12643), .ZN(
        P3_U3165) );
  XNOR2_X1 U14932 ( .A(n12645), .B(n12646), .ZN(n12652) );
  NAND2_X1 U14933 ( .A1(n12696), .A2(n12995), .ZN(n12648) );
  AOI22_X1 U14934 ( .A1(n12964), .A2(n12692), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12647) );
  OAI211_X1 U14935 ( .C1(n12990), .C2(n12694), .A(n12648), .B(n12647), .ZN(
        n12649) );
  AOI21_X1 U14936 ( .B1(n12650), .B2(n15186), .A(n12649), .ZN(n12651) );
  OAI21_X1 U14937 ( .B1(n12652), .B2(n15172), .A(n12651), .ZN(P3_U3168) );
  INV_X1 U14938 ( .A(n12653), .ZN(n12655) );
  NOR3_X1 U14939 ( .A1(n12656), .A2(n12655), .A3(n12654), .ZN(n12658) );
  OAI21_X1 U14940 ( .B1(n12658), .B2(n12657), .A(n15180), .ZN(n12665) );
  OR2_X1 U14941 ( .A1(n12659), .A2(n15302), .ZN(n12661) );
  OR2_X1 U14942 ( .A1(n12865), .A2(n15303), .ZN(n12660) );
  AND2_X1 U14943 ( .A1(n12661), .A2(n12660), .ZN(n12888) );
  INV_X1 U14944 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12662) );
  OAI22_X1 U14945 ( .A1(n12888), .A2(n15189), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12662), .ZN(n12663) );
  AOI21_X1 U14946 ( .B1(n12896), .B2(n12696), .A(n12663), .ZN(n12664) );
  OAI211_X1 U14947 ( .C1(n12898), .C2(n15170), .A(n12665), .B(n12664), .ZN(
        P3_U3169) );
  XNOR2_X1 U14948 ( .A(n12667), .B(n12666), .ZN(n12672) );
  NAND2_X1 U14949 ( .A1(n12696), .A2(n12945), .ZN(n12669) );
  AOI22_X1 U14950 ( .A1(n12705), .A2(n12692), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12668) );
  OAI211_X1 U14951 ( .C1(n12979), .C2(n12694), .A(n12669), .B(n12668), .ZN(
        n12670) );
  AOI21_X1 U14952 ( .B1(n12950), .B2(n15186), .A(n12670), .ZN(n12671) );
  OAI21_X1 U14953 ( .B1(n12672), .B2(n15172), .A(n12671), .ZN(P3_U3173) );
  AOI21_X1 U14954 ( .B1(n12909), .B2(n12673), .A(n6565), .ZN(n12679) );
  AOI22_X1 U14955 ( .A1(n12704), .A2(n12962), .B1(n12963), .B2(n12705), .ZN(
        n12920) );
  OAI22_X1 U14956 ( .A1(n12920), .A2(n15189), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12674), .ZN(n12677) );
  INV_X1 U14957 ( .A(n12675), .ZN(n13084) );
  NOR2_X1 U14958 ( .A1(n13084), .A2(n15170), .ZN(n12676) );
  AOI211_X1 U14959 ( .C1(n12924), .C2(n12696), .A(n12677), .B(n12676), .ZN(
        n12678) );
  OAI21_X1 U14960 ( .B1(n12679), .B2(n15172), .A(n12678), .ZN(P3_U3175) );
  XNOR2_X1 U14961 ( .A(n12681), .B(n12680), .ZN(n12687) );
  NAND2_X1 U14962 ( .A1(n12706), .A2(n12692), .ZN(n12682) );
  NAND2_X1 U14963 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12796)
         );
  OAI211_X1 U14964 ( .C1(n12978), .C2(n12694), .A(n12682), .B(n12796), .ZN(
        n12685) );
  INV_X1 U14965 ( .A(n12683), .ZN(n13101) );
  NOR2_X1 U14966 ( .A1(n13101), .A2(n15170), .ZN(n12684) );
  AOI211_X1 U14967 ( .C1(n12982), .C2(n12696), .A(n12685), .B(n12684), .ZN(
        n12686) );
  OAI21_X1 U14968 ( .B1(n12687), .B2(n15172), .A(n12686), .ZN(P3_U3178) );
  OAI21_X1 U14969 ( .B1(n12690), .B2(n12689), .A(n12688), .ZN(n12691) );
  NAND2_X1 U14970 ( .A1(n12691), .A2(n15180), .ZN(n12698) );
  AOI22_X1 U14971 ( .A1(n12701), .A2(n12692), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12693) );
  OAI21_X1 U14972 ( .B1(n12865), .B2(n12694), .A(n12693), .ZN(n12695) );
  AOI21_X1 U14973 ( .B1(n12869), .B2(n12696), .A(n12695), .ZN(n12697) );
  OAI211_X1 U14974 ( .C1(n13071), .C2(n15170), .A(n12698), .B(n12697), .ZN(
        P3_U3180) );
  MUX2_X1 U14975 ( .A(n14603), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12720), .Z(
        P3_U3522) );
  MUX2_X1 U14976 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12699), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14977 ( .A(n12700), .B(P3_DATAO_REG_28__SCAN_IN), .S(n12720), .Z(
        P3_U3519) );
  MUX2_X1 U14978 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12701), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14979 ( .A(n12702), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12720), .Z(
        P3_U3517) );
  MUX2_X1 U14980 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12703), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14981 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12908), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14982 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12704), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14983 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12909), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14984 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12705), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14985 ( .A(n12961), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12720), .Z(
        P3_U3511) );
  MUX2_X1 U14986 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12706), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14987 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12964), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14988 ( .A(n12707), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12720), .Z(
        P3_U3508) );
  MUX2_X1 U14989 ( .A(n12708), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12720), .Z(
        P3_U3507) );
  MUX2_X1 U14990 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12709), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14991 ( .A(n12710), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12720), .Z(
        P3_U3505) );
  MUX2_X1 U14992 ( .A(n12711), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12720), .Z(
        P3_U3504) );
  MUX2_X1 U14993 ( .A(n12712), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12720), .Z(
        P3_U3503) );
  MUX2_X1 U14994 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12713), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14995 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12714), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14996 ( .A(n12715), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12720), .Z(
        P3_U3500) );
  MUX2_X1 U14997 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12716), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14998 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n11810), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14999 ( .A(n12717), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12720), .Z(
        P3_U3497) );
  MUX2_X1 U15000 ( .A(n12718), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12720), .Z(
        P3_U3496) );
  MUX2_X1 U15001 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12719), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15002 ( .A(n12721), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12720), .Z(
        P3_U3494) );
  MUX2_X1 U15003 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12722), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15004 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12723), .S(P3_U3897), .Z(
        P3_U3492) );
  INV_X1 U15005 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12726) );
  OR2_X1 U15006 ( .A1(n12735), .A2(n12726), .ZN(n12760) );
  NAND2_X1 U15007 ( .A1(n12735), .A2(n12726), .ZN(n12727) );
  AND2_X1 U15008 ( .A1(n12760), .A2(n12727), .ZN(n12742) );
  INV_X1 U15009 ( .A(n12742), .ZN(n12729) );
  INV_X1 U15010 ( .A(n12753), .ZN(n12728) );
  AOI21_X1 U15011 ( .B1(n12730), .B2(n12729), .A(n12728), .ZN(n12752) );
  NAND2_X1 U15012 ( .A1(n12732), .A2(n12731), .ZN(n12734) );
  XNOR2_X1 U15013 ( .A(n12735), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12741) );
  OAI21_X1 U15014 ( .B1(n12736), .B2(n12741), .A(n12757), .ZN(n12750) );
  NAND2_X1 U15015 ( .A1(n15245), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n12737) );
  OAI211_X1 U15016 ( .C1(n15285), .C2(n12756), .A(n12738), .B(n12737), .ZN(
        n12749) );
  INV_X1 U15017 ( .A(n12739), .ZN(n12740) );
  NAND2_X1 U15018 ( .A1(n12740), .A2(n12257), .ZN(n12744) );
  MUX2_X1 U15019 ( .A(n12742), .B(n12741), .S(n12823), .Z(n12743) );
  NAND3_X1 U15020 ( .A1(n12745), .A2(n12744), .A3(n12743), .ZN(n12762) );
  INV_X1 U15021 ( .A(n12762), .ZN(n12747) );
  AOI21_X1 U15022 ( .B1(n12745), .B2(n12744), .A(n12743), .ZN(n12746) );
  NOR3_X1 U15023 ( .A1(n12747), .A2(n12746), .A3(n15241), .ZN(n12748) );
  AOI211_X1 U15024 ( .C1(n15287), .C2(n12750), .A(n12749), .B(n12748), .ZN(
        n12751) );
  OAI21_X1 U15025 ( .B1(n12752), .B2(n15291), .A(n12751), .ZN(P3_U3196) );
  INV_X1 U15026 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12755) );
  AOI21_X1 U15027 ( .B1(n12755), .B2(n12754), .A(n12786), .ZN(n12774) );
  NAND2_X1 U15028 ( .A1(n12756), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12759) );
  OAI21_X1 U15029 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12758), .A(n12799), 
        .ZN(n12772) );
  MUX2_X1 U15030 ( .A(n12760), .B(n12759), .S(n12823), .Z(n12761) );
  NAND2_X1 U15031 ( .A1(n12762), .A2(n12761), .ZN(n12775) );
  XNOR2_X1 U15032 ( .A(n12775), .B(n12798), .ZN(n12764) );
  MUX2_X1 U15033 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12823), .Z(n12763) );
  NOR2_X1 U15034 ( .A1(n12764), .A2(n12763), .ZN(n12776) );
  AOI21_X1 U15035 ( .B1(n12764), .B2(n12763), .A(n12776), .ZN(n12770) );
  NOR2_X1 U15036 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12765), .ZN(n12768) );
  NOR2_X1 U15037 ( .A1(n15296), .A2(n12766), .ZN(n12767) );
  AOI211_X1 U15038 ( .C1(n14584), .C2(n12785), .A(n12768), .B(n12767), .ZN(
        n12769) );
  OAI21_X1 U15039 ( .B1(n12770), .B2(n15241), .A(n12769), .ZN(n12771) );
  AOI21_X1 U15040 ( .B1(n15287), .B2(n12772), .A(n12771), .ZN(n12773) );
  OAI21_X1 U15041 ( .B1(n12774), .B2(n15291), .A(n12773), .ZN(P3_U3197) );
  MUX2_X1 U15042 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12823), .Z(n12782) );
  MUX2_X1 U15043 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12823), .Z(n12780) );
  INV_X1 U15044 ( .A(n12775), .ZN(n12777) );
  AOI21_X1 U15045 ( .B1(n12777), .B2(n12785), .A(n12776), .ZN(n14573) );
  INV_X1 U15046 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12788) );
  INV_X1 U15047 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12778) );
  MUX2_X1 U15048 ( .A(n12788), .B(n12778), .S(n12823), .Z(n12779) );
  INV_X1 U15049 ( .A(n12801), .ZN(n14566) );
  NOR2_X1 U15050 ( .A1(n12779), .A2(n14566), .ZN(n14569) );
  NAND2_X1 U15051 ( .A1(n12779), .A2(n14566), .ZN(n14570) );
  OAI21_X1 U15052 ( .B1(n14573), .B2(n14569), .A(n14570), .ZN(n14588) );
  XNOR2_X1 U15053 ( .A(n12780), .B(n12803), .ZN(n14589) );
  NOR2_X1 U15054 ( .A1(n14588), .A2(n14589), .ZN(n14587) );
  XOR2_X1 U15055 ( .A(n12818), .B(n12828), .Z(n12781) );
  NOR2_X1 U15056 ( .A1(n12781), .A2(n12782), .ZN(n12826) );
  AOI21_X1 U15057 ( .B1(n12782), .B2(n12781), .A(n12826), .ZN(n12813) );
  INV_X1 U15058 ( .A(n12818), .ZN(n12827) );
  INV_X1 U15059 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12783) );
  AND2_X1 U15060 ( .A1(n12818), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12814) );
  AOI21_X1 U15061 ( .B1(n12827), .B2(n12783), .A(n12814), .ZN(n12794) );
  NOR2_X1 U15062 ( .A1(n12787), .A2(n12786), .ZN(n14577) );
  OR2_X1 U15063 ( .A1(n12801), .A2(n12788), .ZN(n12790) );
  NAND2_X1 U15064 ( .A1(n12801), .A2(n12788), .ZN(n12789) );
  AND2_X1 U15065 ( .A1(n12790), .A2(n12789), .ZN(n14576) );
  INV_X1 U15066 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14595) );
  OAI21_X1 U15067 ( .B1(n12794), .B2(n12793), .A(n12816), .ZN(n12795) );
  NAND2_X1 U15068 ( .A1(n12795), .A2(n14593), .ZN(n12812) );
  OAI21_X1 U15069 ( .B1(n15296), .B2(n8553), .A(n12796), .ZN(n12810) );
  NAND2_X1 U15070 ( .A1(n12798), .A2(n12797), .ZN(n12800) );
  XOR2_X1 U15071 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12801), .Z(n14567) );
  AOI22_X1 U15072 ( .A1(n14568), .A2(n14567), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n12801), .ZN(n12802) );
  NAND2_X1 U15073 ( .A1(n12804), .A2(n12803), .ZN(n12805) );
  XNOR2_X1 U15074 ( .A(n12818), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12806) );
  INV_X1 U15075 ( .A(n12817), .ZN(n12808) );
  NAND3_X1 U15076 ( .A1(n14585), .A2(n12806), .A3(n12805), .ZN(n12807) );
  AOI21_X1 U15077 ( .B1(n12808), .B2(n12807), .A(n15257), .ZN(n12809) );
  AOI211_X1 U15078 ( .C1(n14584), .C2(n12827), .A(n12810), .B(n12809), .ZN(
        n12811) );
  OAI211_X1 U15079 ( .C1(n12813), .C2(n15241), .A(n12812), .B(n12811), .ZN(
        P3_U3200) );
  INV_X1 U15080 ( .A(n12814), .ZN(n12815) );
  XNOR2_X1 U15081 ( .A(n12822), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12825) );
  AOI21_X1 U15082 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n12818), .A(n12817), 
        .ZN(n12819) );
  XNOR2_X1 U15083 ( .A(n12822), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12824) );
  AOI21_X1 U15084 ( .B1(n15245), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12820), 
        .ZN(n12821) );
  OAI21_X1 U15085 ( .B1(n15285), .B2(n12822), .A(n12821), .ZN(n12832) );
  MUX2_X1 U15086 ( .A(n12825), .B(n12824), .S(n12823), .Z(n12830) );
  AOI21_X1 U15087 ( .B1(n12828), .B2(n12827), .A(n12826), .ZN(n12829) );
  XOR2_X1 U15088 ( .A(n12830), .B(n12829), .Z(n12831) );
  OAI21_X1 U15089 ( .B1(n12834), .B2(n15291), .A(n12833), .ZN(P3_U3201) );
  NOR2_X1 U15090 ( .A1(n12835), .A2(n15308), .ZN(n12840) );
  OAI21_X1 U15091 ( .B1(n12849), .B2(n12836), .A(n12842), .ZN(n12839) );
  OAI22_X1 U15092 ( .A1(n12866), .A2(n15302), .B1(n12837), .B2(n15303), .ZN(
        n12838) );
  OAI21_X1 U15093 ( .B1(n12843), .B2(n12842), .A(n12841), .ZN(n13004) );
  INV_X1 U15094 ( .A(n13003), .ZN(n12846) );
  AOI22_X1 U15095 ( .A1(n13001), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15331), 
        .B2(n12844), .ZN(n12845) );
  OAI21_X1 U15096 ( .B1(n12846), .B2(n12997), .A(n12845), .ZN(n12847) );
  AOI21_X1 U15097 ( .B1(n13004), .B2(n12999), .A(n12847), .ZN(n12848) );
  OAI21_X1 U15098 ( .B1(n13006), .B2(n13001), .A(n12848), .ZN(P3_U3205) );
  AOI21_X1 U15099 ( .B1(n12852), .B2(n12850), .A(n12849), .ZN(n12856) );
  OAI21_X1 U15100 ( .B1(n12853), .B2(n12852), .A(n12851), .ZN(n13008) );
  AOI21_X1 U15101 ( .B1(n13008), .B2(n15324), .A(n12854), .ZN(n12855) );
  OAI21_X1 U15102 ( .B1(n12856), .B2(n15308), .A(n12855), .ZN(n13007) );
  INV_X1 U15103 ( .A(n13007), .ZN(n12862) );
  INV_X1 U15104 ( .A(n12857), .ZN(n13067) );
  AOI22_X1 U15105 ( .A1(n13001), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15331), 
        .B2(n12858), .ZN(n12859) );
  OAI21_X1 U15106 ( .B1(n13067), .B2(n12997), .A(n12859), .ZN(n12860) );
  AOI21_X1 U15107 ( .B1(n13008), .B2(n15332), .A(n12860), .ZN(n12861) );
  OAI21_X1 U15108 ( .B1(n12862), .B2(n13001), .A(n12861), .ZN(P3_U3206) );
  XOR2_X1 U15109 ( .A(n12868), .B(n12863), .Z(n12864) );
  INV_X1 U15110 ( .A(n13011), .ZN(n12873) );
  XOR2_X1 U15111 ( .A(n12868), .B(n12867), .Z(n13012) );
  AOI22_X1 U15112 ( .A1(n13001), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15331), 
        .B2(n12869), .ZN(n12870) );
  OAI21_X1 U15113 ( .B1(n13071), .B2(n12997), .A(n12870), .ZN(n12871) );
  AOI21_X1 U15114 ( .B1(n13012), .B2(n12999), .A(n12871), .ZN(n12872) );
  OAI21_X1 U15115 ( .B1(n12873), .B2(n13001), .A(n12872), .ZN(P3_U3207) );
  XNOR2_X1 U15116 ( .A(n12874), .B(n12876), .ZN(n12880) );
  OAI211_X1 U15117 ( .C1(n12877), .C2(n12876), .A(n12875), .B(n15317), .ZN(
        n12879) );
  OAI211_X1 U15118 ( .C1(n12912), .C2(n12880), .A(n12879), .B(n12878), .ZN(
        n13015) );
  INV_X1 U15119 ( .A(n13015), .ZN(n12885) );
  INV_X1 U15120 ( .A(n12880), .ZN(n13016) );
  AOI22_X1 U15121 ( .A1(n13001), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15331), 
        .B2(n12881), .ZN(n12882) );
  OAI21_X1 U15122 ( .B1(n13075), .B2(n12997), .A(n12882), .ZN(n12883) );
  AOI21_X1 U15123 ( .B1(n13016), .B2(n15332), .A(n12883), .ZN(n12884) );
  OAI21_X1 U15124 ( .B1(n12885), .B2(n13001), .A(n12884), .ZN(P3_U3208) );
  OAI211_X1 U15125 ( .C1(n12887), .C2(n12892), .A(n12886), .B(n15317), .ZN(
        n12889) );
  NAND2_X1 U15126 ( .A1(n12889), .A2(n12888), .ZN(n13023) );
  INV_X1 U15127 ( .A(n13023), .ZN(n12901) );
  INV_X1 U15128 ( .A(n12890), .ZN(n12891) );
  NAND2_X1 U15129 ( .A1(n12905), .A2(n12891), .ZN(n12893) );
  NAND2_X1 U15130 ( .A1(n12893), .A2(n12892), .ZN(n12895) );
  NAND2_X1 U15131 ( .A1(n12895), .A2(n12894), .ZN(n13020) );
  AOI22_X1 U15132 ( .A1(n13001), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15331), 
        .B2(n12896), .ZN(n12897) );
  OAI21_X1 U15133 ( .B1(n12898), .B2(n12997), .A(n12897), .ZN(n12899) );
  AOI21_X1 U15134 ( .B1(n13020), .B2(n12999), .A(n12899), .ZN(n12900) );
  OAI21_X1 U15135 ( .B1(n12901), .B2(n13001), .A(n12900), .ZN(P3_U3209) );
  OR2_X1 U15136 ( .A1(n12903), .A2(n12902), .ZN(n12904) );
  NAND2_X1 U15137 ( .A1(n12905), .A2(n12904), .ZN(n12913) );
  OAI211_X1 U15138 ( .C1(n6609), .C2(n12907), .A(n12906), .B(n15317), .ZN(
        n12911) );
  AOI22_X1 U15139 ( .A1(n12909), .A2(n12963), .B1(n12962), .B2(n12908), .ZN(
        n12910) );
  OAI211_X1 U15140 ( .C1(n12912), .C2(n12913), .A(n12911), .B(n12910), .ZN(
        n13024) );
  INV_X1 U15141 ( .A(n13024), .ZN(n12918) );
  INV_X1 U15142 ( .A(n12913), .ZN(n13025) );
  AOI22_X1 U15143 ( .A1(n13001), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12914), 
        .B2(n15331), .ZN(n12915) );
  OAI21_X1 U15144 ( .B1(n13080), .B2(n12997), .A(n12915), .ZN(n12916) );
  AOI21_X1 U15145 ( .B1(n13025), .B2(n15332), .A(n12916), .ZN(n12917) );
  OAI21_X1 U15146 ( .B1(n12918), .B2(n13001), .A(n12917), .ZN(P3_U3210) );
  XNOR2_X1 U15147 ( .A(n12919), .B(n12923), .ZN(n12921) );
  OAI21_X1 U15148 ( .B1(n12921), .B2(n15308), .A(n12920), .ZN(n13028) );
  INV_X1 U15149 ( .A(n13028), .ZN(n12928) );
  XOR2_X1 U15150 ( .A(n12923), .B(n12922), .Z(n13029) );
  AOI22_X1 U15151 ( .A1(n13001), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15331), 
        .B2(n12924), .ZN(n12925) );
  OAI21_X1 U15152 ( .B1(n13084), .B2(n12997), .A(n12925), .ZN(n12926) );
  AOI21_X1 U15153 ( .B1(n13029), .B2(n12999), .A(n12926), .ZN(n12927) );
  OAI21_X1 U15154 ( .B1(n12928), .B2(n13001), .A(n12927), .ZN(P3_U3211) );
  INV_X1 U15155 ( .A(n12929), .ZN(n12930) );
  AOI21_X1 U15156 ( .B1(n12936), .B2(n12931), .A(n12930), .ZN(n12932) );
  OAI222_X1 U15157 ( .A1(n15302), .A2(n12934), .B1(n15303), .B2(n12933), .C1(
        n15308), .C2(n12932), .ZN(n13032) );
  INV_X1 U15158 ( .A(n13032), .ZN(n12941) );
  XOR2_X1 U15159 ( .A(n12936), .B(n12935), .Z(n13033) );
  AOI22_X1 U15160 ( .A1(n13001), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15331), 
        .B2(n12937), .ZN(n12938) );
  OAI21_X1 U15161 ( .B1(n13088), .B2(n12997), .A(n12938), .ZN(n12939) );
  AOI21_X1 U15162 ( .B1(n13033), .B2(n12999), .A(n12939), .ZN(n12940) );
  OAI21_X1 U15163 ( .B1(n12941), .B2(n13001), .A(n12940), .ZN(P3_U3212) );
  XNOR2_X1 U15164 ( .A(n12942), .B(n12951), .ZN(n12943) );
  OAI222_X1 U15165 ( .A1(n15302), .A2(n12979), .B1(n15303), .B2(n12944), .C1(
        n12943), .C2(n15308), .ZN(n13036) );
  INV_X1 U15166 ( .A(n13036), .ZN(n12957) );
  INV_X1 U15167 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12948) );
  INV_X1 U15168 ( .A(n12945), .ZN(n12947) );
  OAI22_X1 U15169 ( .A1(n15334), .A2(n12948), .B1(n12947), .B2(n12946), .ZN(
        n12949) );
  AOI21_X1 U15170 ( .B1(n12950), .B2(n14607), .A(n12949), .ZN(n12956) );
  NAND2_X1 U15171 ( .A1(n12952), .A2(n12951), .ZN(n12953) );
  NAND2_X1 U15172 ( .A1(n13037), .A2(n12999), .ZN(n12955) );
  OAI211_X1 U15173 ( .C1(n12957), .C2(n13001), .A(n12956), .B(n12955), .ZN(
        P3_U3213) );
  NAND2_X1 U15174 ( .A1(n12958), .A2(n7029), .ZN(n12959) );
  NAND3_X1 U15175 ( .A1(n12960), .A2(n15317), .A3(n12959), .ZN(n12966) );
  AOI22_X1 U15176 ( .A1(n12964), .A2(n12963), .B1(n12962), .B2(n12961), .ZN(
        n12965) );
  XNOR2_X1 U15177 ( .A(n12968), .B(n12967), .ZN(n13040) );
  INV_X1 U15178 ( .A(n13095), .ZN(n12971) );
  AOI22_X1 U15179 ( .A1(n13001), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15331), 
        .B2(n12969), .ZN(n12970) );
  OAI21_X1 U15180 ( .B1(n12971), .B2(n12997), .A(n12970), .ZN(n12972) );
  AOI21_X1 U15181 ( .B1(n13040), .B2(n12999), .A(n12972), .ZN(n12973) );
  OAI21_X1 U15182 ( .B1(n13042), .B2(n13001), .A(n12973), .ZN(P3_U3214) );
  INV_X1 U15183 ( .A(n12974), .ZN(n12975) );
  AOI21_X1 U15184 ( .B1(n12980), .B2(n12976), .A(n12975), .ZN(n12977) );
  OAI222_X1 U15185 ( .A1(n15303), .A2(n12979), .B1(n15302), .B2(n12978), .C1(
        n15308), .C2(n12977), .ZN(n13046) );
  INV_X1 U15186 ( .A(n13046), .ZN(n12986) );
  XNOR2_X1 U15187 ( .A(n12981), .B(n12980), .ZN(n13047) );
  AOI22_X1 U15188 ( .A1(n13001), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15331), 
        .B2(n12982), .ZN(n12983) );
  OAI21_X1 U15189 ( .B1(n13101), .B2(n12997), .A(n12983), .ZN(n12984) );
  AOI21_X1 U15190 ( .B1(n13047), .B2(n12999), .A(n12984), .ZN(n12985) );
  OAI21_X1 U15191 ( .B1(n12986), .B2(n13001), .A(n12985), .ZN(P3_U3215) );
  XNOR2_X1 U15192 ( .A(n12987), .B(n12988), .ZN(n12989) );
  OAI222_X1 U15193 ( .A1(n15303), .A2(n12991), .B1(n15302), .B2(n12990), .C1(
        n12989), .C2(n15308), .ZN(n13050) );
  INV_X1 U15194 ( .A(n13050), .ZN(n13002) );
  OAI21_X1 U15195 ( .B1(n12994), .B2(n12993), .A(n12992), .ZN(n13051) );
  AOI22_X1 U15196 ( .A1(n13001), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15331), 
        .B2(n12995), .ZN(n12996) );
  OAI21_X1 U15197 ( .B1(n13105), .B2(n12997), .A(n12996), .ZN(n12998) );
  AOI21_X1 U15198 ( .B1(n13051), .B2(n12999), .A(n12998), .ZN(n13000) );
  OAI21_X1 U15199 ( .B1(n13002), .B2(n13001), .A(n13000), .ZN(P3_U3216) );
  AOI22_X1 U15200 ( .A1(n13004), .A2(n15339), .B1(n15325), .B2(n13003), .ZN(
        n13005) );
  NAND2_X1 U15201 ( .A1(n13006), .A2(n13005), .ZN(n13063) );
  MUX2_X1 U15202 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13063), .S(n15374), .Z(
        P3_U3487) );
  INV_X1 U15203 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13009) );
  INV_X1 U15204 ( .A(n15359), .ZN(n15355) );
  AOI21_X1 U15205 ( .B1(n15355), .B2(n13008), .A(n13007), .ZN(n13064) );
  MUX2_X1 U15206 ( .A(n13009), .B(n13064), .S(n15374), .Z(n13010) );
  OAI21_X1 U15207 ( .B1(n13067), .B2(n13062), .A(n13010), .ZN(P3_U3486) );
  INV_X1 U15208 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13013) );
  MUX2_X1 U15209 ( .A(n13013), .B(n13068), .S(n15374), .Z(n13014) );
  OAI21_X1 U15210 ( .B1(n13071), .B2(n13062), .A(n13014), .ZN(P3_U3485) );
  INV_X1 U15211 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13017) );
  AOI21_X1 U15212 ( .B1(n15355), .B2(n13016), .A(n13015), .ZN(n13072) );
  MUX2_X1 U15213 ( .A(n13017), .B(n13072), .S(n15374), .Z(n13018) );
  OAI21_X1 U15214 ( .B1(n13075), .B2(n13062), .A(n13018), .ZN(P3_U3484) );
  AND2_X1 U15215 ( .A1(n13019), .A2(n15325), .ZN(n13022) );
  AND2_X1 U15216 ( .A1(n13020), .A2(n15339), .ZN(n13021) );
  MUX2_X1 U15217 ( .A(n13076), .B(P3_REG1_REG_24__SCAN_IN), .S(n15371), .Z(
        P3_U3483) );
  INV_X1 U15218 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13026) );
  AOI21_X1 U15219 ( .B1(n15355), .B2(n13025), .A(n13024), .ZN(n13077) );
  MUX2_X1 U15220 ( .A(n13026), .B(n13077), .S(n15374), .Z(n13027) );
  OAI21_X1 U15221 ( .B1(n13080), .B2(n13062), .A(n13027), .ZN(P3_U3482) );
  INV_X1 U15222 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13030) );
  AOI21_X1 U15223 ( .B1(n15339), .B2(n13029), .A(n13028), .ZN(n13081) );
  MUX2_X1 U15224 ( .A(n13030), .B(n13081), .S(n15374), .Z(n13031) );
  OAI21_X1 U15225 ( .B1(n13084), .B2(n13062), .A(n13031), .ZN(P3_U3481) );
  INV_X1 U15226 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13034) );
  AOI21_X1 U15227 ( .B1(n15339), .B2(n13033), .A(n13032), .ZN(n13085) );
  MUX2_X1 U15228 ( .A(n13034), .B(n13085), .S(n15374), .Z(n13035) );
  OAI21_X1 U15229 ( .B1(n13088), .B2(n13062), .A(n13035), .ZN(P3_U3480) );
  INV_X1 U15230 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13038) );
  AOI21_X1 U15231 ( .B1(n13037), .B2(n15339), .A(n13036), .ZN(n13089) );
  MUX2_X1 U15232 ( .A(n13038), .B(n13089), .S(n15374), .Z(n13039) );
  OAI21_X1 U15233 ( .B1(n13092), .B2(n13062), .A(n13039), .ZN(P3_U3479) );
  NAND2_X1 U15234 ( .A1(n13040), .A2(n15339), .ZN(n13041) );
  NAND2_X1 U15235 ( .A1(n13042), .A2(n13041), .ZN(n13093) );
  MUX2_X1 U15236 ( .A(n13093), .B(P3_REG1_REG_19__SCAN_IN), .S(n15371), .Z(
        n13043) );
  AOI21_X1 U15237 ( .B1(n13044), .B2(n13095), .A(n13043), .ZN(n13045) );
  INV_X1 U15238 ( .A(n13045), .ZN(P3_U3478) );
  INV_X1 U15239 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13048) );
  AOI21_X1 U15240 ( .B1(n13047), .B2(n15339), .A(n13046), .ZN(n13098) );
  MUX2_X1 U15241 ( .A(n13048), .B(n13098), .S(n15374), .Z(n13049) );
  OAI21_X1 U15242 ( .B1(n13101), .B2(n13062), .A(n13049), .ZN(P3_U3477) );
  INV_X1 U15243 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13052) );
  AOI21_X1 U15244 ( .B1(n15339), .B2(n13051), .A(n13050), .ZN(n13102) );
  MUX2_X1 U15245 ( .A(n13052), .B(n13102), .S(n15374), .Z(n13053) );
  OAI21_X1 U15246 ( .B1(n13105), .B2(n13062), .A(n13053), .ZN(P3_U3476) );
  AOI22_X1 U15247 ( .A1(n13055), .A2(n15339), .B1(n15325), .B2(n13054), .ZN(
        n13056) );
  NAND2_X1 U15248 ( .A1(n13057), .A2(n13056), .ZN(n13106) );
  MUX2_X1 U15249 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13106), .S(n15374), .Z(
        P3_U3475) );
  INV_X1 U15250 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13060) );
  AOI21_X1 U15251 ( .B1(n15339), .B2(n13059), .A(n13058), .ZN(n13107) );
  MUX2_X1 U15252 ( .A(n13060), .B(n13107), .S(n15374), .Z(n13061) );
  OAI21_X1 U15253 ( .B1(n13111), .B2(n13062), .A(n13061), .ZN(P3_U3474) );
  MUX2_X1 U15254 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13063), .S(n15365), .Z(
        P3_U3455) );
  INV_X1 U15255 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13065) );
  MUX2_X1 U15256 ( .A(n13065), .B(n13064), .S(n15365), .Z(n13066) );
  OAI21_X1 U15257 ( .B1(n13067), .B2(n13110), .A(n13066), .ZN(P3_U3454) );
  INV_X1 U15258 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13069) );
  MUX2_X1 U15259 ( .A(n13069), .B(n13068), .S(n15365), .Z(n13070) );
  OAI21_X1 U15260 ( .B1(n13071), .B2(n13110), .A(n13070), .ZN(P3_U3453) );
  INV_X1 U15261 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13073) );
  MUX2_X1 U15262 ( .A(n13073), .B(n13072), .S(n15365), .Z(n13074) );
  OAI21_X1 U15263 ( .B1(n13075), .B2(n13110), .A(n13074), .ZN(P3_U3452) );
  MUX2_X1 U15264 ( .A(n13076), .B(P3_REG0_REG_24__SCAN_IN), .S(n15363), .Z(
        P3_U3451) );
  INV_X1 U15265 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13078) );
  MUX2_X1 U15266 ( .A(n13078), .B(n13077), .S(n15365), .Z(n13079) );
  OAI21_X1 U15267 ( .B1(n13080), .B2(n13110), .A(n13079), .ZN(P3_U3450) );
  INV_X1 U15268 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13082) );
  MUX2_X1 U15269 ( .A(n13082), .B(n13081), .S(n15365), .Z(n13083) );
  OAI21_X1 U15270 ( .B1(n13084), .B2(n13110), .A(n13083), .ZN(P3_U3449) );
  INV_X1 U15271 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13086) );
  MUX2_X1 U15272 ( .A(n13086), .B(n13085), .S(n15365), .Z(n13087) );
  OAI21_X1 U15273 ( .B1(n13088), .B2(n13110), .A(n13087), .ZN(P3_U3448) );
  INV_X1 U15274 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13090) );
  MUX2_X1 U15275 ( .A(n13090), .B(n13089), .S(n15365), .Z(n13091) );
  OAI21_X1 U15276 ( .B1(n13092), .B2(n13110), .A(n13091), .ZN(P3_U3447) );
  INV_X1 U15277 ( .A(n13110), .ZN(n13096) );
  MUX2_X1 U15278 ( .A(n13093), .B(P3_REG0_REG_19__SCAN_IN), .S(n15363), .Z(
        n13094) );
  AOI21_X1 U15279 ( .B1(n13096), .B2(n13095), .A(n13094), .ZN(n13097) );
  INV_X1 U15280 ( .A(n13097), .ZN(P3_U3446) );
  INV_X1 U15281 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13099) );
  MUX2_X1 U15282 ( .A(n13099), .B(n13098), .S(n15365), .Z(n13100) );
  OAI21_X1 U15283 ( .B1(n13101), .B2(n13110), .A(n13100), .ZN(P3_U3444) );
  INV_X1 U15284 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13103) );
  MUX2_X1 U15285 ( .A(n13103), .B(n13102), .S(n15365), .Z(n13104) );
  OAI21_X1 U15286 ( .B1(n13105), .B2(n13110), .A(n13104), .ZN(P3_U3441) );
  MUX2_X1 U15287 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13106), .S(n15365), .Z(
        P3_U3438) );
  INV_X1 U15288 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13108) );
  MUX2_X1 U15289 ( .A(n13108), .B(n13107), .S(n15365), .Z(n13109) );
  OAI21_X1 U15290 ( .B1(n13111), .B2(n13110), .A(n13109), .ZN(P3_U3435) );
  NAND2_X1 U15291 ( .A1(n13113), .A2(n13112), .ZN(n13118) );
  INV_X1 U15292 ( .A(n13114), .ZN(n13116) );
  NAND4_X1 U15293 ( .A1(n13116), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n13115), .ZN(n13117) );
  OAI211_X1 U15294 ( .C1(n13125), .C2(n13119), .A(n13118), .B(n13117), .ZN(
        P3_U3264) );
  INV_X1 U15295 ( .A(n13120), .ZN(n13122) );
  OAI222_X1 U15296 ( .A1(n13125), .A2(n13124), .B1(n13123), .B2(n13122), .C1(
        P3_U3151), .C2(n13121), .ZN(P3_U3266) );
  INV_X1 U15297 ( .A(n13126), .ZN(n13129) );
  OAI222_X1 U15298 ( .A1(n13130), .A2(n13129), .B1(n6501), .B2(P3_U3151), .C1(
        n13128), .C2(n13125), .ZN(P3_U3267) );
  AOI21_X1 U15299 ( .B1(n13131), .B2(n13132), .A(n14926), .ZN(n13134) );
  NAND2_X1 U15300 ( .A1(n13134), .A2(n13133), .ZN(n13141) );
  OAI22_X1 U15301 ( .A1(n13461), .A2(n14921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13135), .ZN(n13136) );
  AOI21_X1 U15302 ( .B1(n13430), .B2(n13235), .A(n13136), .ZN(n13137) );
  OAI21_X1 U15303 ( .B1(n13138), .B2(n14920), .A(n13137), .ZN(n13139) );
  AOI21_X1 U15304 ( .B1(n13656), .B2(n14930), .A(n13139), .ZN(n13140) );
  NAND2_X1 U15305 ( .A1(n13141), .A2(n13140), .ZN(P2_U3186) );
  INV_X1 U15306 ( .A(n13505), .ZN(n13745) );
  OAI21_X1 U15307 ( .B1(n13142), .B2(n13145), .A(n13144), .ZN(n13146) );
  NAND2_X1 U15308 ( .A1(n13146), .A2(n13243), .ZN(n13151) );
  OAI22_X1 U15309 ( .A1(n13460), .A2(n13537), .B1(n13536), .B2(n13539), .ZN(
        n13497) );
  INV_X1 U15310 ( .A(n13504), .ZN(n13148) );
  OAI22_X1 U15311 ( .A1(n13148), .A2(n14934), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13147), .ZN(n13149) );
  AOI21_X1 U15312 ( .B1(n13497), .B2(n13249), .A(n13149), .ZN(n13150) );
  OAI211_X1 U15313 ( .C1(n13745), .C2(n13252), .A(n13151), .B(n13150), .ZN(
        P2_U3188) );
  INV_X1 U15314 ( .A(n13154), .ZN(n13155) );
  AOI21_X1 U15315 ( .B1(n13156), .B2(n13152), .A(n13155), .ZN(n13160) );
  AOI22_X1 U15316 ( .A1(n13565), .A2(n13219), .B1(n13220), .B2(n13564), .ZN(
        n13157) );
  NAND2_X1 U15317 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13381)
         );
  OAI211_X1 U15318 ( .C1(n14934), .C2(n13568), .A(n13157), .B(n13381), .ZN(
        n13158) );
  AOI21_X1 U15319 ( .B1(n13702), .B2(n14930), .A(n13158), .ZN(n13159) );
  OAI21_X1 U15320 ( .B1(n13160), .B2(n14926), .A(n13159), .ZN(P2_U3191) );
  AOI21_X1 U15321 ( .B1(n13161), .B2(n13162), .A(n14926), .ZN(n13164) );
  NAND2_X1 U15322 ( .A1(n13164), .A2(n13163), .ZN(n13170) );
  INV_X1 U15323 ( .A(n13165), .ZN(n13542) );
  AOI22_X1 U15324 ( .A1(n13542), .A2(n13235), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13166) );
  OAI21_X1 U15325 ( .B1(n13538), .B2(n14921), .A(n13166), .ZN(n13167) );
  AOI21_X1 U15326 ( .B1(n13168), .B2(n13219), .A(n13167), .ZN(n13169) );
  OAI211_X1 U15327 ( .C1(n13755), .C2(n13252), .A(n13170), .B(n13169), .ZN(
        P2_U3195) );
  OAI211_X1 U15328 ( .C1(n13171), .C2(n13173), .A(n13172), .B(n13243), .ZN(
        n13178) );
  INV_X1 U15329 ( .A(n13461), .ZN(n13428) );
  INV_X1 U15330 ( .A(n13174), .ZN(n13470) );
  AOI22_X1 U15331 ( .A1(n13470), .A2(n13235), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13175) );
  OAI21_X1 U15332 ( .B1(n13460), .B2(n14921), .A(n13175), .ZN(n13176) );
  AOI21_X1 U15333 ( .B1(n13428), .B2(n13219), .A(n13176), .ZN(n13177) );
  OAI211_X1 U15334 ( .C1(n13179), .C2(n13252), .A(n13178), .B(n13177), .ZN(
        P2_U3197) );
  INV_X1 U15335 ( .A(n13712), .ZN(n13607) );
  INV_X1 U15336 ( .A(n13181), .ZN(n14639) );
  INV_X1 U15337 ( .A(n13182), .ZN(n13184) );
  NOR3_X1 U15338 ( .A1(n14639), .A2(n13184), .A3(n13183), .ZN(n13186) );
  OAI21_X1 U15339 ( .B1(n13186), .B2(n13185), .A(n13243), .ZN(n13191) );
  NAND2_X1 U15340 ( .A1(n13564), .A2(n13614), .ZN(n13188) );
  NAND2_X1 U15341 ( .A1(n13256), .A2(n13612), .ZN(n13187) );
  NAND2_X1 U15342 ( .A1(n13188), .A2(n13187), .ZN(n13595) );
  OAI22_X1 U15343 ( .A1(n14934), .A2(n13603), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15024), .ZN(n13189) );
  AOI21_X1 U15344 ( .B1(n13595), .B2(n13249), .A(n13189), .ZN(n13190) );
  OAI211_X1 U15345 ( .C1(n13607), .C2(n13252), .A(n13191), .B(n13190), .ZN(
        P2_U3200) );
  AOI21_X1 U15346 ( .B1(n13192), .B2(n13193), .A(n14926), .ZN(n13195) );
  NAND2_X1 U15347 ( .A1(n13195), .A2(n13194), .ZN(n13200) );
  INV_X1 U15348 ( .A(n13196), .ZN(n13488) );
  AOI22_X1 U15349 ( .A1(n13488), .A2(n13235), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13197) );
  OAI21_X1 U15350 ( .B1(n13483), .B2(n14921), .A(n13197), .ZN(n13198) );
  AOI21_X1 U15351 ( .B1(n13219), .B2(n13481), .A(n13198), .ZN(n13199) );
  OAI211_X1 U15352 ( .C1(n13490), .C2(n13252), .A(n13200), .B(n13199), .ZN(
        P2_U3201) );
  INV_X1 U15353 ( .A(n13203), .ZN(n13205) );
  NAND3_X1 U15354 ( .A1(n13154), .A2(n13205), .A3(n13204), .ZN(n13206) );
  AOI21_X1 U15355 ( .B1(n13201), .B2(n13206), .A(n14926), .ZN(n13210) );
  AOI22_X1 U15356 ( .A1(n13552), .A2(n13235), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13208) );
  AOI22_X1 U15357 ( .A1(n13558), .A2(n13219), .B1(n13220), .B2(n13579), .ZN(
        n13207) );
  OAI211_X1 U15358 ( .C1(n13554), .C2(n13252), .A(n13208), .B(n13207), .ZN(
        n13209) );
  OR2_X1 U15359 ( .A1(n13210), .A2(n13209), .ZN(P2_U3205) );
  OAI211_X1 U15360 ( .C1(n13213), .C2(n13212), .A(n13211), .B(n13243), .ZN(
        n13218) );
  OAI22_X1 U15361 ( .A1(n13514), .A2(n14921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13214), .ZN(n13216) );
  NOR2_X1 U15362 ( .A1(n13483), .A2(n14920), .ZN(n13215) );
  AOI211_X1 U15363 ( .C1(n13235), .C2(n13522), .A(n13216), .B(n13215), .ZN(
        n13217) );
  OAI211_X1 U15364 ( .C1(n13521), .C2(n13252), .A(n13218), .B(n13217), .ZN(
        P2_U3207) );
  AOI22_X1 U15365 ( .A1(n13220), .A2(n13615), .B1(n13219), .B2(n13579), .ZN(
        n13221) );
  NAND2_X1 U15366 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15046)
         );
  OAI211_X1 U15367 ( .C1(n14934), .C2(n13583), .A(n13221), .B(n15046), .ZN(
        n13228) );
  INV_X1 U15368 ( .A(n13224), .ZN(n13225) );
  AOI211_X1 U15369 ( .C1(n13707), .C2(n14930), .A(n13228), .B(n13227), .ZN(
        n13229) );
  INV_X1 U15370 ( .A(n13229), .ZN(P2_U3210) );
  AOI21_X1 U15372 ( .B1(n13233), .B2(n13230), .A(n15400), .ZN(n13240) );
  NOR2_X1 U15373 ( .A1(n13234), .A2(n14920), .ZN(n13238) );
  AOI22_X1 U15374 ( .A1(n13449), .A2(n13235), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13236) );
  OAI21_X1 U15375 ( .B1(n13443), .B2(n14921), .A(n13236), .ZN(n13237) );
  AOI211_X1 U15376 ( .C1(n13661), .C2(n14930), .A(n13238), .B(n13237), .ZN(
        n13239) );
  OAI21_X1 U15377 ( .B1(n13240), .B2(n14926), .A(n13239), .ZN(P2_U3212) );
  INV_X1 U15378 ( .A(n13721), .ZN(n13637) );
  OAI211_X1 U15379 ( .C1(n13245), .C2(n13244), .A(n13242), .B(n13243), .ZN(
        n13251) );
  OAI22_X1 U15380 ( .A1(n13247), .A2(n13539), .B1(n13246), .B2(n13537), .ZN(
        n13630) );
  NAND2_X1 U15381 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15019)
         );
  OAI21_X1 U15382 ( .B1(n14934), .B2(n13633), .A(n15019), .ZN(n13248) );
  AOI21_X1 U15383 ( .B1(n13630), .B2(n13249), .A(n13248), .ZN(n13250) );
  OAI211_X1 U15384 ( .C1(n13637), .C2(n13252), .A(n13251), .B(n13250), .ZN(
        P2_U3213) );
  MUX2_X1 U15385 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13388), .S(P2_U3947), .Z(
        P2_U3562) );
  MUX2_X1 U15386 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13253), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15387 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13254), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15388 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13427), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15389 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13441), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15390 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13428), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15391 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13481), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15392 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13255), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15393 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13512), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15394 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13558), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15395 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13565), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15396 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13579), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15397 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13564), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15398 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13615), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15399 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13256), .S(P2_U3947), .Z(
        P2_U3547) );
  MUX2_X1 U15400 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13613), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U15401 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13257), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U15402 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13258), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U15403 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13259), .S(P2_U3947), .Z(
        P2_U3543) );
  MUX2_X1 U15404 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13260), .S(P2_U3947), .Z(
        P2_U3542) );
  MUX2_X1 U15405 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13261), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U15406 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13262), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U15407 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13263), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15408 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13264), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15409 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13265), .S(P2_U3947), .Z(
        P2_U3537) );
  MUX2_X1 U15410 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13266), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U15411 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13267), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15412 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13268), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U15413 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n10668), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U15414 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13269), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U15415 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13270), .S(P2_U3947), .Z(
        P2_U3531) );
  NOR2_X1 U15416 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13271), .ZN(n13274) );
  NOR2_X1 U15417 ( .A1(n15048), .A2(n13272), .ZN(n13273) );
  AOI211_X1 U15418 ( .C1(n15051), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n13274), .B(
        n13273), .ZN(n13284) );
  OAI211_X1 U15419 ( .C1(n13277), .C2(n13276), .A(n15021), .B(n13275), .ZN(
        n13283) );
  INV_X1 U15420 ( .A(n13294), .ZN(n13281) );
  NAND3_X1 U15421 ( .A1(n14965), .A2(n13279), .A3(n13278), .ZN(n13280) );
  NAND3_X1 U15422 ( .A1(n15033), .A2(n13281), .A3(n13280), .ZN(n13282) );
  NAND3_X1 U15423 ( .A1(n13284), .A2(n13283), .A3(n13282), .ZN(P2_U3217) );
  INV_X1 U15424 ( .A(n13285), .ZN(n13288) );
  NOR2_X1 U15425 ( .A1(n15048), .A2(n13286), .ZN(n13287) );
  AOI211_X1 U15426 ( .C1(n15051), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n13288), .B(
        n13287), .ZN(n13298) );
  OAI211_X1 U15427 ( .C1(n13291), .C2(n13290), .A(n15021), .B(n13289), .ZN(
        n13297) );
  OR3_X1 U15428 ( .A1(n13294), .A2(n13293), .A3(n13292), .ZN(n13295) );
  NAND3_X1 U15429 ( .A1(n15033), .A2(n13309), .A3(n13295), .ZN(n13296) );
  NAND3_X1 U15430 ( .A1(n13298), .A2(n13297), .A3(n13296), .ZN(P2_U3218) );
  INV_X1 U15431 ( .A(n13299), .ZN(n13302) );
  NOR2_X1 U15432 ( .A1(n15048), .A2(n13300), .ZN(n13301) );
  AOI211_X1 U15433 ( .C1(n15051), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n13302), .B(
        n13301), .ZN(n13314) );
  OAI211_X1 U15434 ( .C1(n13305), .C2(n13304), .A(n15021), .B(n13303), .ZN(
        n13313) );
  INV_X1 U15435 ( .A(n13306), .ZN(n13311) );
  NAND3_X1 U15436 ( .A1(n13309), .A2(n13308), .A3(n13307), .ZN(n13310) );
  NAND3_X1 U15437 ( .A1(n15033), .A2(n13311), .A3(n13310), .ZN(n13312) );
  NAND3_X1 U15438 ( .A1(n13314), .A2(n13313), .A3(n13312), .ZN(P2_U3219) );
  NAND2_X1 U15439 ( .A1(n13315), .A2(n8985), .ZN(n14987) );
  MUX2_X1 U15440 ( .A(n13316), .B(P2_REG2_REG_12__SCAN_IN), .S(n14994), .Z(
        n14988) );
  AOI21_X1 U15441 ( .B1(n14989), .B2(n14987), .A(n14988), .ZN(n14986) );
  AOI21_X1 U15442 ( .B1(n13316), .B2(n13317), .A(n14986), .ZN(n13320) );
  AOI22_X1 U15443 ( .A1(n13343), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11911), 
        .B2(n13318), .ZN(n13319) );
  NAND2_X1 U15444 ( .A1(n13319), .A2(n13320), .ZN(n13333) );
  OAI211_X1 U15445 ( .C1(n13320), .C2(n13319), .A(n15033), .B(n13333), .ZN(
        n13332) );
  INV_X1 U15446 ( .A(n13321), .ZN(n13322) );
  AOI21_X1 U15447 ( .B1(n15051), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n13322), 
        .ZN(n13331) );
  NAND2_X1 U15448 ( .A1(n13323), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U15449 ( .A1(n13325), .A2(n13324), .ZN(n14983) );
  INV_X1 U15450 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14680) );
  MUX2_X1 U15451 ( .A(n14680), .B(P2_REG1_REG_12__SCAN_IN), .S(n14994), .Z(
        n14982) );
  OR2_X1 U15452 ( .A1(n14994), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n13326) );
  MUX2_X1 U15453 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9020), .S(n13343), .Z(
        n13327) );
  NAND2_X1 U15454 ( .A1(n13328), .A2(n13327), .ZN(n13345) );
  OAI211_X1 U15455 ( .C1(n13328), .C2(n13327), .A(n13345), .B(n15021), .ZN(
        n13330) );
  NAND2_X1 U15456 ( .A1(n15027), .A2(n13343), .ZN(n13329) );
  NAND4_X1 U15457 ( .A1(n13332), .A2(n13331), .A3(n13330), .A4(n13329), .ZN(
        P2_U3227) );
  NAND2_X1 U15458 ( .A1(n13343), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n13334) );
  NAND2_X1 U15459 ( .A1(n13334), .A2(n13333), .ZN(n13335) );
  NOR2_X1 U15460 ( .A1(n13335), .A2(n13349), .ZN(n13336) );
  NOR2_X1 U15461 ( .A1(n13336), .A2(n14998), .ZN(n13337) );
  NAND2_X1 U15462 ( .A1(n15016), .A2(n13337), .ZN(n13338) );
  XOR2_X1 U15463 ( .A(n15016), .B(n13337), .Z(n15015) );
  NAND2_X1 U15464 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15015), .ZN(n15014) );
  NAND2_X1 U15465 ( .A1(n13338), .A2(n15014), .ZN(n13341) );
  INV_X1 U15466 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13362) );
  NAND2_X1 U15467 ( .A1(n13368), .A2(n13362), .ZN(n13339) );
  OAI21_X1 U15468 ( .B1(n13368), .B2(n13362), .A(n13339), .ZN(n13340) );
  OAI211_X1 U15469 ( .C1(n13341), .C2(n13340), .A(n13360), .B(n15033), .ZN(
        n13359) );
  NAND2_X1 U15470 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14645)
         );
  INV_X1 U15471 ( .A(n14645), .ZN(n13342) );
  AOI21_X1 U15472 ( .B1(n15051), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n13342), 
        .ZN(n13358) );
  NAND2_X1 U15473 ( .A1(n13343), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n13344) );
  NAND2_X1 U15474 ( .A1(n13345), .A2(n13344), .ZN(n15001) );
  OR2_X1 U15475 ( .A1(n13349), .A2(n13346), .ZN(n13348) );
  NAND2_X1 U15476 ( .A1(n13349), .A2(n13346), .ZN(n13347) );
  NAND2_X1 U15477 ( .A1(n13348), .A2(n13347), .ZN(n15000) );
  AOI21_X1 U15478 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n13349), .A(n15002), 
        .ZN(n13351) );
  NOR2_X1 U15479 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  XNOR2_X1 U15480 ( .A(n13351), .B(n13350), .ZN(n15012) );
  NOR2_X1 U15481 ( .A1(n15011), .A2(n15012), .ZN(n15010) );
  NOR2_X1 U15482 ( .A1(n13352), .A2(n15010), .ZN(n13354) );
  XNOR2_X1 U15483 ( .A(n13368), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13353) );
  AOI21_X1 U15484 ( .B1(n13354), .B2(n13353), .A(n15042), .ZN(n13355) );
  NAND2_X1 U15485 ( .A1(n13355), .A2(n13370), .ZN(n13357) );
  NAND2_X1 U15486 ( .A1(n15027), .A2(n13368), .ZN(n13356) );
  NAND4_X1 U15487 ( .A1(n13359), .A2(n13358), .A3(n13357), .A4(n13356), .ZN(
        P2_U3230) );
  AOI22_X1 U15488 ( .A1(n15026), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9074), 
        .B2(n13363), .ZN(n15035) );
  NAND2_X1 U15489 ( .A1(n15035), .A2(n15034), .ZN(n15032) );
  XNOR2_X1 U15490 ( .A(n13364), .B(n13365), .ZN(n15041) );
  NOR2_X1 U15491 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15041), .ZN(n15040) );
  NOR2_X1 U15492 ( .A1(n13365), .A2(n13364), .ZN(n13366) );
  XOR2_X1 U15493 ( .A(n13367), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13378) );
  INV_X1 U15494 ( .A(n13378), .ZN(n13376) );
  NAND2_X1 U15495 ( .A1(n13368), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n13369) );
  NAND2_X1 U15496 ( .A1(n13370), .A2(n13369), .ZN(n15023) );
  XNOR2_X1 U15497 ( .A(n15026), .B(n13371), .ZN(n15022) );
  AOI21_X1 U15498 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n15026), .A(n15029), 
        .ZN(n13372) );
  XNOR2_X1 U15499 ( .A(n15047), .B(n13372), .ZN(n15045) );
  NOR2_X1 U15500 ( .A1(n15044), .A2(n15045), .ZN(n15043) );
  NOR2_X1 U15501 ( .A1(n13372), .A2(n15047), .ZN(n13373) );
  NOR2_X1 U15502 ( .A1(n15043), .A2(n13373), .ZN(n13374) );
  XNOR2_X1 U15503 ( .A(n13374), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13377) );
  NOR2_X1 U15504 ( .A1(n13377), .A2(n15042), .ZN(n13375) );
  AOI22_X1 U15505 ( .A1(n13378), .A2(n15033), .B1(n15021), .B2(n13377), .ZN(
        n13380) );
  OAI211_X1 U15506 ( .C1(n13383), .C2(n15039), .A(n13382), .B(n13381), .ZN(
        P2_U3233) );
  NAND2_X1 U15507 ( .A1(n13731), .A2(n13392), .ZN(n13391) );
  XNOR2_X1 U15508 ( .A(n13391), .B(n13728), .ZN(n13385) );
  NAND2_X1 U15509 ( .A1(n13385), .A2(n6483), .ZN(n13645) );
  INV_X1 U15510 ( .A(n13386), .ZN(n13387) );
  NAND2_X1 U15511 ( .A1(n13388), .A2(n13387), .ZN(n13648) );
  NOR2_X1 U15512 ( .A1(n13648), .A2(n14668), .ZN(n13394) );
  NOR2_X1 U15513 ( .A1(n13728), .A2(n13636), .ZN(n13389) );
  AOI211_X1 U15514 ( .C1(n14668), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13394), 
        .B(n13389), .ZN(n13390) );
  OAI21_X1 U15515 ( .B1(n13645), .B2(n13525), .A(n13390), .ZN(P2_U3234) );
  OAI211_X1 U15516 ( .C1(n13731), .C2(n13392), .A(n6483), .B(n13391), .ZN(
        n13649) );
  NOR2_X1 U15517 ( .A1(n7490), .A2(n13393), .ZN(n13395) );
  AOI211_X1 U15518 ( .C1(n13396), .C2(n14655), .A(n13395), .B(n13394), .ZN(
        n13397) );
  OAI21_X1 U15519 ( .B1(n13649), .B2(n13525), .A(n13397), .ZN(P2_U3235) );
  INV_X1 U15520 ( .A(n13398), .ZN(n13406) );
  INV_X1 U15521 ( .A(n13399), .ZN(n13400) );
  AOI22_X1 U15522 ( .A1(n13400), .A2(n14654), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14668), .ZN(n13403) );
  NAND2_X1 U15523 ( .A1(n13401), .A2(n14655), .ZN(n13402) );
  OAI211_X1 U15524 ( .C1(n13404), .C2(n13525), .A(n13403), .B(n13402), .ZN(
        n13405) );
  NAND3_X1 U15525 ( .A1(n13411), .A2(n9268), .A3(n13410), .ZN(n13414) );
  INV_X1 U15526 ( .A(n13412), .ZN(n13413) );
  INV_X1 U15527 ( .A(n13653), .ZN(n13424) );
  OAI211_X1 U15528 ( .C1(n9255), .C2(n13429), .A(n6483), .B(n13417), .ZN(
        n13651) );
  INV_X1 U15529 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13418) );
  OAI22_X1 U15530 ( .A1(n13420), .A2(n13419), .B1(n13418), .B2(n7490), .ZN(
        n13421) );
  AOI21_X1 U15531 ( .B1(n13733), .B2(n14655), .A(n13421), .ZN(n13422) );
  OAI21_X1 U15532 ( .B1(n13651), .B2(n13525), .A(n13422), .ZN(n13423) );
  AOI21_X1 U15533 ( .B1(n13424), .B2(n14665), .A(n13423), .ZN(n13425) );
  OAI21_X1 U15534 ( .B1(n13652), .B2(n14668), .A(n13425), .ZN(P2_U3237) );
  AOI211_X1 U15535 ( .C1(n13656), .C2(n13446), .A(n12562), .B(n13429), .ZN(
        n13655) );
  AOI22_X1 U15536 ( .A1(n13430), .A2(n14654), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14668), .ZN(n13431) );
  OAI21_X1 U15537 ( .B1(n13432), .B2(n13636), .A(n13431), .ZN(n13438) );
  NAND2_X1 U15538 ( .A1(n13434), .A2(n9190), .ZN(n13435) );
  NAND2_X1 U15539 ( .A1(n13436), .A2(n13435), .ZN(n13659) );
  NOR2_X1 U15540 ( .A1(n13659), .A2(n13641), .ZN(n13437) );
  AOI211_X1 U15541 ( .C1(n13655), .C2(n14664), .A(n13438), .B(n13437), .ZN(
        n13439) );
  OAI21_X1 U15542 ( .B1(n14668), .B2(n13657), .A(n13439), .ZN(P2_U3238) );
  XNOR2_X1 U15543 ( .A(n13440), .B(n13452), .ZN(n13445) );
  NAND2_X1 U15544 ( .A1(n13441), .A2(n13614), .ZN(n13442) );
  OAI21_X1 U15545 ( .B1(n13443), .B2(n13539), .A(n13442), .ZN(n13444) );
  AOI21_X1 U15546 ( .B1(n13445), .B2(n9268), .A(n13444), .ZN(n13662) );
  INV_X1 U15547 ( .A(n13469), .ZN(n13448) );
  INV_X1 U15548 ( .A(n13446), .ZN(n13447) );
  AOI211_X1 U15549 ( .C1(n13661), .C2(n13448), .A(n12562), .B(n13447), .ZN(
        n13660) );
  AOI22_X1 U15550 ( .A1(n13449), .A2(n14654), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14668), .ZN(n13450) );
  OAI21_X1 U15551 ( .B1(n13451), .B2(n13636), .A(n13450), .ZN(n13455) );
  XNOR2_X1 U15552 ( .A(n13453), .B(n13452), .ZN(n13664) );
  NOR2_X1 U15553 ( .A1(n13664), .A2(n13641), .ZN(n13454) );
  AOI211_X1 U15554 ( .C1(n13660), .C2(n14664), .A(n13455), .B(n13454), .ZN(
        n13456) );
  OAI21_X1 U15555 ( .B1(n14668), .B2(n13662), .A(n13456), .ZN(P2_U3239) );
  OAI21_X1 U15556 ( .B1(n13459), .B2(n13458), .A(n13457), .ZN(n13463) );
  OAI22_X1 U15557 ( .A1(n13461), .A2(n13537), .B1(n13460), .B2(n13539), .ZN(
        n13462) );
  AOI21_X1 U15558 ( .B1(n13463), .B2(n9268), .A(n13462), .ZN(n13667) );
  OAI21_X1 U15559 ( .B1(n13466), .B2(n13465), .A(n13464), .ZN(n13665) );
  NAND2_X1 U15560 ( .A1(n13739), .A2(n13487), .ZN(n13467) );
  NAND2_X1 U15561 ( .A1(n13467), .A2(n6483), .ZN(n13468) );
  OR2_X1 U15562 ( .A1(n13469), .A2(n13468), .ZN(n13666) );
  AOI22_X1 U15563 ( .A1(n13470), .A2(n14654), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14668), .ZN(n13472) );
  NAND2_X1 U15564 ( .A1(n13739), .A2(n14655), .ZN(n13471) );
  OAI211_X1 U15565 ( .C1(n13666), .C2(n13525), .A(n13472), .B(n13471), .ZN(
        n13473) );
  AOI21_X1 U15566 ( .B1(n13665), .B2(n14665), .A(n13473), .ZN(n13474) );
  OAI21_X1 U15567 ( .B1(n14668), .B2(n13667), .A(n13474), .ZN(P2_U3240) );
  OAI21_X1 U15568 ( .B1(n13476), .B2(n13478), .A(n13475), .ZN(n13674) );
  NAND2_X1 U15569 ( .A1(n13478), .A2(n13477), .ZN(n13479) );
  NAND2_X1 U15570 ( .A1(n13480), .A2(n13479), .ZN(n13485) );
  NAND2_X1 U15571 ( .A1(n13481), .A2(n13614), .ZN(n13482) );
  OAI21_X1 U15572 ( .B1(n13483), .B2(n13539), .A(n13482), .ZN(n13484) );
  AOI21_X1 U15573 ( .B1(n13485), .B2(n9268), .A(n13484), .ZN(n13486) );
  OAI21_X1 U15574 ( .B1(n13674), .B2(n9219), .A(n13486), .ZN(n13676) );
  NAND2_X1 U15575 ( .A1(n13676), .A2(n7490), .ZN(n13494) );
  OAI211_X1 U15576 ( .C1(n13490), .C2(n13503), .A(n6483), .B(n13487), .ZN(
        n13672) );
  INV_X1 U15577 ( .A(n13672), .ZN(n13492) );
  AOI22_X1 U15578 ( .A1(n13488), .A2(n14654), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14668), .ZN(n13489) );
  OAI21_X1 U15579 ( .B1(n13490), .B2(n13636), .A(n13489), .ZN(n13491) );
  AOI21_X1 U15580 ( .B1(n13492), .B2(n14664), .A(n13491), .ZN(n13493) );
  OAI211_X1 U15581 ( .C1(n13674), .C2(n13495), .A(n13494), .B(n13493), .ZN(
        P2_U3241) );
  XNOR2_X1 U15582 ( .A(n6538), .B(n13496), .ZN(n13498) );
  AOI21_X1 U15583 ( .B1(n13498), .B2(n9268), .A(n13497), .ZN(n13679) );
  XNOR2_X1 U15584 ( .A(n13500), .B(n13499), .ZN(n13677) );
  NAND2_X1 U15585 ( .A1(n13505), .A2(n13520), .ZN(n13501) );
  NAND2_X1 U15586 ( .A1(n13501), .A2(n6483), .ZN(n13502) );
  OR2_X1 U15587 ( .A1(n13503), .A2(n13502), .ZN(n13678) );
  AOI22_X1 U15588 ( .A1(n13504), .A2(n14654), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14668), .ZN(n13507) );
  NAND2_X1 U15589 ( .A1(n13505), .A2(n14655), .ZN(n13506) );
  OAI211_X1 U15590 ( .C1(n13678), .C2(n13525), .A(n13507), .B(n13506), .ZN(
        n13508) );
  AOI21_X1 U15591 ( .B1(n13677), .B2(n14665), .A(n13508), .ZN(n13509) );
  OAI21_X1 U15592 ( .B1(n14668), .B2(n13679), .A(n13509), .ZN(P2_U3242) );
  XNOR2_X1 U15593 ( .A(n13511), .B(n13510), .ZN(n13516) );
  NAND2_X1 U15594 ( .A1(n13512), .A2(n13614), .ZN(n13513) );
  OAI21_X1 U15595 ( .B1(n13514), .B2(n13539), .A(n13513), .ZN(n13515) );
  AOI21_X1 U15596 ( .B1(n13516), .B2(n9268), .A(n13515), .ZN(n13685) );
  OAI21_X1 U15597 ( .B1(n13519), .B2(n13518), .A(n13517), .ZN(n13683) );
  INV_X1 U15598 ( .A(n13683), .ZN(n13527) );
  OAI211_X1 U15599 ( .C1(n13521), .C2(n13540), .A(n6483), .B(n13520), .ZN(
        n13684) );
  AOI22_X1 U15600 ( .A1(n13522), .A2(n14654), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n14668), .ZN(n13524) );
  NAND2_X1 U15601 ( .A1(n13748), .A2(n14655), .ZN(n13523) );
  OAI211_X1 U15602 ( .C1(n13684), .C2(n13525), .A(n13524), .B(n13523), .ZN(
        n13526) );
  AOI21_X1 U15603 ( .B1(n13527), .B2(n14665), .A(n13526), .ZN(n13528) );
  OAI21_X1 U15604 ( .B1(n14668), .B2(n13685), .A(n13528), .ZN(P2_U3243) );
  XNOR2_X1 U15605 ( .A(n13529), .B(n13534), .ZN(n13692) );
  INV_X1 U15606 ( .A(n13692), .ZN(n13547) );
  AOI21_X1 U15607 ( .B1(n13563), .B2(n13531), .A(n13530), .ZN(n13556) );
  INV_X1 U15608 ( .A(n13548), .ZN(n13557) );
  NAND2_X1 U15609 ( .A1(n13556), .A2(n13557), .ZN(n13555) );
  NAND2_X1 U15610 ( .A1(n13555), .A2(n13532), .ZN(n13533) );
  XOR2_X1 U15611 ( .A(n13534), .B(n13533), .Z(n13535) );
  OAI222_X1 U15612 ( .A1(n13539), .A2(n13538), .B1(n13537), .B2(n13536), .C1(
        n13593), .C2(n13535), .ZN(n13690) );
  AOI211_X1 U15613 ( .C1(n13541), .C2(n13550), .A(n12562), .B(n13540), .ZN(
        n13691) );
  NAND2_X1 U15614 ( .A1(n13691), .A2(n14664), .ZN(n13544) );
  AOI22_X1 U15615 ( .A1(n13542), .A2(n14654), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14668), .ZN(n13543) );
  OAI211_X1 U15616 ( .C1(n13755), .C2(n13636), .A(n13544), .B(n13543), .ZN(
        n13545) );
  AOI21_X1 U15617 ( .B1(n13690), .B2(n7490), .A(n13545), .ZN(n13546) );
  OAI21_X1 U15618 ( .B1(n13547), .B2(n13641), .A(n13546), .ZN(P2_U3244) );
  XNOR2_X1 U15619 ( .A(n13549), .B(n13548), .ZN(n13700) );
  INV_X1 U15620 ( .A(n13550), .ZN(n13551) );
  AOI211_X1 U15621 ( .C1(n13697), .C2(n13567), .A(n12562), .B(n13551), .ZN(
        n13696) );
  AOI22_X1 U15622 ( .A1(n13552), .A2(n14654), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n14668), .ZN(n13553) );
  OAI21_X1 U15623 ( .B1(n13554), .B2(n13636), .A(n13553), .ZN(n13561) );
  OAI21_X1 U15624 ( .B1(n13557), .B2(n13556), .A(n13555), .ZN(n13559) );
  AOI222_X1 U15625 ( .A1(n9268), .A2(n13559), .B1(n13558), .B2(n13614), .C1(
        n13579), .C2(n13612), .ZN(n13699) );
  NOR2_X1 U15626 ( .A1(n13699), .A2(n14668), .ZN(n13560) );
  AOI211_X1 U15627 ( .C1(n13696), .C2(n14664), .A(n13561), .B(n13560), .ZN(
        n13562) );
  OAI21_X1 U15628 ( .B1(n13641), .B2(n13700), .A(n13562), .ZN(P2_U3245) );
  XOR2_X1 U15629 ( .A(n13572), .B(n13563), .Z(n13566) );
  AOI222_X1 U15630 ( .A1(n9268), .A2(n13566), .B1(n13565), .B2(n13614), .C1(
        n13564), .C2(n13612), .ZN(n13704) );
  AOI211_X1 U15631 ( .C1(n13702), .C2(n13581), .A(n12562), .B(n6933), .ZN(
        n13701) );
  INV_X1 U15632 ( .A(n13568), .ZN(n13569) );
  AOI22_X1 U15633 ( .A1(n13569), .A2(n14654), .B1(n14668), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n13570) );
  OAI21_X1 U15634 ( .B1(n13571), .B2(n13636), .A(n13570), .ZN(n13575) );
  XNOR2_X1 U15635 ( .A(n13573), .B(n13572), .ZN(n13705) );
  NOR2_X1 U15636 ( .A1(n13705), .A2(n13641), .ZN(n13574) );
  AOI211_X1 U15637 ( .C1(n13701), .C2(n14664), .A(n13575), .B(n13574), .ZN(
        n13576) );
  OAI21_X1 U15638 ( .B1(n14668), .B2(n13704), .A(n13576), .ZN(P2_U3246) );
  XNOR2_X1 U15639 ( .A(n13578), .B(n13577), .ZN(n13580) );
  AOI222_X1 U15640 ( .A1(n9268), .A2(n13580), .B1(n13579), .B2(n13614), .C1(
        n13615), .C2(n13612), .ZN(n13709) );
  INV_X1 U15641 ( .A(n13581), .ZN(n13582) );
  AOI211_X1 U15642 ( .C1(n13707), .C2(n13601), .A(n12562), .B(n13582), .ZN(
        n13706) );
  INV_X1 U15643 ( .A(n13583), .ZN(n13584) );
  AOI22_X1 U15644 ( .A1(n14668), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14654), 
        .B2(n13584), .ZN(n13585) );
  OAI21_X1 U15645 ( .B1(n6934), .B2(n13636), .A(n13585), .ZN(n13591) );
  INV_X1 U15646 ( .A(n13586), .ZN(n13587) );
  AOI21_X1 U15647 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(n13710) );
  NOR2_X1 U15648 ( .A1(n13710), .A2(n13641), .ZN(n13590) );
  AOI211_X1 U15649 ( .C1(n13706), .C2(n14664), .A(n13591), .B(n13590), .ZN(
        n13592) );
  OAI21_X1 U15650 ( .B1(n14668), .B2(n13709), .A(n13592), .ZN(P2_U3247) );
  AOI21_X1 U15651 ( .B1(n13594), .B2(n13599), .A(n13593), .ZN(n13597) );
  AOI21_X1 U15652 ( .B1(n13597), .B2(n13596), .A(n13595), .ZN(n13714) );
  OAI21_X1 U15653 ( .B1(n13600), .B2(n13599), .A(n13598), .ZN(n13715) );
  INV_X1 U15654 ( .A(n13715), .ZN(n13609) );
  AOI21_X1 U15655 ( .B1(n13621), .B2(n13712), .A(n12562), .ZN(n13602) );
  AND2_X1 U15656 ( .A1(n13602), .A2(n13601), .ZN(n13711) );
  NAND2_X1 U15657 ( .A1(n13711), .A2(n14664), .ZN(n13606) );
  INV_X1 U15658 ( .A(n13603), .ZN(n13604) );
  AOI22_X1 U15659 ( .A1(n14668), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14654), 
        .B2(n13604), .ZN(n13605) );
  OAI211_X1 U15660 ( .C1(n13607), .C2(n13636), .A(n13606), .B(n13605), .ZN(
        n13608) );
  AOI21_X1 U15661 ( .B1(n13609), .B2(n14665), .A(n13608), .ZN(n13610) );
  OAI21_X1 U15662 ( .B1(n14668), .B2(n13714), .A(n13610), .ZN(P2_U3248) );
  XNOR2_X1 U15663 ( .A(n13611), .B(n13618), .ZN(n13616) );
  AOI222_X1 U15664 ( .A1(n9268), .A2(n13616), .B1(n13615), .B2(n13614), .C1(
        n13613), .C2(n13612), .ZN(n13718) );
  OAI21_X1 U15665 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n13719) );
  INV_X1 U15666 ( .A(n13719), .ZN(n13627) );
  OR2_X1 U15667 ( .A1(n13625), .A2(n13632), .ZN(n13620) );
  AND3_X1 U15668 ( .A1(n13621), .A2(n13620), .A3(n6483), .ZN(n13716) );
  NAND2_X1 U15669 ( .A1(n13716), .A2(n14664), .ZN(n13624) );
  INV_X1 U15670 ( .A(n14647), .ZN(n13622) );
  AOI22_X1 U15671 ( .A1(n14668), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n14654), 
        .B2(n13622), .ZN(n13623) );
  OAI211_X1 U15672 ( .C1(n13625), .C2(n13636), .A(n13624), .B(n13623), .ZN(
        n13626) );
  AOI21_X1 U15673 ( .B1(n13627), .B2(n14665), .A(n13626), .ZN(n13628) );
  OAI21_X1 U15674 ( .B1(n13718), .B2(n14668), .A(n13628), .ZN(P2_U3249) );
  XNOR2_X1 U15675 ( .A(n13629), .B(n7152), .ZN(n13631) );
  AOI21_X1 U15676 ( .B1(n13631), .B2(n9268), .A(n13630), .ZN(n13723) );
  AOI211_X1 U15677 ( .C1(n13721), .C2(n14661), .A(n12562), .B(n13632), .ZN(
        n13720) );
  INV_X1 U15678 ( .A(n13633), .ZN(n13634) );
  AOI22_X1 U15679 ( .A1(n14668), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14654), 
        .B2(n13634), .ZN(n13635) );
  OAI21_X1 U15680 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13643) );
  INV_X1 U15681 ( .A(n13638), .ZN(n13639) );
  AOI21_X1 U15682 ( .B1(n7152), .B2(n13640), .A(n13639), .ZN(n13725) );
  NOR2_X1 U15683 ( .A1(n13725), .A2(n13641), .ZN(n13642) );
  AOI211_X1 U15684 ( .C1(n13720), .C2(n14664), .A(n13643), .B(n13642), .ZN(
        n13644) );
  OAI21_X1 U15685 ( .B1(n14668), .B2(n13723), .A(n13644), .ZN(P2_U3250) );
  INV_X1 U15686 ( .A(n13688), .ZN(n13695) );
  OAI21_X1 U15687 ( .B1(n13728), .B2(n13695), .A(n13647), .ZN(P2_U3530) );
  AND2_X1 U15688 ( .A1(n13649), .A2(n13648), .ZN(n13729) );
  INV_X1 U15689 ( .A(n13654), .ZN(P2_U3527) );
  AOI21_X1 U15690 ( .B1(n15100), .B2(n13656), .A(n13655), .ZN(n13658) );
  OAI211_X1 U15691 ( .C1(n13724), .C2(n13659), .A(n13658), .B(n13657), .ZN(
        n13735) );
  MUX2_X1 U15692 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13735), .S(n15156), .Z(
        P2_U3526) );
  AOI21_X1 U15693 ( .B1(n15100), .B2(n13661), .A(n13660), .ZN(n13663) );
  OAI211_X1 U15694 ( .C1(n13724), .C2(n13664), .A(n13663), .B(n13662), .ZN(
        n13736) );
  MUX2_X1 U15695 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13736), .S(n15156), .Z(
        P2_U3525) );
  NAND2_X1 U15696 ( .A1(n13665), .A2(n15137), .ZN(n13668) );
  NAND3_X1 U15697 ( .A1(n13668), .A2(n13667), .A3(n13666), .ZN(n13737) );
  MUX2_X1 U15698 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13737), .S(n15156), .Z(
        n13669) );
  AOI21_X1 U15699 ( .B1(n13688), .B2(n13739), .A(n13669), .ZN(n13670) );
  INV_X1 U15700 ( .A(n13670), .ZN(P2_U3524) );
  NAND2_X1 U15701 ( .A1(n13671), .A2(n15100), .ZN(n13673) );
  OAI211_X1 U15702 ( .C1(n13674), .C2(n15123), .A(n13673), .B(n13672), .ZN(
        n13675) );
  OR2_X1 U15703 ( .A1(n13676), .A2(n13675), .ZN(n13741) );
  MUX2_X1 U15704 ( .A(n13741), .B(P2_REG1_REG_24__SCAN_IN), .S(n15154), .Z(
        P2_U3523) );
  NAND2_X1 U15705 ( .A1(n13677), .A2(n15137), .ZN(n13680) );
  AND3_X1 U15706 ( .A1(n13680), .A2(n13679), .A3(n13678), .ZN(n13742) );
  MUX2_X1 U15707 ( .A(n13681), .B(n13742), .S(n15156), .Z(n13682) );
  OAI21_X1 U15708 ( .B1(n13745), .B2(n13695), .A(n13682), .ZN(P2_U3522) );
  OR2_X1 U15709 ( .A1(n13683), .A2(n13724), .ZN(n13686) );
  NAND3_X1 U15710 ( .A1(n13686), .A2(n13685), .A3(n13684), .ZN(n13746) );
  MUX2_X1 U15711 ( .A(n13746), .B(P2_REG1_REG_22__SCAN_IN), .S(n15154), .Z(
        n13687) );
  AOI21_X1 U15712 ( .B1(n13688), .B2(n13748), .A(n13687), .ZN(n13689) );
  INV_X1 U15713 ( .A(n13689), .ZN(P2_U3521) );
  AOI211_X1 U15714 ( .C1(n15137), .C2(n13692), .A(n13691), .B(n13690), .ZN(
        n13751) );
  MUX2_X1 U15715 ( .A(n13693), .B(n13751), .S(n15156), .Z(n13694) );
  OAI21_X1 U15716 ( .B1(n13755), .B2(n13695), .A(n13694), .ZN(P2_U3520) );
  AOI21_X1 U15717 ( .B1(n15100), .B2(n13697), .A(n13696), .ZN(n13698) );
  OAI211_X1 U15718 ( .C1(n13724), .C2(n13700), .A(n13699), .B(n13698), .ZN(
        n13756) );
  MUX2_X1 U15719 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13756), .S(n15156), .Z(
        P2_U3519) );
  AOI21_X1 U15720 ( .B1(n15100), .B2(n13702), .A(n13701), .ZN(n13703) );
  OAI211_X1 U15721 ( .C1(n13724), .C2(n13705), .A(n13704), .B(n13703), .ZN(
        n13757) );
  MUX2_X1 U15722 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13757), .S(n15156), .Z(
        P2_U3518) );
  AOI21_X1 U15723 ( .B1(n15100), .B2(n13707), .A(n13706), .ZN(n13708) );
  OAI211_X1 U15724 ( .C1(n13710), .C2(n13724), .A(n13709), .B(n13708), .ZN(
        n13758) );
  MUX2_X1 U15725 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13758), .S(n15156), .Z(
        P2_U3517) );
  AOI21_X1 U15726 ( .B1(n15100), .B2(n13712), .A(n13711), .ZN(n13713) );
  OAI211_X1 U15727 ( .C1(n13715), .C2(n13724), .A(n13714), .B(n13713), .ZN(
        n13759) );
  MUX2_X1 U15728 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13759), .S(n15156), .Z(
        P2_U3516) );
  AOI21_X1 U15729 ( .B1(n15100), .B2(n14644), .A(n13716), .ZN(n13717) );
  OAI211_X1 U15730 ( .C1(n13724), .C2(n13719), .A(n13718), .B(n13717), .ZN(
        n13760) );
  MUX2_X1 U15731 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13760), .S(n15156), .Z(
        P2_U3515) );
  AOI21_X1 U15732 ( .B1(n15100), .B2(n13721), .A(n13720), .ZN(n13722) );
  OAI211_X1 U15733 ( .C1(n13725), .C2(n13724), .A(n13723), .B(n13722), .ZN(
        n13761) );
  MUX2_X1 U15734 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13761), .S(n15156), .Z(
        P2_U3514) );
  OAI21_X1 U15735 ( .B1(n13728), .B2(n13754), .A(n13727), .ZN(P2_U3498) );
  INV_X1 U15736 ( .A(n13734), .ZN(P2_U3495) );
  MUX2_X1 U15737 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13735), .S(n15147), .Z(
        P2_U3494) );
  MUX2_X1 U15738 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13736), .S(n15147), .Z(
        P2_U3493) );
  MUX2_X1 U15739 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13737), .S(n15147), .Z(
        n13738) );
  AOI21_X1 U15740 ( .B1(n13749), .B2(n13739), .A(n13738), .ZN(n13740) );
  INV_X1 U15741 ( .A(n13740), .ZN(P2_U3492) );
  MUX2_X1 U15742 ( .A(n13741), .B(P2_REG0_REG_24__SCAN_IN), .S(n15145), .Z(
        P2_U3491) );
  INV_X1 U15743 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13743) );
  MUX2_X1 U15744 ( .A(n13743), .B(n13742), .S(n15147), .Z(n13744) );
  OAI21_X1 U15745 ( .B1(n13745), .B2(n13754), .A(n13744), .ZN(P2_U3490) );
  MUX2_X1 U15746 ( .A(n13746), .B(P2_REG0_REG_22__SCAN_IN), .S(n15145), .Z(
        n13747) );
  AOI21_X1 U15747 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13750) );
  INV_X1 U15748 ( .A(n13750), .ZN(P2_U3489) );
  INV_X1 U15749 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13752) );
  MUX2_X1 U15750 ( .A(n13752), .B(n13751), .S(n15147), .Z(n13753) );
  OAI21_X1 U15751 ( .B1(n13755), .B2(n13754), .A(n13753), .ZN(P2_U3488) );
  MUX2_X1 U15752 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13756), .S(n15147), .Z(
        P2_U3487) );
  MUX2_X1 U15753 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13757), .S(n15147), .Z(
        P2_U3486) );
  MUX2_X1 U15754 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13758), .S(n15147), .Z(
        P2_U3484) );
  MUX2_X1 U15755 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13759), .S(n15147), .Z(
        P2_U3481) );
  MUX2_X1 U15756 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13760), .S(n15147), .Z(
        P2_U3478) );
  MUX2_X1 U15757 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13761), .S(n15147), .Z(
        P2_U3475) );
  INV_X1 U15758 ( .A(n13762), .ZN(n14511) );
  NOR4_X1 U15759 ( .A1(n13763), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8741), .A4(
        P2_U3088), .ZN(n13764) );
  AOI21_X1 U15760 ( .B1(n13770), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13764), 
        .ZN(n13765) );
  OAI21_X1 U15761 ( .B1(n14511), .B2(n13781), .A(n13765), .ZN(P2_U3296) );
  INV_X1 U15762 ( .A(n13766), .ZN(n14512) );
  OAI222_X1 U15763 ( .A1(n13781), .A2(n14512), .B1(P2_U3088), .B2(n13768), 
        .C1(n13767), .C2(n13783), .ZN(P2_U3298) );
  AOI21_X1 U15764 ( .B1(n13770), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13769), 
        .ZN(n13771) );
  OAI21_X1 U15765 ( .B1(n13772), .B2(n13781), .A(n13771), .ZN(P2_U3299) );
  INV_X1 U15766 ( .A(n13773), .ZN(n14517) );
  OAI222_X1 U15767 ( .A1(n13783), .A2(n13775), .B1(n13781), .B2(n14517), .C1(
        n13774), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15768 ( .A(n13776), .ZN(n14520) );
  OAI222_X1 U15769 ( .A1(P2_U3088), .A2(n13778), .B1(n13781), .B2(n14520), 
        .C1(n13777), .C2(n13783), .ZN(P2_U3301) );
  INV_X1 U15770 ( .A(n13779), .ZN(n14524) );
  OAI222_X1 U15771 ( .A1(n13783), .A2(n13782), .B1(n13781), .B2(n14524), .C1(
        P2_U3088), .C2(n13780), .ZN(P2_U3302) );
  MUX2_X1 U15772 ( .A(n13784), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U15773 ( .A1(n14205), .A2(n11847), .B1(n13932), .B2(n14069), .ZN(
        n13928) );
  NAND2_X1 U15774 ( .A1(n14205), .A2(n13935), .ZN(n13786) );
  NAND2_X1 U15775 ( .A1(n14069), .A2(n11847), .ZN(n13785) );
  NAND2_X1 U15776 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  XOR2_X1 U15777 ( .A(n13928), .B(n13929), .Z(n13930) );
  INV_X1 U15778 ( .A(n13788), .ZN(n13791) );
  NAND2_X1 U15779 ( .A1(n13793), .A2(n13792), .ZN(n14017) );
  NOR2_X1 U15780 ( .A1(n13854), .A2(n13794), .ZN(n13795) );
  AOI21_X1 U15781 ( .B1(n14710), .B2(n13933), .A(n13795), .ZN(n13798) );
  AOI22_X1 U15782 ( .A1(n14710), .A2(n13935), .B1(n13933), .B2(n14075), .ZN(
        n13796) );
  XNOR2_X1 U15783 ( .A(n13796), .B(n12151), .ZN(n13797) );
  XOR2_X1 U15784 ( .A(n13798), .B(n13797), .Z(n14016) );
  NAND2_X1 U15785 ( .A1(n14017), .A2(n14016), .ZN(n13802) );
  INV_X1 U15786 ( .A(n13797), .ZN(n13800) );
  INV_X1 U15787 ( .A(n13798), .ZN(n13799) );
  NAND2_X1 U15788 ( .A1(n13800), .A2(n13799), .ZN(n13801) );
  NAND2_X1 U15789 ( .A1(n13802), .A2(n13801), .ZN(n14684) );
  INV_X1 U15790 ( .A(n14684), .ZN(n13810) );
  NAND2_X1 U15791 ( .A1(n14688), .A2(n13935), .ZN(n13804) );
  NAND2_X1 U15792 ( .A1(n14074), .A2(n13933), .ZN(n13803) );
  NAND2_X1 U15793 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  XNOR2_X1 U15794 ( .A(n13805), .B(n7488), .ZN(n13808) );
  NOR2_X1 U15795 ( .A1(n13854), .A2(n14058), .ZN(n13806) );
  AOI21_X1 U15796 ( .B1(n14688), .B2(n13933), .A(n13806), .ZN(n13807) );
  NAND2_X1 U15797 ( .A1(n13808), .A2(n13807), .ZN(n13811) );
  OAI21_X1 U15798 ( .B1(n13808), .B2(n13807), .A(n13811), .ZN(n14683) );
  INV_X1 U15799 ( .A(n14683), .ZN(n13809) );
  OAI22_X1 U15800 ( .A1(n14697), .A2(n13838), .B1(n13977), .B2(n13855), .ZN(
        n13813) );
  XOR2_X1 U15801 ( .A(n12151), .B(n13813), .Z(n13814) );
  OAI22_X1 U15802 ( .A1(n14697), .A2(n13855), .B1(n13977), .B2(n13854), .ZN(
        n14054) );
  NAND2_X1 U15803 ( .A1(n14480), .A2(n13935), .ZN(n13816) );
  NAND2_X1 U15804 ( .A1(n14365), .A2(n13933), .ZN(n13815) );
  NAND2_X1 U15805 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  XNOR2_X1 U15806 ( .A(n13817), .B(n12151), .ZN(n13818) );
  AOI22_X1 U15807 ( .A1(n14480), .A2(n13933), .B1(n13932), .B2(n14365), .ZN(
        n13819) );
  XNOR2_X1 U15808 ( .A(n13818), .B(n13819), .ZN(n13975) );
  NAND2_X1 U15809 ( .A1(n13974), .A2(n13975), .ZN(n13973) );
  INV_X1 U15810 ( .A(n13818), .ZN(n13820) );
  NAND2_X1 U15811 ( .A1(n13820), .A2(n13819), .ZN(n13821) );
  NAND2_X1 U15812 ( .A1(n13973), .A2(n13821), .ZN(n13986) );
  NAND2_X1 U15813 ( .A1(n14475), .A2(n13935), .ZN(n13823) );
  NAND2_X1 U15814 ( .A1(n14072), .A2(n13933), .ZN(n13822) );
  NAND2_X1 U15815 ( .A1(n13823), .A2(n13822), .ZN(n13824) );
  XNOR2_X1 U15816 ( .A(n13824), .B(n12151), .ZN(n13827) );
  NAND2_X1 U15817 ( .A1(n14475), .A2(n11847), .ZN(n13826) );
  NAND2_X1 U15818 ( .A1(n13932), .A2(n14072), .ZN(n13825) );
  NAND2_X1 U15819 ( .A1(n13826), .A2(n13825), .ZN(n13828) );
  NAND2_X1 U15820 ( .A1(n13827), .A2(n13828), .ZN(n13988) );
  NAND2_X1 U15821 ( .A1(n13986), .A2(n13988), .ZN(n13985) );
  INV_X1 U15822 ( .A(n13827), .ZN(n13830) );
  INV_X1 U15823 ( .A(n13828), .ZN(n13829) );
  NAND2_X1 U15824 ( .A1(n13830), .A2(n13829), .ZN(n13987) );
  NAND2_X1 U15825 ( .A1(n13985), .A2(n13987), .ZN(n14037) );
  NOR2_X1 U15826 ( .A1(n13833), .A2(n13855), .ZN(n13831) );
  AOI21_X1 U15827 ( .B1(n14470), .B2(n13935), .A(n13831), .ZN(n13832) );
  XNOR2_X1 U15828 ( .A(n13832), .B(n12151), .ZN(n13836) );
  INV_X1 U15829 ( .A(n14470), .ZN(n14347) );
  OAI22_X1 U15830 ( .A1(n14347), .A2(n13855), .B1(n13833), .B2(n13854), .ZN(
        n13834) );
  XNOR2_X1 U15831 ( .A(n13836), .B(n13834), .ZN(n14038) );
  INV_X1 U15832 ( .A(n13834), .ZN(n13835) );
  NAND2_X1 U15833 ( .A1(n13836), .A2(n13835), .ZN(n13837) );
  OAI22_X1 U15834 ( .A1(n14335), .A2(n13838), .B1(n14352), .B2(n13855), .ZN(
        n13839) );
  XNOR2_X1 U15835 ( .A(n13839), .B(n12151), .ZN(n13841) );
  OAI22_X1 U15836 ( .A1(n14335), .A2(n13855), .B1(n14352), .B2(n13854), .ZN(
        n13840) );
  XNOR2_X1 U15837 ( .A(n13841), .B(n13840), .ZN(n13921) );
  NAND2_X1 U15838 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  NAND2_X1 U15839 ( .A1(n13923), .A2(n13842), .ZN(n14009) );
  NOR2_X1 U15840 ( .A1(n13843), .A2(n13854), .ZN(n13844) );
  AOI21_X1 U15841 ( .B1(n14455), .B2(n13933), .A(n13844), .ZN(n13846) );
  AOI22_X1 U15842 ( .A1(n14455), .A2(n13935), .B1(n11847), .B2(n14292), .ZN(
        n13845) );
  XNOR2_X1 U15843 ( .A(n13845), .B(n12151), .ZN(n13847) );
  XOR2_X1 U15844 ( .A(n13846), .B(n13847), .Z(n14008) );
  OR2_X1 U15845 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  AOI22_X1 U15846 ( .A1(n14449), .A2(n13935), .B1(n11847), .B2(n14285), .ZN(
        n13849) );
  XNOR2_X1 U15847 ( .A(n13849), .B(n12151), .ZN(n13852) );
  AOI22_X1 U15848 ( .A1(n14449), .A2(n13933), .B1(n13932), .B2(n14285), .ZN(
        n13851) );
  XNOR2_X1 U15849 ( .A(n13852), .B(n13851), .ZN(n13952) );
  NAND2_X1 U15850 ( .A1(n13852), .A2(n13851), .ZN(n13853) );
  NAND2_X2 U15851 ( .A1(n13949), .A2(n13853), .ZN(n13960) );
  OAI22_X1 U15852 ( .A1(n14281), .A2(n13855), .B1(n13954), .B2(n13854), .ZN(
        n13883) );
  NAND2_X1 U15853 ( .A1(n14444), .A2(n13935), .ZN(n13857) );
  NAND2_X1 U15854 ( .A1(n14293), .A2(n13933), .ZN(n13856) );
  NAND2_X1 U15855 ( .A1(n13857), .A2(n13856), .ZN(n13858) );
  XNOR2_X1 U15856 ( .A(n13858), .B(n12151), .ZN(n13882) );
  XOR2_X1 U15857 ( .A(n13883), .B(n13882), .Z(n14026) );
  NAND2_X1 U15858 ( .A1(n14438), .A2(n13935), .ZN(n13860) );
  NAND2_X1 U15859 ( .A1(n14284), .A2(n13933), .ZN(n13859) );
  NAND2_X1 U15860 ( .A1(n13860), .A2(n13859), .ZN(n13861) );
  XNOR2_X1 U15861 ( .A(n13861), .B(n12151), .ZN(n13864) );
  INV_X1 U15862 ( .A(n13864), .ZN(n13862) );
  AOI22_X1 U15863 ( .A1(n14438), .A2(n13933), .B1(n13932), .B2(n14284), .ZN(
        n13863) );
  NAND2_X1 U15864 ( .A1(n13862), .A2(n13863), .ZN(n13886) );
  INV_X1 U15865 ( .A(n13886), .ZN(n13865) );
  XNOR2_X1 U15866 ( .A(n13864), .B(n13863), .ZN(n13907) );
  NAND2_X1 U15867 ( .A1(n14433), .A2(n13935), .ZN(n13867) );
  NAND2_X1 U15868 ( .A1(n14228), .A2(n13933), .ZN(n13866) );
  NAND2_X1 U15869 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  AOI22_X1 U15870 ( .A1(n14433), .A2(n13933), .B1(n13932), .B2(n14228), .ZN(
        n13878) );
  AND2_X1 U15871 ( .A1(n14026), .A2(n13881), .ZN(n13961) );
  NAND2_X1 U15872 ( .A1(n14427), .A2(n13935), .ZN(n13870) );
  NAND2_X1 U15873 ( .A1(n14070), .A2(n11847), .ZN(n13869) );
  NAND2_X1 U15874 ( .A1(n13870), .A2(n13869), .ZN(n13871) );
  XNOR2_X1 U15875 ( .A(n13871), .B(n12151), .ZN(n13874) );
  INV_X1 U15876 ( .A(n13874), .ZN(n13872) );
  AOI22_X1 U15877 ( .A1(n14427), .A2(n13933), .B1(n13932), .B2(n14070), .ZN(
        n13873) );
  NAND2_X1 U15878 ( .A1(n13872), .A2(n13873), .ZN(n13880) );
  XNOR2_X1 U15879 ( .A(n13874), .B(n13873), .ZN(n13967) );
  AND2_X1 U15880 ( .A1(n13961), .A2(n13876), .ZN(n13875) );
  INV_X1 U15881 ( .A(n13877), .ZN(n13879) );
  NAND2_X1 U15882 ( .A1(n13879), .A2(n13878), .ZN(n13964) );
  AND2_X1 U15883 ( .A1(n13964), .A2(n13880), .ZN(n13888) );
  INV_X1 U15884 ( .A(n13882), .ZN(n13885) );
  INV_X1 U15885 ( .A(n13883), .ZN(n13884) );
  NAND2_X1 U15886 ( .A1(n13885), .A2(n13884), .ZN(n13905) );
  AND2_X1 U15887 ( .A1(n13905), .A2(n13886), .ZN(n13997) );
  AND2_X1 U15888 ( .A1(n13962), .A2(n13888), .ZN(n13889) );
  NAND2_X1 U15889 ( .A1(n14420), .A2(n13935), .ZN(n13893) );
  NAND2_X1 U15890 ( .A1(n14229), .A2(n11847), .ZN(n13892) );
  NAND2_X1 U15891 ( .A1(n13893), .A2(n13892), .ZN(n13894) );
  XNOR2_X1 U15892 ( .A(n13894), .B(n12151), .ZN(n13897) );
  AOI22_X1 U15893 ( .A1(n14420), .A2(n13933), .B1(n13932), .B2(n14229), .ZN(
        n13895) );
  XNOR2_X1 U15894 ( .A(n13897), .B(n13895), .ZN(n14046) );
  INV_X1 U15895 ( .A(n13895), .ZN(n13896) );
  NOR2_X1 U15896 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  XOR2_X1 U15897 ( .A(n13931), .B(n13930), .Z(n13904) );
  NOR2_X1 U15898 ( .A1(n13899), .A2(n14030), .ZN(n13902) );
  INV_X1 U15899 ( .A(n14057), .ZN(n14033) );
  AOI22_X1 U15900 ( .A1(n14229), .A2(n14033), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13900) );
  OAI21_X1 U15901 ( .B1(n14203), .B2(n14696), .A(n13900), .ZN(n13901) );
  AOI211_X1 U15902 ( .C1(n14205), .C2(n14687), .A(n13902), .B(n13901), .ZN(
        n13903) );
  OAI21_X1 U15903 ( .B1(n13904), .B2(n14065), .A(n13903), .ZN(P1_U3214) );
  NAND2_X1 U15904 ( .A1(n13960), .A2(n14026), .ZN(n14025) );
  NAND2_X1 U15905 ( .A1(n14025), .A2(n13905), .ZN(n13906) );
  XOR2_X1 U15906 ( .A(n13907), .B(n13906), .Z(n13912) );
  AOI22_X1 U15907 ( .A1(n14228), .A2(n14362), .B1(n14364), .B2(n14293), .ZN(
        n14260) );
  OAI22_X1 U15908 ( .A1(n14260), .A2(n14049), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13908), .ZN(n13909) );
  AOI21_X1 U15909 ( .B1(n14262), .B2(n14063), .A(n13909), .ZN(n13911) );
  NAND2_X1 U15910 ( .A1(n14438), .A2(n14687), .ZN(n13910) );
  OAI211_X1 U15911 ( .C1(n13912), .C2(n14065), .A(n13911), .B(n13910), .ZN(
        P1_U3216) );
  OAI211_X1 U15912 ( .C1(n13915), .C2(n13914), .A(n13913), .B(n14689), .ZN(
        n13920) );
  AOI22_X1 U15913 ( .A1(n14055), .A2(n14084), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13919) );
  AOI22_X1 U15914 ( .A1(n7859), .A2(n14063), .B1(n14687), .B2(n13916), .ZN(
        n13918) );
  NAND2_X1 U15915 ( .A1(n14033), .A2(n14086), .ZN(n13917) );
  NAND4_X1 U15916 ( .A1(n13920), .A2(n13919), .A3(n13918), .A4(n13917), .ZN(
        P1_U3218) );
  AOI21_X1 U15917 ( .B1(n13922), .B2(n13921), .A(n14065), .ZN(n13924) );
  NAND2_X1 U15918 ( .A1(n13924), .A2(n13923), .ZN(n13927) );
  AOI22_X1 U15919 ( .A1(n14363), .A2(n14364), .B1(n14362), .B2(n14292), .ZN(
        n14338) );
  NAND2_X1 U15920 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14175)
         );
  OAI21_X1 U15921 ( .B1(n14338), .B2(n14049), .A(n14175), .ZN(n13925) );
  AOI21_X1 U15922 ( .B1(n14333), .B2(n14063), .A(n13925), .ZN(n13926) );
  OAI211_X1 U15923 ( .C1(n14335), .C2(n14059), .A(n13927), .B(n13926), .ZN(
        P1_U3219) );
  AOI22_X1 U15924 ( .A1(n14409), .A2(n13933), .B1(n13932), .B2(n14193), .ZN(
        n13934) );
  XNOR2_X1 U15925 ( .A(n13934), .B(n12151), .ZN(n13937) );
  AOI22_X1 U15926 ( .A1(n14409), .A2(n13935), .B1(n11847), .B2(n14193), .ZN(
        n13936) );
  XNOR2_X1 U15927 ( .A(n13937), .B(n13936), .ZN(n13938) );
  XNOR2_X1 U15928 ( .A(n13939), .B(n13938), .ZN(n13948) );
  OAI22_X1 U15929 ( .A1(n13941), .A2(n14057), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13940), .ZN(n13946) );
  INV_X1 U15930 ( .A(n13942), .ZN(n13943) );
  OAI22_X1 U15931 ( .A1(n13944), .A2(n14030), .B1(n13943), .B2(n14696), .ZN(
        n13945) );
  AOI211_X1 U15932 ( .C1(n14409), .C2(n14687), .A(n13946), .B(n13945), .ZN(
        n13947) );
  OAI21_X1 U15933 ( .B1(n13948), .B2(n14065), .A(n13947), .ZN(P1_U3220) );
  INV_X1 U15934 ( .A(n13949), .ZN(n13950) );
  AOI21_X1 U15935 ( .B1(n13952), .B2(n13951), .A(n13950), .ZN(n13959) );
  OAI22_X1 U15936 ( .A1(n14030), .A2(n13954), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13953), .ZN(n13955) );
  AOI21_X1 U15937 ( .B1(n14033), .B2(n14292), .A(n13955), .ZN(n13956) );
  OAI21_X1 U15938 ( .B1(n14299), .B2(n14696), .A(n13956), .ZN(n13957) );
  AOI21_X1 U15939 ( .B1(n14449), .B2(n14687), .A(n13957), .ZN(n13958) );
  OAI21_X1 U15940 ( .B1(n13959), .B2(n14065), .A(n13958), .ZN(P1_U3223) );
  NAND2_X1 U15941 ( .A1(n13960), .A2(n13961), .ZN(n13963) );
  AND2_X1 U15942 ( .A1(n13963), .A2(n13962), .ZN(n13965) );
  NAND2_X1 U15943 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  XOR2_X1 U15944 ( .A(n13967), .B(n13966), .Z(n13972) );
  AOI22_X1 U15945 ( .A1(n14229), .A2(n14055), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13969) );
  NAND2_X1 U15946 ( .A1(n14033), .A2(n14228), .ZN(n13968) );
  OAI211_X1 U15947 ( .C1(n14696), .C2(n14232), .A(n13969), .B(n13968), .ZN(
        n13970) );
  AOI21_X1 U15948 ( .B1(n6805), .B2(n14687), .A(n13970), .ZN(n13971) );
  OAI21_X1 U15949 ( .B1(n13972), .B2(n14065), .A(n13971), .ZN(P1_U3225) );
  OAI21_X1 U15950 ( .B1(n13975), .B2(n13974), .A(n13973), .ZN(n13976) );
  NAND2_X1 U15951 ( .A1(n13976), .A2(n14689), .ZN(n13983) );
  OR2_X1 U15952 ( .A1(n13977), .A2(n14353), .ZN(n13979) );
  NAND2_X1 U15953 ( .A1(n14072), .A2(n14362), .ZN(n13978) );
  AND2_X1 U15954 ( .A1(n13979), .A2(n13978), .ZN(n14382) );
  OAI21_X1 U15955 ( .B1(n14382), .B2(n14049), .A(n13980), .ZN(n13981) );
  AOI21_X1 U15956 ( .B1(n14379), .B2(n14063), .A(n13981), .ZN(n13982) );
  OAI211_X1 U15957 ( .C1(n14395), .C2(n14059), .A(n13983), .B(n13982), .ZN(
        P1_U3226) );
  INV_X1 U15958 ( .A(n13987), .ZN(n13984) );
  NOR2_X1 U15959 ( .A1(n13985), .A2(n13984), .ZN(n13990) );
  AOI21_X1 U15960 ( .B1(n13988), .B2(n13987), .A(n13986), .ZN(n13989) );
  OAI21_X1 U15961 ( .B1(n13990), .B2(n13989), .A(n14689), .ZN(n13996) );
  NAND2_X1 U15962 ( .A1(n14055), .A2(n14363), .ZN(n13992) );
  OAI211_X1 U15963 ( .C1(n13993), .C2(n14057), .A(n13992), .B(n13991), .ZN(
        n13994) );
  AOI21_X1 U15964 ( .B1(n14370), .B2(n14063), .A(n13994), .ZN(n13995) );
  OAI211_X1 U15965 ( .C1(n6809), .C2(n14059), .A(n13996), .B(n13995), .ZN(
        P1_U3228) );
  NAND2_X1 U15966 ( .A1(n14025), .A2(n13997), .ZN(n13999) );
  XOR2_X1 U15967 ( .A(n14001), .B(n14000), .Z(n14006) );
  AOI22_X1 U15968 ( .A1(n14070), .A2(n14362), .B1(n14364), .B2(n14284), .ZN(
        n14247) );
  INV_X1 U15969 ( .A(n14253), .ZN(n14002) );
  AOI22_X1 U15970 ( .A1(n14063), .A2(n14002), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14003) );
  OAI21_X1 U15971 ( .B1(n14247), .B2(n14049), .A(n14003), .ZN(n14004) );
  AOI21_X1 U15972 ( .B1(n14433), .B2(n14687), .A(n14004), .ZN(n14005) );
  OAI21_X1 U15973 ( .B1(n14006), .B2(n14065), .A(n14005), .ZN(P1_U3229) );
  OAI211_X1 U15974 ( .C1(n14009), .C2(n14008), .A(n14007), .B(n14689), .ZN(
        n14015) );
  NAND2_X1 U15975 ( .A1(n14285), .A2(n14362), .ZN(n14011) );
  OR2_X1 U15976 ( .A1(n14352), .A2(n14353), .ZN(n14010) );
  NAND2_X1 U15977 ( .A1(n14011), .A2(n14010), .ZN(n14314) );
  AOI22_X1 U15978 ( .A1(n14691), .A2(n14314), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14012) );
  OAI21_X1 U15979 ( .B1(n14317), .B2(n14696), .A(n14012), .ZN(n14013) );
  AOI21_X1 U15980 ( .B1(n14455), .B2(n14687), .A(n14013), .ZN(n14014) );
  NAND2_X1 U15981 ( .A1(n14015), .A2(n14014), .ZN(P1_U3233) );
  XNOR2_X1 U15982 ( .A(n14017), .B(n14016), .ZN(n14024) );
  OAI22_X1 U15983 ( .A1(n14049), .A2(n14019), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14018), .ZN(n14020) );
  AOI21_X1 U15984 ( .B1(n14021), .B2(n14063), .A(n14020), .ZN(n14023) );
  NAND2_X1 U15985 ( .A1(n14710), .A2(n14687), .ZN(n14022) );
  OAI211_X1 U15986 ( .C1(n14024), .C2(n14065), .A(n14023), .B(n14022), .ZN(
        P1_U3234) );
  OAI21_X1 U15987 ( .B1(n14026), .B2(n13960), .A(n14025), .ZN(n14027) );
  NAND2_X1 U15988 ( .A1(n14027), .A2(n14689), .ZN(n14035) );
  NOR2_X1 U15989 ( .A1(n14696), .A2(n14278), .ZN(n14032) );
  OAI22_X1 U15990 ( .A1(n14030), .A2(n14029), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14028), .ZN(n14031) );
  AOI211_X1 U15991 ( .C1(n14033), .C2(n14285), .A(n14032), .B(n14031), .ZN(
        n14034) );
  OAI211_X1 U15992 ( .C1(n14059), .C2(n14281), .A(n14035), .B(n14034), .ZN(
        P1_U3235) );
  OAI21_X1 U15993 ( .B1(n14038), .B2(n14037), .A(n14036), .ZN(n14039) );
  NAND2_X1 U15994 ( .A1(n14039), .A2(n14689), .ZN(n14044) );
  NAND2_X1 U15995 ( .A1(n14055), .A2(n14071), .ZN(n14041) );
  OAI211_X1 U15996 ( .C1(n14354), .C2(n14057), .A(n14041), .B(n14040), .ZN(
        n14042) );
  AOI21_X1 U15997 ( .B1(n14345), .B2(n14063), .A(n14042), .ZN(n14043) );
  OAI211_X1 U15998 ( .C1(n14347), .C2(n14059), .A(n14044), .B(n14043), .ZN(
        P1_U3238) );
  XOR2_X1 U15999 ( .A(n14046), .B(n14045), .Z(n14052) );
  AND2_X1 U16000 ( .A1(n14070), .A2(n14364), .ZN(n14047) );
  AOI21_X1 U16001 ( .B1(n14069), .B2(n14362), .A(n14047), .ZN(n14215) );
  AOI22_X1 U16002 ( .A1(n14220), .A2(n14063), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14048) );
  OAI21_X1 U16003 ( .B1(n14215), .B2(n14049), .A(n14048), .ZN(n14050) );
  AOI21_X1 U16004 ( .B1(n14420), .B2(n14687), .A(n14050), .ZN(n14051) );
  OAI21_X1 U16005 ( .B1(n14052), .B2(n14065), .A(n14051), .ZN(P1_U3240) );
  AOI21_X1 U16006 ( .B1(n14054), .B2(n14053), .A(n6516), .ZN(n14066) );
  NAND2_X1 U16007 ( .A1(n14055), .A2(n14365), .ZN(n14056) );
  NAND2_X1 U16008 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14810)
         );
  OAI211_X1 U16009 ( .C1(n14058), .C2(n14057), .A(n14056), .B(n14810), .ZN(
        n14061) );
  NOR2_X1 U16010 ( .A1(n14697), .A2(n14059), .ZN(n14060) );
  AOI211_X1 U16011 ( .C1(n14063), .C2(n14062), .A(n14061), .B(n14060), .ZN(
        n14064) );
  OAI21_X1 U16012 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(P1_U3241) );
  MUX2_X1 U16013 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14067), .S(n14102), .Z(
        P1_U3590) );
  MUX2_X1 U16014 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14068), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16015 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14193), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16016 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14069), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16017 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14229), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16018 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14070), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16019 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14228), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16020 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14284), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16021 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14293), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16022 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14285), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16023 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14292), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16024 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14071), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16025 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14363), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16026 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14072), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16027 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14365), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16028 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14073), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16029 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14074), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16030 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14075), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16031 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14076), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16032 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14077), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16033 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14078), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16034 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14079), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16035 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14080), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16036 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14081), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16037 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14082), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16038 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14083), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16039 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14084), .S(n14102), .Z(
        P1_U3564) );
  MUX2_X1 U16040 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14085), .S(n14102), .Z(
        P1_U3563) );
  MUX2_X1 U16041 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14086), .S(n14102), .Z(
        P1_U3562) );
  MUX2_X1 U16042 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7088), .S(n14102), .Z(
        P1_U3561) );
  MUX2_X1 U16043 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8099), .S(n14102), .Z(
        P1_U3560) );
  OAI211_X1 U16044 ( .C1(n14089), .C2(n14088), .A(n14801), .B(n14087), .ZN(
        n14097) );
  AOI22_X1 U16045 ( .A1(n14757), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14096) );
  NAND2_X1 U16046 ( .A1(n14804), .A2(n14090), .ZN(n14095) );
  NAND2_X1 U16047 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14098) );
  INV_X1 U16048 ( .A(n14098), .ZN(n14093) );
  MUX2_X1 U16049 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n11710), .S(n14090), .Z(
        n14092) );
  OAI211_X1 U16050 ( .C1(n14093), .C2(n14092), .A(n14771), .B(n14091), .ZN(
        n14094) );
  NAND4_X1 U16051 ( .A1(n14097), .A2(n14096), .A3(n14095), .A4(n14094), .ZN(
        P1_U3244) );
  MUX2_X1 U16052 ( .A(n14099), .B(n14098), .S(n14749), .Z(n14103) );
  OR2_X1 U16053 ( .A1(n14516), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14100) );
  NAND2_X1 U16054 ( .A1(n14101), .A2(n14100), .ZN(n14750) );
  NAND2_X1 U16055 ( .A1(n14750), .A2(n14752), .ZN(n14755) );
  OAI211_X1 U16056 ( .C1(n14103), .C2(n7828), .A(n14102), .B(n14755), .ZN(
        n14778) );
  AOI22_X1 U16057 ( .A1(n14757), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14116) );
  OAI211_X1 U16058 ( .C1(n14106), .C2(n14105), .A(n14801), .B(n14104), .ZN(
        n14112) );
  INV_X1 U16059 ( .A(n14107), .ZN(n14108) );
  XNOR2_X1 U16060 ( .A(n14109), .B(n14108), .ZN(n14110) );
  NAND2_X1 U16061 ( .A1(n14771), .A2(n14110), .ZN(n14111) );
  AND2_X1 U16062 ( .A1(n14112), .A2(n14111), .ZN(n14115) );
  NAND2_X1 U16063 ( .A1(n14804), .A2(n14113), .ZN(n14114) );
  NAND4_X1 U16064 ( .A1(n14778), .A2(n14116), .A3(n14115), .A4(n14114), .ZN(
        P1_U3245) );
  OAI211_X1 U16065 ( .C1(n14118), .C2(n14117), .A(n14801), .B(n14761), .ZN(
        n14126) );
  NOR2_X1 U16066 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7859), .ZN(n14119) );
  AOI21_X1 U16067 ( .B1(n14757), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14119), .ZN(
        n14125) );
  NAND2_X1 U16068 ( .A1(n14804), .A2(n14120), .ZN(n14124) );
  OAI211_X1 U16069 ( .C1(n14122), .C2(n14121), .A(n14771), .B(n14767), .ZN(
        n14123) );
  NAND4_X1 U16070 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        P1_U3246) );
  OAI21_X1 U16071 ( .B1(n14129), .B2(n14128), .A(n14127), .ZN(n14130) );
  NAND2_X1 U16072 ( .A1(n14130), .A2(n14801), .ZN(n14142) );
  AOI21_X1 U16073 ( .B1(n14757), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14131), .ZN(
        n14141) );
  MUX2_X1 U16074 ( .A(n10749), .B(P1_REG2_REG_9__SCAN_IN), .S(n14138), .Z(
        n14134) );
  INV_X1 U16075 ( .A(n14132), .ZN(n14133) );
  NAND2_X1 U16076 ( .A1(n14134), .A2(n14133), .ZN(n14136) );
  OAI211_X1 U16077 ( .C1(n14137), .C2(n14136), .A(n14135), .B(n14771), .ZN(
        n14140) );
  NAND2_X1 U16078 ( .A1(n14804), .A2(n14138), .ZN(n14139) );
  NAND4_X1 U16079 ( .A1(n14142), .A2(n14141), .A3(n14140), .A4(n14139), .ZN(
        P1_U3252) );
  OAI211_X1 U16080 ( .C1(n14145), .C2(n14144), .A(n14771), .B(n14143), .ZN(
        n14155) );
  NAND2_X1 U16081 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14693)
         );
  INV_X1 U16082 ( .A(n14693), .ZN(n14146) );
  AOI21_X1 U16083 ( .B1(n14757), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n14146), 
        .ZN(n14154) );
  OAI21_X1 U16084 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14150) );
  NAND2_X1 U16085 ( .A1(n14150), .A2(n14801), .ZN(n14153) );
  NAND2_X1 U16086 ( .A1(n14804), .A2(n14151), .ZN(n14152) );
  NAND4_X1 U16087 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        P1_U3257) );
  INV_X1 U16088 ( .A(n14757), .ZN(n14812) );
  NOR2_X1 U16089 ( .A1(n14157), .A2(n14156), .ZN(n14158) );
  NOR2_X1 U16090 ( .A1(n14159), .A2(n14158), .ZN(n14160) );
  XNOR2_X1 U16091 ( .A(n14160), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14171) );
  NAND2_X1 U16092 ( .A1(n14162), .A2(n14161), .ZN(n14163) );
  NAND2_X1 U16093 ( .A1(n14164), .A2(n14163), .ZN(n14165) );
  XOR2_X1 U16094 ( .A(n14165), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14170) );
  INV_X1 U16095 ( .A(n14170), .ZN(n14166) );
  NAND2_X1 U16096 ( .A1(n14166), .A2(n14771), .ZN(n14167) );
  OAI211_X1 U16097 ( .C1(n14171), .C2(n14168), .A(n14775), .B(n14167), .ZN(
        n14169) );
  INV_X1 U16098 ( .A(n14169), .ZN(n14174) );
  AOI22_X1 U16099 ( .A1(n14171), .A2(n14801), .B1(n14771), .B2(n14170), .ZN(
        n14173) );
  OAI211_X1 U16100 ( .C1(n14177), .C2(n14812), .A(n14176), .B(n14175), .ZN(
        P1_U3262) );
  NAND2_X1 U16101 ( .A1(n14179), .A2(n14178), .ZN(n14405) );
  NOR2_X1 U16102 ( .A1(n14377), .A2(n14405), .ZN(n14185) );
  AOI21_X1 U16103 ( .B1(n14377), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14185), 
        .ZN(n14181) );
  NAND2_X1 U16104 ( .A1(n8424), .A2(n14322), .ZN(n14180) );
  OAI211_X1 U16105 ( .C1(n14402), .C2(n14319), .A(n14181), .B(n14180), .ZN(
        P1_U3263) );
  INV_X1 U16106 ( .A(n14182), .ZN(n14183) );
  NAND2_X1 U16107 ( .A1(n14184), .A2(n14183), .ZN(n14404) );
  NAND3_X1 U16108 ( .A1(n14404), .A2(n14397), .A3(n14403), .ZN(n14187) );
  AOI21_X1 U16109 ( .B1(n14377), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14185), 
        .ZN(n14186) );
  OAI211_X1 U16110 ( .C1(n14407), .C2(n14394), .A(n14187), .B(n14186), .ZN(
        P1_U3264) );
  AND2_X1 U16111 ( .A1(n14219), .A2(n14205), .ZN(n14189) );
  XNOR2_X1 U16112 ( .A(n14191), .B(n14190), .ZN(n14192) );
  NAND2_X1 U16113 ( .A1(n14192), .A2(n14384), .ZN(n14201) );
  AOI22_X1 U16114 ( .A1(n14193), .A2(n14362), .B1(n14364), .B2(n14229), .ZN(
        n14200) );
  NAND2_X1 U16115 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  NAND2_X1 U16116 ( .A1(n14197), .A2(n14196), .ZN(n14198) );
  NAND2_X1 U16117 ( .A1(n14198), .A2(n14879), .ZN(n14199) );
  NAND3_X1 U16118 ( .A1(n14201), .A2(n14200), .A3(n14199), .ZN(n14417) );
  NAND2_X1 U16119 ( .A1(n14417), .A2(n14393), .ZN(n14207) );
  INV_X1 U16120 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14202) );
  OAI22_X1 U16121 ( .A1(n14203), .A2(n14386), .B1(n14202), .B2(n14393), .ZN(
        n14204) );
  AOI21_X1 U16122 ( .B1(n14205), .B2(n14322), .A(n14204), .ZN(n14206) );
  OAI211_X1 U16123 ( .C1(n14415), .C2(n14319), .A(n14207), .B(n14206), .ZN(
        P1_U3266) );
  OR2_X1 U16124 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U16125 ( .A1(n14211), .A2(n14210), .ZN(n14423) );
  XNOR2_X1 U16126 ( .A(n14213), .B(n14212), .ZN(n14214) );
  NAND2_X1 U16127 ( .A1(n14214), .A2(n14384), .ZN(n14216) );
  NAND2_X1 U16128 ( .A1(n14216), .A2(n14215), .ZN(n14424) );
  NAND2_X1 U16129 ( .A1(n14424), .A2(n14393), .ZN(n14224) );
  NAND2_X1 U16130 ( .A1(n14217), .A2(n14420), .ZN(n14218) );
  AND2_X1 U16131 ( .A1(n14219), .A2(n14218), .ZN(n14421) );
  AOI22_X1 U16132 ( .A1(n14220), .A2(n14369), .B1(n14377), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n14221) );
  OAI21_X1 U16133 ( .B1(n6801), .B2(n14394), .A(n14221), .ZN(n14222) );
  AOI21_X1 U16134 ( .B1(n14397), .B2(n14421), .A(n14222), .ZN(n14223) );
  OAI211_X1 U16135 ( .C1(n14423), .C2(n14400), .A(n14224), .B(n14223), .ZN(
        P1_U3267) );
  OAI21_X1 U16136 ( .B1(n14226), .B2(n14237), .A(n14225), .ZN(n14227) );
  NAND2_X1 U16137 ( .A1(n14227), .A2(n14384), .ZN(n14231) );
  AOI22_X1 U16138 ( .A1(n14229), .A2(n14362), .B1(n14364), .B2(n14228), .ZN(
        n14230) );
  NAND2_X1 U16139 ( .A1(n14231), .A2(n14230), .ZN(n14432) );
  INV_X1 U16140 ( .A(n14432), .ZN(n14241) );
  XNOR2_X1 U16141 ( .A(n6805), .B(n6529), .ZN(n14428) );
  INV_X1 U16142 ( .A(n14232), .ZN(n14233) );
  AOI22_X1 U16143 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(n14377), .B1(n14233), 
        .B2(n14369), .ZN(n14234) );
  OAI21_X1 U16144 ( .B1(n14235), .B2(n14394), .A(n14234), .ZN(n14236) );
  AOI21_X1 U16145 ( .B1(n14397), .B2(n14428), .A(n14236), .ZN(n14240) );
  NAND2_X1 U16146 ( .A1(n6572), .A2(n14237), .ZN(n14426) );
  NAND3_X1 U16147 ( .A1(n14426), .A2(n14238), .A3(n14325), .ZN(n14239) );
  OAI211_X1 U16148 ( .C1(n14241), .C2(n14377), .A(n14240), .B(n14239), .ZN(
        P1_U3268) );
  INV_X1 U16149 ( .A(n14242), .ZN(n14243) );
  AOI21_X1 U16150 ( .B1(n14245), .B2(n14244), .A(n14243), .ZN(n14437) );
  AOI21_X1 U16151 ( .B1(n14433), .B2(n14264), .A(n6529), .ZN(n14434) );
  INV_X1 U16152 ( .A(n14434), .ZN(n14251) );
  AOI21_X1 U16153 ( .B1(n8137), .B2(n14246), .A(n14348), .ZN(n14250) );
  INV_X1 U16154 ( .A(n14247), .ZN(n14248) );
  AOI21_X1 U16155 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(n14436) );
  OAI21_X1 U16156 ( .B1(n10846), .B2(n14251), .A(n14436), .ZN(n14252) );
  NAND2_X1 U16157 ( .A1(n14252), .A2(n14393), .ZN(n14257) );
  INV_X1 U16158 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14254) );
  OAI22_X1 U16159 ( .A1(n14393), .A2(n14254), .B1(n14253), .B2(n14386), .ZN(
        n14255) );
  AOI21_X1 U16160 ( .B1(n14433), .B2(n14322), .A(n14255), .ZN(n14256) );
  OAI211_X1 U16161 ( .C1(n14437), .C2(n14400), .A(n14257), .B(n14256), .ZN(
        P1_U3269) );
  XNOR2_X1 U16162 ( .A(n14258), .B(n14267), .ZN(n14259) );
  NAND2_X1 U16163 ( .A1(n14259), .A2(n14384), .ZN(n14261) );
  NAND2_X1 U16164 ( .A1(n14261), .A2(n14260), .ZN(n14443) );
  AOI21_X1 U16165 ( .B1(n14262), .B2(n14369), .A(n14443), .ZN(n14274) );
  OR2_X1 U16166 ( .A1(n14266), .A2(n14277), .ZN(n14263) );
  AND2_X1 U16167 ( .A1(n14264), .A2(n14263), .ZN(n14439) );
  INV_X1 U16168 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14265) );
  OAI22_X1 U16169 ( .A1(n14266), .A2(n14394), .B1(n14265), .B2(n14393), .ZN(
        n14272) );
  NAND2_X1 U16170 ( .A1(n14268), .A2(n14267), .ZN(n14269) );
  NAND2_X1 U16171 ( .A1(n14270), .A2(n14269), .ZN(n14441) );
  NOR2_X1 U16172 ( .A1(n14441), .A2(n14400), .ZN(n14271) );
  AOI211_X1 U16173 ( .C1(n14439), .C2(n14397), .A(n14272), .B(n14271), .ZN(
        n14273) );
  OAI21_X1 U16174 ( .B1(n14274), .B2(n14377), .A(n14273), .ZN(P1_U3270) );
  XNOR2_X1 U16175 ( .A(n14275), .B(n14283), .ZN(n14448) );
  AND2_X1 U16176 ( .A1(n14444), .A2(n14296), .ZN(n14276) );
  NOR2_X1 U16177 ( .A1(n14277), .A2(n14276), .ZN(n14445) );
  INV_X1 U16178 ( .A(n14278), .ZN(n14279) );
  AOI22_X1 U16179 ( .A1(n14377), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14279), 
        .B2(n14369), .ZN(n14280) );
  OAI21_X1 U16180 ( .B1(n14281), .B2(n14394), .A(n14280), .ZN(n14288) );
  OAI21_X1 U16181 ( .B1(n14283), .B2(n6600), .A(n14282), .ZN(n14286) );
  AOI222_X1 U16182 ( .A1(n14384), .A2(n14286), .B1(n14285), .B2(n14364), .C1(
        n14284), .C2(n14362), .ZN(n14447) );
  NOR2_X1 U16183 ( .A1(n14447), .A2(n14377), .ZN(n14287) );
  AOI211_X1 U16184 ( .C1(n14445), .C2(n14397), .A(n14288), .B(n14287), .ZN(
        n14289) );
  OAI21_X1 U16185 ( .B1(n14448), .B2(n14400), .A(n14289), .ZN(P1_U3271) );
  OAI211_X1 U16186 ( .C1(n14306), .C2(n14291), .A(n14290), .B(n14384), .ZN(
        n14295) );
  AOI22_X1 U16187 ( .A1(n14293), .A2(n14362), .B1(n14364), .B2(n14292), .ZN(
        n14294) );
  AND2_X1 U16188 ( .A1(n14295), .A2(n14294), .ZN(n14452) );
  INV_X1 U16189 ( .A(n14456), .ZN(n14298) );
  INV_X1 U16190 ( .A(n14296), .ZN(n14297) );
  AOI21_X1 U16191 ( .B1(n14449), .B2(n14298), .A(n14297), .ZN(n14450) );
  INV_X1 U16192 ( .A(n14299), .ZN(n14300) );
  AOI22_X1 U16193 ( .A1(n14377), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14300), 
        .B2(n14369), .ZN(n14301) );
  OAI21_X1 U16194 ( .B1(n14302), .B2(n14394), .A(n14301), .ZN(n14308) );
  INV_X1 U16195 ( .A(n14303), .ZN(n14304) );
  AOI21_X1 U16196 ( .B1(n14306), .B2(n6475), .A(n14304), .ZN(n14453) );
  NOR2_X1 U16197 ( .A1(n14453), .A2(n14400), .ZN(n14307) );
  AOI211_X1 U16198 ( .C1(n14450), .C2(n14397), .A(n14308), .B(n14307), .ZN(
        n14309) );
  OAI21_X1 U16199 ( .B1(n14377), .B2(n14452), .A(n14309), .ZN(P1_U3272) );
  NAND2_X1 U16200 ( .A1(n14311), .A2(n14310), .ZN(n14312) );
  NAND3_X1 U16201 ( .A1(n14313), .A2(n14384), .A3(n14312), .ZN(n14316) );
  INV_X1 U16202 ( .A(n14314), .ZN(n14315) );
  NAND2_X1 U16203 ( .A1(n14316), .A2(n14315), .ZN(n14462) );
  INV_X1 U16204 ( .A(n14462), .ZN(n14328) );
  INV_X1 U16205 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14318) );
  OAI22_X1 U16206 ( .A1(n14393), .A2(n14318), .B1(n14317), .B2(n14386), .ZN(
        n14321) );
  AND2_X1 U16207 ( .A1(n14331), .A2(n14455), .ZN(n14457) );
  NOR3_X1 U16208 ( .A1(n14456), .A2(n14457), .A3(n14319), .ZN(n14320) );
  AOI211_X1 U16209 ( .C1(n14322), .C2(n14455), .A(n14321), .B(n14320), .ZN(
        n14327) );
  NAND2_X1 U16210 ( .A1(n14324), .A2(n8007), .ZN(n14454) );
  NAND3_X1 U16211 ( .A1(n14323), .A2(n14454), .A3(n14325), .ZN(n14326) );
  OAI211_X1 U16212 ( .C1(n14328), .C2(n14377), .A(n14327), .B(n14326), .ZN(
        P1_U3273) );
  XNOR2_X1 U16213 ( .A(n14329), .B(n14337), .ZN(n14469) );
  INV_X1 U16214 ( .A(n14331), .ZN(n14332) );
  AOI21_X1 U16215 ( .B1(n14465), .B2(n6810), .A(n14332), .ZN(n14466) );
  AOI22_X1 U16216 ( .A1(n14377), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14333), 
        .B2(n14369), .ZN(n14334) );
  OAI21_X1 U16217 ( .B1(n14335), .B2(n14394), .A(n14334), .ZN(n14342) );
  OAI21_X1 U16218 ( .B1(n7492), .B2(n14337), .A(n14336), .ZN(n14340) );
  INV_X1 U16219 ( .A(n14338), .ZN(n14339) );
  AOI21_X1 U16220 ( .B1(n14340), .B2(n14384), .A(n14339), .ZN(n14468) );
  NOR2_X1 U16221 ( .A1(n14468), .A2(n14377), .ZN(n14341) );
  AOI211_X1 U16222 ( .C1(n14466), .C2(n14397), .A(n14342), .B(n14341), .ZN(
        n14343) );
  OAI21_X1 U16223 ( .B1(n14469), .B2(n14400), .A(n14343), .ZN(P1_U3274) );
  XNOR2_X1 U16224 ( .A(n14344), .B(n14349), .ZN(n14474) );
  AOI21_X1 U16225 ( .B1(n14470), .B2(n14367), .A(n14330), .ZN(n14471) );
  AOI22_X1 U16226 ( .A1(n14377), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14345), 
        .B2(n14369), .ZN(n14346) );
  OAI21_X1 U16227 ( .B1(n14347), .B2(n14394), .A(n14346), .ZN(n14359) );
  AOI21_X1 U16228 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n14357) );
  OAI22_X1 U16229 ( .A1(n14354), .A2(n14353), .B1(n14352), .B2(n14351), .ZN(
        n14355) );
  AOI21_X1 U16230 ( .B1(n14357), .B2(n14356), .A(n14355), .ZN(n14473) );
  NOR2_X1 U16231 ( .A1(n14473), .A2(n14377), .ZN(n14358) );
  AOI211_X1 U16232 ( .C1(n14471), .C2(n14397), .A(n14359), .B(n14358), .ZN(
        n14360) );
  OAI21_X1 U16233 ( .B1(n14474), .B2(n14400), .A(n14360), .ZN(P1_U3275) );
  XNOR2_X1 U16234 ( .A(n14361), .B(n14373), .ZN(n14366) );
  AOI222_X1 U16235 ( .A1(n14384), .A2(n14366), .B1(n14365), .B2(n14364), .C1(
        n14363), .C2(n14362), .ZN(n14478) );
  INV_X1 U16236 ( .A(n14367), .ZN(n14368) );
  AOI21_X1 U16237 ( .B1(n14475), .B2(n14390), .A(n14368), .ZN(n14476) );
  AOI22_X1 U16238 ( .A1(n14377), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14370), 
        .B2(n14369), .ZN(n14371) );
  OAI21_X1 U16239 ( .B1(n6809), .B2(n14394), .A(n14371), .ZN(n14375) );
  XNOR2_X1 U16240 ( .A(n14372), .B(n14373), .ZN(n14479) );
  NOR2_X1 U16241 ( .A1(n14479), .A2(n14400), .ZN(n14374) );
  AOI211_X1 U16242 ( .C1(n14476), .C2(n14397), .A(n14375), .B(n14374), .ZN(
        n14376) );
  OAI21_X1 U16243 ( .B1(n14478), .B2(n14377), .A(n14376), .ZN(P1_U3276) );
  XNOR2_X1 U16244 ( .A(n14378), .B(n14381), .ZN(n14484) );
  INV_X1 U16245 ( .A(n14379), .ZN(n14387) );
  OAI21_X1 U16246 ( .B1(n6629), .B2(n14381), .A(n14380), .ZN(n14385) );
  INV_X1 U16247 ( .A(n14382), .ZN(n14383) );
  AOI21_X1 U16248 ( .B1(n14385), .B2(n14384), .A(n14383), .ZN(n14483) );
  OAI21_X1 U16249 ( .B1(n14387), .B2(n14386), .A(n14483), .ZN(n14388) );
  NAND2_X1 U16250 ( .A1(n14388), .A2(n14393), .ZN(n14399) );
  INV_X1 U16251 ( .A(n14389), .ZN(n14392) );
  INV_X1 U16252 ( .A(n14390), .ZN(n14391) );
  AOI21_X1 U16253 ( .B1(n14480), .B2(n14392), .A(n14391), .ZN(n14481) );
  OAI22_X1 U16254 ( .A1(n14395), .A2(n14394), .B1(n14393), .B2(n11766), .ZN(
        n14396) );
  AOI21_X1 U16255 ( .B1(n14481), .B2(n14397), .A(n14396), .ZN(n14398) );
  OAI211_X1 U16256 ( .C1(n14484), .C2(n14400), .A(n14399), .B(n14398), .ZN(
        P1_U3277) );
  NAND2_X1 U16257 ( .A1(n8424), .A2(n14882), .ZN(n14401) );
  OAI211_X1 U16258 ( .C1(n14402), .C2(n10323), .A(n14401), .B(n14405), .ZN(
        n14486) );
  MUX2_X1 U16259 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14486), .S(n14916), .Z(
        P1_U3559) );
  NAND3_X1 U16260 ( .A1(n14404), .A2(n14883), .A3(n14403), .ZN(n14406) );
  OAI211_X1 U16261 ( .C1(n14407), .C2(n14875), .A(n14406), .B(n14405), .ZN(
        n14487) );
  MUX2_X1 U16262 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14487), .S(n14916), .Z(
        P1_U3558) );
  NAND3_X1 U16263 ( .A1(n6495), .A2(n14904), .A3(n14408), .ZN(n14413) );
  AOI22_X1 U16264 ( .A1(n14410), .A2(n14883), .B1(n14882), .B2(n14409), .ZN(
        n14411) );
  NAND3_X1 U16265 ( .A1(n14413), .A2(n14412), .A3(n14411), .ZN(n14488) );
  MUX2_X1 U16266 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14488), .S(n14916), .Z(
        P1_U3556) );
  OAI22_X1 U16267 ( .A1(n14415), .A2(n10323), .B1(n14414), .B2(n14875), .ZN(
        n14416) );
  NOR2_X1 U16268 ( .A1(n14417), .A2(n14416), .ZN(n14489) );
  MUX2_X1 U16269 ( .A(n14418), .B(n14489), .S(n14916), .Z(n14419) );
  INV_X1 U16270 ( .A(n14419), .ZN(P1_U3555) );
  AOI22_X1 U16271 ( .A1(n14421), .A2(n14883), .B1(n14882), .B2(n14420), .ZN(
        n14422) );
  OAI21_X1 U16272 ( .B1(n14423), .B2(n14888), .A(n14422), .ZN(n14425) );
  MUX2_X1 U16273 ( .A(n14492), .B(P1_REG1_REG_26__SCAN_IN), .S(n14917), .Z(
        P1_U3554) );
  NAND3_X1 U16274 ( .A1(n14426), .A2(n14238), .A3(n14904), .ZN(n14430) );
  AOI22_X1 U16275 ( .A1(n14428), .A2(n14883), .B1(n14882), .B2(n14427), .ZN(
        n14429) );
  NAND2_X1 U16276 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  MUX2_X1 U16277 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14493), .S(n14916), .Z(
        P1_U3553) );
  AOI22_X1 U16278 ( .A1(n14434), .A2(n14883), .B1(n14882), .B2(n14433), .ZN(
        n14435) );
  OAI211_X1 U16279 ( .C1(n14437), .C2(n14888), .A(n14436), .B(n14435), .ZN(
        n14494) );
  MUX2_X1 U16280 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14494), .S(n14916), .Z(
        P1_U3552) );
  AOI22_X1 U16281 ( .A1(n14439), .A2(n14883), .B1(n14882), .B2(n14438), .ZN(
        n14440) );
  OAI21_X1 U16282 ( .B1(n14441), .B2(n14888), .A(n14440), .ZN(n14442) );
  MUX2_X1 U16283 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14495), .S(n14916), .Z(
        P1_U3551) );
  AOI22_X1 U16284 ( .A1(n14445), .A2(n14883), .B1(n14444), .B2(n14882), .ZN(
        n14446) );
  OAI211_X1 U16285 ( .C1(n14888), .C2(n14448), .A(n14447), .B(n14446), .ZN(
        n14496) );
  MUX2_X1 U16286 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14496), .S(n14916), .Z(
        P1_U3550) );
  AOI22_X1 U16287 ( .A1(n14450), .A2(n14883), .B1(n14882), .B2(n14449), .ZN(
        n14451) );
  OAI211_X1 U16288 ( .C1(n14453), .C2(n14888), .A(n14452), .B(n14451), .ZN(
        n14497) );
  MUX2_X1 U16289 ( .A(n14497), .B(P1_REG1_REG_21__SCAN_IN), .S(n14917), .Z(
        P1_U3549) );
  NAND3_X1 U16290 ( .A1(n14323), .A2(n14454), .A3(n14904), .ZN(n14460) );
  NAND2_X1 U16291 ( .A1(n14455), .A2(n14882), .ZN(n14459) );
  OR3_X1 U16292 ( .A1(n14457), .A2(n14456), .A3(n10323), .ZN(n14458) );
  NAND3_X1 U16293 ( .A1(n14460), .A2(n14459), .A3(n14458), .ZN(n14461) );
  NOR2_X1 U16294 ( .A1(n14462), .A2(n14461), .ZN(n14499) );
  INV_X1 U16295 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14463) );
  MUX2_X1 U16296 ( .A(n14499), .B(n14463), .S(n14917), .Z(n14464) );
  INV_X1 U16297 ( .A(n14464), .ZN(P1_U3548) );
  AOI22_X1 U16298 ( .A1(n14466), .A2(n14883), .B1(n14882), .B2(n14465), .ZN(
        n14467) );
  OAI211_X1 U16299 ( .C1(n14888), .C2(n14469), .A(n14468), .B(n14467), .ZN(
        n14501) );
  MUX2_X1 U16300 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14501), .S(n14916), .Z(
        P1_U3547) );
  AOI22_X1 U16301 ( .A1(n14471), .A2(n14883), .B1(n14882), .B2(n14470), .ZN(
        n14472) );
  OAI211_X1 U16302 ( .C1(n14888), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        n14502) );
  MUX2_X1 U16303 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14502), .S(n14916), .Z(
        P1_U3546) );
  AOI22_X1 U16304 ( .A1(n14476), .A2(n14883), .B1(n14882), .B2(n14475), .ZN(
        n14477) );
  OAI211_X1 U16305 ( .C1(n14888), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n14503) );
  MUX2_X1 U16306 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14503), .S(n14916), .Z(
        P1_U3545) );
  AOI22_X1 U16307 ( .A1(n14481), .A2(n14883), .B1(n14882), .B2(n14480), .ZN(
        n14482) );
  OAI211_X1 U16308 ( .C1(n14888), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14505) );
  MUX2_X1 U16309 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14505), .S(n14916), .Z(
        P1_U3544) );
  MUX2_X1 U16310 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14485), .S(n14916), .Z(
        P1_U3528) );
  MUX2_X1 U16311 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14486), .S(n14504), .Z(
        P1_U3527) );
  MUX2_X1 U16312 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14487), .S(n14504), .Z(
        P1_U3526) );
  MUX2_X1 U16313 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14488), .S(n14504), .Z(
        P1_U3524) );
  INV_X1 U16314 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14490) );
  MUX2_X1 U16315 ( .A(n14490), .B(n14489), .S(n14504), .Z(n14491) );
  INV_X1 U16316 ( .A(n14491), .ZN(P1_U3523) );
  MUX2_X1 U16317 ( .A(n14492), .B(P1_REG0_REG_26__SCAN_IN), .S(n14905), .Z(
        P1_U3522) );
  MUX2_X1 U16318 ( .A(n14493), .B(P1_REG0_REG_25__SCAN_IN), .S(n14905), .Z(
        P1_U3521) );
  MUX2_X1 U16319 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14494), .S(n14504), .Z(
        P1_U3520) );
  MUX2_X1 U16320 ( .A(n14495), .B(P1_REG0_REG_23__SCAN_IN), .S(n14905), .Z(
        P1_U3519) );
  MUX2_X1 U16321 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14496), .S(n14504), .Z(
        P1_U3518) );
  MUX2_X1 U16322 ( .A(n14497), .B(P1_REG0_REG_21__SCAN_IN), .S(n14905), .Z(
        P1_U3517) );
  INV_X1 U16323 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14498) );
  MUX2_X1 U16324 ( .A(n14499), .B(n14498), .S(n14905), .Z(n14500) );
  INV_X1 U16325 ( .A(n14500), .ZN(P1_U3516) );
  MUX2_X1 U16326 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14501), .S(n14504), .Z(
        P1_U3515) );
  MUX2_X1 U16327 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14502), .S(n14504), .Z(
        P1_U3513) );
  MUX2_X1 U16328 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14503), .S(n14504), .Z(
        P1_U3510) );
  MUX2_X1 U16329 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14505), .S(n14504), .Z(
        P1_U3507) );
  INV_X1 U16330 ( .A(n14506), .ZN(n14507) );
  NOR4_X1 U16331 ( .A1(n14507), .A2(P1_IR_REG_30__SCAN_IN), .A3(n7832), .A4(
        P1_U3086), .ZN(n14508) );
  AOI21_X1 U16332 ( .B1(n14509), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14508), 
        .ZN(n14510) );
  OAI21_X1 U16333 ( .B1(n14511), .B2(n14521), .A(n14510), .ZN(P1_U3324) );
  OAI222_X1 U16334 ( .A1(n14527), .A2(n14515), .B1(P1_U3086), .B2(n14513), 
        .C1(n14521), .C2(n14512), .ZN(P1_U3326) );
  OAI222_X1 U16335 ( .A1(n14527), .A2(n14518), .B1(n14525), .B2(n14517), .C1(
        n14516), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16336 ( .A1(n14522), .A2(P1_U3086), .B1(n14521), .B2(n14520), 
        .C1(n14519), .C2(n14527), .ZN(P1_U3329) );
  OAI222_X1 U16337 ( .A1(n14527), .A2(n14526), .B1(n14525), .B2(n14524), .C1(
        n14523), .C2(P1_U3086), .ZN(P1_U3330) );
  MUX2_X1 U16338 ( .A(n14528), .B(n8194), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16339 ( .A(n14529), .ZN(n14530) );
  MUX2_X1 U16340 ( .A(n14530), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U16341 ( .A1(n14532), .A2(n14531), .ZN(n14533) );
  XOR2_X1 U16342 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14533), .Z(SUB_1596_U62)
         );
  AOI21_X1 U16343 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14534) );
  OAI21_X1 U16344 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14534), 
        .ZN(U28) );
  OAI221_X1 U16345 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7499), .C2(n14536), .A(n14535), .ZN(U29) );
  OAI21_X1 U16346 ( .B1(n14539), .B2(n14538), .A(n14537), .ZN(n14540) );
  XNOR2_X1 U16347 ( .A(n14540), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16348 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(SUB_1596_U57) );
  OAI222_X1 U16349 ( .A1(n14548), .A2(n14547), .B1(n14548), .B2(n14546), .C1(
        n14545), .C2(n14544), .ZN(SUB_1596_U55) );
  AOI21_X1 U16350 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(SUB_1596_U54) );
  AOI21_X1 U16351 ( .B1(n14554), .B2(n14553), .A(n14552), .ZN(n14555) );
  XOR2_X1 U16352 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14555), .Z(SUB_1596_U70)
         );
  OAI22_X1 U16353 ( .A1(n14557), .A2(n10323), .B1(n14556), .B2(n14875), .ZN(
        n14559) );
  NOR2_X1 U16354 ( .A1(n14559), .A2(n14558), .ZN(n14562) );
  INV_X1 U16355 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14560) );
  AOI22_X1 U16356 ( .A1(n14504), .A2(n14562), .B1(n14560), .B2(n14905), .ZN(
        P1_U3495) );
  AOI22_X1 U16357 ( .A1(n14916), .A2(n14562), .B1(n14561), .B2(n14917), .ZN(
        P1_U3540) );
  AOI21_X1 U16358 ( .B1(n14564), .B2(n14563), .A(n6602), .ZN(n14565) );
  XNOR2_X1 U16359 ( .A(n14565), .B(n15038), .ZN(SUB_1596_U63) );
  AOI22_X1 U16360 ( .A1(n14584), .A2(n14566), .B1(n15245), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14582) );
  XNOR2_X1 U16361 ( .A(n14568), .B(n14567), .ZN(n14575) );
  INV_X1 U16362 ( .A(n14569), .ZN(n14571) );
  NAND2_X1 U16363 ( .A1(n14571), .A2(n14570), .ZN(n14572) );
  XNOR2_X1 U16364 ( .A(n14573), .B(n14572), .ZN(n14574) );
  AOI22_X1 U16365 ( .A1(n14575), .A2(n15287), .B1(n14574), .B2(n15280), .ZN(
        n14581) );
  NAND2_X1 U16366 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14580)
         );
  OAI221_X1 U16367 ( .B1(n14578), .B2(n14577), .C1(n14578), .C2(n14576), .A(
        n14593), .ZN(n14579) );
  NAND4_X1 U16368 ( .A1(n14582), .A2(n14581), .A3(n14580), .A4(n14579), .ZN(
        P3_U3198) );
  AOI22_X1 U16369 ( .A1(n14584), .A2(n14583), .B1(n15245), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14600) );
  OAI21_X1 U16370 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14586), .A(n14585), 
        .ZN(n14591) );
  AOI211_X1 U16371 ( .C1(n14589), .C2(n14588), .A(n15241), .B(n14587), .ZN(
        n14590) );
  AOI21_X1 U16372 ( .B1(n15287), .B2(n14591), .A(n14590), .ZN(n14599) );
  NAND2_X1 U16373 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14598)
         );
  OAI221_X1 U16374 ( .B1(n14596), .B2(n14595), .C1(n14596), .C2(n14594), .A(
        n14593), .ZN(n14597) );
  NAND4_X1 U16375 ( .A1(n14600), .A2(n14599), .A3(n14598), .A4(n14597), .ZN(
        P3_U3199) );
  INV_X1 U16376 ( .A(n14601), .ZN(n14602) );
  AOI22_X1 U16377 ( .A1(n14604), .A2(n15331), .B1(n14614), .B2(n15334), .ZN(
        n14609) );
  AOI22_X1 U16378 ( .A1(n14605), .A2(n14607), .B1(P3_REG2_REG_31__SCAN_IN), 
        .B2(n13001), .ZN(n14606) );
  NAND2_X1 U16379 ( .A1(n14609), .A2(n14606), .ZN(P3_U3202) );
  AOI22_X1 U16380 ( .A1(n14615), .A2(n14607), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n13001), .ZN(n14608) );
  NAND2_X1 U16381 ( .A1(n14609), .A2(n14608), .ZN(P3_U3203) );
  OR2_X1 U16382 ( .A1(n14610), .A2(n15357), .ZN(n14612) );
  INV_X1 U16383 ( .A(n14614), .ZN(n14611) );
  INV_X1 U16384 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U16385 ( .A1(n15374), .A2(n14629), .B1(n14613), .B2(n15371), .ZN(
        P3_U3490) );
  AOI21_X1 U16386 ( .B1(n14615), .B2(n15325), .A(n14614), .ZN(n14631) );
  INV_X1 U16387 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14616) );
  AOI22_X1 U16388 ( .A1(n15374), .A2(n14631), .B1(n14616), .B2(n15371), .ZN(
        P3_U3489) );
  NOR2_X1 U16389 ( .A1(n14617), .A2(n15357), .ZN(n14619) );
  AOI211_X1 U16390 ( .C1(n15339), .C2(n14620), .A(n14619), .B(n14618), .ZN(
        n14633) );
  AOI22_X1 U16391 ( .A1(n15374), .A2(n14633), .B1(n14621), .B2(n15371), .ZN(
        P3_U3471) );
  OAI22_X1 U16392 ( .A1(n14624), .A2(n14623), .B1(n14622), .B2(n15357), .ZN(
        n14625) );
  NOR2_X1 U16393 ( .A1(n14626), .A2(n14625), .ZN(n14635) );
  INV_X1 U16394 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14627) );
  AOI22_X1 U16395 ( .A1(n15374), .A2(n14635), .B1(n14627), .B2(n15371), .ZN(
        P3_U3470) );
  INV_X1 U16396 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14628) );
  AOI22_X1 U16397 ( .A1(n15365), .A2(n14629), .B1(n14628), .B2(n15363), .ZN(
        P3_U3458) );
  INV_X1 U16398 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14630) );
  AOI22_X1 U16399 ( .A1(n15365), .A2(n14631), .B1(n14630), .B2(n15363), .ZN(
        P3_U3457) );
  INV_X1 U16400 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U16401 ( .A1(n15365), .A2(n14633), .B1(n14632), .B2(n15363), .ZN(
        P3_U3426) );
  INV_X1 U16402 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U16403 ( .A1(n15365), .A2(n14635), .B1(n14634), .B2(n15363), .ZN(
        P3_U3423) );
  OAI22_X1 U16404 ( .A1(n14637), .A2(n14921), .B1(n14920), .B2(n14636), .ZN(
        n14643) );
  AOI21_X1 U16405 ( .B1(n14640), .B2(n14638), .A(n14639), .ZN(n14641) );
  NOR2_X1 U16406 ( .A1(n14641), .A2(n14926), .ZN(n14642) );
  AOI211_X1 U16407 ( .C1(n14644), .C2(n14930), .A(n14643), .B(n14642), .ZN(
        n14646) );
  OAI211_X1 U16408 ( .C1(n14934), .C2(n14647), .A(n14646), .B(n14645), .ZN(
        P2_U3198) );
  XNOR2_X1 U16409 ( .A(n14649), .B(n14648), .ZN(n14651) );
  AOI21_X1 U16410 ( .B1(n14651), .B2(n9268), .A(n14650), .ZN(n14670) );
  INV_X1 U16411 ( .A(n14652), .ZN(n14653) );
  AOI222_X1 U16412 ( .A1(n14656), .A2(n14655), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14668), .C1(n14654), .C2(n14653), .ZN(n14667) );
  INV_X1 U16413 ( .A(n14657), .ZN(n14658) );
  AOI21_X1 U16414 ( .B1(n14660), .B2(n14659), .A(n14658), .ZN(n14673) );
  OAI211_X1 U16415 ( .C1(n6678), .C2(n6632), .A(n6483), .B(n14661), .ZN(n14669) );
  INV_X1 U16416 ( .A(n14669), .ZN(n14663) );
  AOI22_X1 U16417 ( .A1(n14673), .A2(n14665), .B1(n14664), .B2(n14663), .ZN(
        n14666) );
  OAI211_X1 U16418 ( .C1(n14668), .C2(n14670), .A(n14667), .B(n14666), .ZN(
        P2_U3251) );
  OAI21_X1 U16419 ( .B1(n6678), .B2(n15140), .A(n14669), .ZN(n14672) );
  INV_X1 U16420 ( .A(n14670), .ZN(n14671) );
  AOI211_X1 U16421 ( .C1(n14673), .C2(n15137), .A(n14672), .B(n14671), .ZN(
        n14681) );
  AOI22_X1 U16422 ( .A1(n15156), .A2(n14681), .B1(n13346), .B2(n15154), .ZN(
        P2_U3513) );
  INV_X1 U16423 ( .A(n14674), .ZN(n14679) );
  OAI21_X1 U16424 ( .B1(n14676), .B2(n15140), .A(n14675), .ZN(n14678) );
  AOI211_X1 U16425 ( .C1(n15135), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        n14682) );
  AOI22_X1 U16426 ( .A1(n15156), .A2(n14682), .B1(n14680), .B2(n15154), .ZN(
        P2_U3511) );
  AOI22_X1 U16427 ( .A1(n15147), .A2(n14681), .B1(n9036), .B2(n15145), .ZN(
        P2_U3472) );
  AOI22_X1 U16428 ( .A1(n15147), .A2(n14682), .B1(n9006), .B2(n15145), .ZN(
        P2_U3466) );
  NAND2_X1 U16429 ( .A1(n14684), .A2(n14683), .ZN(n14685) );
  NAND2_X1 U16430 ( .A1(n14686), .A2(n14685), .ZN(n14690) );
  AOI222_X1 U16431 ( .A1(n14692), .A2(n14691), .B1(n14690), .B2(n14689), .C1(
        n14688), .C2(n14687), .ZN(n14694) );
  OAI211_X1 U16432 ( .C1(n14696), .C2(n14695), .A(n14694), .B(n14693), .ZN(
        P1_U3215) );
  OAI22_X1 U16433 ( .A1(n14698), .A2(n10323), .B1(n14697), .B2(n14875), .ZN(
        n14699) );
  AOI21_X1 U16434 ( .B1(n14700), .B2(n14904), .A(n14699), .ZN(n14701) );
  AOI22_X1 U16435 ( .A1(n14916), .A2(n14722), .B1(n14799), .B2(n14917), .ZN(
        P1_U3543) );
  OAI22_X1 U16436 ( .A1(n14704), .A2(n10323), .B1(n14703), .B2(n14875), .ZN(
        n14707) );
  INV_X1 U16437 ( .A(n14705), .ZN(n14706) );
  AOI211_X1 U16438 ( .C1(n14708), .C2(n14904), .A(n14707), .B(n14706), .ZN(
        n14724) );
  AOI22_X1 U16439 ( .A1(n14916), .A2(n14724), .B1(n11773), .B2(n14917), .ZN(
        P1_U3542) );
  AND2_X1 U16440 ( .A1(n14709), .A2(n14904), .ZN(n14713) );
  OAI22_X1 U16441 ( .A1(n14711), .A2(n10323), .B1(n6816), .B2(n14875), .ZN(
        n14712) );
  NOR3_X1 U16442 ( .A1(n14714), .A2(n14713), .A3(n14712), .ZN(n14726) );
  AOI22_X1 U16443 ( .A1(n14916), .A2(n14726), .B1(n11127), .B2(n14917), .ZN(
        P1_U3541) );
  AND2_X1 U16444 ( .A1(n14715), .A2(n14904), .ZN(n14719) );
  OAI22_X1 U16445 ( .A1(n14717), .A2(n10323), .B1(n14716), .B2(n14875), .ZN(
        n14718) );
  NOR3_X1 U16446 ( .A1(n14720), .A2(n14719), .A3(n14718), .ZN(n14728) );
  AOI22_X1 U16447 ( .A1(n14916), .A2(n14728), .B1(n10755), .B2(n14917), .ZN(
        P1_U3539) );
  INV_X1 U16448 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14721) );
  AOI22_X1 U16449 ( .A1(n14504), .A2(n14722), .B1(n14721), .B2(n14905), .ZN(
        P1_U3504) );
  INV_X1 U16450 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U16451 ( .A1(n14504), .A2(n14724), .B1(n14723), .B2(n14905), .ZN(
        P1_U3501) );
  INV_X1 U16452 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14725) );
  AOI22_X1 U16453 ( .A1(n14504), .A2(n14726), .B1(n14725), .B2(n14905), .ZN(
        P1_U3498) );
  INV_X1 U16454 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U16455 ( .A1(n14504), .A2(n14728), .B1(n14727), .B2(n14905), .ZN(
        P1_U3492) );
  OAI21_X1 U16456 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(SUB_1596_U69) );
  OAI21_X1 U16457 ( .B1(n14733), .B2(n14997), .A(n14732), .ZN(SUB_1596_U68) );
  OAI21_X1 U16458 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n14737) );
  XNOR2_X1 U16459 ( .A(n14737), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16460 ( .B1(n14740), .B2(n14739), .A(n14738), .ZN(n14741) );
  XNOR2_X1 U16461 ( .A(n14741), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16462 ( .B1(n14744), .B2(n14743), .A(n14742), .ZN(n14745) );
  XOR2_X1 U16463 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14745), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16464 ( .A1(n14747), .A2(n14746), .ZN(n14748) );
  XOR2_X1 U16465 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14748), .Z(SUB_1596_U64)
         );
  NOR2_X1 U16466 ( .A1(n14749), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14751) );
  OR2_X1 U16467 ( .A1(n14750), .A2(n14751), .ZN(n14754) );
  INV_X1 U16468 ( .A(n14751), .ZN(n14753) );
  MUX2_X1 U16469 ( .A(n14754), .B(n14753), .S(n14752), .Z(n14756) );
  NAND2_X1 U16470 ( .A1(n14756), .A2(n14755), .ZN(n14759) );
  AOI22_X1 U16471 ( .A1(n14757), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14758) );
  OAI21_X1 U16472 ( .B1(n14760), .B2(n14759), .A(n14758), .ZN(P1_U3243) );
  NAND3_X1 U16473 ( .A1(n14763), .A2(n14762), .A3(n14761), .ZN(n14764) );
  NAND3_X1 U16474 ( .A1(n14801), .A2(n14765), .A3(n14764), .ZN(n14773) );
  MUX2_X1 U16475 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10606), .S(n14774), .Z(
        n14768) );
  NAND3_X1 U16476 ( .A1(n14768), .A2(n14767), .A3(n14766), .ZN(n14769) );
  NAND3_X1 U16477 ( .A1(n14771), .A2(n14770), .A3(n14769), .ZN(n14772) );
  OAI211_X1 U16478 ( .C1(n14775), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        n14776) );
  INV_X1 U16479 ( .A(n14776), .ZN(n14777) );
  AND2_X1 U16480 ( .A1(n14778), .A2(n14777), .ZN(n14780) );
  OAI211_X1 U16481 ( .C1(n14812), .C2(n8494), .A(n14780), .B(n14779), .ZN(
        P1_U3247) );
  INV_X1 U16482 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14795) );
  AOI21_X1 U16483 ( .B1(n14783), .B2(n14782), .A(n14781), .ZN(n14791) );
  OAI21_X1 U16484 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(n14787) );
  NAND2_X1 U16485 ( .A1(n14787), .A2(n14801), .ZN(n14790) );
  NAND2_X1 U16486 ( .A1(n14804), .A2(n14788), .ZN(n14789) );
  OAI211_X1 U16487 ( .C1(n14791), .C2(n14807), .A(n14790), .B(n14789), .ZN(
        n14792) );
  INV_X1 U16488 ( .A(n14792), .ZN(n14794) );
  OAI211_X1 U16489 ( .C1(n14795), .C2(n14812), .A(n14794), .B(n14793), .ZN(
        P1_U3255) );
  AOI21_X1 U16490 ( .B1(n14797), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14796), 
        .ZN(n14808) );
  OAI21_X1 U16491 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n14802) );
  NAND2_X1 U16492 ( .A1(n14802), .A2(n14801), .ZN(n14806) );
  NAND2_X1 U16493 ( .A1(n14804), .A2(n14803), .ZN(n14805) );
  OAI211_X1 U16494 ( .C1(n14808), .C2(n14807), .A(n14806), .B(n14805), .ZN(
        n14809) );
  INV_X1 U16495 ( .A(n14809), .ZN(n14811) );
  OAI211_X1 U16496 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        P1_U3258) );
  INV_X1 U16497 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14814) );
  NOR2_X1 U16498 ( .A1(n14844), .A2(n14814), .ZN(P1_U3294) );
  INV_X1 U16499 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14815) );
  NOR2_X1 U16500 ( .A1(n14844), .A2(n14815), .ZN(P1_U3295) );
  INV_X1 U16501 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14816) );
  NOR2_X1 U16502 ( .A1(n14844), .A2(n14816), .ZN(P1_U3296) );
  INV_X1 U16503 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14817) );
  NOR2_X1 U16504 ( .A1(n14844), .A2(n14817), .ZN(P1_U3297) );
  INV_X1 U16505 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14818) );
  NOR2_X1 U16506 ( .A1(n14844), .A2(n14818), .ZN(P1_U3298) );
  INV_X1 U16507 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14819) );
  NOR2_X1 U16508 ( .A1(n14844), .A2(n14819), .ZN(P1_U3299) );
  INV_X1 U16509 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14820) );
  NOR2_X1 U16510 ( .A1(n14844), .A2(n14820), .ZN(P1_U3300) );
  INV_X1 U16511 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14821) );
  NOR2_X1 U16512 ( .A1(n14844), .A2(n14821), .ZN(P1_U3301) );
  INV_X1 U16513 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14822) );
  NOR2_X1 U16514 ( .A1(n14844), .A2(n14822), .ZN(P1_U3302) );
  INV_X1 U16515 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14823) );
  NOR2_X1 U16516 ( .A1(n14844), .A2(n14823), .ZN(P1_U3303) );
  INV_X1 U16517 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14824) );
  NOR2_X1 U16518 ( .A1(n14844), .A2(n14824), .ZN(P1_U3304) );
  INV_X1 U16519 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14825) );
  NOR2_X1 U16520 ( .A1(n14844), .A2(n14825), .ZN(P1_U3305) );
  INV_X1 U16521 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14826) );
  NOR2_X1 U16522 ( .A1(n14844), .A2(n14826), .ZN(P1_U3306) );
  INV_X1 U16523 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14827) );
  NOR2_X1 U16524 ( .A1(n14844), .A2(n14827), .ZN(P1_U3307) );
  INV_X1 U16525 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14828) );
  NOR2_X1 U16526 ( .A1(n14844), .A2(n14828), .ZN(P1_U3308) );
  INV_X1 U16527 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14829) );
  NOR2_X1 U16528 ( .A1(n14844), .A2(n14829), .ZN(P1_U3309) );
  INV_X1 U16529 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14830) );
  NOR2_X1 U16530 ( .A1(n14844), .A2(n14830), .ZN(P1_U3310) );
  INV_X1 U16531 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14831) );
  NOR2_X1 U16532 ( .A1(n14844), .A2(n14831), .ZN(P1_U3311) );
  INV_X1 U16533 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14832) );
  NOR2_X1 U16534 ( .A1(n14844), .A2(n14832), .ZN(P1_U3312) );
  INV_X1 U16535 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14833) );
  NOR2_X1 U16536 ( .A1(n14844), .A2(n14833), .ZN(P1_U3313) );
  INV_X1 U16537 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14834) );
  NOR2_X1 U16538 ( .A1(n14844), .A2(n14834), .ZN(P1_U3314) );
  INV_X1 U16539 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14835) );
  NOR2_X1 U16540 ( .A1(n14844), .A2(n14835), .ZN(P1_U3315) );
  INV_X1 U16541 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14836) );
  NOR2_X1 U16542 ( .A1(n14844), .A2(n14836), .ZN(P1_U3316) );
  INV_X1 U16543 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14837) );
  NOR2_X1 U16544 ( .A1(n14844), .A2(n14837), .ZN(P1_U3317) );
  INV_X1 U16545 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14838) );
  NOR2_X1 U16546 ( .A1(n14844), .A2(n14838), .ZN(P1_U3318) );
  INV_X1 U16547 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14839) );
  NOR2_X1 U16548 ( .A1(n14844), .A2(n14839), .ZN(P1_U3319) );
  NOR2_X1 U16549 ( .A1(n14844), .A2(n14840), .ZN(P1_U3320) );
  NOR2_X1 U16550 ( .A1(n14844), .A2(n14841), .ZN(P1_U3321) );
  NOR2_X1 U16551 ( .A1(n14844), .A2(n14842), .ZN(P1_U3322) );
  NOR2_X1 U16552 ( .A1(n14844), .A2(n14843), .ZN(P1_U3323) );
  OAI22_X1 U16553 ( .A1(n14846), .A2(n10323), .B1(n14845), .B2(n14875), .ZN(
        n14848) );
  NOR2_X1 U16554 ( .A1(n14848), .A2(n14847), .ZN(n14907) );
  INV_X1 U16555 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14849) );
  AOI22_X1 U16556 ( .A1(n14504), .A2(n14907), .B1(n14849), .B2(n14905), .ZN(
        P1_U3465) );
  OAI22_X1 U16557 ( .A1(n14851), .A2(n10323), .B1(n14850), .B2(n14875), .ZN(
        n14853) );
  AOI211_X1 U16558 ( .C1(n14854), .C2(n14904), .A(n14853), .B(n14852), .ZN(
        n14908) );
  INV_X1 U16559 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U16560 ( .A1(n14504), .A2(n14908), .B1(n14855), .B2(n14905), .ZN(
        P1_U3471) );
  AOI211_X1 U16561 ( .C1(n14883), .C2(n14858), .A(n14857), .B(n14856), .ZN(
        n14859) );
  OAI21_X1 U16562 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n14862) );
  INV_X1 U16563 ( .A(n14862), .ZN(n14910) );
  INV_X1 U16564 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14863) );
  AOI22_X1 U16565 ( .A1(n14504), .A2(n14910), .B1(n14863), .B2(n14905), .ZN(
        P1_U3474) );
  AOI22_X1 U16566 ( .A1(n14865), .A2(n14883), .B1(n14882), .B2(n14864), .ZN(
        n14866) );
  OAI211_X1 U16567 ( .C1(n14888), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14869) );
  INV_X1 U16568 ( .A(n14869), .ZN(n14911) );
  INV_X1 U16569 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U16570 ( .A1(n14504), .A2(n14911), .B1(n14870), .B2(n14905), .ZN(
        P1_U3477) );
  INV_X1 U16571 ( .A(n14871), .ZN(n14878) );
  NAND2_X1 U16572 ( .A1(n14872), .A2(n14883), .ZN(n14873) );
  OAI211_X1 U16573 ( .C1(n14876), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        n14877) );
  AOI21_X1 U16574 ( .B1(n14879), .B2(n14878), .A(n14877), .ZN(n14912) );
  INV_X1 U16575 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14880) );
  AOI22_X1 U16576 ( .A1(n14504), .A2(n14912), .B1(n14880), .B2(n14905), .ZN(
        P1_U3480) );
  AOI22_X1 U16577 ( .A1(n14884), .A2(n14883), .B1(n14882), .B2(n14881), .ZN(
        n14885) );
  OAI211_X1 U16578 ( .C1(n14888), .C2(n14887), .A(n14886), .B(n14885), .ZN(
        n14889) );
  INV_X1 U16579 ( .A(n14889), .ZN(n14913) );
  INV_X1 U16580 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U16581 ( .A1(n14504), .A2(n14913), .B1(n14890), .B2(n14905), .ZN(
        P1_U3483) );
  AND2_X1 U16582 ( .A1(n14891), .A2(n14904), .ZN(n14895) );
  OAI21_X1 U16583 ( .B1(n14893), .B2(n10323), .A(n14892), .ZN(n14894) );
  NOR3_X1 U16584 ( .A1(n14896), .A2(n14895), .A3(n14894), .ZN(n14915) );
  INV_X1 U16585 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14897) );
  AOI22_X1 U16586 ( .A1(n14504), .A2(n14915), .B1(n14897), .B2(n14905), .ZN(
        P1_U3486) );
  INV_X1 U16587 ( .A(n14898), .ZN(n14903) );
  NAND3_X1 U16588 ( .A1(n14901), .A2(n14900), .A3(n14899), .ZN(n14902) );
  AOI21_X1 U16589 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n14918) );
  INV_X1 U16590 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14906) );
  AOI22_X1 U16591 ( .A1(n14504), .A2(n14918), .B1(n14906), .B2(n14905), .ZN(
        P1_U3489) );
  AOI22_X1 U16592 ( .A1(n14916), .A2(n14907), .B1(n10622), .B2(n14917), .ZN(
        P1_U3530) );
  AOI22_X1 U16593 ( .A1(n14916), .A2(n14908), .B1(n10624), .B2(n14917), .ZN(
        P1_U3532) );
  INV_X1 U16594 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14909) );
  AOI22_X1 U16595 ( .A1(n14916), .A2(n14910), .B1(n14909), .B2(n14917), .ZN(
        P1_U3533) );
  AOI22_X1 U16596 ( .A1(n14916), .A2(n14911), .B1(n10619), .B2(n14917), .ZN(
        P1_U3534) );
  AOI22_X1 U16597 ( .A1(n14916), .A2(n14912), .B1(n10651), .B2(n14917), .ZN(
        P1_U3535) );
  AOI22_X1 U16598 ( .A1(n14916), .A2(n14913), .B1(n10653), .B2(n14917), .ZN(
        P1_U3536) );
  INV_X1 U16599 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14914) );
  AOI22_X1 U16600 ( .A1(n14916), .A2(n14915), .B1(n14914), .B2(n14917), .ZN(
        P1_U3537) );
  AOI22_X1 U16601 ( .A1(n14916), .A2(n14918), .B1(n10754), .B2(n14917), .ZN(
        P1_U3538) );
  OAI22_X1 U16602 ( .A1(n14922), .A2(n14921), .B1(n14920), .B2(n14919), .ZN(
        n14929) );
  NAND2_X1 U16603 ( .A1(n14925), .A2(n14924), .ZN(n14927) );
  AOI21_X1 U16604 ( .B1(n14923), .B2(n14927), .A(n14926), .ZN(n14928) );
  AOI211_X1 U16605 ( .C1(n14931), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14932) );
  NAND2_X1 U16606 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14995)
         );
  OAI211_X1 U16607 ( .C1(n14934), .C2(n14933), .A(n14932), .B(n14995), .ZN(
        P2_U3196) );
  AOI22_X1 U16608 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15033), .B1(n15021), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14938) );
  AOI22_X1 U16609 ( .A1(n15051), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14937) );
  OAI22_X1 U16610 ( .A1(n15053), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n15042), .ZN(n14935) );
  OAI21_X1 U16611 ( .B1(n15027), .B2(n14935), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14936) );
  OAI211_X1 U16612 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14938), .A(n14937), .B(
        n14936), .ZN(P2_U3214) );
  OAI21_X1 U16613 ( .B1(n14941), .B2(n14940), .A(n14939), .ZN(n14947) );
  NOR2_X1 U16614 ( .A1(n14942), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14943) );
  AOI21_X1 U16615 ( .B1(n15027), .B2(n14944), .A(n14943), .ZN(n14946) );
  NAND2_X1 U16616 ( .A1(n15051), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n14945) );
  OAI211_X1 U16617 ( .C1(n15042), .C2(n14947), .A(n14946), .B(n14945), .ZN(
        n14948) );
  INV_X1 U16618 ( .A(n14948), .ZN(n14954) );
  AOI211_X1 U16619 ( .C1(n14951), .C2(n14950), .A(n14949), .B(n15053), .ZN(
        n14952) );
  INV_X1 U16620 ( .A(n14952), .ZN(n14953) );
  NAND2_X1 U16621 ( .A1(n14954), .A2(n14953), .ZN(P2_U3215) );
  AOI22_X1 U16622 ( .A1(n15051), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14968) );
  OAI21_X1 U16623 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14960) );
  NAND2_X1 U16624 ( .A1(n15027), .A2(n14958), .ZN(n14959) );
  OAI21_X1 U16625 ( .B1(n15042), .B2(n14960), .A(n14959), .ZN(n14961) );
  INV_X1 U16626 ( .A(n14961), .ZN(n14967) );
  NAND2_X1 U16627 ( .A1(n14963), .A2(n14962), .ZN(n14964) );
  NAND3_X1 U16628 ( .A1(n15033), .A2(n14965), .A3(n14964), .ZN(n14966) );
  NAND3_X1 U16629 ( .A1(n14968), .A2(n14967), .A3(n14966), .ZN(P2_U3216) );
  OAI21_X1 U16630 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n14972) );
  INV_X1 U16631 ( .A(n14972), .ZN(n14981) );
  AOI22_X1 U16632 ( .A1(n15051), .A2(P2_ADDR_REG_9__SCAN_IN), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(P2_U3088), .ZN(n14980) );
  NAND2_X1 U16633 ( .A1(n14974), .A2(n14973), .ZN(n14975) );
  AOI21_X1 U16634 ( .B1(n14976), .B2(n14975), .A(n15042), .ZN(n14977) );
  AOI21_X1 U16635 ( .B1(n15027), .B2(n14978), .A(n14977), .ZN(n14979) );
  OAI211_X1 U16636 ( .C1(n14981), .C2(n15053), .A(n14980), .B(n14979), .ZN(
        P2_U3223) );
  NAND2_X1 U16637 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  AOI21_X1 U16638 ( .B1(n14985), .B2(n14984), .A(n15042), .ZN(n14993) );
  INV_X1 U16639 ( .A(n14986), .ZN(n14991) );
  NAND3_X1 U16640 ( .A1(n14989), .A2(n14988), .A3(n14987), .ZN(n14990) );
  AOI21_X1 U16641 ( .B1(n14991), .B2(n14990), .A(n15053), .ZN(n14992) );
  AOI211_X1 U16642 ( .C1(n15027), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        n14996) );
  OAI211_X1 U16643 ( .C1(n14997), .C2(n15039), .A(n14996), .B(n14995), .ZN(
        P2_U3226) );
  AOI21_X1 U16644 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n14999), .A(n14998), 
        .ZN(n15009) );
  OAI21_X1 U16645 ( .B1(n15001), .B2(n15000), .A(n15021), .ZN(n15003) );
  NOR2_X1 U16646 ( .A1(n15003), .A2(n15002), .ZN(n15007) );
  OAI21_X1 U16647 ( .B1(n15048), .B2(n15005), .A(n15004), .ZN(n15006) );
  AOI211_X1 U16648 ( .C1(n15051), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n15007), 
        .B(n15006), .ZN(n15008) );
  OAI21_X1 U16649 ( .B1(n15009), .B2(n15053), .A(n15008), .ZN(P2_U3228) );
  AOI211_X1 U16650 ( .C1(n15012), .C2(n15011), .A(n15010), .B(n15042), .ZN(
        n15013) );
  AOI21_X1 U16651 ( .B1(n15051), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n15013), 
        .ZN(n15020) );
  OAI211_X1 U16652 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15015), .A(n15033), 
        .B(n15014), .ZN(n15018) );
  NAND2_X1 U16653 ( .A1(n15027), .A2(n15016), .ZN(n15017) );
  NAND4_X1 U16654 ( .A1(n15020), .A2(n15019), .A3(n15018), .A4(n15017), .ZN(
        P2_U3229) );
  OAI21_X1 U16655 ( .B1(n15023), .B2(n15022), .A(n15021), .ZN(n15030) );
  NOR2_X1 U16656 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15024), .ZN(n15025) );
  AOI21_X1 U16657 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15028) );
  OAI21_X1 U16658 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(n15031) );
  INV_X1 U16659 ( .A(n15031), .ZN(n15037) );
  OAI211_X1 U16660 ( .C1(n15035), .C2(n15034), .A(n15033), .B(n15032), .ZN(
        n15036) );
  OAI211_X1 U16661 ( .C1(n15039), .C2(n15038), .A(n15037), .B(n15036), .ZN(
        P2_U3231) );
  AOI21_X1 U16662 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n15041), .A(n15040), 
        .ZN(n15054) );
  AOI211_X1 U16663 ( .C1(n15045), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        n15050) );
  OAI21_X1 U16664 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(n15049) );
  AOI211_X1 U16665 ( .C1(n15051), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n15050), 
        .B(n15049), .ZN(n15052) );
  OAI21_X1 U16666 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(P2_U3232) );
  NOR2_X1 U16667 ( .A1(n15055), .A2(n15093), .ZN(n15083) );
  CLKBUF_X1 U16668 ( .A(n15083), .Z(n15087) );
  INV_X1 U16669 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15056) );
  NOR2_X1 U16670 ( .A1(n15087), .A2(n15056), .ZN(P2_U3266) );
  INV_X1 U16671 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15057) );
  NOR2_X1 U16672 ( .A1(n15087), .A2(n15057), .ZN(P2_U3267) );
  INV_X1 U16673 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15058) );
  NOR2_X1 U16674 ( .A1(n15087), .A2(n15058), .ZN(P2_U3268) );
  INV_X1 U16675 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15059) );
  NOR2_X1 U16676 ( .A1(n15083), .A2(n15059), .ZN(P2_U3269) );
  INV_X1 U16677 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15060) );
  NOR2_X1 U16678 ( .A1(n15083), .A2(n15060), .ZN(P2_U3270) );
  INV_X1 U16679 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15061) );
  NOR2_X1 U16680 ( .A1(n15083), .A2(n15061), .ZN(P2_U3271) );
  INV_X1 U16681 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15062) );
  NOR2_X1 U16682 ( .A1(n15083), .A2(n15062), .ZN(P2_U3272) );
  INV_X1 U16683 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15063) );
  NOR2_X1 U16684 ( .A1(n15083), .A2(n15063), .ZN(P2_U3273) );
  INV_X1 U16685 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15064) );
  NOR2_X1 U16686 ( .A1(n15083), .A2(n15064), .ZN(P2_U3274) );
  INV_X1 U16687 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15065) );
  NOR2_X1 U16688 ( .A1(n15083), .A2(n15065), .ZN(P2_U3275) );
  INV_X1 U16689 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15066) );
  NOR2_X1 U16690 ( .A1(n15083), .A2(n15066), .ZN(P2_U3276) );
  INV_X1 U16691 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15067) );
  NOR2_X1 U16692 ( .A1(n15083), .A2(n15067), .ZN(P2_U3277) );
  INV_X1 U16693 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15068) );
  NOR2_X1 U16694 ( .A1(n15087), .A2(n15068), .ZN(P2_U3278) );
  INV_X1 U16695 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15069) );
  NOR2_X1 U16696 ( .A1(n15087), .A2(n15069), .ZN(P2_U3279) );
  INV_X1 U16697 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15070) );
  NOR2_X1 U16698 ( .A1(n15087), .A2(n15070), .ZN(P2_U3280) );
  INV_X1 U16699 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15071) );
  NOR2_X1 U16700 ( .A1(n15087), .A2(n15071), .ZN(P2_U3281) );
  INV_X1 U16701 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U16702 ( .A1(n15087), .A2(n15072), .ZN(P2_U3282) );
  INV_X1 U16703 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15073) );
  NOR2_X1 U16704 ( .A1(n15087), .A2(n15073), .ZN(P2_U3283) );
  INV_X1 U16705 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15074) );
  NOR2_X1 U16706 ( .A1(n15087), .A2(n15074), .ZN(P2_U3284) );
  INV_X1 U16707 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15075) );
  NOR2_X1 U16708 ( .A1(n15087), .A2(n15075), .ZN(P2_U3285) );
  INV_X1 U16709 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15076) );
  NOR2_X1 U16710 ( .A1(n15087), .A2(n15076), .ZN(P2_U3286) );
  INV_X1 U16711 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15077) );
  NOR2_X1 U16712 ( .A1(n15087), .A2(n15077), .ZN(P2_U3287) );
  INV_X1 U16713 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15078) );
  NOR2_X1 U16714 ( .A1(n15087), .A2(n15078), .ZN(P2_U3288) );
  INV_X1 U16715 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15079) );
  NOR2_X1 U16716 ( .A1(n15087), .A2(n15079), .ZN(P2_U3289) );
  INV_X1 U16717 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15080) );
  NOR2_X1 U16718 ( .A1(n15083), .A2(n15080), .ZN(P2_U3290) );
  INV_X1 U16719 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15081) );
  NOR2_X1 U16720 ( .A1(n15087), .A2(n15081), .ZN(P2_U3291) );
  INV_X1 U16721 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15082) );
  NOR2_X1 U16722 ( .A1(n15083), .A2(n15082), .ZN(P2_U3292) );
  INV_X1 U16723 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15084) );
  NOR2_X1 U16724 ( .A1(n15087), .A2(n15084), .ZN(P2_U3293) );
  INV_X1 U16725 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15085) );
  NOR2_X1 U16726 ( .A1(n15087), .A2(n15085), .ZN(P2_U3294) );
  INV_X1 U16727 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15086) );
  NOR2_X1 U16728 ( .A1(n15087), .A2(n15086), .ZN(P2_U3295) );
  AOI22_X1 U16729 ( .A1(n15090), .A2(n15089), .B1(n15088), .B2(n15093), .ZN(
        P2_U3416) );
  AOI21_X1 U16730 ( .B1(n15093), .B2(n15092), .A(n15091), .ZN(P2_U3417) );
  INV_X1 U16731 ( .A(n15094), .ZN(n15097) );
  AOI211_X1 U16732 ( .C1(n15097), .C2(n15135), .A(n15096), .B(n15095), .ZN(
        n15148) );
  AOI22_X1 U16733 ( .A1(n15147), .A2(n15148), .B1(n8838), .B2(n15145), .ZN(
        P2_U3430) );
  INV_X1 U16734 ( .A(n15102), .ZN(n15105) );
  INV_X1 U16735 ( .A(n15098), .ZN(n15104) );
  AOI21_X1 U16736 ( .B1(n15100), .B2(n10663), .A(n15099), .ZN(n15101) );
  OAI21_X1 U16737 ( .B1(n15102), .B2(n15123), .A(n15101), .ZN(n15103) );
  AOI211_X1 U16738 ( .C1(n15106), .C2(n15105), .A(n15104), .B(n15103), .ZN(
        n15149) );
  AOI22_X1 U16739 ( .A1(n15147), .A2(n15149), .B1(n8826), .B2(n15145), .ZN(
        P2_U3433) );
  AOI22_X1 U16740 ( .A1(n15147), .A2(n15107), .B1(n8855), .B2(n15145), .ZN(
        P2_U3436) );
  AOI21_X1 U16741 ( .B1(n9219), .B2(n15123), .A(n15108), .ZN(n15112) );
  OAI211_X1 U16742 ( .C1(n6921), .C2(n15140), .A(n15110), .B(n15109), .ZN(
        n15111) );
  NOR2_X1 U16743 ( .A1(n15112), .A2(n15111), .ZN(n15150) );
  INV_X1 U16744 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U16745 ( .A1(n15147), .A2(n15150), .B1(n15113), .B2(n15145), .ZN(
        P2_U3439) );
  AOI21_X1 U16746 ( .B1(n9219), .B2(n15123), .A(n15114), .ZN(n15120) );
  INV_X1 U16747 ( .A(n15115), .ZN(n15116) );
  OAI211_X1 U16748 ( .C1(n15118), .C2(n15140), .A(n15117), .B(n15116), .ZN(
        n15119) );
  NOR2_X1 U16749 ( .A1(n15120), .A2(n15119), .ZN(n15151) );
  INV_X1 U16750 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U16751 ( .A1(n15147), .A2(n15151), .B1(n15121), .B2(n15145), .ZN(
        P2_U3442) );
  AOI21_X1 U16752 ( .B1(n9219), .B2(n15123), .A(n15122), .ZN(n15129) );
  INV_X1 U16753 ( .A(n15124), .ZN(n15125) );
  OAI211_X1 U16754 ( .C1(n15127), .C2(n15140), .A(n15126), .B(n15125), .ZN(
        n15128) );
  NOR2_X1 U16755 ( .A1(n15129), .A2(n15128), .ZN(n15152) );
  AOI22_X1 U16756 ( .A1(n15147), .A2(n15152), .B1(n8905), .B2(n15145), .ZN(
        P2_U3445) );
  OAI21_X1 U16757 ( .B1(n15131), .B2(n15140), .A(n15130), .ZN(n15133) );
  AOI211_X1 U16758 ( .C1(n15135), .C2(n15134), .A(n15133), .B(n15132), .ZN(
        n15153) );
  INV_X1 U16759 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U16760 ( .A1(n15147), .A2(n15153), .B1(n15136), .B2(n15145), .ZN(
        P2_U3454) );
  AND2_X1 U16761 ( .A1(n15138), .A2(n15137), .ZN(n15144) );
  OAI21_X1 U16762 ( .B1(n15141), .B2(n15140), .A(n15139), .ZN(n15142) );
  NOR3_X1 U16763 ( .A1(n15144), .A2(n15143), .A3(n15142), .ZN(n15155) );
  INV_X1 U16764 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U16765 ( .A1(n15147), .A2(n15155), .B1(n15146), .B2(n15145), .ZN(
        P2_U3460) );
  AOI22_X1 U16766 ( .A1(n15156), .A2(n15148), .B1(n8845), .B2(n15154), .ZN(
        P2_U3499) );
  AOI22_X1 U16767 ( .A1(n15156), .A2(n15149), .B1(n10460), .B2(n15154), .ZN(
        P2_U3500) );
  AOI22_X1 U16768 ( .A1(n15156), .A2(n15150), .B1(n10464), .B2(n15154), .ZN(
        P2_U3502) );
  AOI22_X1 U16769 ( .A1(n15156), .A2(n15151), .B1(n10466), .B2(n15154), .ZN(
        P2_U3503) );
  AOI22_X1 U16770 ( .A1(n15156), .A2(n15152), .B1(n10468), .B2(n15154), .ZN(
        P2_U3504) );
  AOI22_X1 U16771 ( .A1(n15156), .A2(n15153), .B1(n8945), .B2(n15154), .ZN(
        P2_U3507) );
  AOI22_X1 U16772 ( .A1(n15156), .A2(n15155), .B1(n10527), .B2(n15154), .ZN(
        P2_U3509) );
  NOR2_X1 U16773 ( .A1(P3_U3897), .A2(n15245), .ZN(P3_U3150) );
  OAI211_X1 U16774 ( .C1(n15159), .C2(n15158), .A(n15157), .B(n15180), .ZN(
        n15164) );
  NOR2_X1 U16775 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15160), .ZN(n15161) );
  AOI21_X1 U16776 ( .B1(n15186), .B2(n15162), .A(n15161), .ZN(n15163) );
  OAI211_X1 U16777 ( .C1(n15165), .C2(n15189), .A(n15164), .B(n15163), .ZN(
        n15166) );
  INV_X1 U16778 ( .A(n15166), .ZN(n15167) );
  OAI21_X1 U16779 ( .B1(n15168), .B2(n15193), .A(n15167), .ZN(P3_U3153) );
  OAI22_X1 U16780 ( .A1(n15170), .A2(n15169), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15203), .ZN(n15176) );
  AOI211_X1 U16781 ( .C1(n15174), .C2(n15173), .A(n15172), .B(n15171), .ZN(
        n15175) );
  AOI211_X1 U16782 ( .C1(n15178), .C2(n15177), .A(n15176), .B(n15175), .ZN(
        n15179) );
  OAI21_X1 U16783 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15193), .A(n15179), .ZN(
        P3_U3158) );
  OAI211_X1 U16784 ( .C1(n15183), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15188) );
  AOI21_X1 U16785 ( .B1(n15186), .B2(n15185), .A(n15184), .ZN(n15187) );
  OAI211_X1 U16786 ( .C1(n15190), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15191) );
  INV_X1 U16787 ( .A(n15191), .ZN(n15192) );
  OAI21_X1 U16788 ( .B1(n15194), .B2(n15193), .A(n15192), .ZN(P3_U3179) );
  AOI21_X1 U16789 ( .B1(n10919), .B2(n15196), .A(n15195), .ZN(n15213) );
  INV_X1 U16790 ( .A(n15197), .ZN(n15198) );
  NAND3_X1 U16791 ( .A1(n15200), .A2(n15199), .A3(n15198), .ZN(n15201) );
  AOI21_X1 U16792 ( .B1(n15202), .B2(n15201), .A(n15241), .ZN(n15208) );
  NOR2_X1 U16793 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15203), .ZN(n15204) );
  AOI21_X1 U16794 ( .B1(n15245), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n15204), .ZN(
        n15205) );
  OAI21_X1 U16795 ( .B1(n15285), .B2(n15206), .A(n15205), .ZN(n15207) );
  NOR2_X1 U16796 ( .A1(n15208), .A2(n15207), .ZN(n15212) );
  XNOR2_X1 U16797 ( .A(n15209), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U16798 ( .A1(n15287), .A2(n15210), .ZN(n15211) );
  OAI211_X1 U16799 ( .C1(n15213), .C2(n15291), .A(n15212), .B(n15211), .ZN(
        P3_U3185) );
  AOI21_X1 U16800 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15232) );
  OAI21_X1 U16801 ( .B1(n15219), .B2(n15218), .A(n15217), .ZN(n15225) );
  NOR2_X1 U16802 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15220), .ZN(n15221) );
  AOI21_X1 U16803 ( .B1(n15245), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n15221), .ZN(
        n15222) );
  OAI21_X1 U16804 ( .B1(n15285), .B2(n15223), .A(n15222), .ZN(n15224) );
  AOI21_X1 U16805 ( .B1(n15225), .B2(n15280), .A(n15224), .ZN(n15231) );
  AOI21_X1 U16806 ( .B1(n15228), .B2(n15227), .A(n15226), .ZN(n15229) );
  OR2_X1 U16807 ( .A1(n15257), .A2(n15229), .ZN(n15230) );
  OAI211_X1 U16808 ( .C1(n15232), .C2(n15291), .A(n15231), .B(n15230), .ZN(
        P3_U3186) );
  AOI21_X1 U16809 ( .B1(n15235), .B2(n15234), .A(n15233), .ZN(n15251) );
  AND2_X1 U16810 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n15244) );
  NAND2_X1 U16811 ( .A1(n15237), .A2(n15236), .ZN(n15238) );
  XNOR2_X1 U16812 ( .A(n15239), .B(n15238), .ZN(n15242) );
  OAI22_X1 U16813 ( .A1(n15242), .A2(n15241), .B1(n15240), .B2(n15285), .ZN(
        n15243) );
  AOI211_X1 U16814 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15245), .A(n15244), .B(
        n15243), .ZN(n15250) );
  OAI21_X1 U16815 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15247), .A(n15246), .ZN(
        n15248) );
  NAND2_X1 U16816 ( .A1(n15287), .A2(n15248), .ZN(n15249) );
  OAI211_X1 U16817 ( .C1(n15251), .C2(n15291), .A(n15250), .B(n15249), .ZN(
        P3_U3187) );
  XNOR2_X1 U16818 ( .A(n15253), .B(n15252), .ZN(n15265) );
  XOR2_X1 U16819 ( .A(n15255), .B(n15254), .Z(n15258) );
  OAI22_X1 U16820 ( .A1(n15258), .A2(n15257), .B1(n15256), .B2(n15285), .ZN(
        n15264) );
  NAND2_X1 U16821 ( .A1(n15260), .A2(n15259), .ZN(n15261) );
  AOI21_X1 U16822 ( .B1(n15262), .B2(n15261), .A(n15291), .ZN(n15263) );
  AOI211_X1 U16823 ( .C1(n15265), .C2(n15280), .A(n15264), .B(n15263), .ZN(
        n15267) );
  OAI211_X1 U16824 ( .C1(n15268), .C2(n15296), .A(n15267), .B(n15266), .ZN(
        P3_U3190) );
  AOI21_X1 U16825 ( .B1(n15271), .B2(n15270), .A(n15269), .ZN(n15292) );
  INV_X1 U16826 ( .A(n15272), .ZN(n15273) );
  NOR2_X1 U16827 ( .A1(n15273), .A2(n15274), .ZN(n15279) );
  INV_X1 U16828 ( .A(n15274), .ZN(n15275) );
  NAND2_X1 U16829 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  OAI21_X1 U16830 ( .B1(n15279), .B2(n15278), .A(n15277), .ZN(n15281) );
  NAND2_X1 U16831 ( .A1(n15281), .A2(n15280), .ZN(n15290) );
  OAI21_X1 U16832 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15283), .A(n15282), .ZN(
        n15288) );
  NOR2_X1 U16833 ( .A1(n15285), .A2(n15284), .ZN(n15286) );
  AOI21_X1 U16834 ( .B1(n15288), .B2(n15287), .A(n15286), .ZN(n15289) );
  OAI211_X1 U16835 ( .C1(n15292), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15293) );
  INV_X1 U16836 ( .A(n15293), .ZN(n15295) );
  NAND2_X1 U16837 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15294) );
  OAI211_X1 U16838 ( .C1(n15297), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        P3_U3191) );
  XNOR2_X1 U16839 ( .A(n15298), .B(n15300), .ZN(n15307) );
  OAI21_X1 U16840 ( .B1(n15301), .B2(n15300), .A(n15299), .ZN(n15343) );
  OAI22_X1 U16841 ( .A1(n15304), .A2(n15303), .B1(n10211), .B2(n15302), .ZN(
        n15305) );
  AOI21_X1 U16842 ( .B1(n15343), .B2(n15324), .A(n15305), .ZN(n15306) );
  OAI21_X1 U16843 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15341) );
  INV_X1 U16844 ( .A(n15343), .ZN(n15313) );
  NOR2_X1 U16845 ( .A1(n15309), .A2(n15357), .ZN(n15342) );
  INV_X1 U16846 ( .A(n15342), .ZN(n15310) );
  OAI22_X1 U16847 ( .A1(n15313), .A2(n15312), .B1(n15311), .B2(n15310), .ZN(
        n15314) );
  AOI211_X1 U16848 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15331), .A(n15341), .B(
        n15314), .ZN(n15315) );
  AOI22_X1 U16849 ( .A1(n13001), .A2(n10960), .B1(n15315), .B2(n15334), .ZN(
        P3_U3231) );
  XNOR2_X1 U16850 ( .A(n15316), .B(n15323), .ZN(n15318) );
  NAND2_X1 U16851 ( .A1(n15318), .A2(n15317), .ZN(n15321) );
  INV_X1 U16852 ( .A(n15319), .ZN(n15320) );
  NAND2_X1 U16853 ( .A1(n15321), .A2(n15320), .ZN(n15336) );
  INV_X1 U16854 ( .A(n15336), .ZN(n15330) );
  XNOR2_X1 U16855 ( .A(n15322), .B(n15323), .ZN(n15338) );
  NAND2_X1 U16856 ( .A1(n15338), .A2(n15324), .ZN(n15329) );
  AND2_X1 U16857 ( .A1(n15326), .A2(n15325), .ZN(n15337) );
  NAND2_X1 U16858 ( .A1(n15337), .A2(n15327), .ZN(n15328) );
  AND3_X1 U16859 ( .A1(n15330), .A2(n15329), .A3(n15328), .ZN(n15335) );
  AOI22_X1 U16860 ( .A1(n15338), .A2(n15332), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15331), .ZN(n15333) );
  OAI221_X1 U16861 ( .B1(n13001), .B2(n15335), .C1(n15334), .C2(n10909), .A(
        n15333), .ZN(P3_U3232) );
  AOI211_X1 U16862 ( .C1(n15339), .C2(n15338), .A(n15337), .B(n15336), .ZN(
        n15366) );
  INV_X1 U16863 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15340) );
  AOI22_X1 U16864 ( .A1(n15365), .A2(n15366), .B1(n15340), .B2(n15363), .ZN(
        P3_U3393) );
  AOI211_X1 U16865 ( .C1(n15355), .C2(n15343), .A(n15342), .B(n15341), .ZN(
        n15367) );
  INV_X1 U16866 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15344) );
  AOI22_X1 U16867 ( .A1(n15365), .A2(n15367), .B1(n15344), .B2(n15363), .ZN(
        P3_U3396) );
  INV_X1 U16868 ( .A(n15345), .ZN(n15349) );
  INV_X1 U16869 ( .A(n15346), .ZN(n15348) );
  AOI211_X1 U16870 ( .C1(n15349), .C2(n15355), .A(n15348), .B(n15347), .ZN(
        n15368) );
  INV_X1 U16871 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15350) );
  AOI22_X1 U16872 ( .A1(n15365), .A2(n15368), .B1(n15350), .B2(n15363), .ZN(
        P3_U3408) );
  NOR2_X1 U16873 ( .A1(n15351), .A2(n15357), .ZN(n15353) );
  AOI211_X1 U16874 ( .C1(n15355), .C2(n15354), .A(n15353), .B(n15352), .ZN(
        n15370) );
  INV_X1 U16875 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15356) );
  AOI22_X1 U16876 ( .A1(n15365), .A2(n15370), .B1(n15356), .B2(n15363), .ZN(
        P3_U3414) );
  OAI22_X1 U16877 ( .A1(n15360), .A2(n15359), .B1(n15358), .B2(n15357), .ZN(
        n15361) );
  NOR2_X1 U16878 ( .A1(n15362), .A2(n15361), .ZN(n15373) );
  INV_X1 U16879 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U16880 ( .A1(n15365), .A2(n15373), .B1(n15364), .B2(n15363), .ZN(
        P3_U3417) );
  AOI22_X1 U16881 ( .A1(n15374), .A2(n15366), .B1(n10908), .B2(n15371), .ZN(
        P3_U3460) );
  AOI22_X1 U16882 ( .A1(n15374), .A2(n15367), .B1(n10945), .B2(n15371), .ZN(
        P3_U3461) );
  AOI22_X1 U16883 ( .A1(n15374), .A2(n15368), .B1(n10942), .B2(n15371), .ZN(
        P3_U3465) );
  INV_X1 U16884 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U16885 ( .A1(n15374), .A2(n15370), .B1(n15369), .B2(n15371), .ZN(
        P3_U3467) );
  INV_X1 U16886 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U16887 ( .A1(n15374), .A2(n15373), .B1(n15372), .B2(n15371), .ZN(
        P3_U3468) );
  AOI21_X1 U16888 ( .B1(n15377), .B2(n15376), .A(n15375), .ZN(SUB_1596_U59) );
  OAI21_X1 U16889 ( .B1(n15380), .B2(n15379), .A(n15378), .ZN(SUB_1596_U58) );
  XOR2_X1 U16890 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15381), .Z(SUB_1596_U53) );
  AOI21_X1 U16891 ( .B1(n15384), .B2(n15383), .A(n15382), .ZN(SUB_1596_U56) );
  AOI21_X1 U16892 ( .B1(n15387), .B2(n15386), .A(n15385), .ZN(n15388) );
  XOR2_X1 U16893 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15388), .Z(SUB_1596_U60) );
  AOI21_X1 U16894 ( .B1(n15391), .B2(n15390), .A(n15389), .ZN(SUB_1596_U5) );
  NAND4_X1 U10127 ( .A1(n7845), .A2(n7844), .A3(n7843), .A4(n7842), .ZN(n8100)
         );
  CLKBUF_X1 U7221 ( .A(n8787), .Z(n8998) );
  NAND2_X1 U7263 ( .A1(n13211), .A2(n12540), .ZN(n12541) );
  CLKBUF_X1 U7272 ( .A(n13433), .Z(n9190) );
  CLKBUF_X1 U7278 ( .A(n8869), .Z(n9451) );
  AND2_X1 U7291 ( .A1(n13172), .A2(n6603), .ZN(n15400) );
  AND2_X1 U7347 ( .A1(n14323), .A2(n8129), .ZN(n15401) );
endmodule

