

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129;

  OR2_X1 U3546 ( .A1(n5158), .A2(n5157), .ZN(n5612) );
  OR2_X1 U3547 ( .A1(n5090), .A2(n3298), .ZN(n5080) );
  AND2_X1 U3548 ( .A1(n5114), .A2(n4051), .ZN(n5100) );
  AND2_X1 U3549 ( .A1(n5196), .A2(n3149), .ZN(n5114) );
  CLKBUF_X2 U3550 ( .A(n4437), .Z(n4553) );
  OR2_X1 U3551 ( .A1(n6793), .A2(n6698), .ZN(n5718) );
  INV_X1 U3552 ( .A(n4855), .ZN(n3177) );
  INV_X1 U3553 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6956) );
  CLKBUF_X2 U3554 ( .A(n3448), .Z(n3117) );
  AND3_X1 U3555 ( .A1(n3515), .A2(n4585), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4174) );
  OR2_X1 U3556 ( .A1(n4442), .A2(n4325), .ZN(n4332) );
  CLKBUF_X2 U3557 ( .A(n3437), .Z(n5970) );
  INV_X1 U3558 ( .A(n3463), .ZN(n4941) );
  BUF_X2 U3559 ( .A(n4331), .Z(n4585) );
  NAND2_X1 U3560 ( .A1(n3182), .A2(n4932), .ZN(n4334) );
  NAND4_X2 U3561 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3434)
         );
  AND2_X1 U3562 ( .A1(n5025), .A2(n4682), .ZN(n3437) );
  AND2_X1 U3563 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4682) );
  CLKBUF_X2 U3564 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n3112) );
  INV_X1 U3565 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3339) );
  NAND2_X2 U3566 ( .A1(n3186), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3250) );
  XNOR2_X1 U3567 ( .A(n3648), .B(n3649), .ZN(n4215) );
  AND2_X1 U3568 ( .A1(n4682), .A2(n5046), .ZN(n3611) );
  AND2_X1 U3569 ( .A1(n3344), .A2(n5025), .ZN(n3439) );
  OR2_X1 U3570 ( .A1(n3546), .A2(n3545), .ZN(n4276) );
  INV_X1 U3571 ( .A(n4349), .ZN(n3119) );
  XNOR2_X1 U3572 ( .A(n3517), .B(n3516), .ZN(n3649) );
  NAND2_X2 U3573 ( .A1(n4941), .A2(n4585), .ZN(n4343) );
  NAND2_X1 U3574 ( .A1(n4873), .A2(n4249), .ZN(n6523) );
  NAND2_X1 U3576 ( .A1(n3698), .A2(n3697), .ZN(n5346) );
  OR2_X1 U3578 ( .A1(n6693), .A2(n6262), .ZN(n6329) );
  INV_X1 U3579 ( .A(n5415), .ZN(n6473) );
  AND2_X1 U3580 ( .A1(n4993), .A2(n4821), .ZN(n6605) );
  NOR2_X1 U3581 ( .A1(n6175), .A2(n6292), .ZN(n6680) );
  AOI211_X1 U3582 ( .C1(n5725), .C2(n5586), .A(n5585), .B(n5584), .ZN(n5587)
         );
  INV_X2 U3583 ( .A(n4338), .ZN(n4349) );
  AND2_X1 U3584 ( .A1(n4299), .A2(n4298), .ZN(n3098) );
  NAND2_X1 U3585 ( .A1(n3804), .A2(n3803), .ZN(n5265) );
  AND4_X2 U3586 ( .A1(n3339), .A2(n3282), .A3(INSTQUEUERD_ADDR_REG_0__SCAN_IN), 
        .A4(n3112), .ZN(n3099) );
  OAI21_X2 U3588 ( .B1(n5737), .B2(n3258), .A(n5729), .ZN(n3257) );
  XNOR2_X1 U3589 ( .A(n4248), .B(n4352), .ZN(n4870) );
  NOR2_X2 U3590 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  NAND2_X2 U3591 ( .A1(n5627), .A2(n5626), .ZN(n5625) );
  NAND2_X2 U3592 ( .A1(n3381), .A2(n3380), .ZN(n3460) );
  XNOR2_X2 U3593 ( .A(n3690), .B(n3630), .ZN(n4200) );
  AND2_X4 U3594 ( .A1(n3337), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5960)
         );
  CLKBUF_X2 U3596 ( .A(n3505), .Z(n4119) );
  CLKBUF_X2 U3597 ( .A(n3426), .Z(n4120) );
  BUF_X2 U3598 ( .A(n3575), .Z(n3519) );
  BUF_X2 U3599 ( .A(n3611), .Z(n4099) );
  CLKBUF_X2 U3600 ( .A(n3438), .Z(n4118) );
  NOR2_X4 U3601 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4683) );
  OAI211_X1 U3602 ( .C1(n3213), .C2(n3218), .A(n3211), .B(n3210), .ZN(n5778)
         );
  NAND2_X1 U3603 ( .A1(n3212), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3211) );
  XNOR2_X1 U3604 ( .A(n3264), .B(n4514), .ZN(n4540) );
  XNOR2_X1 U3605 ( .A(n3184), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4502)
         );
  NAND2_X1 U3606 ( .A1(n3261), .A2(n3260), .ZN(n3264) );
  AOI21_X1 U3607 ( .B1(n5013), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5012), 
        .ZN(n5014) );
  NOR2_X1 U3608 ( .A1(n5519), .A2(n5718), .ZN(n4537) );
  OR2_X1 U3609 ( .A1(n4533), .A2(n4532), .ZN(n5519) );
  NAND2_X1 U3610 ( .A1(n5102), .A2(n5090), .ZN(n5583) );
  AND2_X1 U3611 ( .A1(n5777), .A2(n5776), .ZN(n3217) );
  CLKBUF_X1 U3612 ( .A(n5114), .Z(n5115) );
  NAND2_X1 U3613 ( .A1(n4552), .A2(n4375), .ZN(n4559) );
  INV_X1 U3614 ( .A(n5265), .ZN(n3178) );
  AND2_X1 U3615 ( .A1(n4437), .A2(n5072), .ZN(n4555) );
  AND2_X1 U3616 ( .A1(n3319), .A2(n4283), .ZN(n3318) );
  NOR2_X1 U3617 ( .A1(n3258), .A2(n3259), .ZN(n3255) );
  NOR2_X1 U3618 ( .A1(n3176), .A2(n4856), .ZN(n3175) );
  AND2_X1 U3619 ( .A1(n6512), .A2(n4214), .ZN(n4260) );
  AND2_X1 U3620 ( .A1(n4240), .A2(n4239), .ZN(n4872) );
  AND2_X1 U3621 ( .A1(n5001), .A2(n3335), .ZN(n3739) );
  NAND2_X1 U3622 ( .A1(n3169), .A2(n4268), .ZN(n4269) );
  NAND2_X1 U3623 ( .A1(n3706), .A2(n3705), .ZN(n5001) );
  NAND2_X1 U3624 ( .A1(n4805), .A2(n3674), .ZN(n4864) );
  NAND2_X1 U3625 ( .A1(n4807), .A2(n4806), .ZN(n4805) );
  NAND3_X1 U3626 ( .A1(n3619), .A2(n3126), .A3(n3630), .ZN(n4271) );
  NAND2_X1 U3627 ( .A1(n3654), .A2(n3653), .ZN(n4807) );
  INV_X2 U3628 ( .A(n6097), .ZN(n4909) );
  NAND2_X1 U3629 ( .A1(n3514), .A2(n3513), .ZN(n3517) );
  NAND2_X1 U3630 ( .A1(n3600), .A2(n3599), .ZN(n4751) );
  CLKBUF_X1 U3631 ( .A(n3662), .Z(n6695) );
  NAND2_X1 U3632 ( .A1(n4995), .A2(n3333), .ZN(n5355) );
  NAND2_X1 U3633 ( .A1(n3230), .A2(n4188), .ZN(n5065) );
  NAND4_X1 U3634 ( .A1(n3249), .A2(n3148), .A3(n3250), .A4(n3247), .ZN(n3495)
         );
  OR2_X1 U3635 ( .A1(n4861), .A2(n3307), .ZN(n3306) );
  OR2_X1 U3636 ( .A1(n4463), .A2(n3484), .ZN(n4459) );
  NOR2_X1 U3637 ( .A1(n5337), .A2(n5357), .ZN(n3310) );
  AND2_X1 U3638 ( .A1(n3562), .A2(n3657), .ZN(n3563) );
  AND2_X1 U3639 ( .A1(n3489), .A2(n3167), .ZN(n3166) );
  BUF_X2 U3640 ( .A(n4348), .Z(n4427) );
  AND2_X1 U3641 ( .A1(n3486), .A2(n4932), .ZN(n3464) );
  NAND2_X1 U3642 ( .A1(n3547), .A2(n4201), .ZN(n3513) );
  NOR2_X1 U3643 ( .A1(n4272), .A2(n3515), .ZN(n4463) );
  NAND2_X1 U3644 ( .A1(n3574), .A2(n3573), .ZN(n4187) );
  AND2_X2 U3645 ( .A1(n4932), .A2(n4331), .ZN(n3487) );
  AND3_X1 U3646 ( .A1(n3182), .A2(n3478), .A3(n4941), .ZN(n4450) );
  INV_X1 U3647 ( .A(n4306), .ZN(n4272) );
  NAND2_X1 U3648 ( .A1(n3558), .A2(n3455), .ZN(n4192) );
  AND2_X2 U3649 ( .A1(n3434), .A2(n4223), .ZN(n4306) );
  OR2_X1 U3650 ( .A1(n3557), .A2(n3556), .ZN(n4228) );
  AND2_X2 U3651 ( .A1(n4331), .A2(n3434), .ZN(n4809) );
  INV_X1 U3652 ( .A(n3434), .ZN(n4932) );
  BUF_X2 U3653 ( .A(n3460), .Z(n3515) );
  CLKBUF_X2 U3654 ( .A(n3458), .Z(n3635) );
  NAND4_X2 U3655 ( .A1(n3421), .A2(n3420), .A3(n3419), .A4(n3418), .ZN(n4331)
         );
  CLKBUF_X1 U3656 ( .A(n3477), .Z(n3478) );
  CLKBUF_X1 U3657 ( .A(n3455), .Z(n4223) );
  AND4_X1 U3658 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n3420)
         );
  AND4_X1 U3659 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3400)
         );
  NAND3_X1 U3660 ( .A1(n3453), .A2(n3332), .A3(n3452), .ZN(n3477) );
  AND4_X1 U3661 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3432)
         );
  AND4_X1 U3662 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3381)
         );
  AND4_X1 U3663 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3431)
         );
  AND4_X1 U3664 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3371)
         );
  AND4_X1 U3665 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(n3399)
         );
  AND4_X1 U3666 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3357)
         );
  AND4_X1 U3667 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3453)
         );
  AND4_X1 U3668 ( .A1(n3413), .A2(n3412), .A3(n3411), .A4(n3410), .ZN(n3419)
         );
  AND4_X1 U3669 ( .A1(n3385), .A2(n3384), .A3(n3383), .A4(n3382), .ZN(n3401)
         );
  AND4_X1 U3670 ( .A1(n3416), .A2(n3417), .A3(n3415), .A4(n3414), .ZN(n3418)
         );
  AND4_X1 U3671 ( .A1(n3342), .A2(n3343), .A3(n3341), .A4(n3340), .ZN(n3136)
         );
  AND4_X1 U3672 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3398)
         );
  AND4_X1 U3673 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3421)
         );
  AND4_X1 U3674 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3380)
         );
  BUF_X2 U3675 ( .A(n3099), .Z(n4094) );
  BUF_X2 U3676 ( .A(n3445), .Z(n4117) );
  AND2_X2 U3677 ( .A1(n5046), .A2(n3344), .ZN(n3121) );
  AND2_X2 U3678 ( .A1(n5050), .A2(n5961), .ZN(n3436) );
  AND2_X2 U3679 ( .A1(n3338), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5050)
         );
  NOR2_X2 U3680 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6691) );
  INV_X2 U3681 ( .A(n4089), .ZN(n3100) );
  INV_X1 U3682 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3337) );
  OR2_X2 U3683 ( .A1(n5633), .A2(n3151), .ZN(n3101) );
  OR2_X1 U3684 ( .A1(n5633), .A2(n3151), .ZN(n4297) );
  NOR2_X4 U3685 ( .A1(n5214), .A2(n5216), .ZN(n5196) );
  AND2_X1 U3687 ( .A1(n3101), .A2(n3140), .ZN(n3102) );
  CLKBUF_X1 U3688 ( .A(n4241), .Z(n3115) );
  INV_X1 U3689 ( .A(n6098), .ZN(n3103) );
  AND2_X2 U3690 ( .A1(n5625), .A2(n3262), .ZN(n5608) );
  CLKBUF_X1 U3691 ( .A(n6532), .Z(n3104) );
  NAND2_X2 U3692 ( .A1(n3371), .A2(n3370), .ZN(n3636) );
  NAND2_X1 U3693 ( .A1(n4220), .A2(n4219), .ZN(n6532) );
  NAND2_X1 U3694 ( .A1(n3101), .A2(n3108), .ZN(n3105) );
  NAND2_X1 U3695 ( .A1(n3105), .A2(n3106), .ZN(n5012) );
  OR2_X1 U3696 ( .A1(n3107), .A2(n4298), .ZN(n3106) );
  INV_X1 U3697 ( .A(n5011), .ZN(n3107) );
  AND2_X1 U3698 ( .A1(n3140), .A2(n5011), .ZN(n3108) );
  NAND2_X1 U3699 ( .A1(n3101), .A2(n3140), .ZN(n3109) );
  NAND2_X1 U3700 ( .A1(n3101), .A2(n3140), .ZN(n3110) );
  NAND3_X1 U3701 ( .A1(n3468), .A2(n3467), .A3(n3484), .ZN(n3111) );
  NAND2_X1 U3702 ( .A1(n4297), .A2(n3140), .ZN(n4299) );
  AND2_X1 U3703 ( .A1(n3339), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5961)
         );
  BUF_X2 U3704 ( .A(n3506), .Z(n4093) );
  NOR2_X2 U3705 ( .A1(n5355), .A2(n3309), .ZN(n5007) );
  OAI21_X2 U3706 ( .B1(n5078), .B2(n4554), .A(n4559), .ZN(n4441) );
  AND2_X1 U3708 ( .A1(n5960), .A2(n5050), .ZN(n3448) );
  AND2_X1 U3709 ( .A1(n5960), .A2(n4683), .ZN(n3506) );
  AND2_X1 U3710 ( .A1(n5046), .A2(n5960), .ZN(n3575) );
  AND2_X2 U3711 ( .A1(n3699), .A2(n4909), .ZN(n3619) );
  NAND2_X2 U3712 ( .A1(n3325), .A2(n4289), .ZN(n3324) );
  INV_X2 U3713 ( .A(n4290), .ZN(n5644) );
  INV_X4 U3714 ( .A(n5644), .ZN(n5720) );
  NOR2_X2 U3715 ( .A1(n3635), .A2(n6956), .ZN(n3813) );
  AND2_X1 U3716 ( .A1(n3636), .A2(n3635), .ZN(n4456) );
  NAND2_X1 U3717 ( .A1(n3434), .A2(n3463), .ZN(n4338) );
  NOR2_X2 U3718 ( .A1(n4880), .A2(n3306), .ZN(n4995) );
  NOR2_X2 U3719 ( .A1(n4541), .A2(n4542), .ZN(n4543) );
  XNOR2_X2 U3720 ( .A(n4441), .B(n4440), .ZN(n5041) );
  CLKBUF_X1 U3721 ( .A(n5690), .Z(n3113) );
  XNOR2_X1 U3723 ( .A(n3518), .B(n3187), .ZN(n3116) );
  XNOR2_X1 U3724 ( .A(n3676), .B(n3677), .ZN(n4241) );
  XNOR2_X1 U3725 ( .A(n3187), .B(n3518), .ZN(n4831) );
  NAND2_X1 U3726 ( .A1(n3482), .A2(n3495), .ZN(n3187) );
  NAND2_X1 U3727 ( .A1(n3101), .A2(n4296), .ZN(n5598) );
  AND2_X1 U3728 ( .A1(n5050), .A2(n4682), .ZN(n3426) );
  AND2_X1 U3729 ( .A1(n5050), .A2(n3344), .ZN(n3445) );
  XNOR2_X2 U3730 ( .A(n4347), .B(n4799), .ZN(n4808) );
  NAND2_X1 U3731 ( .A1(n3110), .A2(n3138), .ZN(n5566) );
  NAND2_X1 U3732 ( .A1(n5642), .A2(n4292), .ZN(n3171) );
  NAND2_X1 U3733 ( .A1(n3647), .A2(n3649), .ZN(n3676) );
  XNOR2_X2 U3734 ( .A(n3571), .B(n3569), .ZN(n3651) );
  INV_X2 U3735 ( .A(n4349), .ZN(n3118) );
  INV_X1 U3736 ( .A(n4349), .ZN(n4402) );
  AND2_X1 U3737 ( .A1(n5046), .A2(n3344), .ZN(n3120) );
  AND2_X2 U3738 ( .A1(n5046), .A2(n3344), .ZN(n3435) );
  NAND2_X4 U3739 ( .A1(n4343), .A2(n3118), .ZN(n4798) );
  OR2_X1 U3740 ( .A1(n3515), .A2(n7091), .ZN(n3573) );
  NAND2_X1 U3741 ( .A1(n3467), .A2(n3248), .ZN(n3247) );
  NOR2_X1 U3742 ( .A1(n3480), .A2(n3476), .ZN(n3248) );
  INV_X1 U3743 ( .A(n4332), .ZN(n3186) );
  AND2_X1 U3744 ( .A1(n5420), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U3745 ( .A1(n3661), .A2(n4941), .ZN(n3167) );
  INV_X1 U3746 ( .A(n3573), .ZN(n3547) );
  AOI22_X1 U3747 ( .A1(n3575), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U3748 ( .A1(n3178), .A2(n3153), .ZN(n5214) );
  INV_X1 U3749 ( .A(n5267), .ZN(n3822) );
  NAND2_X1 U3750 ( .A1(n4263), .A2(n4306), .ZN(n3169) );
  AND2_X1 U3751 ( .A1(n3263), .A2(n4505), .ZN(n3262) );
  INV_X1 U3752 ( .A(n5618), .ZN(n3263) );
  NAND3_X1 U3753 ( .A1(n3468), .A2(n3467), .A3(n3484), .ZN(n3209) );
  NOR2_X1 U3754 ( .A1(n3485), .A2(n3454), .ZN(n3468) );
  AND2_X1 U3755 ( .A1(n4950), .A2(n3460), .ZN(n3841) );
  INV_X1 U3756 ( .A(n3482), .ZN(n3330) );
  AND3_X1 U3757 ( .A1(n3568), .A2(n3567), .A3(n3566), .ZN(n3650) );
  INV_X1 U3758 ( .A(n3618), .ZN(n3172) );
  INV_X1 U3759 ( .A(n4324), .ZN(n4561) );
  OR2_X1 U3760 ( .A1(n5059), .A2(n4565), .ZN(n5420) );
  NOR2_X1 U3761 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  AND2_X1 U3762 ( .A1(n4072), .A2(n4071), .ZN(n5101) );
  OR3_X1 U3763 ( .A1(n4696), .A2(n4328), .A3(n3478), .ZN(n4329) );
  OR2_X1 U3764 ( .A1(n4335), .A2(n4334), .ZN(n5063) );
  NAND2_X1 U3765 ( .A1(n4187), .A2(n4319), .ZN(n4188) );
  NAND2_X1 U3766 ( .A1(n4186), .A2(n4185), .ZN(n3230) );
  NAND2_X1 U3767 ( .A1(n4561), .A2(n3487), .ZN(n6405) );
  NAND2_X1 U3768 ( .A1(n4189), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6788) );
  INV_X1 U3769 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5053) );
  NOR2_X1 U3770 ( .A1(n5065), .A2(n6343), .ZN(n6784) );
  INV_X1 U3771 ( .A(n4175), .ZN(n3235) );
  AND2_X1 U3772 ( .A1(n5183), .A2(n5197), .ZN(n3291) );
  INV_X1 U3773 ( .A(n4287), .ZN(n3326) );
  NAND2_X1 U3774 ( .A1(n4809), .A2(n4402), .ZN(n4348) );
  NAND2_X1 U3775 ( .A1(n3182), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3574) );
  NOR2_X1 U3776 ( .A1(n4151), .A2(n4152), .ZN(n3234) );
  NAND2_X1 U3777 ( .A1(n3547), .A2(n4222), .ZN(n3531) );
  AOI22_X1 U3778 ( .A1(n3611), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U3779 ( .A1(n3435), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U3780 ( .A1(n3206), .A2(n3203), .ZN(n3202) );
  NAND2_X1 U3781 ( .A1(n3207), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U3782 ( .A1(n3205), .A2(n3204), .ZN(n3203) );
  INV_X1 U3783 ( .A(n6436), .ZN(n3207) );
  NOR2_X1 U3784 ( .A1(n5305), .A2(n3289), .ZN(n3288) );
  INV_X1 U3785 ( .A(n3336), .ZN(n3289) );
  NOR3_X2 U3786 ( .A1(n5138), .A2(n5097), .A3(n3302), .ZN(n4437) );
  NAND2_X1 U3787 ( .A1(n3301), .A2(n3300), .ZN(n4541) );
  NOR2_X1 U3788 ( .A1(n3122), .A2(n3161), .ZN(n3300) );
  NOR2_X1 U3789 ( .A1(n5270), .A2(n3314), .ZN(n3313) );
  INV_X1 U3790 ( .A(n5287), .ZN(n3314) );
  NAND2_X1 U3791 ( .A1(n4281), .A2(n3320), .ZN(n3319) );
  INV_X1 U3792 ( .A(n4281), .ZN(n3321) );
  AND2_X1 U3793 ( .A1(n6513), .A2(n4985), .ZN(n4258) );
  NAND2_X1 U3794 ( .A1(n3209), .A2(n3156), .ZN(n3168) );
  NAND2_X1 U3795 ( .A1(n3490), .A2(n3166), .ZN(n3491) );
  AND2_X1 U3796 ( .A1(n4183), .A2(n4182), .ZN(n4319) );
  OR2_X1 U3797 ( .A1(n4181), .A2(n4180), .ZN(n4183) );
  NAND2_X1 U3798 ( .A1(n3500), .A2(n3499), .ZN(n3599) );
  NAND2_X1 U3799 ( .A1(n3127), .A2(n3112), .ZN(n3500) );
  OR2_X1 U3800 ( .A1(n4734), .A2(n4448), .ZN(n5028) );
  INV_X1 U3801 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6417) );
  INV_X1 U3802 ( .A(n3116), .ZN(n5044) );
  AOI21_X1 U3803 ( .B1(n3202), .B2(n6422), .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .ZN(n3200) );
  OAI21_X1 U3804 ( .B1(n3202), .B2(n6422), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n3201) );
  NAND2_X1 U3805 ( .A1(n6477), .A2(n3280), .ZN(n3279) );
  NAND2_X1 U3806 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3280)
         );
  NOR2_X1 U3807 ( .A1(n4570), .A2(n3245), .ZN(n3244) );
  INV_X1 U3808 ( .A(n4569), .ZN(n3245) );
  INV_X1 U3809 ( .A(n4889), .ZN(n6224) );
  AND2_X1 U3810 ( .A1(n4420), .A2(n4419), .ZN(n5135) );
  AOI21_X1 U3811 ( .B1(n4808), .B2(n4809), .A(n4347), .ZN(n4906) );
  INV_X1 U3812 ( .A(n5973), .ZN(n6412) );
  NAND2_X1 U3813 ( .A1(n3270), .A2(n3269), .ZN(n4594) );
  OR2_X1 U3814 ( .A1(n4112), .A2(n6910), .ZN(n3270) );
  NAND2_X1 U3815 ( .A1(n4112), .A2(n3131), .ZN(n4196) );
  OR2_X1 U3816 ( .A1(n4054), .A2(n5582), .ZN(n4111) );
  NOR2_X1 U3817 ( .A1(n4014), .A2(n5139), .ZN(n3266) );
  NAND2_X1 U3818 ( .A1(n3266), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4052)
         );
  NAND2_X1 U3819 ( .A1(n3973), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4014)
         );
  AND3_X1 U3820 ( .A1(n3821), .A2(n3820), .A3(n3819), .ZN(n5267) );
  INV_X1 U3821 ( .A(n5282), .ZN(n3803) );
  NAND2_X1 U3822 ( .A1(n3797), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3834)
         );
  INV_X1 U3823 ( .A(n4856), .ZN(n3174) );
  NAND2_X1 U3824 ( .A1(n3256), .A2(n3185), .ZN(n5728) );
  NAND2_X1 U3825 ( .A1(n6517), .A2(n3255), .ZN(n3185) );
  INV_X1 U3826 ( .A(n4543), .ZN(n5136) );
  OR2_X1 U3827 ( .A1(n5641), .A2(n4504), .ZN(n4505) );
  NOR2_X2 U3828 ( .A1(n5255), .A2(n5242), .ZN(n5241) );
  AND2_X1 U3829 ( .A1(n4395), .A2(n4394), .ZN(n5257) );
  NAND2_X1 U3830 ( .A1(n3310), .A2(n5485), .ZN(n3309) );
  NAND2_X1 U3831 ( .A1(n3246), .A2(n3252), .ZN(n3482) );
  OR2_X1 U3832 ( .A1(n3481), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3252)
         );
  NOR2_X1 U3833 ( .A1(n5983), .A2(n4221), .ZN(n6022) );
  AND2_X1 U3834 ( .A1(n6636), .A2(n6098), .ZN(n6134) );
  OR2_X1 U3835 ( .A1(n6136), .A2(n6135), .ZN(n6138) );
  AND2_X1 U3836 ( .A1(n4837), .A2(n5044), .ZN(n6348) );
  INV_X1 U3837 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6343) );
  XNOR2_X1 U3838 ( .A(n6907), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6372)
         );
  NOR2_X1 U3839 ( .A1(n5030), .A2(n5044), .ZN(n6373) );
  INV_X1 U3840 ( .A(n3477), .ZN(n4950) );
  INV_X1 U3841 ( .A(n3455), .ZN(n4145) );
  INV_X1 U3842 ( .A(n6220), .ZN(n6063) );
  INV_X1 U3843 ( .A(n6809), .ZN(n6338) );
  AND2_X1 U3844 ( .A1(n4835), .A2(n4910), .ZN(n4915) );
  NAND2_X1 U3845 ( .A1(n4697), .A2(n6449), .ZN(n5059) );
  INV_X1 U3846 ( .A(READY_N), .ZN(n6443) );
  NAND2_X1 U3847 ( .A1(n5151), .A2(n3236), .ZN(n5084) );
  AND2_X1 U3848 ( .A1(n3132), .A2(n3237), .ZN(n3236) );
  NOR2_X1 U3849 ( .A1(n7018), .A2(n5109), .ZN(n3237) );
  INV_X1 U3850 ( .A(n3242), .ZN(n3241) );
  OAI21_X1 U3851 ( .B1(n5041), .B2(n5415), .A(n3243), .ZN(n3242) );
  AOI21_X1 U3852 ( .B1(n4621), .B2(REIP_REG_31__SCAN_IN), .A(n4620), .ZN(n3243) );
  AND3_X1 U3853 ( .A1(n5420), .A2(n4594), .A3(STATE2_REG_1__SCAN_IN), .ZN(
        n6488) );
  OAI211_X2 U3854 ( .C1(n4696), .C2(n5063), .A(n4610), .B(n4785), .ZN(n5559)
         );
  AOI21_X1 U3855 ( .B1(n4753), .B2(n4608), .A(n4607), .ZN(n4610) );
  INV_X1 U3856 ( .A(n4502), .ZN(n3170) );
  OAI21_X1 U3857 ( .B1(n5090), .B2(n3294), .A(n3293), .ZN(n3292) );
  INV_X1 U3858 ( .A(n4141), .ZN(n3293) );
  NAND2_X1 U3859 ( .A1(n3909), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3911)
         );
  INV_X1 U3860 ( .A(n6541), .ZN(n5725) );
  NAND2_X1 U3861 ( .A1(n5750), .A2(n4193), .ZN(n5722) );
  INV_X1 U3862 ( .A(n6597), .ZN(n5951) );
  INV_X1 U3863 ( .A(n5957), .ZN(n6602) );
  AND2_X2 U3864 ( .A1(n4475), .A2(n4445), .ZN(n6597) );
  NAND2_X1 U3865 ( .A1(n4475), .A2(n4337), .ZN(n5957) );
  INV_X1 U3866 ( .A(n6691), .ZN(n6698) );
  INV_X1 U3867 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U3868 ( .A1(n3198), .A2(n3197), .ZN(n6416) );
  AOI21_X1 U3869 ( .B1(n5973), .B2(n5053), .A(n5045), .ZN(n3197) );
  NAND2_X1 U3870 ( .A1(n3116), .A2(n3199), .ZN(n3198) );
  INV_X1 U3871 ( .A(n6768), .ZN(n6740) );
  OR2_X1 U3872 ( .A1(n6804), .A2(n3194), .ZN(n3193) );
  INV_X1 U3873 ( .A(n3195), .ZN(n3194) );
  AOI21_X1 U3874 ( .B1(n6784), .B2(n6785), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3195) );
  AND2_X1 U3875 ( .A1(n3192), .A2(n3190), .ZN(n3189) );
  AND2_X1 U3876 ( .A1(n3191), .A2(n6783), .ZN(n3190) );
  NAND2_X1 U3877 ( .A1(n6802), .A2(n6787), .ZN(n3191) );
  NOR2_X1 U3878 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6442) );
  OR2_X1 U3879 ( .A1(n3457), .A2(n3460), .ZN(n3456) );
  AOI22_X1 U3880 ( .A1(n3506), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        INSTQUEUE_REG_0__4__SCAN_IN), .B2(n3438), .ZN(n3379) );
  NAND2_X1 U3881 ( .A1(n6436), .A2(n6421), .ZN(n3205) );
  AND2_X1 U3882 ( .A1(n6420), .A2(n6419), .ZN(n3204) );
  INV_X1 U3883 ( .A(n5691), .ZN(n3225) );
  INV_X1 U3884 ( .A(n4280), .ZN(n3320) );
  OR2_X1 U3885 ( .A1(n3595), .A2(n3594), .ZN(n4208) );
  NAND2_X1 U3886 ( .A1(n3466), .A2(n3182), .ZN(n3484) );
  OR2_X1 U3887 ( .A1(n3512), .A2(n3511), .ZN(n4201) );
  NAND2_X1 U3888 ( .A1(n4836), .A2(n7091), .ZN(n3514) );
  OR2_X1 U3889 ( .A1(n3530), .A2(n3529), .ZN(n4222) );
  OR2_X1 U3890 ( .A1(n3617), .A2(n3616), .ZN(n4242) );
  AOI22_X1 U3891 ( .A1(n3121), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U3892 ( .A1(n3435), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U3893 ( .A1(n3426), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U3894 ( .A1(n3611), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U3895 ( .A1(n3506), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U3896 ( .A1(n3099), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U3897 ( .A1(n3446), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U3898 ( .A1(n3611), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U3899 ( .A1(n3575), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U3900 ( .A1(n3435), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U3901 ( .A1(n3445), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U3902 ( .A1(n3436), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U3903 ( .A1(n5081), .A2(n3299), .ZN(n3298) );
  OR2_X1 U3904 ( .A1(n3961), .A2(n3960), .ZN(n4027) );
  AND2_X1 U3905 ( .A1(n4013), .A2(n3291), .ZN(n3290) );
  NOR2_X1 U3906 ( .A1(n4010), .A2(n5611), .ZN(n3973) );
  OR2_X1 U3907 ( .A1(n5156), .A2(n5172), .ZN(n4530) );
  AND2_X1 U3908 ( .A1(n5196), .A2(n3291), .ZN(n4529) );
  NOR2_X1 U3909 ( .A1(n3910), .A2(n3274), .ZN(n3273) );
  INV_X1 U3910 ( .A(n4109), .ZN(n4136) );
  OR2_X1 U3911 ( .A1(n5043), .A2(n7091), .ZN(n4109) );
  NOR2_X1 U3912 ( .A1(n3286), .A2(n3284), .ZN(n3283) );
  INV_X1 U3913 ( .A(n5240), .ZN(n3284) );
  NAND2_X1 U3914 ( .A1(n3287), .A2(n3822), .ZN(n3286) );
  INV_X1 U3915 ( .A(n5253), .ZN(n3287) );
  NAND2_X1 U3916 ( .A1(n5346), .A2(n3154), .ZN(n3176) );
  AND2_X1 U3917 ( .A1(n3764), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3771)
         );
  XNOR2_X1 U3918 ( .A(n4271), .B(n3634), .ZN(n4263) );
  XNOR2_X1 U3919 ( .A(n3227), .B(n3699), .ZN(n4206) );
  NAND2_X1 U3920 ( .A1(n3126), .A2(n4909), .ZN(n3227) );
  AND2_X1 U3921 ( .A1(n3265), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3642)
         );
  INV_X1 U3922 ( .A(n3666), .ZN(n3265) );
  NOR2_X2 U3923 ( .A1(n3636), .A2(n6956), .ZN(n4140) );
  INV_X1 U3924 ( .A(n3962), .ZN(n4139) );
  AND2_X1 U3925 ( .A1(n4456), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3670) );
  INV_X1 U3926 ( .A(n4140), .ZN(n4134) );
  NAND2_X1 U3927 ( .A1(n5574), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U3928 ( .A1(n3305), .A2(n3303), .ZN(n3302) );
  NOR2_X1 U3929 ( .A1(n5105), .A2(n3304), .ZN(n3303) );
  INV_X1 U3930 ( .A(n5126), .ZN(n3305) );
  INV_X1 U3931 ( .A(n5112), .ZN(n3304) );
  NOR2_X1 U3932 ( .A1(n4273), .A2(n4272), .ZN(n4274) );
  INV_X1 U3933 ( .A(n5355), .ZN(n3311) );
  NAND2_X1 U3934 ( .A1(n3119), .A2(EBX_REG_1__SCAN_IN), .ZN(n4340) );
  NOR2_X1 U3935 ( .A1(n5053), .A2(n7091), .ZN(n3251) );
  OAI21_X1 U3936 ( .B1(n3232), .B2(n3233), .A(n3231), .ZN(n4179) );
  NOR2_X1 U3937 ( .A1(n4325), .A2(n4192), .ZN(n3208) );
  INV_X1 U3938 ( .A(n4835), .ZN(n4887) );
  AOI22_X1 U3939 ( .A1(n3506), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3426), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3452) );
  INV_X1 U3940 ( .A(n3460), .ZN(n3558) );
  AND2_X1 U3941 ( .A1(n6791), .A2(n4686), .ZN(n4687) );
  NAND2_X1 U3942 ( .A1(n3229), .A2(n3228), .ZN(n4697) );
  INV_X1 U3943 ( .A(n5064), .ZN(n3228) );
  INV_X1 U3944 ( .A(n4696), .ZN(n3229) );
  NAND2_X1 U3945 ( .A1(n6442), .A2(n7091), .ZN(n4197) );
  OR2_X1 U3946 ( .A1(n4319), .A2(n4318), .ZN(n5069) );
  NOR2_X1 U3947 ( .A1(n4577), .A2(n3239), .ZN(n3238) );
  INV_X1 U3948 ( .A(n3298), .ZN(n3297) );
  NAND2_X1 U3949 ( .A1(n3297), .A2(n3296), .ZN(n3294) );
  INV_X1 U3950 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5139) );
  OR2_X1 U3951 ( .A1(n4008), .A2(n5621), .ZN(n4010) );
  INV_X1 U3952 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3910) );
  NAND2_X1 U3953 ( .A1(n3909), .A2(n3273), .ZN(n3964) );
  CLKBUF_X1 U3954 ( .A(n5214), .Z(n5215) );
  NOR2_X1 U3955 ( .A1(n3833), .A2(n3277), .ZN(n3276) );
  NAND2_X1 U3956 ( .A1(n3797), .A2(n3123), .ZN(n3873) );
  CLKBUF_X1 U3957 ( .A(n5280), .Z(n5281) );
  NOR2_X1 U3958 ( .A1(n3734), .A2(n7041), .ZN(n3764) );
  NAND2_X1 U3959 ( .A1(n3267), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3734)
         );
  INV_X1 U3960 ( .A(n3732), .ZN(n3267) );
  INV_X1 U3961 ( .A(n4262), .ZN(n3259) );
  NAND2_X1 U3962 ( .A1(n3268), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3732)
         );
  INV_X1 U3963 ( .A(n3694), .ZN(n3268) );
  NOR2_X1 U3964 ( .A1(n3700), .A2(n7111), .ZN(n3701) );
  INV_X1 U3965 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U3966 ( .A1(n3642), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3700)
         );
  AND2_X1 U3967 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5771) );
  AND2_X1 U3968 ( .A1(n3220), .A2(n3219), .ZN(n3215) );
  AND2_X1 U3969 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3220)
         );
  AND2_X1 U3970 ( .A1(n3221), .A2(n3219), .ZN(n3216) );
  INV_X1 U3971 ( .A(n3214), .ZN(n3212) );
  NOR2_X1 U3972 ( .A1(n3222), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3221)
         );
  INV_X1 U3973 ( .A(n5599), .ZN(n3329) );
  NOR2_X1 U3974 ( .A1(n3328), .A2(n5589), .ZN(n3327) );
  INV_X1 U3975 ( .A(n4298), .ZN(n3328) );
  INV_X1 U3976 ( .A(n5135), .ZN(n4421) );
  XNOR2_X1 U3977 ( .A(n5641), .B(n5572), .ZN(n5599) );
  AND2_X1 U3978 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5838) );
  AND2_X1 U3979 ( .A1(n4404), .A2(n4403), .ZN(n5203) );
  INV_X1 U3980 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5878) );
  AND2_X1 U3981 ( .A1(n3313), .A2(n3315), .ZN(n3312) );
  INV_X1 U3982 ( .A(n5257), .ZN(n3315) );
  NAND2_X1 U3983 ( .A1(n5720), .A2(n4286), .ZN(n4287) );
  AOI21_X1 U3984 ( .B1(n3318), .B2(n3321), .A(n3139), .ZN(n3316) );
  NAND2_X1 U3985 ( .A1(n5728), .A2(n3318), .ZN(n3317) );
  AND2_X1 U3986 ( .A1(n4385), .A2(n4384), .ZN(n5307) );
  NAND2_X1 U3987 ( .A1(n4259), .A2(n4260), .ZN(n6517) );
  NAND2_X1 U3988 ( .A1(n4996), .A2(n4358), .ZN(n3307) );
  INV_X1 U3989 ( .A(n4822), .ZN(n5950) );
  CLKBUF_X1 U3990 ( .A(n4983), .Z(n4984) );
  OR2_X1 U3991 ( .A1(n4861), .A2(n4882), .ZN(n3308) );
  NAND2_X1 U3992 ( .A1(n4475), .A2(n5067), .ZN(n6599) );
  OR2_X1 U3993 ( .A1(n4197), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6522) );
  NOR3_X1 U3994 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6421), .A3(n6417), 
        .ZN(n6640) );
  AND2_X1 U3995 ( .A1(n5988), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U3996 ( .A1(n3115), .A2(n4887), .ZN(n6693) );
  AND2_X1 U3997 ( .A1(n4835), .A2(n4886), .ZN(n4963) );
  NAND2_X1 U3998 ( .A1(n4898), .A2(n6803), .ZN(n4951) );
  AND2_X1 U3999 ( .A1(n3201), .A2(n3200), .ZN(n6434) );
  OR2_X1 U4000 ( .A1(n4679), .A2(n6788), .ZN(n6449) );
  INV_X1 U4001 ( .A(n4809), .ZN(n5054) );
  NAND2_X1 U4002 ( .A1(n5420), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6478) );
  INV_X1 U4003 ( .A(n6487), .ZN(n5414) );
  NAND2_X1 U4004 ( .A1(n5151), .A2(n3238), .ZN(n5119) );
  NAND2_X1 U4005 ( .A1(n5151), .A2(REIP_REG_23__SCAN_IN), .ZN(n5144) );
  OR2_X1 U4006 ( .A1(n5222), .A2(n4575), .ZN(n5174) );
  OR2_X1 U4007 ( .A1(n5259), .A2(n4574), .ZN(n5222) );
  NAND2_X1 U4008 ( .A1(n3135), .A2(n4572), .ZN(n5259) );
  AOI21_X1 U4009 ( .B1(n6487), .B2(n3281), .A(n3279), .ZN(n5285) );
  INV_X1 U4010 ( .A(n5686), .ZN(n3281) );
  INV_X1 U4011 ( .A(n6488), .ZN(n5385) );
  AND2_X1 U4012 ( .A1(n5459), .A2(n5363), .ZN(n5379) );
  NAND2_X1 U4013 ( .A1(n5400), .A2(n4569), .ZN(n5429) );
  AND2_X1 U4014 ( .A1(n4583), .A2(n5420), .ZN(n6487) );
  INV_X1 U4015 ( .A(n5449), .ZN(n5462) );
  INV_X1 U4016 ( .A(n5497), .ZN(n6492) );
  INV_X1 U4017 ( .A(n6495), .ZN(n5493) );
  NAND2_X1 U4018 ( .A1(n4601), .A2(n4600), .ZN(n6495) );
  AND2_X1 U4019 ( .A1(n4941), .A2(n3183), .ZN(n4599) );
  NAND2_X1 U4020 ( .A1(n6495), .A2(n4919), .ZN(n5497) );
  NOR2_X2 U4021 ( .A1(n5542), .A2(n4325), .ZN(n5535) );
  AND2_X1 U4022 ( .A1(n5559), .A2(n5021), .ZN(n5536) );
  INV_X1 U4023 ( .A(n5559), .ZN(n5542) );
  NAND2_X1 U4024 ( .A1(n5559), .A2(n4814), .ZN(n5560) );
  OR3_X1 U4025 ( .A1(n4696), .A2(n4692), .A3(n4727), .ZN(n4842) );
  NAND2_X1 U4026 ( .A1(n7091), .A2(n4693), .ZN(n6508) );
  AND2_X1 U4027 ( .A1(n4842), .A2(n6508), .ZN(n6506) );
  INV_X1 U4028 ( .A(n4842), .ZN(n6505) );
  OAI21_X2 U4029 ( .B1(n3487), .B2(n6443), .A(n6448), .ZN(n6825) );
  OR3_X1 U4030 ( .A1(n4696), .A2(READY_N), .A3(n4609), .ZN(n4785) );
  OR2_X1 U4031 ( .A1(n4696), .A2(n6405), .ZN(n6828) );
  INV_X1 U4032 ( .A(n6825), .ZN(n4786) );
  AND2_X1 U4033 ( .A1(n4112), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4113)
         );
  NOR2_X1 U4034 ( .A1(n5079), .A2(n3179), .ZN(n5578) );
  NOR2_X1 U4035 ( .A1(n3180), .A2(n3299), .ZN(n3179) );
  INV_X1 U4036 ( .A(n5090), .ZN(n3180) );
  AND2_X1 U4037 ( .A1(n4111), .A2(n4055), .ZN(n5586) );
  INV_X1 U4038 ( .A(n3266), .ZN(n4015) );
  INV_X1 U4039 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5611) );
  INV_X1 U4040 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5621) );
  OR2_X1 U4041 ( .A1(n5181), .A2(n5198), .ZN(n5635) );
  OR2_X1 U4042 ( .A1(n5306), .A2(n5292), .ZN(n5708) );
  INV_X1 U4043 ( .A(n5004), .ZN(n5482) );
  INV_X1 U4044 ( .A(n5722), .ZN(n6531) );
  INV_X1 U4045 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5751) );
  NOR2_X1 U4046 ( .A1(n4519), .A2(n4518), .ZN(n5811) );
  AND2_X1 U4047 ( .A1(n5641), .A2(n5606), .ZN(n5607) );
  NAND2_X1 U4048 ( .A1(n5625), .A2(n4505), .ZN(n5617) );
  INV_X1 U4049 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7012) );
  CLKBUF_X1 U4050 ( .A(n4870), .Z(n4871) );
  NOR2_X1 U4051 ( .A1(n7079), .A2(n6956), .ZN(n4693) );
  INV_X1 U4052 ( .A(n6140), .ZN(n6214) );
  AND2_X1 U4053 ( .A1(n3103), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6635) );
  CLKBUF_X1 U4054 ( .A(n4836), .Z(n4837) );
  AND2_X1 U4055 ( .A1(n6691), .A2(n7046), .ZN(n6809) );
  INV_X1 U4056 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7079) );
  AND2_X1 U4057 ( .A1(n4309), .A2(n4449), .ZN(n5973) );
  AND2_X1 U4058 ( .A1(n5990), .A2(n5989), .ZN(n6014) );
  AOI22_X1 U4059 ( .A1(n6025), .A2(n6023), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6021), .ZN(n6058) );
  OAI21_X1 U4060 ( .B1(n4893), .B2(n4892), .A(n4891), .ZN(n6626) );
  OAI21_X1 U4061 ( .B1(n6105), .B2(n6343), .A(n6103), .ZN(n6127) );
  AOI22_X1 U4062 ( .A1(n6144), .A2(n6142), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6139), .ZN(n6174) );
  INV_X1 U4063 ( .A(n6179), .ZN(n6211) );
  AND2_X1 U4064 ( .A1(n6299), .A2(n6298), .ZN(n6334) );
  OR2_X1 U4065 ( .A1(n6301), .A2(n6300), .ZN(n6299) );
  INV_X1 U4066 ( .A(n6688), .ZN(n6633) );
  INV_X1 U4067 ( .A(n6708), .ZN(n6611) );
  INV_X1 U4068 ( .A(n6722), .ZN(n6656) );
  INV_X1 U4069 ( .A(n6729), .ZN(n6754) );
  INV_X1 U4070 ( .A(n6665), .ZN(n6755) );
  INV_X1 U4071 ( .A(n6734), .ZN(n6760) );
  INV_X1 U4072 ( .A(n6739), .ZN(n6766) );
  NOR2_X1 U4073 ( .A1(n6907), .A2(n6340), .ZN(n4980) );
  INV_X1 U4074 ( .A(n6745), .ZN(n6772) );
  INV_X1 U4075 ( .A(n6685), .ZN(n6774) );
  AND2_X1 U4076 ( .A1(n4963), .A2(n6140), .ZN(n6776) );
  NOR2_X1 U4077 ( .A1(n5718), .A2(n4930), .ZN(n6646) );
  INV_X1 U4078 ( .A(n6612), .ZN(n6709) );
  NAND2_X1 U4079 ( .A1(n6536), .A2(DATAI_20_), .ZN(n6733) );
  NOR2_X1 U4080 ( .A1(n5718), .A2(n7076), .ZN(n6673) );
  NAND2_X1 U4081 ( .A1(n6536), .A2(DATAI_23_), .ZN(n6752) );
  NOR2_X1 U4082 ( .A1(n5718), .A2(n4911), .ZN(n6681) );
  OR2_X1 U4083 ( .A1(n4951), .A2(n3182), .ZN(n6688) );
  NAND2_X1 U4084 ( .A1(DATAI_1_), .A2(n6063), .ZN(n6649) );
  NAND2_X1 U4085 ( .A1(DATAI_2_), .A2(n6063), .ZN(n6655) );
  OR2_X1 U4086 ( .A1(n4951), .A2(n4950), .ZN(n6715) );
  NAND2_X1 U4087 ( .A1(DATAI_3_), .A2(n6063), .ZN(n6661) );
  OR2_X1 U4088 ( .A1(n4951), .A2(n4941), .ZN(n6722) );
  NAND2_X1 U4089 ( .A1(DATAI_4_), .A2(n6063), .ZN(n6665) );
  NOR2_X1 U4090 ( .A1(n5718), .A2(n4896), .ZN(n6762) );
  NAND2_X1 U4091 ( .A1(DATAI_6_), .A2(n6063), .ZN(n6676) );
  OR2_X1 U4092 ( .A1(n4951), .A2(n4305), .ZN(n6739) );
  NOR2_X1 U4093 ( .A1(n5718), .A2(n4926), .ZN(n6768) );
  NAND2_X1 U4094 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4917), .ZN(n4952) );
  NAND2_X1 U4095 ( .A1(DATAI_7_), .A2(n6063), .ZN(n6685) );
  OR2_X1 U4096 ( .A1(n4951), .A2(n4919), .ZN(n6745) );
  NAND2_X1 U4097 ( .A1(n6638), .A2(n4914), .ZN(n4948) );
  AND2_X1 U4098 ( .A1(n4915), .A2(n6214), .ZN(n6016) );
  INV_X1 U4099 ( .A(n6788), .ZN(n6440) );
  NAND2_X1 U4100 ( .A1(n7079), .A2(n6956), .ZN(n6791) );
  NAND2_X1 U4101 ( .A1(n4313), .A2(n4312), .ZN(n4727) );
  INV_X1 U4102 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4636) );
  INV_X2 U4103 ( .A(n6797), .ZN(n6824) );
  NAND2_X1 U4104 ( .A1(n4622), .A2(n3241), .ZN(n3240) );
  NAND2_X1 U4105 ( .A1(n3170), .A2(n6535), .ZN(n4301) );
  OR2_X1 U4106 ( .A1(n4498), .A2(n3331), .ZN(n4499) );
  AOI211_X1 U4107 ( .C1(n5756), .C2(n6597), .A(n5755), .B(n5754), .ZN(n5757)
         );
  AND2_X1 U4108 ( .A1(n4549), .A2(n4548), .ZN(n4550) );
  OR2_X1 U4109 ( .A1(n5469), .A2(n5951), .ZN(n4549) );
  INV_X1 U4110 ( .A(n6416), .ZN(n6414) );
  NAND2_X1 U4111 ( .A1(n3196), .A2(n3188), .ZN(U3148) );
  NAND2_X1 U4112 ( .A1(n6786), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3196) );
  AND2_X1 U4113 ( .A1(n3193), .A2(n3189), .ZN(n3188) );
  AND3_X1 U4114 ( .A1(n3177), .A2(n3739), .A3(n3145), .ZN(n5004) );
  NAND2_X1 U4115 ( .A1(n4145), .A2(n4950), .ZN(n3476) );
  OR2_X1 U4116 ( .A1(n3128), .A2(n5173), .ZN(n3122) );
  AND2_X1 U4117 ( .A1(n3276), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3123)
         );
  XNOR2_X2 U4118 ( .A(n3651), .B(n3650), .ZN(n4221) );
  NAND2_X1 U4119 ( .A1(n3285), .A2(n3822), .ZN(n5252) );
  NAND2_X1 U4120 ( .A1(n3285), .A2(n3283), .ZN(n5227) );
  NOR2_X1 U4121 ( .A1(n5199), .A2(n3122), .ZN(n5159) );
  OR2_X1 U4122 ( .A1(n5138), .A2(n3302), .ZN(n3124) );
  AND4_X1 U4123 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3125)
         );
  AND3_X1 U4124 ( .A1(n3647), .A2(n3649), .A3(n3226), .ZN(n3126) );
  AND2_X1 U4125 ( .A1(n4145), .A2(n4950), .ZN(n3183) );
  NAND2_X1 U4126 ( .A1(n3467), .A2(n3183), .ZN(n4324) );
  AND2_X1 U4127 ( .A1(n3209), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U4128 ( .A1(n4412), .A2(n4411), .ZN(n3128) );
  OAI211_X1 U4129 ( .C1(n3254), .C2(n3114), .A(n3253), .B(n4270), .ZN(n5727)
         );
  AND2_X1 U4130 ( .A1(n3173), .A2(n3636), .ZN(n3129) );
  NAND2_X2 U4131 ( .A1(n3432), .A2(n3431), .ZN(n3463) );
  NOR2_X1 U4132 ( .A1(n4837), .A2(n3116), .ZN(n3130) );
  NAND2_X1 U4133 ( .A1(n3311), .A2(n4371), .ZN(n5336) );
  OR2_X1 U4134 ( .A1(n4880), .A2(n4882), .ZN(n4860) );
  NAND2_X1 U4135 ( .A1(n4872), .A2(n4870), .ZN(n4873) );
  NAND2_X1 U4136 ( .A1(n4986), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6513)
         );
  AND2_X1 U4137 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3131) );
  AND2_X1 U4138 ( .A1(n3238), .A2(REIP_REG_26__SCAN_IN), .ZN(n3132) );
  AND2_X1 U4139 ( .A1(n3271), .A2(n6910), .ZN(n3133) );
  BUF_X1 U4140 ( .A(n4215), .Z(n4835) );
  NOR2_X1 U4141 ( .A1(n4855), .A2(n4856), .ZN(n4857) );
  AND2_X1 U4142 ( .A1(n5196), .A2(n5197), .ZN(n5181) );
  NAND2_X1 U4143 ( .A1(n5196), .A2(n3290), .ZN(n4521) );
  AND2_X1 U4144 ( .A1(n5004), .A2(n3288), .ZN(n5292) );
  NOR2_X1 U4145 ( .A1(n5265), .A2(n3286), .ZN(n5239) );
  AND2_X1 U4146 ( .A1(n5151), .A2(n3132), .ZN(n3134) );
  AND2_X1 U4147 ( .A1(n5400), .A2(n3244), .ZN(n3135) );
  AND2_X1 U4148 ( .A1(n3208), .A2(n4450), .ZN(n4309) );
  NAND2_X1 U4149 ( .A1(n5004), .A2(n3336), .ZN(n5005) );
  INV_X1 U4150 ( .A(n4456), .ZN(n4325) );
  INV_X1 U4151 ( .A(n3679), .ZN(n3226) );
  NAND2_X1 U4152 ( .A1(n5728), .A2(n4280), .ZN(n5719) );
  NAND2_X1 U4153 ( .A1(n4285), .A2(n5691), .ZN(n5683) );
  NAND2_X1 U4154 ( .A1(n3109), .A2(n3327), .ZN(n3137) );
  NAND2_X1 U4155 ( .A1(n5683), .A2(n5684), .ZN(n5675) );
  AND2_X1 U4156 ( .A1(n3327), .A2(n5771), .ZN(n3138) );
  AND2_X1 U4157 ( .A1(n5641), .A2(n4284), .ZN(n3139) );
  INV_X1 U4158 ( .A(n3165), .ZN(n4462) );
  NAND2_X1 U4159 ( .A1(n3182), .A2(n3463), .ZN(n3165) );
  AND2_X1 U4160 ( .A1(n3329), .A2(n4296), .ZN(n3140) );
  INV_X1 U4161 ( .A(n5265), .ZN(n3285) );
  NOR2_X1 U4162 ( .A1(n5138), .A2(n5126), .ZN(n5111) );
  AND2_X1 U4163 ( .A1(n5719), .A2(n4281), .ZN(n3141) );
  AND2_X1 U4164 ( .A1(n5675), .A2(n4287), .ZN(n3142) );
  AND2_X1 U4165 ( .A1(n5720), .A2(n5875), .ZN(n3143) );
  INV_X1 U4166 ( .A(n5357), .ZN(n4371) );
  INV_X1 U4167 ( .A(n3324), .ZN(n3323) );
  NAND2_X1 U4168 ( .A1(n4305), .A2(n3636), .ZN(n4465) );
  OR3_X1 U4169 ( .A1(n5138), .A2(n5126), .A3(n3304), .ZN(n3144) );
  AND3_X1 U4170 ( .A1(n3174), .A2(n5348), .A3(n5346), .ZN(n3145) );
  BUF_X1 U4171 ( .A(n3558), .Z(n4936) );
  NOR2_X1 U4172 ( .A1(n4173), .A2(n4174), .ZN(n3146) );
  AND2_X1 U4173 ( .A1(n4932), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3147) );
  AND2_X1 U4174 ( .A1(n3479), .A2(n3471), .ZN(n3148) );
  AND2_X1 U4175 ( .A1(n3290), .A2(n4033), .ZN(n3149) );
  NAND2_X1 U4176 ( .A1(n3457), .A2(n3463), .ZN(n3486) );
  NAND3_X1 U4177 ( .A1(n4153), .A2(STATE2_REG_0__SCAN_IN), .A3(n4315), .ZN(
        n3150) );
  AND2_X1 U4178 ( .A1(n5641), .A2(n4294), .ZN(n3151) );
  AND2_X1 U4179 ( .A1(n5241), .A2(n5225), .ZN(n5202) );
  NAND2_X1 U4180 ( .A1(n5294), .A2(n3313), .ZN(n5254) );
  NAND2_X1 U4181 ( .A1(n5294), .A2(n5287), .ZN(n5268) );
  INV_X1 U4182 ( .A(n3458), .ZN(n4305) );
  INV_X1 U4183 ( .A(n5091), .ZN(n3299) );
  INV_X1 U4184 ( .A(n5959), .ZN(n3199) );
  AND2_X1 U4185 ( .A1(n4434), .A2(n4433), .ZN(n5097) );
  INV_X1 U4186 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6413) );
  INV_X1 U4187 ( .A(n4593), .ZN(n3296) );
  OR2_X1 U4188 ( .A1(n5199), .A2(n3128), .ZN(n3152) );
  AND2_X1 U4189 ( .A1(n3283), .A2(n3876), .ZN(n3153) );
  AND2_X1 U4190 ( .A1(n3288), .A2(n5293), .ZN(n3154) );
  AND2_X1 U4191 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3155) );
  AND2_X1 U4192 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3156) );
  INV_X1 U4193 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6909) );
  INV_X1 U4194 ( .A(n3112), .ZN(n5039) );
  INV_X1 U4195 ( .A(n3164), .ZN(n4451) );
  NAND2_X1 U4196 ( .A1(n3463), .A2(n4950), .ZN(n3164) );
  NAND2_X1 U4197 ( .A1(n3797), .A2(n3276), .ZN(n3157) );
  AND2_X1 U4198 ( .A1(n3262), .A2(n5605), .ZN(n3158) );
  AND2_X1 U4199 ( .A1(n3311), .A2(n3310), .ZN(n3159) );
  AND2_X1 U4200 ( .A1(n3123), .A2(n3155), .ZN(n3160) );
  INV_X1 U4201 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3278) );
  INV_X1 U4202 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3277) );
  NOR2_X1 U4203 ( .A1(n4880), .A2(n3308), .ZN(n4859) );
  OR2_X2 U4204 ( .A1(n4696), .A2(n6424), .ZN(n5750) );
  INV_X1 U4205 ( .A(n5750), .ZN(n6535) );
  AND2_X1 U4206 ( .A1(n4415), .A2(n4414), .ZN(n3161) );
  AND2_X1 U4207 ( .A1(n3273), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3162)
         );
  INV_X1 U4208 ( .A(n4334), .ZN(n3181) );
  INV_X1 U4209 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6421) );
  INV_X1 U4210 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7105) );
  INV_X1 U4211 ( .A(n3272), .ZN(n3271) );
  NAND2_X1 U4212 ( .A1(n3131), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3272)
         );
  OR2_X1 U4213 ( .A1(n6791), .A2(n4563), .ZN(n6783) );
  AND2_X1 U4214 ( .A1(n3272), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3163)
         );
  INV_X1 U4215 ( .A(REIP_REG_23__SCAN_IN), .ZN(n3239) );
  INV_X2 U4216 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7091) );
  INV_X1 U4217 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3274) );
  INV_X1 U4218 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3218) );
  INV_X1 U4219 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U4220 ( .A1(n3168), .A2(n3483), .ZN(n3534) );
  NAND2_X1 U4221 ( .A1(n3127), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3605) );
  XNOR2_X2 U4222 ( .A(n4269), .B(n7012), .ZN(n5737) );
  NAND2_X1 U4223 ( .A1(n3129), .A2(n4936), .ZN(n4304) );
  NAND2_X1 U4224 ( .A1(n3456), .A2(n3129), .ZN(n4453) );
  NAND2_X2 U4225 ( .A1(n3171), .A2(n4293), .ZN(n5633) );
  OAI21_X2 U4226 ( .B1(n4285), .B2(n3324), .A(n3223), .ZN(n5642) );
  NAND2_X2 U4227 ( .A1(n5690), .A2(n5692), .ZN(n4285) );
  AOI21_X2 U4228 ( .B1(n4889), .B2(n7091), .A(n3172), .ZN(n6097) );
  XNOR2_X2 U4229 ( .A(n4751), .B(n6337), .ZN(n4889) );
  NAND2_X2 U4230 ( .A1(n3136), .A2(n3125), .ZN(n3455) );
  NAND2_X1 U4231 ( .A1(n4145), .A2(n3458), .ZN(n3173) );
  NAND4_X1 U4232 ( .A1(n3177), .A2(n3739), .A3(n5348), .A4(n3175), .ZN(n5280)
         );
  NAND3_X1 U4233 ( .A1(n3675), .A2(n4864), .A3(n4865), .ZN(n4855) );
  INV_X1 U4234 ( .A(n6532), .ZN(n4238) );
  NAND2_X1 U4235 ( .A1(n6532), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4237)
         );
  NAND3_X1 U4236 ( .A1(n3181), .A2(n4941), .A3(n3183), .ZN(n4442) );
  INV_X2 U4237 ( .A(n4331), .ZN(n3182) );
  OAI21_X2 U4238 ( .B1(n5566), .B2(n4493), .A(n4300), .ZN(n3184) );
  NAND3_X1 U4239 ( .A1(n3494), .A2(n3493), .A3(n4459), .ZN(n3533) );
  AND2_X2 U4240 ( .A1(n3534), .A2(n3533), .ZN(n3518) );
  OR2_X1 U4241 ( .A1(n6789), .A2(n6788), .ZN(n3192) );
  NAND3_X1 U4242 ( .A1(n3208), .A2(n3147), .A3(n4450), .ZN(n3479) );
  NAND2_X1 U4243 ( .A1(n3111), .A2(n3251), .ZN(n3249) );
  OAI21_X1 U4244 ( .B1(n5778), .B2(n5957), .A(n3217), .ZN(U2990) );
  NAND3_X1 U4245 ( .A1(n3214), .A2(n3213), .A3(n3218), .ZN(n3210) );
  NAND2_X1 U4246 ( .A1(n5573), .A2(n3216), .ZN(n3214) );
  NAND2_X1 U4247 ( .A1(n3098), .A2(n3215), .ZN(n3213) );
  NAND2_X1 U4248 ( .A1(n5573), .A2(n3221), .ZN(n5580) );
  INV_X1 U4249 ( .A(n5588), .ZN(n3222) );
  NAND2_X1 U4250 ( .A1(n3323), .A2(n3225), .ZN(n3224) );
  AND2_X2 U4251 ( .A1(n4683), .A2(n3344), .ZN(n3438) );
  NOR2_X4 U4252 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4253 ( .A1(n3126), .A2(n3619), .ZN(n3690) );
  OR2_X2 U4254 ( .A1(n5065), .A2(n6788), .ZN(n4696) );
  AOI21_X1 U4255 ( .B1(n4160), .B2(n3235), .A(n3146), .ZN(n3231) );
  NAND2_X1 U4256 ( .A1(n3235), .A2(n3150), .ZN(n3232) );
  AOI21_X1 U4257 ( .B1(n4150), .B2(n4176), .A(n3234), .ZN(n3233) );
  OR2_X1 U4258 ( .A1(n4619), .A2(n3240), .ZN(U2796) );
  NAND3_X1 U4259 ( .A1(n3250), .A2(n3247), .A3(n3479), .ZN(n3246) );
  NAND2_X1 U4260 ( .A1(n5737), .A2(n3259), .ZN(n3253) );
  INV_X1 U4261 ( .A(n5737), .ZN(n3254) );
  INV_X1 U4262 ( .A(n3257), .ZN(n3256) );
  INV_X1 U4263 ( .A(n4270), .ZN(n3258) );
  NAND2_X1 U4264 ( .A1(n5735), .A2(n5737), .ZN(n5736) );
  NAND2_X1 U4265 ( .A1(n3114), .A2(n4262), .ZN(n5735) );
  AOI21_X2 U4266 ( .B1(n5633), .B2(n5634), .A(n4503), .ZN(n5627) );
  NAND2_X1 U4267 ( .A1(n5625), .A2(n3158), .ZN(n3260) );
  NAND2_X1 U4268 ( .A1(n4527), .A2(n4528), .ZN(n3261) );
  AOI21_X1 U4269 ( .B1(n4112), .B2(n3133), .A(n3163), .ZN(n3269) );
  NAND2_X1 U4270 ( .A1(n3909), .A2(n3162), .ZN(n4008) );
  INV_X1 U4271 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4272 ( .A1(n3797), .A2(n3160), .ZN(n3908) );
  INV_X1 U4273 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3282) );
  AND2_X2 U4274 ( .A1(n3282), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5046)
         );
  INV_X1 U4275 ( .A(n5280), .ZN(n3804) );
  OAI21_X1 U4276 ( .B1(n5090), .B2(n3295), .A(n3292), .ZN(n4614) );
  NOR2_X1 U4277 ( .A1(n5090), .A2(n5091), .ZN(n5079) );
  NAND3_X1 U4278 ( .A1(n3297), .A2(n4141), .A3(n3296), .ZN(n3295) );
  INV_X1 U4279 ( .A(n5199), .ZN(n3301) );
  NAND2_X2 U4280 ( .A1(n5294), .A2(n3312), .ZN(n5255) );
  NAND2_X1 U4281 ( .A1(n3099), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4282 ( .A1(n3317), .A2(n3316), .ZN(n5690) );
  AOI21_X2 U4283 ( .B1(n3323), .B2(n3326), .A(n3143), .ZN(n3322) );
  OR2_X2 U4284 ( .A1(n5684), .A2(n3326), .ZN(n3325) );
  XNOR2_X1 U4285 ( .A(n3598), .B(n3599), .ZN(n4836) );
  OAI21_X2 U4286 ( .B1(n3518), .B2(n3330), .A(n3495), .ZN(n3598) );
  NAND2_X1 U4287 ( .A1(n4212), .A2(n4211), .ZN(n4986) );
  INV_X1 U4288 ( .A(n5020), .ZN(n5024) );
  AOI21_X1 U4289 ( .B1(n5020), .B2(n6493), .A(n4603), .ZN(n4604) );
  NAND2_X1 U4290 ( .A1(n5020), .A2(n6488), .ZN(n4595) );
  XNOR2_X1 U4291 ( .A(n5568), .B(n5765), .ZN(n5759) );
  OAI21_X1 U4292 ( .B1(n3098), .B2(n5567), .A(n5566), .ZN(n5568) );
  NAND2_X1 U4293 ( .A1(n5608), .A2(n4511), .ZN(n4517) );
  INV_X1 U4294 ( .A(n4875), .ZN(n3675) );
  NAND2_X1 U4295 ( .A1(n4206), .A2(n4306), .ZN(n4212) );
  INV_X1 U4296 ( .A(n6493), .ZN(n5490) );
  INV_X1 U4297 ( .A(n5495), .ZN(n6493) );
  NAND2_X2 U4298 ( .A1(n5559), .A2(n4813), .ZN(n5561) );
  OR2_X1 U4299 ( .A1(n4497), .A2(n4496), .ZN(n3331) );
  INV_X2 U4300 ( .A(n5718), .ZN(n6536) );
  INV_X1 U4301 ( .A(n5115), .ZN(n5124) );
  AND2_X1 U4302 ( .A1(n4312), .A2(STATE_REG_1__SCAN_IN), .ZN(n6797) );
  INV_X1 U4303 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5002) );
  INV_X1 U4304 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5552) );
  INV_X1 U4305 ( .A(DATAI_19_), .ZN(n4940) );
  AND3_X1 U4306 ( .A1(n3451), .A2(n3450), .A3(n3449), .ZN(n3332) );
  INV_X1 U4307 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5127) );
  INV_X1 U4308 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3731) );
  AND2_X1 U4309 ( .A1(n4365), .A2(n4364), .ZN(n3333) );
  INV_X1 U4310 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6957) );
  INV_X1 U4311 ( .A(REIP_REG_4__SCAN_IN), .ZN(n4670) );
  AND2_X1 U4312 ( .A1(n4351), .A2(n4350), .ZN(n3334) );
  AND2_X1 U4313 ( .A1(n5483), .A2(n5345), .ZN(n3335) );
  OR2_X1 U4314 ( .A1(n3753), .A2(n3752), .ZN(n3336) );
  INV_X1 U4315 ( .A(n3481), .ZN(n3471) );
  OR2_X1 U4316 ( .A1(n3629), .A2(n3628), .ZN(n4265) );
  INV_X1 U4317 ( .A(n3689), .ZN(n3630) );
  OR2_X1 U4318 ( .A1(n3585), .A2(n3584), .ZN(n4251) );
  NAND2_X1 U4319 ( .A1(n4174), .A2(n4306), .ZN(n4176) );
  AOI22_X1 U4320 ( .A1(n3436), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3422) );
  AND2_X1 U4321 ( .A1(n6907), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4155)
         );
  INV_X1 U4322 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n7025) );
  INV_X1 U4323 ( .A(n5229), .ZN(n3876) );
  NAND2_X1 U4324 ( .A1(n3547), .A2(n4276), .ZN(n4273) );
  INV_X1 U4325 ( .A(n4176), .ZN(n4184) );
  NAND2_X1 U4326 ( .A1(n6875), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4182) );
  AND2_X1 U4327 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5313), .ZN(n5296) );
  NAND2_X1 U4328 ( .A1(n3364), .A2(n3363), .ZN(n3369) );
  INV_X1 U4329 ( .A(n5116), .ZN(n4051) );
  NAND2_X1 U4330 ( .A1(n3641), .A2(n3640), .ZN(n5348) );
  OAI21_X1 U4331 ( .B1(n5878), .B2(n4482), .A(n5641), .ZN(n4293) );
  AND2_X1 U4332 ( .A1(n3601), .A2(n4952), .ZN(n6218) );
  OR2_X1 U4333 ( .A1(n4837), .A2(n5044), .ZN(n6295) );
  INV_X1 U4334 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3561) );
  INV_X1 U4335 ( .A(n6478), .ZN(n5454) );
  OR2_X1 U4336 ( .A1(n4375), .A2(EBX_REG_26__SCAN_IN), .ZN(n4425) );
  AND2_X1 U4337 ( .A1(n4010), .A2(n4009), .ZN(n5619) );
  AND2_X1 U4338 ( .A1(n3874), .A2(n3908), .ZN(n5655) );
  AND2_X2 U4339 ( .A1(n4475), .A2(n5973), .ZN(n5917) );
  AND2_X1 U4340 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3496) );
  NOR2_X1 U4341 ( .A1(n6907), .A2(n6143), .ZN(n6169) );
  NAND2_X1 U4342 ( .A1(n3605), .A2(n3604), .ZN(n6337) );
  OAI211_X1 U4343 ( .C1(n3632), .C2(n3561), .A(n3560), .B(n3559), .ZN(n3657)
         );
  INV_X1 U4344 ( .A(n3813), .ZN(n3838) );
  INV_X1 U4345 ( .A(n4033), .ZN(n5125) );
  INV_X1 U4346 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n7041) );
  INV_X1 U4347 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5574) );
  OR2_X1 U4348 ( .A1(n5821), .A2(n4487), .ZN(n4547) );
  AND2_X1 U4349 ( .A1(n5641), .A2(n6995), .ZN(n4503) );
  INV_X1 U4350 ( .A(n4290), .ZN(n5699) );
  OR2_X1 U4351 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5917), .ZN(n4821)
         );
  OR2_X1 U4352 ( .A1(n6784), .A2(n4687), .ZN(n4898) );
  INV_X1 U4353 ( .A(n6695), .ZN(n6135) );
  OR2_X1 U4354 ( .A1(n3115), .A2(n4835), .ZN(n5983) );
  AND2_X1 U4355 ( .A1(n4835), .A2(n6097), .ZN(n6636) );
  NAND2_X1 U4356 ( .A1(n6636), .A2(n6141), .ZN(n6179) );
  INV_X1 U4357 ( .A(n6263), .ZN(n6287) );
  NOR2_X1 U4358 ( .A1(n5988), .A2(n6956), .ZN(n6297) );
  INV_X1 U4359 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6907) );
  OR2_X1 U4360 ( .A1(n4951), .A2(n4932), .ZN(n6708) );
  AOI21_X1 U4361 ( .B1(n6907), .B2(STATE2_REG_3__SCAN_IN), .A(n6220), .ZN(
        n6638) );
  OR2_X1 U4362 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4089) );
  INV_X1 U4363 ( .A(n4697), .ZN(n6448) );
  AND3_X1 U4364 ( .A1(n4809), .A2(EBX_REG_31__SCAN_IN), .A3(n4584), .ZN(n4566)
         );
  INV_X1 U4365 ( .A(n5429), .ZN(n5441) );
  INV_X1 U4366 ( .A(n3636), .ZN(n4919) );
  INV_X1 U4367 ( .A(n6828), .ZN(n6509) );
  INV_X1 U4368 ( .A(n4785), .ZN(n4767) );
  INV_X1 U4369 ( .A(n4535), .ZN(n4536) );
  OR2_X1 U4370 ( .A1(n4335), .A2(n4192), .ZN(n6424) );
  NAND2_X1 U4371 ( .A1(n4517), .A2(n4516), .ZN(n4518) );
  INV_X1 U4372 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5829) );
  AND2_X1 U4373 ( .A1(n5006), .A2(n5009), .ZN(n6543) );
  INV_X1 U4374 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6604) );
  INV_X1 U4375 ( .A(n6522), .ZN(n6586) );
  NAND2_X1 U4376 ( .A1(n4898), .A2(n7091), .ZN(n6220) );
  NAND2_X1 U4377 ( .A1(n5986), .A2(n5985), .ZN(n6012) );
  INV_X1 U4378 ( .A(n6629), .ZN(n6093) );
  OAI221_X1 U4379 ( .B1(n6067), .B2(n6343), .C1(n6067), .C2(n6064), .A(n6304), 
        .ZN(n6089) );
  NOR2_X1 U4380 ( .A1(n6687), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6623)
         );
  NOR2_X2 U4381 ( .A1(n5983), .A2(n6335), .ZN(n6624) );
  INV_X1 U4382 ( .A(n6133), .ZN(n6172) );
  INV_X1 U4383 ( .A(n6677), .ZN(n6666) );
  INV_X1 U4384 ( .A(n6678), .ZN(n6668) );
  OR3_X1 U4385 ( .A1(n6223), .A2(n6222), .A3(n6221), .ZN(n6248) );
  INV_X1 U4386 ( .A(n6746), .ZN(n6331) );
  OAI211_X1 U4387 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6956), .A(n6304), .B(n6303), .ZN(n6327) );
  OAI21_X1 U4388 ( .B1(n6703), .B2(n6700), .A(n6699), .ZN(n6749) );
  OR2_X1 U4389 ( .A1(n6345), .A2(n6344), .ZN(n6778) );
  INV_X1 U4390 ( .A(n6715), .ZN(n6650) );
  INV_X1 U4391 ( .A(n6676), .ZN(n6767) );
  INV_X1 U4392 ( .A(n6721), .ZN(n6651) );
  INV_X1 U4393 ( .A(n6362), .ZN(n6400) );
  NOR2_X1 U4394 ( .A1(n5718), .A2(n4949), .ZN(n6652) );
  AND2_X1 U4395 ( .A1(n7079), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4189) );
  AND2_X1 U4396 ( .A1(n7091), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4564) );
  INV_X1 U4397 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4312) );
  NOR2_X2 U4398 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6824), .ZN(n4666) );
  INV_X1 U4399 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7046) );
  NOR2_X1 U4400 ( .A1(n6466), .A2(n6465), .ZN(n6818) );
  NAND2_X1 U4401 ( .A1(n5400), .A2(n4566), .ZN(n5415) );
  OR2_X1 U4402 ( .A1(n5202), .A2(n5226), .ZN(n5864) );
  NAND2_X1 U4403 ( .A1(n6495), .A2(n3636), .ZN(n5495) );
  INV_X1 U4404 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5547) );
  OR2_X1 U4405 ( .A1(n4858), .A2(n4857), .ZN(n5395) );
  INV_X1 U4406 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6944) );
  INV_X1 U4407 ( .A(n6506), .ZN(n6504) );
  INV_X1 U4408 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6904) );
  INV_X1 U4409 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n7019) );
  INV_X1 U4410 ( .A(DATAI_5_), .ZN(n7066) );
  INV_X1 U4411 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U4412 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  NAND2_X1 U4413 ( .A1(n5722), .A2(n4792), .ZN(n6541) );
  NOR2_X1 U4414 ( .A1(n4500), .A2(n4499), .ZN(n4501) );
  INV_X1 U4415 ( .A(n6812), .ZN(n6814) );
  INV_X1 U4416 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6875) );
  INV_X1 U4417 ( .A(n6056), .ZN(n6019) );
  NAND2_X1 U4418 ( .A1(n6022), .A2(n6214), .ZN(n6096) );
  NAND2_X1 U4419 ( .A1(n4895), .A2(n4894), .ZN(n6629) );
  NAND2_X1 U4420 ( .A1(n6134), .A2(n6140), .ZN(n6133) );
  INV_X1 U4421 ( .A(n6680), .ZN(n6213) );
  OR2_X1 U4422 ( .A1(n6693), .A2(n6215), .ZN(n6291) );
  NAND2_X1 U4423 ( .A1(DATAI_0_), .A2(n6063), .ZN(n6644) );
  NAND2_X1 U4424 ( .A1(DATAI_5_), .A2(n6063), .ZN(n6671) );
  OR2_X1 U4425 ( .A1(n6693), .A2(n6292), .ZN(n6746) );
  OR2_X1 U4426 ( .A1(n6693), .A2(n6335), .ZN(n6781) );
  NAND2_X1 U4427 ( .A1(n4963), .A2(n6214), .ZN(n6362) );
  NAND2_X1 U4428 ( .A1(n6536), .A2(DATAI_16_), .ZN(n6707) );
  INV_X1 U4429 ( .A(n6762), .ZN(n6735) );
  NAND2_X1 U4430 ( .A1(n6536), .A2(DATAI_26_), .ZN(n6721) );
  INV_X1 U4431 ( .A(n6681), .ZN(n6782) );
  INV_X1 U4432 ( .A(n6801), .ZN(n6796) );
  AND2_X1 U4433 ( .A1(n4641), .A2(n6824), .ZN(n6801) );
  INV_X1 U4434 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6888) );
  INV_X1 U4435 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5326) );
  INV_X1 U4436 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5230) );
  INV_X1 U4437 ( .A(n4666), .ZN(n4677) );
  OAI21_X1 U4438 ( .B1(n5811), .B2(n5750), .A(n4526), .ZN(U2962) );
  INV_X1 U4439 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4440 ( .A1(n3575), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3343) );
  AND2_X4 U4441 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5025) );
  AND2_X4 U4442 ( .A1(n5960), .A2(n5025), .ZN(n3446) );
  AND2_X2 U4443 ( .A1(n5961), .A2(n4683), .ZN(n3505) );
  AOI22_X1 U4444 ( .A1(n3505), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3438), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3340) );
  AND2_X2 U4445 ( .A1(n5961), .A2(n5025), .ZN(n3440) );
  AND2_X2 U4446 ( .A1(n4683), .A2(n4682), .ZN(n3447) );
  AOI22_X1 U4447 ( .A1(n3436), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3350) );
  AND4_X2 U4448 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3358)
         );
  AOI22_X1 U4449 ( .A1(n3505), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4450 ( .A1(n3426), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4451 ( .A1(n3506), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3438), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3353) );
  NAND2_X2 U4452 ( .A1(n3358), .A2(n3357), .ZN(n3458) );
  AOI22_X1 U4453 ( .A1(n3506), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3438), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4454 ( .A1(n3505), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4455 ( .A1(n3445), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4456 ( .A1(n3426), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4457 ( .A1(n3121), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4458 ( .A1(n3447), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3367)
         );
  AOI22_X1 U4459 ( .A1(n3575), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4460 ( .A1(n3611), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3365) );
  NAND3_X1 U4461 ( .A1(n3367), .A2(n3366), .A3(n3365), .ZN(n3368) );
  AOI22_X1 U4462 ( .A1(n3435), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4463 ( .A1(n3611), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4464 ( .A1(n3575), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4465 ( .A1(n3436), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4466 ( .A1(n3505), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4467 ( .A1(n3445), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4468 ( .A1(n3426), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4469 ( .A1(n3611), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3385)
         );
  NAND2_X1 U4470 ( .A1(n3446), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3384)
         );
  NAND2_X1 U4471 ( .A1(n3120), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4472 ( .A1(n3575), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4473 ( .A1(n3448), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4474 ( .A1(n3436), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4475 ( .A1(n3447), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3386)
         );
  NAND2_X1 U4476 ( .A1(n3505), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4477 ( .A1(n3440), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3392) );
  NAND2_X1 U4478 ( .A1(n3445), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4479 ( .A1(n3439), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4480 ( .A1(n3506), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3397) );
  NAND2_X1 U4481 ( .A1(n3426), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3396)
         );
  NAND2_X1 U4482 ( .A1(n3438), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4483 ( .A1(n3437), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3394)
         );
  NAND2_X1 U4484 ( .A1(n3611), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3405)
         );
  NAND2_X1 U4485 ( .A1(n3446), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3404)
         );
  NAND2_X1 U4486 ( .A1(n3575), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4487 ( .A1(n3099), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4488 ( .A1(n3448), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3409)
         );
  NAND2_X1 U4489 ( .A1(n3435), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4490 ( .A1(n3436), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3407) );
  NAND2_X1 U4491 ( .A1(n3447), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3406)
         );
  NAND2_X1 U4492 ( .A1(n3506), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4493 ( .A1(n3426), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3412)
         );
  NAND2_X1 U4494 ( .A1(n3440), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4495 ( .A1(n3439), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4496 ( .A1(n3445), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3417) );
  NAND2_X1 U4497 ( .A1(n3505), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3416) );
  NAND2_X1 U4498 ( .A1(n3438), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4499 ( .A1(n3437), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3414)
         );
  NAND2_X1 U4500 ( .A1(n4304), .A2(n3487), .ZN(n3433) );
  AOI22_X1 U4501 ( .A1(n3611), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4502 ( .A1(n3575), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4503 ( .A1(n3505), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4504 ( .A1(n3506), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3438), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4505 ( .A1(n3445), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4506 ( .A1(n3437), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        INSTQUEUE_REG_14__3__SCAN_IN), .B2(n3426), .ZN(n3427) );
  OR2_X1 U4507 ( .A1(n4192), .A2(n4338), .ZN(n4737) );
  NAND2_X1 U4508 ( .A1(n3433), .A2(n4737), .ZN(n3485) );
  XNOR2_X1 U4509 ( .A(n4636), .B(STATE_REG_1__SCAN_IN), .ZN(n4313) );
  NOR2_X1 U4510 ( .A1(n3434), .A2(n4313), .ZN(n3473) );
  AOI22_X1 U4511 ( .A1(n3438), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4512 ( .A1(n3440), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4513 ( .A1(n3505), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4514 ( .A1(n3448), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3449) );
  OAI21_X1 U4515 ( .B1(n3473), .B2(n4223), .A(n4950), .ZN(n3454) );
  NAND2_X1 U4516 ( .A1(n3455), .A2(n4305), .ZN(n3457) );
  NOR2_X2 U4517 ( .A1(n4453), .A2(n4941), .ZN(n4190) );
  NAND2_X1 U4518 ( .A1(n4812), .A2(n3515), .ZN(n3472) );
  AND2_X2 U4519 ( .A1(n4190), .A2(n3472), .ZN(n3467) );
  OAI21_X1 U4520 ( .B1(n4192), .B2(n4950), .A(n3476), .ZN(n3459) );
  NAND2_X1 U4521 ( .A1(n3459), .A2(n4456), .ZN(n3462) );
  INV_X1 U4522 ( .A(n4465), .ZN(n3661) );
  NAND2_X1 U4523 ( .A1(n3661), .A2(n3841), .ZN(n3461) );
  NAND2_X1 U4524 ( .A1(n3462), .A2(n3461), .ZN(n3465) );
  NAND2_X1 U4525 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  INV_X1 U4526 ( .A(n4197), .ZN(n3603) );
  NAND2_X1 U4527 ( .A1(n3603), .A2(n6372), .ZN(n3470) );
  INV_X1 U4528 ( .A(n4189), .ZN(n3602) );
  NAND2_X1 U4529 ( .A1(n3602), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4530 ( .A1(n3470), .A2(n3469), .ZN(n3481) );
  NAND2_X1 U4531 ( .A1(n4190), .A2(n3472), .ZN(n3492) );
  INV_X1 U4532 ( .A(n3473), .ZN(n3475) );
  NAND2_X1 U4533 ( .A1(n4585), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4144) );
  INV_X1 U4534 ( .A(n4144), .ZN(n3474) );
  NAND2_X1 U4535 ( .A1(n3475), .A2(n3474), .ZN(n3480) );
  MUX2_X1 U4536 ( .A(n4189), .B(n4197), .S(n6907), .Z(n3483) );
  NAND2_X1 U4537 ( .A1(n3486), .A2(n3487), .ZN(n3490) );
  NAND2_X1 U4538 ( .A1(n6442), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3488) );
  AOI21_X1 U4539 ( .B1(n3478), .B2(n4585), .A(n3488), .ZN(n3489) );
  NOR2_X1 U4540 ( .A1(n3485), .A2(n3491), .ZN(n3494) );
  NAND2_X1 U4541 ( .A1(n3492), .A2(n4449), .ZN(n3493) );
  NAND2_X1 U4542 ( .A1(n3496), .A2(n6421), .ZN(n6687) );
  INV_X1 U4543 ( .A(n3496), .ZN(n3497) );
  NAND2_X1 U4544 ( .A1(n3497), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3498) );
  NAND2_X1 U4545 ( .A1(n6687), .A2(n3498), .ZN(n5988) );
  AOI22_X1 U4546 ( .A1(n3603), .A2(n5988), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3602), .ZN(n3499) );
  AOI22_X1 U4547 ( .A1(n4099), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4548 ( .A1(n3121), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4549 ( .A1(n3519), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3502) );
  CLKBUF_X2 U4550 ( .A(n3436), .Z(n3606) );
  BUF_X1 U4551 ( .A(n3447), .Z(n3536) );
  AOI22_X1 U4552 ( .A1(n3606), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4553 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3512)
         );
  INV_X1 U4554 ( .A(n3440), .ZN(n3524) );
  INV_X2 U4555 ( .A(n3524), .ZN(n4092) );
  AOI22_X1 U4556 ( .A1(n4119), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3510) );
  INV_X1 U4557 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n7098) );
  AOI22_X1 U4558 ( .A1(n4093), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3509) );
  INV_X1 U4559 ( .A(n3439), .ZN(n5963) );
  INV_X2 U4560 ( .A(n5963), .ZN(n4100) );
  AOI22_X1 U4561 ( .A1(n4117), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4562 ( .A1(n4120), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4563 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3511)
         );
  INV_X1 U4564 ( .A(n3574), .ZN(n3565) );
  AOI22_X1 U4565 ( .A1(n4174), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3565), 
        .B2(n4201), .ZN(n3516) );
  NAND2_X1 U4566 ( .A1(n4831), .A2(n7091), .ZN(n3532) );
  AOI22_X1 U4567 ( .A1(n4099), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4568 ( .A1(n3121), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4569 ( .A1(n3519), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4570 ( .A1(n3606), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4571 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3530)
         );
  AOI22_X1 U4572 ( .A1(n4119), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4573 ( .A1(n4093), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4574 ( .A1(n4117), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4575 ( .A1(n4120), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3525) );
  NAND4_X1 U4576 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3529)
         );
  NAND2_X2 U4577 ( .A1(n3532), .A2(n3531), .ZN(n3571) );
  INV_X1 U4578 ( .A(n3533), .ZN(n3535) );
  XNOR2_X1 U4579 ( .A(n3535), .B(n3534), .ZN(n3662) );
  AOI22_X1 U4580 ( .A1(n4099), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4581 ( .A1(n3435), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4582 ( .A1(n3519), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4583 ( .A1(n3606), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3537) );
  NAND4_X1 U4584 ( .A1(n3540), .A2(n3539), .A3(n3538), .A4(n3537), .ZN(n3546)
         );
  AOI22_X1 U4585 ( .A1(n3505), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4586 ( .A1(n4093), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3438), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4587 ( .A1(n4117), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4588 ( .A1(n3426), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3541) );
  NAND4_X1 U4589 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3545)
         );
  AOI22_X1 U4590 ( .A1(n4093), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4591 ( .A1(n3519), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4592 ( .A1(n3121), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4593 ( .A1(n3438), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3437), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4594 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3557)
         );
  AOI22_X1 U4595 ( .A1(n4099), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4596 ( .A1(n3426), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4597 ( .A1(n3446), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4598 ( .A1(n3448), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4599 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3556)
         );
  NOR2_X1 U4600 ( .A1(n3573), .A2(n4276), .ZN(n3564) );
  NAND2_X1 U4601 ( .A1(n3564), .A2(n4228), .ZN(n3656) );
  OAI21_X1 U4602 ( .B1(n4273), .B2(n4228), .A(n3656), .ZN(n3562) );
  INV_X1 U4603 ( .A(n4174), .ZN(n3632) );
  AOI21_X1 U4604 ( .B1(n4936), .B2(n4276), .A(n7091), .ZN(n3560) );
  NAND2_X1 U4605 ( .A1(n3182), .A2(n4228), .ZN(n3559) );
  AOI21_X2 U4606 ( .B1(n3662), .B2(n7091), .A(n3563), .ZN(n3655) );
  AND2_X2 U4607 ( .A1(n3655), .A2(n4273), .ZN(n3569) );
  INV_X1 U4608 ( .A(n3564), .ZN(n3568) );
  NAND2_X1 U4609 ( .A1(n4174), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4610 ( .A1(n3565), .A2(n4222), .ZN(n3566) );
  INV_X1 U4611 ( .A(n3569), .ZN(n3570) );
  NOR2_X1 U4612 ( .A1(n3571), .A2(n3570), .ZN(n3572) );
  AOI21_X2 U4613 ( .B1(n3651), .B2(n3650), .A(n3572), .ZN(n3647) );
  AOI22_X1 U4614 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4099), .B1(n3446), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4615 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3121), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4616 ( .A1(n3519), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4617 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3606), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3576) );
  NAND4_X1 U4618 ( .A1(n3579), .A2(n3578), .A3(n3577), .A4(n3576), .ZN(n3585)
         );
  AOI22_X1 U4619 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4092), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4620 ( .A1(n4093), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4621 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4117), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4622 ( .A1(n4120), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3580) );
  NAND4_X1 U4623 ( .A1(n3583), .A2(n3582), .A3(n3581), .A4(n3580), .ZN(n3584)
         );
  AOI22_X1 U4624 ( .A1(n4187), .A2(n4251), .B1(n4174), .B2(
        INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4625 ( .A1(n4099), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4626 ( .A1(n3519), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4627 ( .A1(n4093), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4628 ( .A1(n4117), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4629 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3595)
         );
  AOI22_X1 U4630 ( .A1(n3435), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4631 ( .A1(n4092), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4632 ( .A1(n3117), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4633 ( .A1(n4120), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3590) );
  NAND4_X1 U4634 ( .A1(n3593), .A2(n3592), .A3(n3591), .A4(n3590), .ZN(n3594)
         );
  NAND2_X1 U4635 ( .A1(n4187), .A2(n4208), .ZN(n3597) );
  NAND2_X1 U4636 ( .A1(n4174), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4637 ( .A1(n3597), .A2(n3596), .ZN(n3699) );
  INV_X1 U4638 ( .A(n3598), .ZN(n3600) );
  NAND2_X1 U4639 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6640), .ZN(n6677) );
  NAND2_X1 U4640 ( .A1(n6982), .A2(n6677), .ZN(n3601) );
  NAND3_X1 U4641 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6366) );
  INV_X1 U4642 ( .A(n6366), .ZN(n4917) );
  AOI22_X1 U4643 ( .A1(n3603), .A2(n6218), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3602), .ZN(n3604) );
  AOI22_X1 U4644 ( .A1(n3446), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4645 ( .A1(n3519), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4646 ( .A1(n4120), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4647 ( .A1(n3606), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3607) );
  NAND4_X1 U4648 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3617)
         );
  AOI22_X1 U4649 ( .A1(n4099), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4650 ( .A1(n4119), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4651 ( .A1(n4093), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4652 ( .A1(n4117), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4653 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3616)
         );
  AOI22_X1 U4654 ( .A1(n4187), .A2(n4242), .B1(n4174), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4655 ( .A1(n4099), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4656 ( .A1(n3121), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4657 ( .A1(n3519), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4658 ( .A1(n3606), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3620) );
  NAND4_X1 U4659 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3629)
         );
  AOI22_X1 U4660 ( .A1(n4119), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3627) );
  INV_X1 U4661 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U4662 ( .A1(n4093), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4663 ( .A1(n4117), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4664 ( .A1(n4120), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4665 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3628)
         );
  AOI22_X1 U4666 ( .A1(n4187), .A2(n4265), .B1(n4174), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3689) );
  INV_X1 U4667 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3633) );
  NAND2_X1 U4668 ( .A1(n4187), .A2(n4276), .ZN(n3631) );
  OAI21_X1 U4669 ( .B1(n3633), .B2(n3632), .A(n3631), .ZN(n3634) );
  NAND2_X1 U4670 ( .A1(n4263), .A2(n3813), .ZN(n3641) );
  NAND2_X1 U4671 ( .A1(n6956), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3962) );
  NAND2_X1 U4672 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4673 ( .A1(n3701), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3694)
         );
  NAND2_X1 U4674 ( .A1(n3694), .A2(n6909), .ZN(n3637) );
  NAND2_X1 U4675 ( .A1(n3732), .A2(n3637), .ZN(n5739) );
  NAND2_X1 U4676 ( .A1(n5739), .A2(n3100), .ZN(n3638) );
  OAI21_X1 U4677 ( .B1(n6909), .B2(n3962), .A(n3638), .ZN(n3639) );
  AOI21_X1 U4678 ( .B1(n4140), .B2(EAX_REG_7__SCAN_IN), .A(n3639), .ZN(n3640)
         );
  INV_X1 U4679 ( .A(n3670), .ZN(n3683) );
  INV_X1 U4680 ( .A(n3642), .ZN(n3684) );
  INV_X1 U4681 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U4682 ( .A1(n5412), .A2(n3666), .ZN(n3643) );
  NAND2_X1 U4683 ( .A1(n3684), .A2(n3643), .ZN(n5413) );
  AOI22_X1 U4684 ( .A1(n5413), .A2(n3100), .B1(n4139), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4685 ( .A1(n4140), .A2(EAX_REG_3__SCAN_IN), .ZN(n3644) );
  OAI211_X1 U4686 ( .C1(n3683), .C2(n3339), .A(n3645), .B(n3644), .ZN(n3646)
         );
  AOI21_X1 U4687 ( .B1(n3115), .B2(n3813), .A(n3646), .ZN(n4875) );
  INV_X1 U4688 ( .A(n3647), .ZN(n3648) );
  AOI21_X1 U4689 ( .B1(n4835), .B2(n3813), .A(n4139), .ZN(n4867) );
  NAND2_X1 U4690 ( .A1(n4221), .A2(n3813), .ZN(n3654) );
  INV_X1 U4691 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4780) );
  INV_X1 U4692 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5443) );
  OAI22_X1 U4693 ( .A1(n4134), .A2(n4780), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5443), .ZN(n3652) );
  AOI21_X1 U4694 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3670), .A(n3652), 
        .ZN(n3653) );
  INV_X1 U4695 ( .A(n3655), .ZN(n3660) );
  INV_X1 U4696 ( .A(n3656), .ZN(n3658) );
  NOR2_X1 U4697 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  OR2_X2 U4698 ( .A1(n3660), .A2(n3659), .ZN(n6140) );
  AOI21_X1 U4699 ( .B1(n6140), .B2(n3661), .A(n6956), .ZN(n4790) );
  NAND2_X1 U4700 ( .A1(n6695), .A2(n3813), .ZN(n3665) );
  INV_X1 U4701 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4776) );
  INV_X1 U4702 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4793) );
  OAI22_X1 U4703 ( .A1(n4134), .A2(n4776), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4793), .ZN(n3663) );
  AOI21_X1 U4704 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3670), .A(n3663), 
        .ZN(n3664) );
  NAND2_X1 U4705 ( .A1(n3665), .A2(n3664), .ZN(n4789) );
  MUX2_X1 U4706 ( .A(n3100), .B(n4790), .S(n4789), .Z(n4806) );
  INV_X1 U4707 ( .A(n4805), .ZN(n3672) );
  INV_X1 U4708 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3668) );
  OAI21_X1 U4709 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3666), .ZN(n6540) );
  AOI22_X1 U4710 ( .A1(n4139), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3100), 
        .B2(n6540), .ZN(n3667) );
  OAI21_X1 U4711 ( .B1(n4134), .B2(n3668), .A(n3667), .ZN(n3669) );
  AOI21_X1 U4712 ( .B1(n3112), .B2(n3670), .A(n3669), .ZN(n3674) );
  INV_X1 U4713 ( .A(n3674), .ZN(n3671) );
  NAND2_X1 U4714 ( .A1(n3672), .A2(n3671), .ZN(n3673) );
  NAND2_X1 U4715 ( .A1(n4867), .A2(n3673), .ZN(n4865) );
  INV_X1 U4716 ( .A(n4864), .ZN(n4868) );
  INV_X1 U4717 ( .A(n3676), .ZN(n3678) );
  INV_X1 U4718 ( .A(n6097), .ZN(n3677) );
  NAND2_X1 U4719 ( .A1(n3678), .A2(n3677), .ZN(n3680) );
  XNOR2_X1 U4720 ( .A(n3680), .B(n3226), .ZN(n4250) );
  NAND2_X1 U4721 ( .A1(n6956), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3682)
         );
  NAND2_X1 U4722 ( .A1(n4140), .A2(EAX_REG_4__SCAN_IN), .ZN(n3681) );
  OAI211_X1 U4723 ( .C1(n3683), .C2(n6875), .A(n3682), .B(n3681), .ZN(n3687)
         );
  INV_X1 U4724 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3685) );
  NAND2_X1 U4725 ( .A1(n3685), .A2(n3684), .ZN(n3686) );
  NAND2_X1 U4726 ( .A1(n3700), .A2(n3686), .ZN(n6529) );
  MUX2_X1 U4727 ( .A(n3687), .B(n6529), .S(n3100), .Z(n3688) );
  AOI21_X1 U4728 ( .B1(n4250), .B2(n3813), .A(n3688), .ZN(n4856) );
  NAND2_X1 U4729 ( .A1(n4200), .A2(n3813), .ZN(n3698) );
  INV_X1 U4730 ( .A(n3701), .ZN(n3692) );
  INV_X1 U4731 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3691) );
  NAND2_X1 U4732 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  NAND2_X1 U4733 ( .A1(n3694), .A2(n3693), .ZN(n6521) );
  AOI22_X1 U4734 ( .A1(n6521), .A2(n3100), .B1(n4139), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3695) );
  OAI21_X1 U4735 ( .B1(n4134), .B2(n5002), .A(n3695), .ZN(n3696) );
  INV_X1 U4736 ( .A(n3696), .ZN(n3697) );
  NAND2_X1 U4737 ( .A1(n4206), .A2(n3813), .ZN(n3706) );
  AND2_X1 U4738 ( .A1(n3700), .A2(n7111), .ZN(n3702) );
  OR2_X1 U4739 ( .A1(n3702), .A2(n3701), .ZN(n5745) );
  NAND2_X1 U4740 ( .A1(n5745), .A2(n3100), .ZN(n3703) );
  OAI21_X1 U4741 ( .B1(n7111), .B2(n3962), .A(n3703), .ZN(n3704) );
  AOI21_X1 U4742 ( .B1(n4140), .B2(EAX_REG_5__SCAN_IN), .A(n3704), .ZN(n3705)
         );
  AOI22_X1 U4743 ( .A1(n4099), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4744 ( .A1(n3519), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4745 ( .A1(n4093), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4746 ( .A1(n4119), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4747 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3716)
         );
  AOI22_X1 U4748 ( .A1(n3446), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4749 ( .A1(n4092), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4750 ( .A1(n4120), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4751 ( .A1(n3606), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3711) );
  NAND4_X1 U4752 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3715)
         );
  NOR2_X1 U4753 ( .A1(n3716), .A2(n3715), .ZN(n3720) );
  NAND2_X1 U4754 ( .A1(n4140), .A2(EAX_REG_9__SCAN_IN), .ZN(n3719) );
  AOI21_X1 U4755 ( .B1(n7041), .B2(n3734), .A(n3764), .ZN(n6486) );
  INV_X1 U4756 ( .A(n6486), .ZN(n3717) );
  AOI22_X1 U4757 ( .A1(n4139), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n3100), 
        .B2(n3717), .ZN(n3718) );
  OAI211_X1 U4758 ( .C1(n3720), .C2(n3838), .A(n3719), .B(n3718), .ZN(n5483)
         );
  AOI22_X1 U4759 ( .A1(n4099), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4760 ( .A1(n4094), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4761 ( .A1(n4119), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4762 ( .A1(n4120), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4763 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3730)
         );
  AOI22_X1 U4764 ( .A1(n3435), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4765 ( .A1(n4092), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4766 ( .A1(n3519), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4767 ( .A1(n4093), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4768 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  OAI21_X1 U4769 ( .B1(n3730), .B2(n3729), .A(n3813), .ZN(n3738) );
  NAND2_X1 U4770 ( .A1(n4140), .A2(EAX_REG_8__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4771 ( .A1(n4139), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3736)
         );
  NAND2_X1 U4772 ( .A1(n3732), .A2(n3731), .ZN(n3733) );
  NAND2_X1 U4773 ( .A1(n3734), .A2(n3733), .ZN(n5731) );
  NAND2_X1 U4774 ( .A1(n5731), .A2(n3100), .ZN(n3735) );
  NAND4_X1 U4775 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n5345)
         );
  INV_X1 U4776 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5554) );
  XNOR2_X1 U4777 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3764), .ZN(n5713)
         );
  AOI22_X1 U4778 ( .A1(n3100), .A2(n5713), .B1(n4139), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3740) );
  OAI21_X1 U4779 ( .B1(n4134), .B2(n5554), .A(n3740), .ZN(n3753) );
  AOI22_X1 U4780 ( .A1(n4099), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4781 ( .A1(n3435), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4782 ( .A1(n3519), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4783 ( .A1(n4120), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4784 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3750)
         );
  AOI22_X1 U4785 ( .A1(n4093), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4786 ( .A1(n4117), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4787 ( .A1(n3446), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4788 ( .A1(n4118), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4789 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  NOR2_X1 U4790 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  NOR2_X1 U4791 ( .A1(n3838), .A2(n3751), .ZN(n3752) );
  AOI22_X1 U4792 ( .A1(n3446), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4793 ( .A1(n3519), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4794 ( .A1(n4119), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4795 ( .A1(n4118), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4796 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3763)
         );
  AOI22_X1 U4797 ( .A1(n4099), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4798 ( .A1(n4093), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4799 ( .A1(n4092), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4800 ( .A1(n3606), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4801 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  NOR2_X1 U4802 ( .A1(n3763), .A2(n3762), .ZN(n3766) );
  XNOR2_X1 U4803 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3771), .ZN(n5705)
         );
  AOI22_X1 U4804 ( .A1(n3100), .A2(n5705), .B1(n4139), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3765) );
  OAI21_X1 U4805 ( .B1(n3838), .B2(n3766), .A(n3765), .ZN(n3768) );
  NOR2_X1 U4806 ( .A1(n4134), .A2(n5552), .ZN(n3767) );
  NOR2_X1 U4807 ( .A1(n3768), .A2(n3767), .ZN(n5305) );
  INV_X1 U4808 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5550) );
  AOI21_X1 U4809 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3277), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3769) );
  INV_X1 U4810 ( .A(n3769), .ZN(n3770) );
  OAI21_X1 U4811 ( .B1(n4134), .B2(n5550), .A(n3770), .ZN(n3773) );
  NAND2_X1 U4812 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n3771), .ZN(n3796)
         );
  XNOR2_X1 U4813 ( .A(n3796), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5697)
         );
  NAND2_X1 U4814 ( .A1(n5697), .A2(n3100), .ZN(n3772) );
  NAND2_X1 U4815 ( .A1(n3773), .A2(n3772), .ZN(n3785) );
  AOI22_X1 U4816 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4094), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4817 ( .A1(n4093), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4818 ( .A1(n4120), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4819 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3606), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4820 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3783)
         );
  AOI22_X1 U4821 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4099), .B1(n3446), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4822 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3519), .B1(n3121), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4823 ( .A1(n4119), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4824 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n4117), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4825 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3782)
         );
  OAI21_X1 U4826 ( .B1(n3783), .B2(n3782), .A(n3813), .ZN(n3784) );
  NAND2_X1 U4827 ( .A1(n3785), .A2(n3784), .ZN(n5293) );
  AOI22_X1 U4828 ( .A1(n3446), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4829 ( .A1(n3519), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4830 ( .A1(n4093), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4831 ( .A1(n4118), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4832 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3795)
         );
  AOI22_X1 U4833 ( .A1(n4099), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4834 ( .A1(n4120), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4835 ( .A1(n4117), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4836 ( .A1(n3606), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4837 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3794)
         );
  NOR2_X1 U4838 ( .A1(n3795), .A2(n3794), .ZN(n3800) );
  INV_X1 U4839 ( .A(n3796), .ZN(n3797) );
  INV_X1 U4840 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3798) );
  XNOR2_X1 U4841 ( .A(n3834), .B(n3798), .ZN(n5686) );
  AOI22_X1 U4842 ( .A1(n5686), .A2(n3100), .B1(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .B2(n4139), .ZN(n3799) );
  OAI21_X1 U4843 ( .B1(n3838), .B2(n3800), .A(n3799), .ZN(n3802) );
  NOR2_X1 U4844 ( .A1(n4134), .A2(n5547), .ZN(n3801) );
  NOR2_X1 U4845 ( .A1(n3802), .A2(n3801), .ZN(n5282) );
  AOI22_X1 U4846 ( .A1(n4099), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4847 ( .A1(n4120), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4848 ( .A1(n3446), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4849 ( .A1(n3519), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4850 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3815)
         );
  AOI22_X1 U4851 ( .A1(n4093), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4852 ( .A1(n3117), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4853 ( .A1(n3121), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4854 ( .A1(n4118), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4855 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3814)
         );
  OAI21_X1 U4856 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(n3821) );
  INV_X1 U4857 ( .A(n3834), .ZN(n3816) );
  NAND2_X1 U4858 ( .A1(n3816), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3818)
         );
  INV_X1 U4859 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3817) );
  XNOR2_X1 U4860 ( .A(n3818), .B(n3817), .ZN(n5679) );
  AOI22_X1 U4861 ( .A1(n5679), .A2(n3100), .B1(PHYADDRPOINTER_REG_14__SCAN_IN), 
        .B2(n4139), .ZN(n3820) );
  NAND2_X1 U4862 ( .A1(n4140), .A2(EAX_REG_14__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4863 ( .A1(n4099), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4864 ( .A1(n3435), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4865 ( .A1(n4120), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4866 ( .A1(n4119), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4867 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3832)
         );
  AOI22_X1 U4868 ( .A1(n3519), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4869 ( .A1(n4093), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4870 ( .A1(n4118), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4871 ( .A1(n3606), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3827) );
  NAND4_X1 U4872 ( .A1(n3830), .A2(n3829), .A3(n3828), .A4(n3827), .ZN(n3831)
         );
  NOR2_X1 U4873 ( .A1(n3832), .A2(n3831), .ZN(n3837) );
  NAND2_X1 U4874 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3833) );
  NAND2_X1 U4875 ( .A1(n3157), .A2(n3278), .ZN(n3835) );
  NAND2_X1 U4876 ( .A1(n3873), .A2(n3835), .ZN(n5671) );
  AOI22_X1 U4877 ( .A1(n5671), .A2(n3100), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .B2(n4139), .ZN(n3836) );
  OAI21_X1 U4878 ( .B1(n3838), .B2(n3837), .A(n3836), .ZN(n3840) );
  INV_X1 U4879 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U4880 ( .A1(n4134), .A2(n5540), .ZN(n3839) );
  NOR2_X1 U4881 ( .A1(n3840), .A2(n3839), .ZN(n5253) );
  INV_X1 U4882 ( .A(n4812), .ZN(n3842) );
  NAND3_X1 U4883 ( .A1(n3842), .A2(n3841), .A3(n3636), .ZN(n5043) );
  AOI22_X1 U4884 ( .A1(n3435), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4885 ( .A1(n3117), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4886 ( .A1(n4120), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4887 ( .A1(n4117), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4888 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3852)
         );
  AOI22_X1 U4889 ( .A1(n4099), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4890 ( .A1(n4093), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4891 ( .A1(n4118), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4892 ( .A1(n3519), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4893 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3851)
         );
  NOR2_X1 U4894 ( .A1(n3852), .A2(n3851), .ZN(n3858) );
  INV_X1 U4895 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3855) );
  INV_X1 U4896 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3872) );
  XNOR2_X1 U4897 ( .A(n3873), .B(n3872), .ZN(n5663) );
  NAND2_X1 U4898 ( .A1(n5663), .A2(n3100), .ZN(n3854) );
  NAND2_X1 U4899 ( .A1(n4139), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3853)
         );
  OAI211_X1 U4900 ( .C1(n4134), .C2(n3855), .A(n3854), .B(n3853), .ZN(n3856)
         );
  INV_X1 U4901 ( .A(n3856), .ZN(n3857) );
  OAI21_X1 U4902 ( .B1(n4109), .B2(n3858), .A(n3857), .ZN(n5240) );
  AOI22_X1 U4903 ( .A1(n4099), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4904 ( .A1(n3519), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4905 ( .A1(n3446), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4906 ( .A1(n4120), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4907 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3868)
         );
  AOI22_X1 U4908 ( .A1(n4092), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4909 ( .A1(n4093), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4910 ( .A1(n3121), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4911 ( .A1(n3606), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4912 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3867)
         );
  OR2_X1 U4913 ( .A1(n3868), .A2(n3867), .ZN(n3871) );
  INV_X1 U4914 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3869) );
  INV_X1 U4915 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5657) );
  OAI22_X1 U4916 ( .A1(n4134), .A2(n3869), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5657), .ZN(n3870) );
  AOI21_X1 U4917 ( .B1(n4136), .B2(n3871), .A(n3870), .ZN(n3875) );
  OAI21_X1 U4918 ( .B1(n3873), .B2(n3872), .A(n5657), .ZN(n3874) );
  MUX2_X1 U4919 ( .A(n3875), .B(n5655), .S(n3100), .Z(n5229) );
  AOI22_X1 U4920 ( .A1(n3121), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4921 ( .A1(n3117), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4922 ( .A1(n3519), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4923 ( .A1(n4100), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4924 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3888)
         );
  AOI22_X1 U4925 ( .A1(n4120), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4926 ( .A1(n3446), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4927 ( .A1(n4099), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3884) );
  NAND2_X1 U4928 ( .A1(n4093), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3882)
         );
  NAND2_X1 U4929 ( .A1(n3447), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3881)
         );
  AND3_X1 U4930 ( .A1(n3882), .A2(n4089), .A3(n3881), .ZN(n3883) );
  NAND4_X1 U4931 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3887)
         );
  NAND2_X1 U4932 ( .A1(n4109), .A2(n4089), .ZN(n3987) );
  OAI21_X1 U4933 ( .B1(n3888), .B2(n3887), .A(n3987), .ZN(n3891) );
  NAND2_X1 U4934 ( .A1(n4140), .A2(EAX_REG_18__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4935 ( .A1(n6956), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3889)
         );
  NAND3_X1 U4936 ( .A1(n3891), .A2(n3890), .A3(n3889), .ZN(n3893) );
  XNOR2_X1 U4937 ( .A(n3908), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5648)
         );
  NAND2_X1 U4938 ( .A1(n5648), .A2(n3100), .ZN(n3892) );
  NAND2_X1 U4939 ( .A1(n3893), .A2(n3892), .ZN(n5216) );
  AOI22_X1 U4940 ( .A1(n3121), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4941 ( .A1(n4099), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4942 ( .A1(n4093), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4943 ( .A1(n3606), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4944 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3903)
         );
  AOI22_X1 U4945 ( .A1(n3519), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4946 ( .A1(n4119), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4947 ( .A1(n4120), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4948 ( .A1(n3446), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4949 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3902)
         );
  NOR2_X1 U4950 ( .A1(n3903), .A2(n3902), .ZN(n3907) );
  INV_X1 U4951 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3904) );
  OAI22_X1 U4952 ( .A1(n4134), .A2(n3904), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3910), .ZN(n3905) );
  INV_X1 U4953 ( .A(n3905), .ZN(n3906) );
  OAI21_X1 U4954 ( .B1(n4109), .B2(n3907), .A(n3906), .ZN(n3913) );
  INV_X1 U4955 ( .A(n3908), .ZN(n3909) );
  NAND2_X1 U4956 ( .A1(n3911), .A2(n3910), .ZN(n3912) );
  NAND2_X1 U4957 ( .A1(n3964), .A2(n3912), .ZN(n5637) );
  MUX2_X1 U4958 ( .A(n3913), .B(n5637), .S(n3100), .Z(n5197) );
  AOI22_X1 U4959 ( .A1(n3519), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3919) );
  NAND2_X1 U4960 ( .A1(n4093), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3915)
         );
  NAND2_X1 U4961 ( .A1(n3606), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3914) );
  AND3_X1 U4962 ( .A1(n3915), .A2(n3914), .A3(n4089), .ZN(n3918) );
  AOI22_X1 U4963 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3446), .B1(n4120), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4964 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3120), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4965 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3925)
         );
  AOI22_X1 U4966 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4099), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4967 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3117), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4968 ( .A1(n4117), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4969 ( .A1(n4119), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4970 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3924)
         );
  OR2_X1 U4971 ( .A1(n3925), .A2(n3924), .ZN(n3926) );
  NAND2_X1 U4972 ( .A1(n3987), .A2(n3926), .ZN(n3931) );
  INV_X1 U4973 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3927) );
  OAI22_X1 U4974 ( .A1(n4134), .A2(n3927), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3275), .ZN(n3928) );
  INV_X1 U4975 ( .A(n3928), .ZN(n3930) );
  XNOR2_X1 U4976 ( .A(n3964), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5631)
         );
  AND2_X1 U4977 ( .A1(n5631), .A2(n3100), .ZN(n3929) );
  AOI21_X1 U4978 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n5183) );
  AOI22_X1 U4979 ( .A1(n4099), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4980 ( .A1(n3117), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4981 ( .A1(n4093), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4982 ( .A1(n4119), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4983 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3941)
         );
  AOI22_X1 U4984 ( .A1(n3435), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4985 ( .A1(n4092), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4986 ( .A1(n4118), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4987 ( .A1(n3519), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4988 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3940)
         );
  NOR2_X1 U4989 ( .A1(n3941), .A2(n3940), .ZN(n3968) );
  AOI22_X1 U4990 ( .A1(n4099), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4991 ( .A1(n3446), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4992 ( .A1(n4093), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4993 ( .A1(n3117), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4994 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3951)
         );
  AOI22_X1 U4995 ( .A1(n3519), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4996 ( .A1(n4119), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4997 ( .A1(n4120), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4998 ( .A1(n3121), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4999 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3950)
         );
  NOR2_X1 U5000 ( .A1(n3951), .A2(n3950), .ZN(n3969) );
  NOR2_X1 U5001 ( .A1(n3968), .A2(n3969), .ZN(n4028) );
  AOI22_X1 U5002 ( .A1(n4099), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U5003 ( .A1(n3121), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U5004 ( .A1(n3519), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U5005 ( .A1(n3606), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U5006 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3961)
         );
  AOI22_X1 U5007 ( .A1(n4119), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U5008 ( .A1(n4093), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U5009 ( .A1(n4117), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U5010 ( .A1(n4120), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U5011 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3960)
         );
  XNOR2_X1 U5012 ( .A(n4028), .B(n4027), .ZN(n3967) );
  INV_X1 U5013 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4712) );
  OAI22_X1 U5014 ( .A1(n4134), .A2(n4712), .B1(n5139), .B2(n3962), .ZN(n3963)
         );
  INV_X1 U5015 ( .A(n3963), .ZN(n3966) );
  XNOR2_X1 U5016 ( .A(n4014), .B(n5139), .ZN(n5140) );
  NAND2_X1 U5017 ( .A1(n5140), .A2(n3100), .ZN(n3965) );
  OAI211_X1 U5018 ( .C1(n3967), .C2(n4109), .A(n3966), .B(n3965), .ZN(n4522)
         );
  XNOR2_X1 U5019 ( .A(n3969), .B(n3968), .ZN(n3972) );
  INV_X1 U5020 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4699) );
  INV_X1 U5021 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5147) );
  OAI22_X1 U5022 ( .A1(n4134), .A2(n4699), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5147), .ZN(n3970) );
  INV_X1 U5023 ( .A(n3970), .ZN(n3971) );
  OAI21_X1 U5024 ( .B1(n3972), .B2(n4109), .A(n3971), .ZN(n3976) );
  INV_X1 U5025 ( .A(n3973), .ZN(n3974) );
  NAND2_X1 U5026 ( .A1(n3974), .A2(n5147), .ZN(n3975) );
  NAND2_X1 U5027 ( .A1(n4014), .A2(n3975), .ZN(n5148) );
  MUX2_X1 U5028 ( .A(n3976), .B(n5148), .S(n3100), .Z(n4531) );
  INV_X1 U5029 ( .A(n4531), .ZN(n4012) );
  AOI22_X1 U5030 ( .A1(n3446), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U5031 ( .A1(n4094), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U5032 ( .A1(n4099), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5033 ( .A1(n3117), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3977) );
  NAND4_X1 U5034 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3989)
         );
  AOI22_X1 U5035 ( .A1(n3519), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U5036 ( .A1(n4119), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3982) );
  NAND2_X1 U5037 ( .A1(n3447), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3981)
         );
  AND3_X1 U5038 ( .A1(n3982), .A2(n4089), .A3(n3981), .ZN(n3985) );
  AOI22_X1 U5039 ( .A1(n4092), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U5040 ( .A1(n4093), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U5041 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3988)
         );
  OAI21_X1 U5042 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n3992) );
  NAND2_X1 U5043 ( .A1(n4140), .A2(EAX_REG_22__SCAN_IN), .ZN(n3991) );
  NAND2_X1 U5044 ( .A1(n6956), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3990)
         );
  NAND3_X1 U5045 ( .A1(n3992), .A2(n3991), .A3(n3990), .ZN(n3994) );
  XNOR2_X1 U5046 ( .A(n4010), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5615)
         );
  NAND2_X1 U5047 ( .A1(n5615), .A2(n3100), .ZN(n3993) );
  NAND2_X1 U5048 ( .A1(n3994), .A2(n3993), .ZN(n5156) );
  AOI22_X1 U5049 ( .A1(n4099), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5050 ( .A1(n3121), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5051 ( .A1(n3519), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U5052 ( .A1(n4119), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U5053 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n4004)
         );
  AOI22_X1 U5054 ( .A1(n4093), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5055 ( .A1(n4120), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U5056 ( .A1(n4117), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U5057 ( .A1(n3117), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U5058 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4003)
         );
  OR2_X1 U5059 ( .A1(n4004), .A2(n4003), .ZN(n4007) );
  INV_X1 U5060 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4005) );
  OAI22_X1 U5061 ( .A1(n4134), .A2(n4005), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5621), .ZN(n4006) );
  AOI21_X1 U5062 ( .B1(n4136), .B2(n4007), .A(n4006), .ZN(n4011) );
  NAND2_X1 U5063 ( .A1(n4008), .A2(n5621), .ZN(n4009) );
  MUX2_X1 U5064 ( .A(n4011), .B(n5619), .S(n3100), .Z(n5172) );
  NOR2_X1 U5065 ( .A1(n4012), .A2(n4530), .ZN(n4520) );
  AND2_X1 U5066 ( .A1(n4522), .A2(n4520), .ZN(n4013) );
  NAND2_X1 U5067 ( .A1(n4015), .A2(n5127), .ZN(n4016) );
  NAND2_X1 U5068 ( .A1(n4052), .A2(n4016), .ZN(n5601) );
  AOI22_X1 U5069 ( .A1(n4119), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5070 ( .A1(n4093), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5071 ( .A1(n4117), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5072 ( .A1(n4120), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4017) );
  NAND4_X1 U5073 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4026)
         );
  AOI22_X1 U5074 ( .A1(n4099), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5075 ( .A1(n3435), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5076 ( .A1(n3519), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5077 ( .A1(n3606), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4021) );
  NAND4_X1 U5078 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4025)
         );
  NOR2_X1 U5079 ( .A1(n4026), .A2(n4025), .ZN(n4035) );
  NAND2_X1 U5080 ( .A1(n4028), .A2(n4027), .ZN(n4034) );
  XNOR2_X1 U5081 ( .A(n4035), .B(n4034), .ZN(n4031) );
  INV_X1 U5082 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4704) );
  OAI22_X1 U5083 ( .A1(n4134), .A2(n4704), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5127), .ZN(n4029) );
  INV_X1 U5084 ( .A(n4029), .ZN(n4030) );
  OAI21_X1 U5085 ( .B1(n4031), .B2(n4109), .A(n4030), .ZN(n4032) );
  MUX2_X1 U5086 ( .A(n5601), .B(n4032), .S(n4089), .Z(n4033) );
  NOR2_X1 U5087 ( .A1(n4035), .A2(n4034), .ZN(n4057) );
  AOI22_X1 U5088 ( .A1(n4099), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5089 ( .A1(n3121), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5090 ( .A1(n3519), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5091 ( .A1(n3606), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U5092 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4045)
         );
  AOI22_X1 U5093 ( .A1(n4119), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5094 ( .A1(n4093), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5095 ( .A1(n4117), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5096 ( .A1(n4120), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U5097 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  OR2_X1 U5098 ( .A1(n4045), .A2(n4044), .ZN(n4056) );
  INV_X1 U5099 ( .A(n4056), .ZN(n4046) );
  XNOR2_X1 U5100 ( .A(n4057), .B(n4046), .ZN(n4049) );
  INV_X1 U5101 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4047) );
  INV_X1 U5102 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5593) );
  OAI22_X1 U5103 ( .A1(n4134), .A2(n4047), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5593), .ZN(n4048) );
  AOI21_X1 U5104 ( .B1(n4049), .B2(n4136), .A(n4048), .ZN(n4050) );
  XNOR2_X1 U5105 ( .A(n4052), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5591)
         );
  MUX2_X1 U5106 ( .A(n4050), .B(n5591), .S(n3100), .Z(n5116) );
  INV_X1 U5107 ( .A(n4052), .ZN(n4053) );
  NAND2_X1 U5108 ( .A1(n4053), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4054)
         );
  INV_X1 U5109 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U5110 ( .A1(n4054), .A2(n5582), .ZN(n4055) );
  NAND2_X1 U5111 ( .A1(n5586), .A2(n3100), .ZN(n4072) );
  NAND2_X1 U5112 ( .A1(n4057), .A2(n4056), .ZN(n4073) );
  AOI22_X1 U5113 ( .A1(n4099), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5114 ( .A1(n4093), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5115 ( .A1(n3446), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5116 ( .A1(n3117), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5117 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4067)
         );
  AOI22_X1 U5118 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3519), .B1(n3606), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5119 ( .A1(n4094), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5120 ( .A1(n4092), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5121 ( .A1(n4120), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5122 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4066)
         );
  NOR2_X1 U5123 ( .A1(n4067), .A2(n4066), .ZN(n4074) );
  XNOR2_X1 U5124 ( .A(n4073), .B(n4074), .ZN(n4070) );
  OAI21_X1 U5125 ( .B1(n7046), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6956), 
        .ZN(n4069) );
  NAND2_X1 U5126 ( .A1(n4140), .A2(EAX_REG_27__SCAN_IN), .ZN(n4068) );
  OAI211_X1 U5127 ( .C1(n4070), .C2(n4109), .A(n4069), .B(n4068), .ZN(n4071)
         );
  XOR2_X1 U5128 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n4111), .Z(n5576) );
  NOR2_X1 U5129 ( .A1(n4074), .A2(n4073), .ZN(n4091) );
  AOI22_X1 U5130 ( .A1(n4099), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5131 ( .A1(n3121), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3099), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5132 ( .A1(n3519), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5133 ( .A1(n3606), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5134 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4084)
         );
  AOI22_X1 U5135 ( .A1(n4119), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5136 ( .A1(n4093), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5137 ( .A1(n4117), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5138 ( .A1(n4120), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U5139 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4083)
         );
  OR2_X1 U5140 ( .A1(n4084), .A2(n4083), .ZN(n4090) );
  XNOR2_X1 U5141 ( .A(n4091), .B(n4090), .ZN(n4087) );
  NAND2_X1 U5142 ( .A1(n4140), .A2(EAX_REG_28__SCAN_IN), .ZN(n4086) );
  OAI21_X1 U5143 ( .B1(n7046), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6956), 
        .ZN(n4085) );
  OAI211_X1 U5144 ( .C1(n4087), .C2(n4109), .A(n4086), .B(n4085), .ZN(n4088)
         );
  OAI21_X1 U5145 ( .B1(n5576), .B2(n4089), .A(n4088), .ZN(n5091) );
  NAND2_X1 U5146 ( .A1(n4091), .A2(n4090), .ZN(n4115) );
  AOI22_X1 U5147 ( .A1(n4093), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5148 ( .A1(n4094), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5149 ( .A1(n4118), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5150 ( .A1(n3606), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4095) );
  NAND4_X1 U5151 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4106)
         );
  AOI22_X1 U5152 ( .A1(n4099), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5153 ( .A1(n3519), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5154 ( .A1(n4120), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5155 ( .A1(n3446), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5156 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  NOR2_X1 U5157 ( .A1(n4106), .A2(n4105), .ZN(n4116) );
  XNOR2_X1 U5158 ( .A(n4115), .B(n4116), .ZN(n4110) );
  NAND2_X1 U5159 ( .A1(n6956), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4108)
         );
  NAND2_X1 U5160 ( .A1(n4140), .A2(EAX_REG_29__SCAN_IN), .ZN(n4107) );
  OAI211_X1 U5161 ( .C1(n4110), .C2(n4109), .A(n4108), .B(n4107), .ZN(n4114)
         );
  INV_X1 U5162 ( .A(n4111), .ZN(n4112) );
  OAI21_X1 U5163 ( .B1(n4113), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4196), 
        .ZN(n5564) );
  MUX2_X1 U5164 ( .A(n4114), .B(n5564), .S(n3100), .Z(n5081) );
  NOR2_X1 U5165 ( .A1(n4116), .A2(n4115), .ZN(n4132) );
  AOI22_X1 U5166 ( .A1(n4099), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5167 ( .A1(n3446), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5168 ( .A1(n4119), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5169 ( .A1(n4120), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5970), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5170 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4130)
         );
  AOI22_X1 U5171 ( .A1(n3435), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5172 ( .A1(n4093), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5173 ( .A1(n3099), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4100), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5174 ( .A1(n3519), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4125) );
  NAND4_X1 U5175 ( .A1(n4128), .A2(n4127), .A3(n4126), .A4(n4125), .ZN(n4129)
         );
  NOR2_X1 U5176 ( .A1(n4130), .A2(n4129), .ZN(n4131) );
  XNOR2_X1 U5177 ( .A(n4132), .B(n4131), .ZN(n4137) );
  INV_X1 U5178 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4133) );
  INV_X1 U5179 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5017) );
  OAI22_X1 U5180 ( .A1(n4134), .A2(n4133), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5017), .ZN(n4135) );
  AOI21_X1 U5181 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4138) );
  XNOR2_X1 U5182 ( .A(n4196), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5015)
         );
  MUX2_X1 U5183 ( .A(n4138), .B(n5015), .S(n3100), .Z(n4593) );
  AOI22_X1 U5184 ( .A1(n4140), .A2(EAX_REG_31__SCAN_IN), .B1(n4139), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4141) );
  NAND2_X1 U5185 ( .A1(n4564), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6793) );
  XNOR2_X1 U5186 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4154) );
  INV_X1 U5187 ( .A(n4154), .ZN(n4142) );
  XNOR2_X1 U5188 ( .A(n4142), .B(n4155), .ZN(n4315) );
  INV_X1 U5189 ( .A(n4315), .ZN(n4152) );
  AND2_X1 U5190 ( .A1(n6413), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4143)
         );
  NOR2_X1 U5191 ( .A1(n4155), .A2(n4143), .ZN(n4148) );
  AOI21_X1 U5192 ( .B1(n4192), .B2(n4148), .A(n4144), .ZN(n4146) );
  AOI21_X1 U5193 ( .B1(n4145), .B2(n4585), .A(n4449), .ZN(n4166) );
  OR2_X1 U5194 ( .A1(n4146), .A2(n4166), .ZN(n4151) );
  NAND2_X1 U5195 ( .A1(n4187), .A2(n4449), .ZN(n4147) );
  NAND2_X1 U5196 ( .A1(n4147), .A2(n4223), .ZN(n4153) );
  AND2_X1 U5197 ( .A1(n4187), .A2(n4148), .ZN(n4149) );
  OAI211_X1 U5198 ( .C1(n4153), .C2(n4315), .A(n4149), .B(n4151), .ZN(n4150)
         );
  NAND2_X1 U5199 ( .A1(n4155), .A2(n4154), .ZN(n4157) );
  NAND2_X1 U5200 ( .A1(n6417), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U5201 ( .A1(n4157), .A2(n4156), .ZN(n4163) );
  NAND2_X1 U5202 ( .A1(n6421), .A2(n3112), .ZN(n4164) );
  NAND2_X1 U5203 ( .A1(n5039), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4158) );
  NAND2_X1 U5204 ( .A1(n4164), .A2(n4158), .ZN(n4161) );
  XNOR2_X1 U5205 ( .A(n4163), .B(n4161), .ZN(n4316) );
  MUX2_X1 U5206 ( .A(n4174), .B(n4187), .S(n4316), .Z(n4159) );
  NOR2_X1 U5207 ( .A1(n4159), .A2(n4166), .ZN(n4160) );
  INV_X1 U5208 ( .A(n4161), .ZN(n4162) );
  NAND2_X1 U5209 ( .A1(n4163), .A2(n4162), .ZN(n4165) );
  NAND2_X1 U5210 ( .A1(n4165), .A2(n4164), .ZN(n4170) );
  XNOR2_X1 U5211 ( .A(n3339), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4168)
         );
  XNOR2_X1 U5212 ( .A(n4170), .B(n4168), .ZN(n4317) );
  NAND3_X1 U5213 ( .A1(n4166), .A2(n4187), .A3(n4316), .ZN(n4167) );
  OAI21_X1 U5214 ( .B1(n4317), .B2(n4272), .A(n4167), .ZN(n4175) );
  INV_X1 U5215 ( .A(n4168), .ZN(n4169) );
  NAND2_X1 U5216 ( .A1(n4170), .A2(n4169), .ZN(n4172) );
  NAND2_X1 U5217 ( .A1(n6982), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4171) );
  NAND2_X1 U5218 ( .A1(n4172), .A2(n4171), .ZN(n4181) );
  OR2_X1 U5219 ( .A1(n4181), .A2(n4182), .ZN(n4314) );
  AND2_X1 U5220 ( .A1(n4314), .A2(n4317), .ZN(n4173) );
  INV_X1 U5221 ( .A(n4314), .ZN(n4177) );
  AOI22_X1 U5222 ( .A1(n4184), .A2(n4177), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7091), .ZN(n4178) );
  NAND2_X1 U5223 ( .A1(n4179), .A2(n4178), .ZN(n4186) );
  NOR2_X1 U5224 ( .A1(n6875), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4180)
         );
  NAND2_X1 U5225 ( .A1(n4184), .A2(n4319), .ZN(n4185) );
  OAI21_X1 U5226 ( .B1(n3182), .B2(n3478), .A(n5043), .ZN(n4191) );
  NAND2_X1 U5227 ( .A1(n4190), .A2(n4191), .ZN(n4335) );
  NAND2_X1 U5228 ( .A1(n6698), .A2(n4197), .ZN(n5060) );
  NAND2_X1 U5229 ( .A1(n5060), .A2(n7091), .ZN(n4193) );
  INV_X1 U5230 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U5231 ( .A1(n7091), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U5232 ( .A1(n7046), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U5233 ( .A1(n4195), .A2(n4194), .ZN(n4792) );
  NAND2_X1 U5234 ( .A1(n5725), .A2(n4594), .ZN(n4198) );
  NAND2_X1 U5235 ( .A1(n6586), .A2(REIP_REG_31__SCAN_IN), .ZN(n4495) );
  OAI211_X1 U5236 ( .C1(n5722), .C2(n6910), .A(n4198), .B(n4495), .ZN(n4199)
         );
  AOI21_X1 U5237 ( .B1(n4614), .B2(n6536), .A(n4199), .ZN(n4302) );
  NAND2_X1 U5238 ( .A1(n4200), .A2(n4306), .ZN(n4205) );
  NAND2_X1 U5239 ( .A1(n4222), .A2(n4228), .ZN(n4217) );
  INV_X1 U5240 ( .A(n4201), .ZN(n4216) );
  NAND2_X1 U5241 ( .A1(n4217), .A2(n4216), .ZN(n4244) );
  NAND2_X1 U5242 ( .A1(n4244), .A2(n4242), .ZN(n4252) );
  NAND2_X1 U5243 ( .A1(n4251), .A2(n4208), .ZN(n4202) );
  OR2_X1 U5244 ( .A1(n4252), .A2(n4202), .ZN(n4264) );
  XNOR2_X1 U5245 ( .A(n4264), .B(n4265), .ZN(n4203) );
  NAND2_X1 U5246 ( .A1(n4203), .A2(n3487), .ZN(n4204) );
  NAND2_X1 U5247 ( .A1(n4205), .A2(n4204), .ZN(n4261) );
  INV_X1 U5248 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6574) );
  XNOR2_X1 U5249 ( .A(n4261), .B(n6574), .ZN(n6512) );
  INV_X1 U5250 ( .A(n4251), .ZN(n4207) );
  OR2_X1 U5251 ( .A1(n4252), .A2(n4207), .ZN(n4209) );
  XNOR2_X1 U5252 ( .A(n4209), .B(n4208), .ZN(n4210) );
  NAND2_X1 U5253 ( .A1(n4210), .A2(n3487), .ZN(n4211) );
  INV_X1 U5254 ( .A(n4986), .ZN(n4213) );
  INV_X1 U5255 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U5256 ( .A1(n4213), .A2(n4989), .ZN(n4214) );
  NAND2_X1 U5257 ( .A1(n4215), .A2(n4306), .ZN(n4220) );
  XNOR2_X1 U5258 ( .A(n4217), .B(n4216), .ZN(n4218) );
  AOI21_X1 U5259 ( .B1(n4218), .B2(n3487), .A(n4462), .ZN(n4219) );
  NAND2_X1 U5260 ( .A1(n4221), .A2(n4449), .ZN(n4227) );
  XNOR2_X1 U5261 ( .A(n4222), .B(n4228), .ZN(n4224) );
  INV_X1 U5262 ( .A(n3487), .ZN(n4229) );
  OAI211_X1 U5263 ( .C1(n4224), .C2(n4229), .A(n4451), .B(n4223), .ZN(n4225)
         );
  INV_X1 U5264 ( .A(n4225), .ZN(n4226) );
  NAND2_X1 U5265 ( .A1(n4227), .A2(n4226), .ZN(n4817) );
  OAI21_X1 U5266 ( .B1(n4229), .B2(n4228), .A(n3165), .ZN(n4230) );
  INV_X1 U5267 ( .A(n4230), .ZN(n4231) );
  OAI21_X2 U5268 ( .B1(n6140), .B2(n4272), .A(n4231), .ZN(n4791) );
  NAND2_X1 U5269 ( .A1(n4791), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4232)
         );
  INV_X1 U5270 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U5271 ( .A1(n4232), .A2(n5027), .ZN(n4234) );
  AND2_X1 U5272 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4233) );
  NAND2_X1 U5273 ( .A1(n4791), .A2(n4233), .ZN(n4235) );
  AND2_X1 U5274 ( .A1(n4234), .A2(n4235), .ZN(n4816) );
  INV_X1 U5275 ( .A(n4235), .ZN(n4236) );
  AOI21_X2 U5276 ( .B1(n4817), .B2(n4816), .A(n4236), .ZN(n6533) );
  NAND2_X1 U5277 ( .A1(n4237), .A2(n6533), .ZN(n4240) );
  NAND2_X1 U5278 ( .A1(n4238), .A2(n6604), .ZN(n4239) );
  NAND2_X1 U5279 ( .A1(n4241), .A2(n4306), .ZN(n4247) );
  INV_X1 U5280 ( .A(n4242), .ZN(n4243) );
  XNOR2_X1 U5281 ( .A(n4244), .B(n4243), .ZN(n4245) );
  NAND2_X1 U5282 ( .A1(n4245), .A2(n3487), .ZN(n4246) );
  INV_X1 U5283 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4352) );
  NAND2_X1 U5284 ( .A1(n4248), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4249)
         );
  NAND2_X1 U5285 ( .A1(n4250), .A2(n4306), .ZN(n4255) );
  XNOR2_X1 U5286 ( .A(n4252), .B(n4251), .ZN(n4253) );
  NAND2_X1 U5287 ( .A1(n4253), .A2(n3487), .ZN(n4254) );
  NAND2_X1 U5288 ( .A1(n4255), .A2(n4254), .ZN(n4257) );
  INV_X1 U5289 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4256) );
  XNOR2_X1 U5290 ( .A(n4257), .B(n4256), .ZN(n6524) );
  NAND2_X1 U5291 ( .A1(n6523), .A2(n6524), .ZN(n4983) );
  NAND2_X1 U5292 ( .A1(n4257), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4985)
         );
  NAND2_X1 U5293 ( .A1(n4983), .A2(n4258), .ZN(n4259) );
  NAND2_X1 U5294 ( .A1(n4261), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4262)
         );
  INV_X1 U5295 ( .A(n4264), .ZN(n4266) );
  NAND2_X1 U5296 ( .A1(n4266), .A2(n4265), .ZN(n4275) );
  XNOR2_X1 U5297 ( .A(n4275), .B(n4276), .ZN(n4267) );
  NAND2_X1 U5298 ( .A1(n4267), .A2(n3487), .ZN(n4268) );
  NAND2_X1 U5299 ( .A1(n4269), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4270)
         );
  NAND2_X2 U5300 ( .A1(n4271), .A2(n4274), .ZN(n4290) );
  INV_X1 U5301 ( .A(n4275), .ZN(n4277) );
  NAND3_X1 U5302 ( .A1(n4277), .A2(n3487), .A3(n4276), .ZN(n4278) );
  NAND2_X1 U5303 ( .A1(n4290), .A2(n4278), .ZN(n4279) );
  INV_X1 U5304 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6559) );
  XNOR2_X1 U5305 ( .A(n4279), .B(n6559), .ZN(n5729) );
  NAND2_X1 U5306 ( .A1(n4279), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4280)
         );
  INV_X2 U5307 ( .A(n5644), .ZN(n5641) );
  INV_X1 U5308 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5309 ( .A1(n5641), .A2(n4373), .ZN(n4281) );
  INV_X1 U5310 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5700) );
  INV_X1 U5311 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5940) );
  AND3_X1 U5312 ( .A1(n5700), .A2(n4373), .A3(n5940), .ZN(n4282) );
  OR2_X1 U5313 ( .A1(n5641), .A2(n4282), .ZN(n4283) );
  NAND2_X1 U5314 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4284) );
  INV_X1 U5315 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5928) );
  OR2_X1 U5316 ( .A1(n5641), .A2(n5928), .ZN(n5692) );
  NAND2_X1 U5317 ( .A1(n5720), .A2(n5928), .ZN(n5691) );
  XNOR2_X1 U5318 ( .A(n5720), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5684)
         );
  NAND2_X1 U5319 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4286) );
  NOR2_X1 U5320 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4288) );
  OR2_X1 U5321 ( .A1(n5641), .A2(n4288), .ZN(n4289) );
  INV_X1 U5322 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5875) );
  INV_X1 U5323 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5856) );
  NAND3_X1 U5324 ( .A1(n5829), .A2(n5856), .A3(n5878), .ZN(n4291) );
  NAND2_X1 U5325 ( .A1(n5699), .A2(n4291), .ZN(n4292) );
  NAND2_X1 U5326 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4482) );
  AND2_X1 U5327 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5813) );
  AND2_X1 U5328 ( .A1(n5838), .A2(n5813), .ZN(n4528) );
  AND2_X1 U5329 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5330 ( .A1(n4528), .A2(n4488), .ZN(n4294) );
  NOR2_X1 U5331 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5805) );
  NOR2_X1 U5332 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U5333 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5812) );
  AND3_X1 U5334 ( .A1(n5805), .A2(n5837), .A3(n5812), .ZN(n4295) );
  OR2_X1 U5335 ( .A1(n5641), .A2(n4295), .ZN(n4296) );
  NAND2_X1 U5336 ( .A1(n5720), .A2(n5572), .ZN(n4298) );
  NAND2_X1 U5337 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U5338 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4493) );
  INV_X1 U5339 ( .A(n3109), .ZN(n5597) );
  NOR2_X1 U5340 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5588)
         );
  NOR2_X1 U5341 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U5342 ( .A1(n5588), .A2(n5772), .ZN(n5567) );
  NOR2_X1 U5343 ( .A1(n5567), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5011)
         );
  NAND3_X1 U5344 ( .A1(n3102), .A2(n5011), .A3(n5751), .ZN(n4300) );
  NAND2_X1 U5345 ( .A1(n4302), .A2(n4301), .ZN(U2955) );
  INV_X1 U5346 ( .A(n5043), .ZN(n4303) );
  NAND3_X1 U5347 ( .A1(n5065), .A2(n4303), .A3(n4449), .ZN(n4322) );
  INV_X1 U5348 ( .A(n4304), .ZN(n4308) );
  NAND2_X1 U5349 ( .A1(n4306), .A2(n4305), .ZN(n4448) );
  NAND2_X1 U5350 ( .A1(n4448), .A2(n4585), .ZN(n4307) );
  AOI21_X1 U5351 ( .B1(n4308), .B2(n4812), .A(n4307), .ZN(n4458) );
  OR2_X1 U5352 ( .A1(n4335), .A2(n4458), .ZN(n4311) );
  INV_X1 U5353 ( .A(n4309), .ZN(n4310) );
  NAND2_X1 U5354 ( .A1(n4311), .A2(n4310), .ZN(n4447) );
  NAND2_X1 U5355 ( .A1(n4449), .A2(n4727), .ZN(n4320) );
  AND4_X1 U5356 ( .A1(n4317), .A2(n4316), .A3(n4315), .A4(n4314), .ZN(n4318)
         );
  NOR2_X1 U5357 ( .A1(READY_N), .A2(n5069), .ZN(n4732) );
  NAND3_X1 U5358 ( .A1(n4320), .A2(n4732), .A3(n3478), .ZN(n4321) );
  NAND3_X1 U5359 ( .A1(n4322), .A2(n4447), .A3(n4321), .ZN(n4323) );
  NAND2_X1 U5360 ( .A1(n4323), .A2(n6440), .ZN(n4330) );
  NAND2_X1 U5361 ( .A1(n4932), .A2(n4727), .ZN(n4568) );
  NAND2_X1 U5362 ( .A1(n4568), .A2(n6443), .ZN(n4326) );
  OAI211_X1 U5363 ( .C1(n4324), .C2(n4326), .A(n4585), .B(n4325), .ZN(n4327)
         );
  INV_X1 U5364 ( .A(n4327), .ZN(n4328) );
  NAND2_X2 U5365 ( .A1(n4330), .A2(n4329), .ZN(n4475) );
  NAND2_X1 U5366 ( .A1(n4561), .A2(n4809), .ZN(n4609) );
  AND2_X1 U5367 ( .A1(n4309), .A2(n4932), .ZN(n4753) );
  INV_X1 U5368 ( .A(n4753), .ZN(n6432) );
  OAI211_X1 U5369 ( .C1(n4936), .C2(n4332), .A(n6424), .B(n6432), .ZN(n4333)
         );
  INV_X1 U5370 ( .A(n4333), .ZN(n4336) );
  NAND3_X1 U5371 ( .A1(n4609), .A2(n4336), .A3(n5063), .ZN(n4337) );
  INV_X1 U5372 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U5373 ( .A1(n4348), .A2(n4339), .ZN(n4341) );
  INV_X1 U5374 ( .A(n4349), .ZN(n4375) );
  NAND2_X1 U5375 ( .A1(n4341), .A2(n4340), .ZN(n4342) );
  OAI21_X2 U5376 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n4798), .A(n4342), 
        .ZN(n4347) );
  INV_X1 U5377 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4344) );
  OR2_X1 U5378 ( .A1(n4343), .A2(n4344), .ZN(n4346) );
  INV_X1 U5379 ( .A(n4375), .ZN(n5184) );
  NAND2_X1 U5380 ( .A1(n4349), .A2(n4344), .ZN(n4345) );
  NAND2_X1 U5381 ( .A1(n4346), .A2(n4345), .ZN(n4799) );
  MUX2_X1 U5382 ( .A(n4427), .B(n3119), .S(EBX_REG_2__SCAN_IN), .Z(n4351) );
  OR2_X1 U5383 ( .A1(n4798), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4350)
         );
  NAND2_X1 U5384 ( .A1(n4906), .A2(n3334), .ZN(n4880) );
  NAND2_X1 U5385 ( .A1(n4343), .A2(n4352), .ZN(n4354) );
  INV_X1 U5386 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4355) );
  NAND2_X1 U5387 ( .A1(n4809), .A2(n4355), .ZN(n4353) );
  NAND3_X1 U5388 ( .A1(n4354), .A2(n3119), .A3(n4353), .ZN(n4357) );
  NAND2_X1 U5389 ( .A1(n4349), .A2(n4355), .ZN(n4356) );
  AND2_X1 U5390 ( .A1(n4357), .A2(n4356), .ZN(n4882) );
  INV_X1 U5391 ( .A(n4882), .ZN(n4358) );
  MUX2_X1 U5392 ( .A(n4427), .B(n3119), .S(EBX_REG_4__SCAN_IN), .Z(n4359) );
  OAI21_X1 U5393 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4798), .A(n4359), 
        .ZN(n4861) );
  NAND2_X1 U5394 ( .A1(n4429), .A2(n4989), .ZN(n4361) );
  INV_X1 U5395 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5396 ( .A1(n4809), .A2(n5496), .ZN(n4360) );
  NAND3_X1 U5397 ( .A1(n4361), .A2(n3119), .A3(n4360), .ZN(n4363) );
  NAND2_X1 U5398 ( .A1(n4349), .A2(n5496), .ZN(n4362) );
  NAND2_X1 U5399 ( .A1(n4363), .A2(n4362), .ZN(n4996) );
  MUX2_X1 U5400 ( .A(n4427), .B(n3119), .S(EBX_REG_6__SCAN_IN), .Z(n4365) );
  OR2_X1 U5401 ( .A1(n4798), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4364)
         );
  NAND2_X1 U5402 ( .A1(n4343), .A2(n7012), .ZN(n4367) );
  INV_X1 U5403 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U5404 ( .A1(n4809), .A2(n4368), .ZN(n4366) );
  NAND3_X1 U5405 ( .A1(n4367), .A2(n3119), .A3(n4366), .ZN(n4370) );
  NAND2_X1 U5406 ( .A1(n5184), .A2(n4368), .ZN(n4369) );
  AND2_X1 U5407 ( .A1(n4370), .A2(n4369), .ZN(n5357) );
  MUX2_X1 U5408 ( .A(n4427), .B(n3119), .S(EBX_REG_8__SCAN_IN), .Z(n4372) );
  OAI21_X1 U5409 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n4798), .A(n4372), 
        .ZN(n5337) );
  NAND2_X1 U5410 ( .A1(n4429), .A2(n4373), .ZN(n4376) );
  INV_X1 U5411 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U5412 ( .A1(n4809), .A2(n5487), .ZN(n4374) );
  NAND3_X1 U5413 ( .A1(n4376), .A2(n3119), .A3(n4374), .ZN(n4378) );
  NAND2_X1 U5414 ( .A1(n5184), .A2(n5487), .ZN(n4377) );
  NAND2_X1 U5415 ( .A1(n4378), .A2(n4377), .ZN(n5485) );
  INV_X1 U5416 ( .A(n4427), .ZN(n4379) );
  INV_X1 U5417 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U5418 ( .A1(n4379), .A2(n6922), .ZN(n4383) );
  NAND2_X1 U5419 ( .A1(n4809), .A2(n6922), .ZN(n4381) );
  NAND2_X1 U5420 ( .A1(n3118), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4380) );
  NAND3_X1 U5421 ( .A1(n4429), .A2(n4381), .A3(n4380), .ZN(n4382) );
  AND2_X1 U5422 ( .A1(n4383), .A2(n4382), .ZN(n5008) );
  NAND2_X1 U5423 ( .A1(n5007), .A2(n5008), .ZN(n5006) );
  MUX2_X1 U5424 ( .A(n3119), .B(n4343), .S(EBX_REG_11__SCAN_IN), .Z(n4385) );
  NAND2_X1 U5425 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4384) );
  OR2_X2 U5426 ( .A1(n5006), .A2(n5307), .ZN(n5309) );
  INV_X1 U5427 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U5428 ( .A1(n4809), .A2(n5298), .ZN(n4387) );
  NAND2_X1 U5429 ( .A1(n3118), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4386) );
  NAND3_X1 U5430 ( .A1(n4343), .A2(n4387), .A3(n4386), .ZN(n4388) );
  OAI21_X1 U5431 ( .B1(n4427), .B2(EBX_REG_12__SCAN_IN), .A(n4388), .ZN(n5295)
         );
  NOR2_X4 U5432 ( .A1(n5309), .A2(n5295), .ZN(n5294) );
  MUX2_X1 U5433 ( .A(n3118), .B(n4429), .S(EBX_REG_13__SCAN_IN), .Z(n4390) );
  NAND2_X1 U5434 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U5435 ( .A1(n4390), .A2(n4389), .ZN(n5287) );
  INV_X1 U5436 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U5437 ( .A1(n4809), .A2(n5276), .ZN(n4392) );
  NAND2_X1 U5438 ( .A1(n3118), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4391) );
  NAND3_X1 U5439 ( .A1(n4429), .A2(n4392), .A3(n4391), .ZN(n4393) );
  OAI21_X1 U5440 ( .B1(n4427), .B2(EBX_REG_14__SCAN_IN), .A(n4393), .ZN(n5270)
         );
  MUX2_X1 U5441 ( .A(n3119), .B(n4343), .S(EBX_REG_15__SCAN_IN), .Z(n4395) );
  NAND2_X1 U5442 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4394) );
  INV_X1 U5443 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5444 ( .A1(n4809), .A2(n4396), .ZN(n4398) );
  NAND2_X1 U5445 ( .A1(n3118), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4397) );
  NAND3_X1 U5446 ( .A1(n4343), .A2(n4398), .A3(n4397), .ZN(n4399) );
  OAI21_X1 U5447 ( .B1(n4427), .B2(EBX_REG_16__SCAN_IN), .A(n4399), .ZN(n5242)
         );
  MUX2_X1 U5448 ( .A(n3118), .B(n4429), .S(EBX_REG_17__SCAN_IN), .Z(n4401) );
  NAND2_X1 U5449 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5450 ( .A1(n4401), .A2(n4400), .ZN(n5225) );
  MUX2_X1 U5451 ( .A(n4427), .B(n4375), .S(EBX_REG_19__SCAN_IN), .Z(n4404) );
  OR2_X1 U5452 ( .A1(n4798), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4403)
         );
  NAND2_X1 U5453 ( .A1(n5202), .A2(n5203), .ZN(n5199) );
  NAND2_X1 U5454 ( .A1(n4798), .A2(EBX_REG_18__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5455 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U5456 ( .A1(n4406), .A2(n4405), .ZN(n5185) );
  OR2_X1 U5457 ( .A1(n5185), .A2(n3119), .ZN(n5201) );
  OR2_X1 U5458 ( .A1(n4798), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4409)
         );
  INV_X1 U5459 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U5460 ( .A1(n4809), .A2(n4407), .ZN(n4408) );
  NAND2_X1 U5461 ( .A1(n4409), .A2(n4408), .ZN(n5186) );
  NAND2_X1 U5462 ( .A1(n5201), .A2(n5186), .ZN(n4412) );
  NAND2_X1 U5463 ( .A1(n5185), .A2(n4402), .ZN(n5200) );
  INV_X1 U5464 ( .A(n5186), .ZN(n4410) );
  NAND2_X1 U5465 ( .A1(n5200), .A2(n4410), .ZN(n4411) );
  MUX2_X1 U5466 ( .A(n4427), .B(n3118), .S(EBX_REG_21__SCAN_IN), .Z(n4413) );
  OAI21_X1 U5467 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4798), .A(n4413), 
        .ZN(n5173) );
  MUX2_X1 U5468 ( .A(n4375), .B(n4343), .S(EBX_REG_22__SCAN_IN), .Z(n4415) );
  NAND2_X1 U5469 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4414) );
  INV_X1 U5470 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U5471 ( .A1(n4809), .A2(n5470), .ZN(n4417) );
  NAND2_X1 U5472 ( .A1(n4375), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4416) );
  NAND3_X1 U5473 ( .A1(n4429), .A2(n4417), .A3(n4416), .ZN(n4418) );
  OAI21_X1 U5474 ( .B1(n4427), .B2(EBX_REG_23__SCAN_IN), .A(n4418), .ZN(n4542)
         );
  MUX2_X1 U5475 ( .A(n4375), .B(n4343), .S(EBX_REG_24__SCAN_IN), .Z(n4420) );
  NAND2_X1 U5476 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4419) );
  NAND2_X2 U5477 ( .A1(n4543), .A2(n4421), .ZN(n5138) );
  MUX2_X1 U5478 ( .A(n4427), .B(n4375), .S(EBX_REG_25__SCAN_IN), .Z(n4422) );
  OAI21_X1 U5479 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4798), .A(n4422), 
        .ZN(n5126) );
  NAND2_X1 U5480 ( .A1(n4343), .A2(n5574), .ZN(n4424) );
  INV_X1 U5481 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U5482 ( .A1(n4809), .A2(n5466), .ZN(n4423) );
  NAND3_X1 U5483 ( .A1(n4424), .A2(n4375), .A3(n4423), .ZN(n4426) );
  NAND2_X1 U5484 ( .A1(n4426), .A2(n4425), .ZN(n5112) );
  MUX2_X1 U5485 ( .A(n4427), .B(n4375), .S(EBX_REG_27__SCAN_IN), .Z(n4428) );
  OAI21_X1 U5486 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4798), .A(n4428), 
        .ZN(n5105) );
  NAND2_X1 U5487 ( .A1(n4429), .A2(n3218), .ZN(n4432) );
  INV_X1 U5488 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U5489 ( .A1(n4809), .A2(n4430), .ZN(n4431) );
  NAND3_X1 U5490 ( .A1(n4432), .A2(n4375), .A3(n4431), .ZN(n4434) );
  OR2_X1 U5491 ( .A1(n4375), .A2(EBX_REG_28__SCAN_IN), .ZN(n4433) );
  OR2_X1 U5492 ( .A1(n4798), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4436)
         );
  INV_X1 U5493 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U5494 ( .A1(n4809), .A2(n5463), .ZN(n4435) );
  AND2_X1 U5495 ( .A1(n4436), .A2(n4435), .ZN(n5072) );
  NOR2_X1 U5496 ( .A1(n4375), .A2(EBX_REG_29__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U5497 ( .A1(n4555), .A2(n4375), .B1(n5073), .B2(n4553), .ZN(n5078)
         );
  NAND2_X1 U5498 ( .A1(n4798), .A2(EBX_REG_30__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U5499 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U5500 ( .A1(n4439), .A2(n4438), .ZN(n4554) );
  INV_X1 U5501 ( .A(n4555), .ZN(n4552) );
  OAI22_X1 U5502 ( .A1(n4798), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5054), .B2(EBX_REG_31__SCAN_IN), .ZN(n4440) );
  INV_X1 U5503 ( .A(n4442), .ZN(n4443) );
  NAND3_X1 U5504 ( .A1(n4443), .A2(n4936), .A3(n4456), .ZN(n4444) );
  NAND2_X1 U5505 ( .A1(n6405), .A2(n4444), .ZN(n4445) );
  NOR2_X1 U5506 ( .A1(n5041), .A2(n5951), .ZN(n4500) );
  NAND2_X1 U5507 ( .A1(n3182), .A2(n4449), .ZN(n5398) );
  OR2_X1 U5508 ( .A1(n5398), .A2(n3478), .ZN(n4446) );
  NAND2_X1 U5509 ( .A1(n4447), .A2(n4446), .ZN(n4734) );
  INV_X1 U5510 ( .A(n5028), .ZN(n5067) );
  NAND3_X1 U5511 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n4991) );
  NOR2_X1 U5512 ( .A1(n6574), .A2(n4991), .ZN(n5946) );
  NOR2_X1 U5513 ( .A1(n7012), .A2(n6559), .ZN(n6554) );
  NAND4_X1 U5514 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5946), .A4(n6554), .ZN(n4477)
         );
  INV_X1 U5515 ( .A(n4477), .ZN(n4469) );
  NAND2_X1 U5516 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U5517 ( .A1(n6604), .A2(n6600), .ZN(n4990) );
  NAND2_X1 U5518 ( .A1(n4469), .A2(n4990), .ZN(n5871) );
  OR2_X1 U5519 ( .A1(n6599), .A2(n5871), .ZN(n5896) );
  INV_X1 U5520 ( .A(n4450), .ZN(n4452) );
  NAND3_X1 U5521 ( .A1(n4452), .A2(n4334), .A3(n3164), .ZN(n4455) );
  NAND2_X1 U5522 ( .A1(n4453), .A2(n5184), .ZN(n4454) );
  OAI211_X1 U5523 ( .C1(n4950), .C2(n4456), .A(n4455), .B(n4454), .ZN(n4457)
         );
  NOR2_X1 U5524 ( .A1(n4458), .A2(n4457), .ZN(n4460) );
  NAND2_X1 U5525 ( .A1(n4460), .A2(n4459), .ZN(n4741) );
  NAND2_X1 U5526 ( .A1(n4941), .A2(n3182), .ZN(n4461) );
  OR2_X1 U5527 ( .A1(n5043), .A2(n4461), .ZN(n5969) );
  NAND2_X1 U5528 ( .A1(n4463), .A2(n4462), .ZN(n4464) );
  OAI211_X1 U5529 ( .C1(n4442), .C2(n4465), .A(n5969), .B(n4464), .ZN(n4466)
         );
  OR2_X1 U5530 ( .A1(n4741), .A2(n4466), .ZN(n4467) );
  AND2_X2 U5531 ( .A1(n4475), .A2(n4467), .ZN(n5894) );
  OR2_X2 U5532 ( .A1(n5917), .A2(n5894), .ZN(n4993) );
  NAND3_X1 U5533 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6605), .ZN(n5833) );
  INV_X1 U5534 ( .A(n5833), .ZN(n4468) );
  NAND2_X1 U5535 ( .A1(n4469), .A2(n4468), .ZN(n4470) );
  NAND2_X1 U5536 ( .A1(n5896), .A2(n4470), .ZN(n5938) );
  AND3_X1 U5537 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5904) );
  AND2_X1 U5538 ( .A1(n5904), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5879)
         );
  AND2_X1 U5539 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5540 ( .A1(n5879), .A2(n4471), .ZN(n4481) );
  INV_X1 U5541 ( .A(n4481), .ZN(n4472) );
  NAND2_X1 U5542 ( .A1(n5938), .A2(n4472), .ZN(n5863) );
  NOR2_X1 U5543 ( .A1(n5863), .A2(n4482), .ZN(n5836) );
  NAND2_X1 U5544 ( .A1(n5836), .A2(n5838), .ZN(n5824) );
  INV_X1 U5545 ( .A(n5813), .ZN(n4486) );
  OR2_X2 U5546 ( .A1(n5824), .A2(n4486), .ZN(n5806) );
  INV_X1 U5547 ( .A(n4488), .ZN(n4508) );
  OR2_X2 U5548 ( .A1(n5806), .A2(n4508), .ZN(n5799) );
  NOR2_X1 U5549 ( .A1(n5572), .A2(n5574), .ZN(n4491) );
  INV_X1 U5550 ( .A(n4491), .ZN(n4473) );
  NOR2_X1 U5551 ( .A1(n5799), .A2(n4473), .ZN(n5770) );
  NAND2_X1 U5552 ( .A1(n5770), .A2(n5771), .ZN(n5760) );
  NOR3_X1 U5553 ( .A1(n5760), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4493), 
        .ZN(n4498) );
  INV_X1 U5554 ( .A(n4993), .ZN(n4474) );
  NAND2_X1 U5555 ( .A1(n4474), .A2(n6599), .ZN(n4822) );
  INV_X1 U5556 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U5557 ( .A1(n5894), .A2(n7015), .ZN(n4476) );
  OR2_X1 U5558 ( .A1(n4475), .A2(n6586), .ZN(n4819) );
  NAND2_X1 U5559 ( .A1(n4476), .A2(n4819), .ZN(n4992) );
  INV_X1 U5560 ( .A(n4992), .ZN(n5926) );
  NAND2_X1 U5561 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4994) );
  NOR2_X1 U5562 ( .A1(n4994), .A2(n4477), .ZN(n5916) );
  INV_X1 U5563 ( .A(n5916), .ZN(n4478) );
  NAND2_X1 U5564 ( .A1(n4993), .A2(n4478), .ZN(n4479) );
  NAND2_X1 U5565 ( .A1(n5926), .A2(n4479), .ZN(n5874) );
  AND2_X1 U5566 ( .A1(n4993), .A2(n4481), .ZN(n4480) );
  NOR2_X1 U5567 ( .A1(n5874), .A2(n4480), .ZN(n5831) );
  OR2_X1 U5568 ( .A1(n5871), .A2(n4481), .ZN(n5830) );
  NOR2_X1 U5569 ( .A1(n5830), .A2(n4482), .ZN(n4483) );
  NAND2_X1 U5570 ( .A1(n5838), .A2(n4483), .ZN(n4484) );
  NAND2_X1 U5571 ( .A1(n4822), .A2(n4484), .ZN(n4485) );
  NAND2_X1 U5572 ( .A1(n5831), .A2(n4485), .ZN(n5821) );
  AND2_X1 U5573 ( .A1(n4822), .A2(n4486), .ZN(n4487) );
  INV_X1 U5574 ( .A(n6605), .ZN(n4489) );
  AOI21_X1 U5575 ( .B1(n4489), .B2(n6599), .A(n4488), .ZN(n4490) );
  NOR2_X1 U5576 ( .A1(n4547), .A2(n4490), .ZN(n5804) );
  OAI21_X1 U5577 ( .B1(n5950), .B2(n4491), .A(n5804), .ZN(n5780) );
  INV_X1 U5578 ( .A(n5771), .ZN(n4492) );
  NOR2_X1 U5579 ( .A1(n5780), .A2(n4492), .ZN(n5762) );
  INV_X1 U5580 ( .A(n4493), .ZN(n4494) );
  INV_X1 U5581 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5026) );
  INV_X1 U5582 ( .A(n5804), .ZN(n5796) );
  NOR2_X1 U5583 ( .A1(n5796), .A2(n4822), .ZN(n5761) );
  AOI211_X1 U5584 ( .C1(n5762), .C2(n4494), .A(n5026), .B(n5761), .ZN(n4497)
         );
  INV_X1 U5585 ( .A(n4495), .ZN(n4496) );
  OAI21_X1 U5586 ( .B1(n4502), .B2(n5957), .A(n4501), .ZN(U2987) );
  XNOR2_X1 U5587 ( .A(n5641), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5634)
         );
  INV_X1 U5588 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6995) );
  XNOR2_X1 U5589 ( .A(n5641), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5626)
         );
  INV_X1 U5590 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4504) );
  XNOR2_X1 U5591 ( .A(n5699), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5618)
         );
  INV_X1 U5592 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4514) );
  INV_X1 U5593 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U5594 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4512) );
  NOR4_X1 U5595 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n7077), 
        .A4(n4512), .ZN(n4506) );
  AOI21_X1 U5596 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4514), .A(n4506), 
        .ZN(n4507) );
  NOR2_X1 U5597 ( .A1(n5608), .A2(n4507), .ZN(n4519) );
  NOR2_X1 U5598 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5605)
         );
  INV_X1 U5599 ( .A(n5605), .ZN(n4510) );
  INV_X1 U5600 ( .A(n5805), .ZN(n4509) );
  OAI21_X1 U5601 ( .B1(n4510), .B2(n4509), .A(n4508), .ZN(n4511) );
  INV_X1 U5602 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7060) );
  NOR3_X1 U5603 ( .A1(n5699), .A2(n7077), .A3(n4512), .ZN(n4513) );
  AOI211_X1 U5604 ( .C1(n5605), .C2(n4514), .A(n7060), .B(n4513), .ZN(n4515)
         );
  INV_X1 U5605 ( .A(n4515), .ZN(n4516) );
  AND2_X1 U5606 ( .A1(n4529), .A2(n4520), .ZN(n4533) );
  OAI21_X1 U5607 ( .B1(n4533), .B2(n4522), .A(n4521), .ZN(n5516) );
  INV_X1 U5608 ( .A(n5516), .ZN(n4525) );
  INV_X1 U5609 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4649) );
  NOR2_X1 U5610 ( .A1(n6522), .A2(n4649), .ZN(n5808) );
  AOI21_X1 U5611 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5808), 
        .ZN(n4523) );
  OAI21_X1 U5612 ( .B1(n5140), .B2(n6541), .A(n4523), .ZN(n4524) );
  AOI21_X1 U5613 ( .B1(n4525), .B2(n6536), .A(n4524), .ZN(n4526) );
  INV_X1 U5614 ( .A(n5625), .ZN(n4527) );
  NAND2_X1 U5615 ( .A1(n4540), .A2(n6535), .ZN(n4539) );
  INV_X1 U5616 ( .A(n4529), .ZN(n5182) );
  NOR2_X1 U5617 ( .A1(n5182), .A2(n4530), .ZN(n5157) );
  NOR2_X1 U5618 ( .A1(n5157), .A2(n4531), .ZN(n4532) );
  NOR2_X1 U5619 ( .A1(n6522), .A2(n3239), .ZN(n4546) );
  NOR2_X1 U5620 ( .A1(n6541), .A2(n5148), .ZN(n4534) );
  AOI211_X1 U5621 ( .C1(n6531), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4546), 
        .B(n4534), .ZN(n4535) );
  NAND2_X1 U5622 ( .A1(n4539), .A2(n4538), .ZN(U2963) );
  NAND2_X1 U5623 ( .A1(n4540), .A2(n6602), .ZN(n4551) );
  INV_X1 U5624 ( .A(n4541), .ZN(n5160) );
  INV_X1 U5625 ( .A(n4542), .ZN(n4544) );
  OAI21_X1 U5626 ( .B1(n5160), .B2(n4544), .A(n5136), .ZN(n5469) );
  NOR2_X1 U5627 ( .A1(n5806), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4545)
         );
  AOI211_X1 U5628 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n4547), .A(n4546), .B(n4545), .ZN(n4548) );
  NAND2_X1 U5629 ( .A1(n4551), .A2(n4550), .ZN(U2995) );
  AOI21_X1 U5630 ( .B1(n4552), .B2(n4553), .A(n4554), .ZN(n4560) );
  INV_X1 U5631 ( .A(n4553), .ZN(n4557) );
  INV_X1 U5632 ( .A(n4554), .ZN(n4556) );
  AOI211_X1 U5633 ( .C1(n5184), .C2(n4557), .A(n4556), .B(n4555), .ZN(n4558)
         );
  AOI21_X1 U5634 ( .B1(n4560), .B2(n4559), .A(n4558), .ZN(n4602) );
  INV_X1 U5635 ( .A(n4602), .ZN(n5756) );
  NAND2_X1 U5636 ( .A1(n4561), .A2(n4585), .ZN(n5064) );
  INV_X1 U5637 ( .A(n5069), .ZN(n4562) );
  NAND2_X1 U5638 ( .A1(n4309), .A2(n4562), .ZN(n4679) );
  NAND2_X1 U5639 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .ZN(n4563) );
  NAND2_X1 U5640 ( .A1(n4564), .A2(n3100), .ZN(n6444) );
  NAND3_X1 U5641 ( .A1(n6522), .A2(n6783), .A3(n6444), .ZN(n4565) );
  NOR2_X1 U5642 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4567) );
  INV_X1 U5643 ( .A(n4567), .ZN(n4584) );
  AND3_X1 U5644 ( .A1(n4568), .A2(n4567), .A3(n4585), .ZN(n4569) );
  INV_X1 U5645 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4667) );
  INV_X1 U5646 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7002) );
  INV_X1 U5647 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6978) );
  NAND3_X1 U5648 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5401) );
  NOR2_X1 U5649 ( .A1(n4670), .A2(n5401), .ZN(n5378) );
  NAND2_X1 U5650 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5378), .ZN(n5362) );
  NOR3_X1 U5651 ( .A1(n7002), .A2(n6978), .A3(n5362), .ZN(n5339) );
  NAND2_X1 U5652 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5339), .ZN(n5340) );
  NOR2_X1 U5653 ( .A1(n4667), .A2(n5340), .ZN(n5325) );
  AND2_X1 U5654 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5325), .ZN(n5313) );
  NAND2_X1 U5655 ( .A1(n5296), .A2(REIP_REG_12__SCAN_IN), .ZN(n4570) );
  AND2_X1 U5656 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n4572) );
  NAND3_X1 U5657 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4574) );
  AND2_X1 U5658 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5188) );
  NAND2_X1 U5659 ( .A1(n5188), .A2(REIP_REG_20__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5660 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n4571) );
  NOR2_X1 U5661 ( .A1(n5174), .A2(n4571), .ZN(n5151) );
  NAND2_X1 U5662 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n4577) );
  INV_X1 U5663 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5563) );
  NOR3_X1 U5664 ( .A1(n5084), .A2(REIP_REG_30__SCAN_IN), .A3(n5563), .ZN(n4592) );
  NAND2_X1 U5665 ( .A1(n5429), .A2(n5420), .ZN(n5459) );
  AND3_X1 U5666 ( .A1(n5296), .A2(REIP_REG_12__SCAN_IN), .A3(n4572), .ZN(n4573) );
  NAND2_X1 U5667 ( .A1(n5420), .A2(n4573), .ZN(n5243) );
  NOR2_X1 U5668 ( .A1(n5243), .A2(n4574), .ZN(n5207) );
  INV_X1 U5669 ( .A(n4575), .ZN(n4576) );
  AND2_X1 U5670 ( .A1(n5207), .A2(n4576), .ZN(n5163) );
  NAND4_X1 U5671 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5163), .ZN(n5129) );
  NOR2_X1 U5672 ( .A1(n4577), .A2(n5129), .ZN(n4578) );
  NAND2_X1 U5673 ( .A1(REIP_REG_26__SCAN_IN), .A2(n4578), .ZN(n4579) );
  NAND2_X1 U5674 ( .A1(n5459), .A2(n4579), .ZN(n5118) );
  NAND2_X1 U5675 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4580) );
  NAND2_X1 U5676 ( .A1(n5441), .A2(n4580), .ZN(n4581) );
  NAND2_X1 U5677 ( .A1(n5118), .A2(n4581), .ZN(n5093) );
  NOR2_X1 U5678 ( .A1(n5429), .A2(REIP_REG_29__SCAN_IN), .ZN(n4582) );
  NOR2_X1 U5679 ( .A1(n5093), .A2(n4582), .ZN(n4615) );
  INV_X1 U5680 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U5681 ( .A1(n4594), .A2(n7079), .ZN(n4583) );
  AOI22_X1 U5682 ( .A1(n6487), .A2(n5015), .B1(n5454), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4590) );
  OR2_X1 U5683 ( .A1(n4727), .A2(n4584), .ZN(n6404) );
  AND2_X1 U5684 ( .A1(n3487), .A2(n6404), .ZN(n4616) );
  INV_X1 U5685 ( .A(n4616), .ZN(n4587) );
  INV_X1 U5686 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5042) );
  NAND3_X1 U5687 ( .A1(n4585), .A2(n5042), .A3(n4584), .ZN(n4586) );
  NAND2_X1 U5688 ( .A1(n4587), .A2(n4586), .ZN(n4588) );
  AND2_X2 U5689 ( .A1(n5400), .A2(n4588), .ZN(n6480) );
  NAND2_X1 U5690 ( .A1(n6480), .A2(EBX_REG_30__SCAN_IN), .ZN(n4589) );
  OAI211_X1 U5691 ( .C1(n4615), .C2(n4675), .A(n4590), .B(n4589), .ZN(n4591)
         );
  AOI211_X1 U5692 ( .C1(n5756), .C2(n6473), .A(n4592), .B(n4591), .ZN(n4596)
         );
  XNOR2_X2 U5693 ( .A(n5080), .B(n3296), .ZN(n5020) );
  NAND2_X1 U5694 ( .A1(n4596), .A2(n4595), .ZN(U2797) );
  NOR2_X1 U5695 ( .A1(n5028), .A2(n6788), .ZN(n4597) );
  NAND2_X1 U5696 ( .A1(n5065), .A2(n4597), .ZN(n4601) );
  NAND4_X1 U5697 ( .A1(n4919), .A2(n4936), .A3(n6440), .A4(n3635), .ZN(n4606)
         );
  INV_X1 U5698 ( .A(n4606), .ZN(n4598) );
  NAND3_X1 U5699 ( .A1(n4599), .A2(n4809), .A3(n4598), .ZN(n4600) );
  INV_X1 U5700 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6923) );
  OAI22_X1 U5701 ( .A1(n4602), .A2(n5497), .B1(n6495), .B2(n6923), .ZN(n4603)
         );
  INV_X1 U5702 ( .A(n4604), .ZN(U2829) );
  INV_X1 U5703 ( .A(n4732), .ZN(n4605) );
  NOR2_X1 U5704 ( .A1(n6788), .A2(n4605), .ZN(n4608) );
  NOR2_X1 U5705 ( .A1(n4442), .A2(n4606), .ZN(n4607) );
  AND2_X1 U5706 ( .A1(n5559), .A2(n4919), .ZN(n4611) );
  NAND2_X1 U5707 ( .A1(n4614), .A2(n4611), .ZN(n4613) );
  AOI22_X1 U5708 ( .A1(n5535), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5542), .ZN(n4612) );
  NAND2_X1 U5709 ( .A1(n4613), .A2(n4612), .ZN(U2860) );
  NAND2_X1 U5710 ( .A1(n4614), .A2(n6488), .ZN(n4622) );
  OAI21_X1 U5711 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5429), .A(n4615), .ZN(n4621) );
  INV_X1 U5712 ( .A(n5400), .ZN(n4618) );
  NAND2_X1 U5713 ( .A1(n4616), .A2(EBX_REG_31__SCAN_IN), .ZN(n4617) );
  OAI22_X1 U5714 ( .A1(n6910), .A2(n6478), .B1(n4618), .B2(n4617), .ZN(n4620)
         );
  NOR4_X1 U5715 ( .A1(n5084), .A2(REIP_REG_31__SCAN_IN), .A3(n4675), .A4(n5563), .ZN(n4619) );
  AOI21_X1 U5716 ( .B1(n4636), .B2(HOLD), .A(READY_N), .ZN(n4626) );
  INV_X1 U5717 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4640) );
  INV_X1 U5718 ( .A(HOLD), .ZN(n4624) );
  INV_X1 U5719 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7033) );
  NOR2_X1 U5720 ( .A1(n4312), .A2(n7033), .ZN(n4623) );
  OAI21_X1 U5721 ( .B1(n4636), .B2(n4624), .A(n4623), .ZN(n4625) );
  OAI211_X1 U5722 ( .C1(n4626), .C2(n4640), .A(n4727), .B(n4625), .ZN(U3182)
         );
  INV_X1 U5723 ( .A(NA_N), .ZN(n4634) );
  AOI22_X1 U5724 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4633) );
  NAND2_X1 U5725 ( .A1(STATE_REG_0__SCAN_IN), .A2(n4633), .ZN(n4635) );
  AOI22_X1 U5726 ( .A1(n4634), .A2(n4312), .B1(STATE_REG_1__SCAN_IN), .B2(
        n4635), .ZN(n4632) );
  NOR2_X1 U5727 ( .A1(NA_N), .A2(n6443), .ZN(n4627) );
  NAND4_X1 U5728 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .A3(
        REQUESTPENDING_REG_SCAN_IN), .A4(n4627), .ZN(n4631) );
  INV_X1 U5729 ( .A(n4627), .ZN(n4628) );
  AOI21_X1 U5730 ( .B1(STATE_REG_1__SCAN_IN), .B2(n4628), .A(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n4629) );
  OAI211_X1 U5731 ( .C1(n4629), .C2(STATE_REG_2__SCAN_IN), .A(HOLD), .B(
        STATE_REG_0__SCAN_IN), .ZN(n4630) );
  OAI211_X1 U5732 ( .C1(n4632), .C2(n4636), .A(n4631), .B(n4630), .ZN(U3183)
         );
  AOI21_X1 U5733 ( .B1(STATE_REG_1__SCAN_IN), .B2(HOLD), .A(n7033), .ZN(n4639)
         );
  OAI21_X1 U5734 ( .B1(n4634), .B2(STATE_REG_0__SCAN_IN), .A(n4633), .ZN(n4637) );
  AOI22_X1 U5735 ( .A1(n4637), .A2(n4640), .B1(n4636), .B2(n4635), .ZN(n4638)
         );
  OAI21_X1 U5736 ( .B1(n4639), .B2(n6797), .A(n4638), .ZN(U3181) );
  INV_X1 U5737 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4642) );
  OAI21_X1 U5738 ( .B1(n4640), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5739 ( .B1(n6797), .B2(n4642), .A(n6796), .ZN(U2789) );
  INV_X1 U5740 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4644) );
  NAND2_X2 U5741 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6797), .ZN(n4678) );
  AOI22_X1 U5742 ( .A1(n4666), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6824), .ZN(n4643) );
  OAI21_X1 U5743 ( .B1(n4644), .B2(n4678), .A(n4643), .ZN(U3188) );
  INV_X1 U5744 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5428) );
  AOI22_X1 U5745 ( .A1(n4666), .A2(REIP_REG_3__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_1__SCAN_IN), .ZN(n4645) );
  OAI21_X1 U5746 ( .B1(n5428), .B2(n4678), .A(n4645), .ZN(U3185) );
  AOI22_X1 U5747 ( .A1(n4666), .A2(REIP_REG_7__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_5__SCAN_IN), .ZN(n4646) );
  OAI21_X1 U5748 ( .B1(n6978), .B2(n4678), .A(n4646), .ZN(U3189) );
  AOI22_X1 U5749 ( .A1(n4666), .A2(REIP_REG_30__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_28__SCAN_IN), .ZN(n4647) );
  OAI21_X1 U5750 ( .B1(n5563), .B2(n4678), .A(n4647), .ZN(U3212) );
  AOI22_X1 U5751 ( .A1(n4666), .A2(REIP_REG_25__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_23__SCAN_IN), .ZN(n4648) );
  OAI21_X1 U5752 ( .B1(n4649), .B2(n4678), .A(n4648), .ZN(U3207) );
  INV_X1 U5753 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U5754 ( .A1(n4666), .A2(REIP_REG_28__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n4650) );
  OAI21_X1 U5755 ( .B1(n5109), .B2(n4678), .A(n4650), .ZN(U3210) );
  AOI22_X1 U5756 ( .A1(n4666), .A2(REIP_REG_2__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n4651) );
  OAI21_X1 U5757 ( .B1(n6888), .B2(n4678), .A(n4651), .ZN(U3184) );
  AOI22_X1 U5758 ( .A1(n4666), .A2(REIP_REG_5__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_3__SCAN_IN), .ZN(n4652) );
  OAI21_X1 U5759 ( .B1(n4670), .B2(n4678), .A(n4652), .ZN(U3187) );
  INV_X1 U5760 ( .A(REIP_REG_18__SCAN_IN), .ZN(n4668) );
  AOI22_X1 U5761 ( .A1(n4666), .A2(REIP_REG_19__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n4653) );
  OAI21_X1 U5762 ( .B1(n4668), .B2(n4678), .A(n4653), .ZN(U3201) );
  AOI22_X1 U5763 ( .A1(n4666), .A2(REIP_REG_24__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n4654) );
  OAI21_X1 U5764 ( .B1(n3239), .B2(n4678), .A(n4654), .ZN(U3206) );
  AOI22_X1 U5765 ( .A1(n4666), .A2(REIP_REG_11__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_9__SCAN_IN), .ZN(n4655) );
  OAI21_X1 U5766 ( .B1(n5326), .B2(n4678), .A(n4655), .ZN(U3193) );
  INV_X1 U5767 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6971) );
  AOI22_X1 U5768 ( .A1(n4666), .A2(REIP_REG_16__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_14__SCAN_IN), .ZN(n4656) );
  OAI21_X1 U5769 ( .B1(n6971), .B2(n4678), .A(n4656), .ZN(U3198) );
  INV_X1 U5770 ( .A(REIP_REG_20__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5771 ( .A1(n4666), .A2(REIP_REG_21__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n4657) );
  OAI21_X1 U5772 ( .B1(n4658), .B2(n4678), .A(n4657), .ZN(U3203) );
  INV_X1 U5773 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6965) );
  AOI22_X1 U5774 ( .A1(n4666), .A2(REIP_REG_14__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_12__SCAN_IN), .ZN(n4659) );
  OAI21_X1 U5775 ( .B1(n6965), .B2(n4678), .A(n4659), .ZN(U3196) );
  INV_X1 U5776 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5302) );
  AOI22_X1 U5777 ( .A1(n4666), .A2(REIP_REG_13__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n4660) );
  OAI21_X1 U5778 ( .B1(n5302), .B2(n4678), .A(n4660), .ZN(U3195) );
  INV_X1 U5779 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5780 ( .A1(n4666), .A2(REIP_REG_12__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_10__SCAN_IN), .ZN(n4661) );
  OAI21_X1 U5781 ( .B1(n4662), .B2(n4678), .A(n4661), .ZN(U3194) );
  INV_X1 U5782 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5783 ( .A1(n4666), .A2(REIP_REG_15__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_13__SCAN_IN), .ZN(n4663) );
  OAI21_X1 U5784 ( .B1(n4664), .B2(n4678), .A(n4663), .ZN(U3197) );
  INV_X1 U5785 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4669) );
  AOI22_X1 U5786 ( .A1(n4666), .A2(REIP_REG_9__SCAN_IN), .B1(n6824), .B2(
        ADDRESS_REG_7__SCAN_IN), .ZN(n4665) );
  OAI21_X1 U5787 ( .B1(n4669), .B2(n4678), .A(n4665), .ZN(U3191) );
  INV_X1 U5788 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7089) );
  OAI222_X1 U5789 ( .A1(n4677), .A2(n5326), .B1(n4678), .B2(n4667), .C1(n6797), 
        .C2(n7089), .ZN(U3192) );
  INV_X1 U5790 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6890) );
  OAI222_X1 U5791 ( .A1(n4677), .A2(n4668), .B1(n6797), .B2(n6890), .C1(n5230), 
        .C2(n4678), .ZN(U3200) );
  INV_X1 U5792 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6939) );
  INV_X1 U5793 ( .A(REIP_REG_22__SCAN_IN), .ZN(n4672) );
  OAI222_X1 U5794 ( .A1(n4677), .A2(n3239), .B1(n6797), .B2(n6939), .C1(n4678), 
        .C2(n4672), .ZN(U3205) );
  INV_X1 U5795 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6945) );
  OAI222_X1 U5796 ( .A1(n4678), .A2(n7002), .B1(n4677), .B2(n4669), .C1(n6945), 
        .C2(n6797), .ZN(U3190) );
  INV_X1 U5797 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6983) );
  INV_X1 U5798 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7082) );
  OAI222_X1 U5799 ( .A1(n4678), .A2(n6983), .B1(n4677), .B2(n4670), .C1(n7082), 
        .C2(n6797), .ZN(U3186) );
  INV_X1 U5800 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5662) );
  INV_X1 U5801 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n4671) );
  OAI222_X1 U5802 ( .A1(n4678), .A2(n5662), .B1(n4677), .B2(n5230), .C1(n6797), 
        .C2(n4671), .ZN(U3199) );
  INV_X1 U5803 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5177) );
  INV_X1 U5804 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6882) );
  OAI222_X1 U5805 ( .A1(n4678), .A2(n5177), .B1(n6797), .B2(n6882), .C1(n4677), 
        .C2(n4672), .ZN(U3204) );
  INV_X1 U5806 ( .A(REIP_REG_19__SCAN_IN), .ZN(n4673) );
  INV_X1 U5807 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7032) );
  OAI222_X1 U5808 ( .A1(n4678), .A2(n4673), .B1(n6797), .B2(n7032), .C1(n4677), 
        .C2(n4658), .ZN(U3202) );
  INV_X1 U5809 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6894) );
  INV_X1 U5810 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4674) );
  OAI222_X1 U5811 ( .A1(n4678), .A2(n4675), .B1(n6797), .B2(n6894), .C1(n4674), 
        .C2(n4677), .ZN(U3213) );
  INV_X1 U5812 ( .A(REIP_REG_25__SCAN_IN), .ZN(n4676) );
  INV_X1 U5813 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7097) );
  OAI222_X1 U5814 ( .A1(n4678), .A2(n4676), .B1(n6797), .B2(n7097), .C1(n7105), 
        .C2(n4677), .ZN(U3208) );
  INV_X1 U5815 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6881) );
  OAI222_X1 U5816 ( .A1(n4678), .A2(n7105), .B1(n6797), .B2(n6881), .C1(n5109), 
        .C2(n4677), .ZN(U3209) );
  INV_X1 U5817 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7018) );
  INV_X1 U5818 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7092) );
  OAI222_X1 U5819 ( .A1(n4678), .A2(n7018), .B1(n6797), .B2(n7092), .C1(n5563), 
        .C2(n4677), .ZN(U3211) );
  AOI22_X1 U5820 ( .A1(n5065), .A2(n4334), .B1(n5064), .B2(n4679), .ZN(n6451)
         );
  NAND3_X1 U5821 ( .A1(n5054), .A2(n4334), .A3(n4727), .ZN(n4680) );
  NAND2_X1 U5822 ( .A1(n4680), .A2(n6443), .ZN(n5057) );
  NAND2_X1 U5823 ( .A1(n6451), .A2(n5057), .ZN(n6426) );
  NAND2_X1 U5824 ( .A1(n6426), .A2(n6440), .ZN(n5070) );
  INV_X1 U5825 ( .A(n5070), .ZN(n4681) );
  OAI21_X1 U5826 ( .B1(n4681), .B2(n6957), .A(n5750), .ZN(U2793) );
  INV_X1 U5827 ( .A(n4682), .ZN(n4684) );
  OAI21_X1 U5828 ( .B1(n4684), .B2(n4683), .A(n6875), .ZN(n4685) );
  NAND2_X1 U5829 ( .A1(n4685), .A2(n6957), .ZN(n6787) );
  NAND2_X1 U5830 ( .A1(n6343), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6810) );
  AOI222_X1 U5831 ( .A1(n6787), .A2(n4693), .B1(n6214), .B2(n6691), .C1(n6695), 
        .C2(n6810), .ZN(n4691) );
  INV_X1 U5832 ( .A(n4693), .ZN(n4686) );
  NAND2_X1 U5833 ( .A1(n6787), .A2(n6957), .ZN(n4688) );
  NAND2_X1 U5834 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4693), .ZN(n6790) );
  INV_X1 U5835 ( .A(n6790), .ZN(n6802) );
  NAND2_X1 U5836 ( .A1(n4688), .A2(n6802), .ZN(n4689) );
  NAND2_X1 U5837 ( .A1(n6220), .A2(n4689), .ZN(n6812) );
  NAND2_X1 U5838 ( .A1(n6814), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4690) );
  OAI21_X1 U5839 ( .B1(n4691), .B2(n6814), .A(n4690), .ZN(U3465) );
  AND2_X1 U5840 ( .A1(n6405), .A2(n6412), .ZN(n4692) );
  NAND2_X1 U5841 ( .A1(n6506), .A2(DATAO_REG_6__SCAN_IN), .ZN(n4695) );
  INV_X2 U5842 ( .A(n6508), .ZN(n6502) );
  NAND2_X1 U5843 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6502), .ZN(n4694) );
  OAI211_X1 U5844 ( .C1(n5002), .C2(n4842), .A(n4695), .B(n4694), .ZN(U2917)
         );
  NAND2_X1 U5845 ( .A1(n6825), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4698) );
  INV_X1 U5846 ( .A(DATAI_7_), .ZN(n5557) );
  OR2_X1 U5847 ( .A1(n4785), .A2(n5557), .ZN(n4705) );
  OAI211_X1 U5848 ( .C1(n6828), .C2(n4699), .A(n4698), .B(n4705), .ZN(U2931)
         );
  INV_X1 U5849 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5850 ( .A1(n6825), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4700) );
  INV_X1 U5851 ( .A(DATAI_9_), .ZN(n5555) );
  OR2_X1 U5852 ( .A1(n4785), .A2(n5555), .ZN(n4702) );
  OAI211_X1 U5853 ( .C1(n6828), .C2(n4701), .A(n4700), .B(n4702), .ZN(U2948)
         );
  NAND2_X1 U5854 ( .A1(n6825), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4703) );
  OAI211_X1 U5855 ( .C1(n6828), .C2(n4704), .A(n4703), .B(n4702), .ZN(U2933)
         );
  INV_X1 U5856 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5857 ( .A1(n6825), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4706) );
  OAI211_X1 U5858 ( .C1(n6828), .C2(n4707), .A(n4706), .B(n4705), .ZN(U2946)
         );
  NAND2_X1 U5859 ( .A1(n6825), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U5860 ( .A1(n4767), .A2(DATAI_10_), .ZN(n4713) );
  OAI211_X1 U5861 ( .C1(n4047), .C2(n6828), .A(n4708), .B(n4713), .ZN(U2934)
         );
  INV_X1 U5862 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5863 ( .A1(n6825), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5864 ( .A1(n4767), .A2(DATAI_11_), .ZN(n4719) );
  OAI211_X1 U5865 ( .C1(n6828), .C2(n4710), .A(n4709), .B(n4719), .ZN(U2935)
         );
  NAND2_X1 U5866 ( .A1(n6825), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U5867 ( .A1(n4767), .A2(DATAI_8_), .ZN(n4721) );
  OAI211_X1 U5868 ( .C1(n6828), .C2(n4712), .A(n4711), .B(n4721), .ZN(U2932)
         );
  NAND2_X1 U5869 ( .A1(n6825), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5870 ( .C1(n5554), .C2(n6828), .A(n4714), .B(n4713), .ZN(U2949)
         );
  INV_X1 U5871 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U5872 ( .A1(n6825), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5873 ( .A1(n4767), .A2(DATAI_2_), .ZN(n6826) );
  OAI211_X1 U5874 ( .C1(n4716), .C2(n6828), .A(n4715), .B(n6826), .ZN(U2926)
         );
  INV_X1 U5875 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U5876 ( .A1(n6825), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5877 ( .A1(n4767), .A2(DATAI_14_), .ZN(n4762) );
  OAI211_X1 U5878 ( .C1(n4718), .C2(n6828), .A(n4717), .B(n4762), .ZN(U2953)
         );
  NAND2_X1 U5879 ( .A1(n6825), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4720) );
  OAI211_X1 U5880 ( .C1(n5552), .C2(n6828), .A(n4720), .B(n4719), .ZN(U2950)
         );
  INV_X1 U5881 ( .A(EAX_REG_8__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U5882 ( .A1(n6825), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4722) );
  OAI211_X1 U5883 ( .C1(n6828), .C2(n4723), .A(n4722), .B(n4721), .ZN(U2947)
         );
  INV_X1 U5884 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U5885 ( .A1(n6825), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U5886 ( .A1(n4767), .A2(DATAI_13_), .ZN(n4760) );
  OAI211_X1 U5887 ( .C1(n4725), .C2(n6828), .A(n4724), .B(n4760), .ZN(U2937)
         );
  INV_X1 U5888 ( .A(n4727), .ZN(n4726) );
  NOR2_X1 U5889 ( .A1(n4809), .A2(n4726), .ZN(n4728) );
  OAI22_X1 U5890 ( .A1(n4324), .A2(n4728), .B1(n6412), .B2(n4727), .ZN(n4730)
         );
  INV_X1 U5891 ( .A(n5063), .ZN(n4729) );
  AOI21_X1 U5892 ( .B1(n4730), .B2(n6443), .A(n4729), .ZN(n4731) );
  MUX2_X1 U5893 ( .A(n4731), .B(n5028), .S(n5065), .Z(n4736) );
  AND2_X1 U5894 ( .A1(n4753), .A2(n4732), .ZN(n4733) );
  NOR2_X1 U5895 ( .A1(n4734), .A2(n4733), .ZN(n4735) );
  NAND2_X1 U5896 ( .A1(n4736), .A2(n4735), .ZN(n6415) );
  AOI22_X1 U5897 ( .A1(n6415), .A2(n6440), .B1(FLUSH_REG_SCAN_IN), .B2(n6802), 
        .ZN(n4755) );
  NAND2_X1 U5898 ( .A1(n7091), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U5899 ( .A1(n4755), .A2(n4897), .ZN(n5981) );
  INV_X1 U5900 ( .A(n5981), .ZN(n5037) );
  AOI21_X1 U5901 ( .B1(n6442), .B2(n5973), .A(n5037), .ZN(n4744) );
  NAND2_X1 U5902 ( .A1(n4442), .A2(n4737), .ZN(n4738) );
  NOR2_X1 U5903 ( .A1(n4753), .A2(n4738), .ZN(n4739) );
  NAND2_X1 U5904 ( .A1(n4324), .A2(n4739), .ZN(n4740) );
  NOR2_X1 U5905 ( .A1(n4741), .A2(n4740), .ZN(n5959) );
  OAI22_X1 U5906 ( .A1(n6135), .A2(n5959), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5043), .ZN(n6410) );
  INV_X1 U5907 ( .A(n6784), .ZN(n5979) );
  OAI22_X1 U5908 ( .A1(n5979), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n7079), .ZN(n4742) );
  AOI21_X1 U5909 ( .B1(n6442), .B2(n6410), .A(n4742), .ZN(n4743) );
  OAI22_X1 U5910 ( .A1(n4744), .A2(n6413), .B1(n4743), .B2(n5037), .ZN(U3461)
         );
  INV_X1 U5911 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4746) );
  AOI22_X1 U5912 ( .A1(n6505), .A2(EAX_REG_9__SCAN_IN), .B1(n6502), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4745) );
  OAI21_X1 U5913 ( .B1(n6504), .B2(n4746), .A(n4745), .ZN(U2914) );
  INV_X1 U5914 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4748) );
  AOI22_X1 U5915 ( .A1(n6505), .A2(EAX_REG_8__SCAN_IN), .B1(n6502), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4747) );
  OAI21_X1 U5916 ( .B1(n6504), .B2(n4748), .A(n4747), .ZN(U2915) );
  INV_X1 U5917 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U5918 ( .A1(n6505), .A2(EAX_REG_1__SCAN_IN), .B1(n6502), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4749) );
  OAI21_X1 U5919 ( .B1(n6504), .B2(n4750), .A(n4749), .ZN(U2922) );
  INV_X1 U5920 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n7065) );
  INV_X1 U5921 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n7028) );
  OAI222_X1 U5922 ( .A1(n4842), .A2(n4707), .B1(n6504), .B2(n7065), .C1(n7028), 
        .C2(n6508), .ZN(U2916) );
  INV_X1 U5923 ( .A(n6337), .ZN(n6178) );
  NOR2_X1 U5924 ( .A1(n4751), .A2(n6178), .ZN(n4752) );
  XNOR2_X1 U5925 ( .A(n4752), .B(n6875), .ZN(n6423) );
  NAND3_X1 U5926 ( .A1(n6423), .A2(n6442), .A3(n4753), .ZN(n4754) );
  OAI22_X1 U5927 ( .A1(n5981), .A2(n6875), .B1(n4755), .B2(n4754), .ZN(U3455)
         );
  AOI222_X1 U5928 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6505), .B1(n6506), .B2(
        DATAO_REG_11__SCAN_IN), .C1(n6502), .C2(LWORD_REG_11__SCAN_IN), .ZN(
        n4756) );
  INV_X1 U5929 ( .A(n4756), .ZN(U2912) );
  AOI222_X1 U5930 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6505), .B1(n6506), .B2(
        DATAO_REG_14__SCAN_IN), .C1(n6502), .C2(LWORD_REG_14__SCAN_IN), .ZN(
        n4757) );
  INV_X1 U5931 ( .A(n4757), .ZN(U2909) );
  AOI222_X1 U5932 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6505), .B1(n6506), .B2(
        DATAO_REG_10__SCAN_IN), .C1(n6502), .C2(LWORD_REG_10__SCAN_IN), .ZN(
        n4758) );
  INV_X1 U5933 ( .A(n4758), .ZN(U2913) );
  NAND2_X1 U5934 ( .A1(n4767), .A2(DATAI_12_), .ZN(n6510) );
  NAND2_X1 U5935 ( .A1(n6509), .A2(EAX_REG_28__SCAN_IN), .ZN(n4759) );
  OAI211_X1 U5936 ( .C1(n4786), .C2(n6904), .A(n6510), .B(n4759), .ZN(U2936)
         );
  NAND2_X1 U5937 ( .A1(n6509), .A2(EAX_REG_13__SCAN_IN), .ZN(n4761) );
  OAI211_X1 U5938 ( .C1(n4786), .C2(n7013), .A(n4761), .B(n4760), .ZN(U2952)
         );
  NAND2_X1 U5939 ( .A1(n6509), .A2(EAX_REG_30__SCAN_IN), .ZN(n4763) );
  OAI211_X1 U5940 ( .C1(n4786), .C2(n7019), .A(n4763), .B(n4762), .ZN(U2938)
         );
  AOI222_X1 U5941 ( .A1(n6825), .A2(UWORD_REG_3__SCAN_IN), .B1(DATAI_3_), .B2(
        n4767), .C1(EAX_REG_19__SCAN_IN), .C2(n6509), .ZN(n4764) );
  INV_X1 U5942 ( .A(n4764), .ZN(U2927) );
  AOI222_X1 U5943 ( .A1(n6825), .A2(UWORD_REG_5__SCAN_IN), .B1(DATAI_5_), .B2(
        n4767), .C1(EAX_REG_21__SCAN_IN), .C2(n6509), .ZN(n4765) );
  INV_X1 U5944 ( .A(n4765), .ZN(U2929) );
  AOI222_X1 U5945 ( .A1(n6825), .A2(UWORD_REG_1__SCAN_IN), .B1(DATAI_1_), .B2(
        n4767), .C1(EAX_REG_17__SCAN_IN), .C2(n6509), .ZN(n4766) );
  INV_X1 U5946 ( .A(n4766), .ZN(U2925) );
  AOI222_X1 U5947 ( .A1(n6825), .A2(UWORD_REG_4__SCAN_IN), .B1(DATAI_4_), .B2(
        n4767), .C1(EAX_REG_20__SCAN_IN), .C2(n6509), .ZN(n4768) );
  INV_X1 U5948 ( .A(n4768), .ZN(U2928) );
  AOI222_X1 U5949 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6505), .B1(
        DATAO_REG_0__SCAN_IN), .B2(n6506), .C1(n6502), .C2(
        LWORD_REG_0__SCAN_IN), .ZN(n4769) );
  INV_X1 U5950 ( .A(n4769), .ZN(U2923) );
  AOI222_X1 U5951 ( .A1(EAX_REG_3__SCAN_IN), .A2(n6505), .B1(
        DATAO_REG_3__SCAN_IN), .B2(n6506), .C1(n6502), .C2(
        LWORD_REG_3__SCAN_IN), .ZN(n4770) );
  INV_X1 U5952 ( .A(n4770), .ZN(U2920) );
  AOI222_X1 U5953 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6505), .B1(
        DATAO_REG_4__SCAN_IN), .B2(n6506), .C1(n6502), .C2(
        LWORD_REG_4__SCAN_IN), .ZN(n4771) );
  INV_X1 U5954 ( .A(n4771), .ZN(U2919) );
  AOI222_X1 U5955 ( .A1(EAX_REG_2__SCAN_IN), .A2(n6505), .B1(
        DATAO_REG_2__SCAN_IN), .B2(n6506), .C1(n6502), .C2(
        LWORD_REG_2__SCAN_IN), .ZN(n4772) );
  INV_X1 U5956 ( .A(n4772), .ZN(U2921) );
  INV_X1 U5957 ( .A(DATAI_6_), .ZN(n5003) );
  INV_X1 U5958 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4774) );
  INV_X1 U5959 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4773) );
  OAI222_X1 U5960 ( .A1(n5003), .A2(n4785), .B1(n6828), .B2(n4774), .C1(n4773), 
        .C2(n4786), .ZN(U2930) );
  INV_X1 U5961 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4775) );
  INV_X1 U5962 ( .A(DATAI_0_), .ZN(n4815) );
  OAI222_X1 U5963 ( .A1(n6828), .A2(n4776), .B1(n4775), .B2(n4786), .C1(n4785), 
        .C2(n4815), .ZN(U2939) );
  INV_X1 U5964 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4778) );
  INV_X1 U5965 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4777) );
  INV_X1 U5966 ( .A(DATAI_4_), .ZN(n4884) );
  OAI222_X1 U5967 ( .A1(n6828), .A2(n4778), .B1(n4777), .B2(n4786), .C1(n4785), 
        .C2(n4884), .ZN(U2943) );
  INV_X1 U5968 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4779) );
  INV_X1 U5969 ( .A(DATAI_1_), .ZN(n6920) );
  OAI222_X1 U5970 ( .A1(n6828), .A2(n4780), .B1(n4779), .B2(n4786), .C1(n4785), 
        .C2(n6920), .ZN(U2940) );
  INV_X1 U5971 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4782) );
  INV_X1 U5972 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4781) );
  OAI222_X1 U5973 ( .A1(n6828), .A2(n4782), .B1(n4781), .B2(n4786), .C1(n4785), 
        .C2(n7066), .ZN(U2944) );
  INV_X1 U5974 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4783) );
  OAI222_X1 U5975 ( .A1(n6828), .A2(n5002), .B1(n4783), .B2(n4786), .C1(n4785), 
        .C2(n5003), .ZN(U2945) );
  INV_X1 U5976 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4784) );
  OAI222_X1 U5977 ( .A1(n4815), .A2(n4785), .B1(n4784), .B2(n4786), .C1(n6828), 
        .C2(n3855), .ZN(U2924) );
  INV_X1 U5978 ( .A(DATAI_15_), .ZN(n5539) );
  OAI222_X1 U5979 ( .A1(n5539), .A2(n4785), .B1(n6944), .B2(n4786), .C1(n5540), 
        .C2(n6828), .ZN(U2954) );
  INV_X1 U5980 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4788) );
  INV_X1 U5981 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4787) );
  INV_X1 U5982 ( .A(DATAI_3_), .ZN(n4885) );
  OAI222_X1 U5983 ( .A1(n6828), .A2(n4788), .B1(n4787), .B2(n4786), .C1(n4785), 
        .C2(n4885), .ZN(U2942) );
  XNOR2_X1 U5984 ( .A(n4790), .B(n4789), .ZN(n5461) );
  XNOR2_X1 U5985 ( .A(n4791), .B(n7015), .ZN(n4797) );
  INV_X1 U5986 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6820) );
  NOR2_X1 U5987 ( .A1(n6522), .A2(n6820), .ZN(n4802) );
  INV_X1 U5988 ( .A(n4792), .ZN(n4794) );
  AOI21_X1 U5989 ( .B1(n5722), .B2(n4794), .A(n4793), .ZN(n4795) );
  AOI211_X1 U5990 ( .C1(n4797), .C2(n6535), .A(n4802), .B(n4795), .ZN(n4796)
         );
  OAI21_X1 U5991 ( .B1(n5461), .B2(n5718), .A(n4796), .ZN(U2986) );
  INV_X1 U5992 ( .A(n4797), .ZN(n4804) );
  INV_X1 U5993 ( .A(n4798), .ZN(n4800) );
  AOI21_X1 U5994 ( .B1(n4800), .B2(n7015), .A(n4799), .ZN(n5453) );
  INV_X1 U5995 ( .A(n5917), .ZN(n5902) );
  AOI21_X1 U5996 ( .B1(n5902), .B2(n4819), .A(n7015), .ZN(n4801) );
  AOI211_X1 U5997 ( .C1(n6597), .C2(n5453), .A(n4802), .B(n4801), .ZN(n4803)
         );
  INV_X1 U5998 ( .A(n6599), .ZN(n5948) );
  OR2_X1 U5999 ( .A1(n5894), .A2(n5948), .ZN(n5900) );
  NAND2_X1 U6000 ( .A1(n5900), .A2(n7015), .ZN(n4820) );
  OAI211_X1 U6001 ( .C1(n4804), .C2(n5957), .A(n4803), .B(n4820), .ZN(U3018)
         );
  OAI21_X1 U6002 ( .B1(n4807), .B2(n4806), .A(n4805), .ZN(n4841) );
  XNOR2_X1 U6003 ( .A(n4808), .B(n4809), .ZN(n4818) );
  AOI22_X1 U6004 ( .A1(n6492), .A2(n4818), .B1(n5493), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4810) );
  OAI21_X1 U6005 ( .B1(n4841), .B2(n5490), .A(n4810), .ZN(U2858) );
  INV_X1 U6006 ( .A(n5453), .ZN(n4811) );
  OAI222_X1 U6007 ( .A1(n4811), .A2(n5497), .B1(n6495), .B2(n4344), .C1(n5490), 
        .C2(n5461), .ZN(U2859) );
  NAND2_X1 U6008 ( .A1(n4812), .A2(n3636), .ZN(n4813) );
  INV_X1 U6009 ( .A(n4813), .ZN(n4814) );
  OAI222_X1 U6010 ( .A1(n5561), .A2(n5461), .B1(n5560), .B2(n4815), .C1(n5559), 
        .C2(n4776), .ZN(U2891) );
  XNOR2_X1 U6011 ( .A(n4817), .B(n4816), .ZN(n4830) );
  AOI22_X1 U6012 ( .A1(n6597), .A2(n4818), .B1(n6586), .B2(REIP_REG_1__SCAN_IN), .ZN(n4826) );
  AND2_X1 U6013 ( .A1(n4820), .A2(n4819), .ZN(n4824) );
  NAND2_X1 U6014 ( .A1(n4822), .A2(n4821), .ZN(n4823) );
  MUX2_X1 U6015 ( .A(n4824), .B(n4823), .S(n5027), .Z(n4825) );
  OAI211_X1 U6016 ( .C1(n4830), .C2(n5957), .A(n4826), .B(n4825), .ZN(U3017)
         );
  INV_X1 U6017 ( .A(n4841), .ZN(n5450) );
  AOI22_X1 U6018 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6586), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4827) );
  OAI21_X1 U6019 ( .B1(n6541), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4827), 
        .ZN(n4828) );
  AOI21_X1 U6020 ( .B1(n5450), .B2(n6536), .A(n4828), .ZN(n4829) );
  OAI21_X1 U6021 ( .B1(n4830), .B2(n5750), .A(n4829), .ZN(U2985) );
  INV_X1 U6022 ( .A(n4221), .ZN(n6098) );
  AOI211_X1 U6023 ( .C1(n6098), .C2(n7046), .A(n6698), .B(n6635), .ZN(n4832)
         );
  AOI21_X1 U6024 ( .B1(n6810), .B2(n3116), .A(n4832), .ZN(n4834) );
  NAND2_X1 U6025 ( .A1(n6814), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4833) );
  OAI21_X1 U6026 ( .B1(n4834), .B2(n6814), .A(n4833), .ZN(U3464) );
  INV_X1 U6027 ( .A(n6635), .ZN(n6692) );
  XNOR2_X1 U6028 ( .A(n6692), .B(n4835), .ZN(n4838) );
  INV_X1 U6029 ( .A(n4837), .ZN(n5030) );
  AOI22_X1 U6030 ( .A1(n4838), .A2(n6691), .B1(n6810), .B2(n4837), .ZN(n4840)
         );
  NAND2_X1 U6031 ( .A1(n6814), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4839) );
  OAI21_X1 U6032 ( .B1(n4840), .B2(n6814), .A(n4839), .ZN(U3463) );
  OAI222_X1 U6033 ( .A1(n4841), .A2(n5561), .B1(n5560), .B2(n6920), .C1(n5559), 
        .C2(n4780), .ZN(U2890) );
  INV_X1 U6034 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4844) );
  NOR2_X2 U6035 ( .A1(n4842), .A2(n3182), .ZN(n6498) );
  AOI22_X1 U6036 ( .A1(n6498), .A2(EAX_REG_25__SCAN_IN), .B1(n6502), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4843) );
  OAI21_X1 U6037 ( .B1(n6504), .B2(n4844), .A(n4843), .ZN(U2898) );
  INV_X1 U6038 ( .A(n6498), .ZN(n4845) );
  INV_X1 U6039 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6925) );
  INV_X1 U6040 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n7043) );
  OAI222_X1 U6041 ( .A1(n4845), .A2(n4047), .B1(n6504), .B2(n6925), .C1(n7043), 
        .C2(n6508), .ZN(U2897) );
  INV_X1 U6042 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n7074) );
  OAI222_X1 U6043 ( .A1(n4845), .A2(n3855), .B1(n6504), .B2(n7074), .C1(n4784), 
        .C2(n6508), .ZN(U2907) );
  AOI222_X1 U6044 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_21__SCAN_IN), .C1(n6502), .C2(UWORD_REG_5__SCAN_IN), .ZN(
        n4846) );
  INV_X1 U6045 ( .A(n4846), .ZN(U2902) );
  AOI222_X1 U6046 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_19__SCAN_IN), .C1(n6502), .C2(UWORD_REG_3__SCAN_IN), .ZN(
        n4847) );
  INV_X1 U6047 ( .A(n4847), .ZN(U2904) );
  AOI222_X1 U6048 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_24__SCAN_IN), .C1(n6502), .C2(UWORD_REG_8__SCAN_IN), .ZN(
        n4848) );
  INV_X1 U6049 ( .A(n4848), .ZN(U2899) );
  AOI222_X1 U6050 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_22__SCAN_IN), .C1(n6502), .C2(UWORD_REG_6__SCAN_IN), .ZN(
        n4849) );
  INV_X1 U6051 ( .A(n4849), .ZN(U2901) );
  AOI222_X1 U6052 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_18__SCAN_IN), .C1(n6502), .C2(UWORD_REG_2__SCAN_IN), .ZN(
        n4850) );
  INV_X1 U6053 ( .A(n4850), .ZN(U2905) );
  AOI222_X1 U6054 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n6502), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4851) );
  INV_X1 U6055 ( .A(n4851), .ZN(U2896) );
  AOI222_X1 U6056 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_20__SCAN_IN), .C1(n6502), .C2(UWORD_REG_4__SCAN_IN), .ZN(
        n4852) );
  INV_X1 U6057 ( .A(n4852), .ZN(U2903) );
  AOI222_X1 U6058 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_29__SCAN_IN), .C1(n6502), .C2(UWORD_REG_13__SCAN_IN), .ZN(
        n4853) );
  INV_X1 U6059 ( .A(n4853), .ZN(U2894) );
  AOI222_X1 U6060 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6498), .B1(n6506), .B2(
        DATAO_REG_17__SCAN_IN), .C1(n6502), .C2(UWORD_REG_1__SCAN_IN), .ZN(
        n4854) );
  INV_X1 U6061 ( .A(n4854), .ZN(U2906) );
  AND2_X1 U6062 ( .A1(n4855), .A2(n4856), .ZN(n4858) );
  AND2_X1 U6063 ( .A1(n4860), .A2(n4861), .ZN(n4862) );
  NOR2_X1 U6064 ( .A1(n4859), .A2(n4862), .ZN(n6581) );
  AOI22_X1 U6065 ( .A1(n6492), .A2(n6581), .B1(n5493), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4863) );
  OAI21_X1 U6066 ( .B1(n5395), .B2(n5490), .A(n4863), .ZN(U2855) );
  NAND2_X1 U6067 ( .A1(n4865), .A2(n4864), .ZN(n4874) );
  INV_X1 U6068 ( .A(n4874), .ZN(n4866) );
  AOI21_X1 U6069 ( .B1(n4868), .B2(n4867), .A(n4866), .ZN(n6537) );
  INV_X1 U6070 ( .A(n6537), .ZN(n5440) );
  INV_X1 U6071 ( .A(DATAI_2_), .ZN(n4869) );
  OAI222_X1 U6072 ( .A1(n5440), .A2(n5561), .B1(n5560), .B2(n4869), .C1(n5559), 
        .C2(n3668), .ZN(U2889) );
  OAI21_X1 U6073 ( .B1(n4871), .B2(n4872), .A(n4873), .ZN(n6588) );
  AOI21_X1 U6074 ( .B1(n4875), .B2(n4874), .A(n3177), .ZN(n4879) );
  AOI22_X1 U6075 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6586), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4876) );
  OAI21_X1 U6076 ( .B1(n5413), .B2(n6541), .A(n4876), .ZN(n4877) );
  AOI21_X1 U6077 ( .B1(n4879), .B2(n6536), .A(n4877), .ZN(n4878) );
  OAI21_X1 U6078 ( .B1(n5750), .B2(n6588), .A(n4878), .ZN(U2983) );
  INV_X1 U6079 ( .A(n4879), .ZN(n5426) );
  INV_X1 U6080 ( .A(n4860), .ZN(n4881) );
  AOI21_X1 U6081 ( .B1(n4882), .B2(n4880), .A(n4881), .ZN(n6587) );
  AOI22_X1 U6082 ( .A1(n6492), .A2(n6587), .B1(n5493), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4883) );
  OAI21_X1 U6083 ( .B1(n5426), .B2(n5495), .A(n4883), .ZN(U2856) );
  OAI222_X1 U6084 ( .A1(n5395), .A2(n5561), .B1(n5560), .B2(n4884), .C1(n5559), 
        .C2(n4778), .ZN(U2887) );
  OAI222_X1 U6085 ( .A1(n5426), .A2(n5561), .B1(n5560), .B2(n4885), .C1(n5559), 
        .C2(n4788), .ZN(U2888) );
  NOR2_X1 U6086 ( .A1(n4221), .A2(n6097), .ZN(n4886) );
  NAND2_X1 U6087 ( .A1(n4963), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4959) );
  NAND2_X1 U6088 ( .A1(n4959), .A2(n6693), .ZN(n6806) );
  NAND2_X1 U6089 ( .A1(n4887), .A2(n6635), .ZN(n4888) );
  OAI21_X1 U6090 ( .B1(n6806), .B2(n4888), .A(n6691), .ZN(n4893) );
  NOR2_X1 U6091 ( .A1(n4889), .A2(n6295), .ZN(n6066) );
  AOI21_X1 U6092 ( .B1(n6066), .B2(n6695), .A(n6623), .ZN(n4890) );
  NAND3_X1 U6093 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6982), .A3(n6421), .ZN(n6059) );
  OAI22_X1 U6094 ( .A1(n4893), .A2(n4890), .B1(n6059), .B2(n6956), .ZN(n6625)
         );
  INV_X1 U6095 ( .A(n6625), .ZN(n4905) );
  INV_X1 U6096 ( .A(n4890), .ZN(n4892) );
  INV_X1 U6097 ( .A(n6638), .ZN(n6697) );
  AOI21_X1 U6098 ( .B1(n6698), .B2(n6059), .A(n6697), .ZN(n4891) );
  NAND2_X1 U6099 ( .A1(n6536), .A2(DATAI_29_), .ZN(n6765) );
  INV_X1 U6100 ( .A(n5983), .ZN(n4895) );
  NAND2_X1 U6101 ( .A1(n4221), .A2(n6140), .ZN(n6292) );
  INV_X1 U6102 ( .A(n6292), .ZN(n4894) );
  NAND2_X1 U6103 ( .A1(n4221), .A2(n6214), .ZN(n6335) );
  INV_X1 U6104 ( .A(DATAI_21_), .ZN(n4896) );
  INV_X1 U6105 ( .A(n4897), .ZN(n6803) );
  OR2_X1 U6106 ( .A1(n4951), .A2(n4145), .ZN(n6734) );
  AOI22_X1 U6107 ( .A1(n6624), .A2(n6762), .B1(n6760), .B2(n6623), .ZN(n4899)
         );
  OAI21_X1 U6108 ( .B1(n6765), .B2(n6629), .A(n4899), .ZN(n4900) );
  AOI21_X1 U6109 ( .B1(n6626), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4900), 
        .ZN(n4901) );
  OAI21_X1 U6110 ( .B1(n4905), .B2(n6671), .A(n4901), .ZN(U3049) );
  NAND2_X1 U6111 ( .A1(n6536), .A2(DATAI_24_), .ZN(n6689) );
  INV_X1 U6112 ( .A(n6707), .ZN(n6641) );
  AOI22_X1 U6113 ( .A1(n6624), .A2(n6641), .B1(n6633), .B2(n6623), .ZN(n4902)
         );
  OAI21_X1 U6114 ( .B1(n6689), .B2(n6629), .A(n4902), .ZN(n4903) );
  AOI21_X1 U6115 ( .B1(n6626), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4903), 
        .ZN(n4904) );
  OAI21_X1 U6116 ( .B1(n4905), .B2(n6644), .A(n4904), .ZN(U3044) );
  OR2_X1 U6117 ( .A1(n4906), .A2(n3334), .ZN(n4907) );
  NAND2_X1 U6118 ( .A1(n4880), .A2(n4907), .ZN(n5431) );
  INV_X1 U6119 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4908) );
  OAI222_X1 U6120 ( .A1(n5431), .A2(n5497), .B1(n4908), .B2(n6495), .C1(n5490), 
        .C2(n5440), .ZN(U2857) );
  AND2_X1 U6121 ( .A1(n4221), .A2(n4909), .ZN(n4910) );
  NAND2_X1 U6122 ( .A1(n4915), .A2(n6140), .ZN(n6403) );
  INV_X1 U6123 ( .A(DATAI_31_), .ZN(n4911) );
  NOR2_X1 U6124 ( .A1(n6224), .A2(n6135), .ZN(n6254) );
  INV_X1 U6125 ( .A(n4952), .ZN(n4912) );
  AOI21_X1 U6126 ( .B1(n6254), .B2(n6373), .A(n4912), .ZN(n4916) );
  OAI21_X1 U6127 ( .B1(n4915), .B2(n5718), .A(n6338), .ZN(n4913) );
  AOI22_X1 U6128 ( .A1(n4916), .A2(n4913), .B1(n6366), .B2(n6698), .ZN(n4914)
         );
  NAND2_X1 U6129 ( .A1(n4948), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4922)
         );
  INV_X1 U6130 ( .A(n6752), .ZN(n6777) );
  INV_X1 U6131 ( .A(n4916), .ZN(n4918) );
  AOI22_X1 U6132 ( .A1(n4918), .A2(n6691), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4917), .ZN(n4953) );
  OAI22_X1 U6133 ( .A1(n4953), .A2(n6685), .B1(n4952), .B2(n6745), .ZN(n4920)
         );
  AOI21_X1 U6134 ( .B1(n6777), .B2(n6016), .A(n4920), .ZN(n4921) );
  OAI211_X1 U6135 ( .C1(n6403), .C2(n6782), .A(n4922), .B(n4921), .ZN(U3147)
         );
  NAND2_X1 U6136 ( .A1(n4948), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4925)
         );
  OAI22_X1 U6137 ( .A1(n4953), .A2(n6671), .B1(n4952), .B2(n6734), .ZN(n4923)
         );
  AOI21_X1 U6138 ( .B1(n6762), .B2(n6016), .A(n4923), .ZN(n4924) );
  OAI211_X1 U6139 ( .C1(n6403), .C2(n6765), .A(n4925), .B(n4924), .ZN(U3145)
         );
  INV_X1 U6140 ( .A(DATAI_30_), .ZN(n7076) );
  INV_X1 U6141 ( .A(n6673), .ZN(n6771) );
  NAND2_X1 U6142 ( .A1(n4948), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4929)
         );
  INV_X1 U6143 ( .A(DATAI_22_), .ZN(n4926) );
  OAI22_X1 U6144 ( .A1(n4953), .A2(n6676), .B1(n4952), .B2(n6739), .ZN(n4927)
         );
  AOI21_X1 U6145 ( .B1(n6768), .B2(n6016), .A(n4927), .ZN(n4928) );
  OAI211_X1 U6146 ( .C1(n6403), .C2(n6771), .A(n4929), .B(n4928), .ZN(U3146)
         );
  INV_X1 U6147 ( .A(DATAI_25_), .ZN(n4930) );
  INV_X1 U6148 ( .A(n6646), .ZN(n6714) );
  NAND2_X1 U6149 ( .A1(n4948), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4935)
         );
  INV_X1 U6150 ( .A(DATAI_17_), .ZN(n4931) );
  NOR2_X1 U6151 ( .A1(n5718), .A2(n4931), .ZN(n6612) );
  OAI22_X1 U6152 ( .A1(n4953), .A2(n6649), .B1(n4952), .B2(n6708), .ZN(n4933)
         );
  AOI21_X1 U6153 ( .B1(n6612), .B2(n6016), .A(n4933), .ZN(n4934) );
  OAI211_X1 U6154 ( .C1(n6403), .C2(n6714), .A(n4935), .B(n4934), .ZN(U3141)
         );
  NAND2_X1 U6155 ( .A1(n6536), .A2(DATAI_28_), .ZN(n6759) );
  NAND2_X1 U6156 ( .A1(n4948), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4939)
         );
  INV_X1 U6157 ( .A(n6733), .ZN(n6756) );
  OR2_X1 U6158 ( .A1(n4951), .A2(n4936), .ZN(n6729) );
  OAI22_X1 U6159 ( .A1(n4953), .A2(n6665), .B1(n4952), .B2(n6729), .ZN(n4937)
         );
  AOI21_X1 U6160 ( .B1(n6756), .B2(n6016), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6161 ( .C1(n6403), .C2(n6759), .A(n4939), .B(n4938), .ZN(U3144)
         );
  NAND2_X1 U6162 ( .A1(n6536), .A2(DATAI_27_), .ZN(n6728) );
  NAND2_X1 U6163 ( .A1(n4948), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4944)
         );
  NOR2_X1 U6164 ( .A1(n5718), .A2(n4940), .ZN(n6658) );
  OAI22_X1 U6165 ( .A1(n4953), .A2(n6661), .B1(n4952), .B2(n6722), .ZN(n4942)
         );
  AOI21_X1 U6166 ( .B1(n6658), .B2(n6016), .A(n4942), .ZN(n4943) );
  OAI211_X1 U6167 ( .C1(n6403), .C2(n6728), .A(n4944), .B(n4943), .ZN(U3143)
         );
  NAND2_X1 U6168 ( .A1(n4948), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4947)
         );
  OAI22_X1 U6169 ( .A1(n4953), .A2(n6644), .B1(n4952), .B2(n6688), .ZN(n4945)
         );
  AOI21_X1 U6170 ( .B1(n6641), .B2(n6016), .A(n4945), .ZN(n4946) );
  OAI211_X1 U6171 ( .C1(n6689), .C2(n6403), .A(n4947), .B(n4946), .ZN(U3140)
         );
  NAND2_X1 U6172 ( .A1(n4948), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4956)
         );
  INV_X1 U6173 ( .A(DATAI_18_), .ZN(n4949) );
  OAI22_X1 U6174 ( .A1(n4953), .A2(n6655), .B1(n4952), .B2(n6715), .ZN(n4954)
         );
  AOI21_X1 U6175 ( .B1(n6652), .B2(n6016), .A(n4954), .ZN(n4955) );
  OAI211_X1 U6176 ( .C1(n6403), .C2(n6721), .A(n4956), .B(n4955), .ZN(U3142)
         );
  NAND2_X1 U6177 ( .A1(n6417), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6099) );
  NOR2_X1 U6178 ( .A1(n6982), .A2(n6099), .ZN(n4958) );
  INV_X1 U6179 ( .A(n4958), .ZN(n6340) );
  AOI21_X1 U6180 ( .B1(n6254), .B2(n6348), .A(n4980), .ZN(n4962) );
  NAND3_X1 U6181 ( .A1(n6691), .A2(n4962), .A3(n4959), .ZN(n4957) );
  OAI211_X1 U6182 ( .C1(n6691), .C2(n4958), .A(n6638), .B(n4957), .ZN(n4979)
         );
  NAND2_X1 U6183 ( .A1(n6691), .A2(n4959), .ZN(n4961) );
  NAND2_X1 U6184 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4960) );
  OAI22_X1 U6185 ( .A1(n4962), .A2(n4961), .B1(n6099), .B2(n4960), .ZN(n4978)
         );
  AOI22_X1 U6186 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4979), .B1(n6774), 
        .B2(n4978), .ZN(n4965) );
  AOI22_X1 U6187 ( .A1(n6776), .A2(n6681), .B1(n6772), .B2(n4980), .ZN(n4964)
         );
  OAI211_X1 U6188 ( .C1(n6752), .C2(n6362), .A(n4965), .B(n4964), .ZN(U3131)
         );
  INV_X1 U6189 ( .A(n6652), .ZN(n6716) );
  INV_X1 U6190 ( .A(n6655), .ZN(n6718) );
  AOI22_X1 U6191 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4979), .B1(n6718), 
        .B2(n4978), .ZN(n4967) );
  AOI22_X1 U6192 ( .A1(n6776), .A2(n6651), .B1(n6650), .B2(n4980), .ZN(n4966)
         );
  OAI211_X1 U6193 ( .C1(n6716), .C2(n6362), .A(n4967), .B(n4966), .ZN(U3126)
         );
  INV_X1 U6194 ( .A(n6658), .ZN(n6723) );
  INV_X1 U6195 ( .A(n6661), .ZN(n6725) );
  AOI22_X1 U6196 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4979), .B1(n6725), 
        .B2(n4978), .ZN(n4969) );
  INV_X1 U6197 ( .A(n6728), .ZN(n6657) );
  AOI22_X1 U6198 ( .A1(n6776), .A2(n6657), .B1(n6656), .B2(n4980), .ZN(n4968)
         );
  OAI211_X1 U6199 ( .C1(n6723), .C2(n6362), .A(n4969), .B(n4968), .ZN(U3127)
         );
  AOI22_X1 U6200 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4979), .B1(n6767), 
        .B2(n4978), .ZN(n4971) );
  AOI22_X1 U6201 ( .A1(n6776), .A2(n6673), .B1(n6766), .B2(n4980), .ZN(n4970)
         );
  OAI211_X1 U6202 ( .C1(n6740), .C2(n6362), .A(n4971), .B(n4970), .ZN(U3130)
         );
  INV_X1 U6203 ( .A(n6671), .ZN(n6761) );
  AOI22_X1 U6204 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4979), .B1(n6761), 
        .B2(n4978), .ZN(n4973) );
  INV_X1 U6205 ( .A(n6765), .ZN(n6667) );
  AOI22_X1 U6206 ( .A1(n6776), .A2(n6667), .B1(n6760), .B2(n4980), .ZN(n4972)
         );
  OAI211_X1 U6207 ( .C1(n6735), .C2(n6362), .A(n4973), .B(n4972), .ZN(U3129)
         );
  AOI22_X1 U6208 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4979), .B1(n6755), 
        .B2(n4978), .ZN(n4975) );
  INV_X1 U6209 ( .A(n6759), .ZN(n6662) );
  AOI22_X1 U6210 ( .A1(n6776), .A2(n6662), .B1(n6754), .B2(n4980), .ZN(n4974)
         );
  OAI211_X1 U6211 ( .C1(n6733), .C2(n6362), .A(n4975), .B(n4974), .ZN(U3128)
         );
  INV_X1 U6212 ( .A(n6649), .ZN(n6711) );
  AOI22_X1 U6213 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4979), .B1(n6711), 
        .B2(n4978), .ZN(n4977) );
  AOI22_X1 U6214 ( .A1(n6776), .A2(n6646), .B1(n6611), .B2(n4980), .ZN(n4976)
         );
  OAI211_X1 U6215 ( .C1(n6709), .C2(n6362), .A(n4977), .B(n4976), .ZN(U3125)
         );
  INV_X1 U6216 ( .A(n6644), .ZN(n6704) );
  AOI22_X1 U6217 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4979), .B1(n6704), 
        .B2(n4978), .ZN(n4982) );
  INV_X1 U6218 ( .A(n6689), .ZN(n6634) );
  AOI22_X1 U6219 ( .A1(n6776), .A2(n6634), .B1(n6633), .B2(n4980), .ZN(n4981)
         );
  OAI211_X1 U6220 ( .C1(n6707), .C2(n6362), .A(n4982), .B(n4981), .ZN(U3124)
         );
  NAND2_X1 U6221 ( .A1(n4984), .A2(n4985), .ZN(n4988) );
  XNOR2_X1 U6222 ( .A(n4986), .B(n4989), .ZN(n4987) );
  NAND2_X1 U6223 ( .A1(n4988), .A2(n4987), .ZN(n6515) );
  OAI21_X1 U6224 ( .B1(n4988), .B2(n4987), .A(n6515), .ZN(n5749) );
  NAND2_X1 U6225 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U6226 ( .A1(n5833), .A2(n6599), .ZN(n6573) );
  NAND2_X1 U6227 ( .A1(n4990), .A2(n6573), .ZN(n6593) );
  OAI21_X1 U6228 ( .B1(n6579), .B2(n6593), .A(n4989), .ZN(n4999) );
  INV_X1 U6229 ( .A(n4990), .ZN(n5947) );
  NOR2_X1 U6230 ( .A1(n5947), .A2(n4991), .ZN(n6575) );
  AOI21_X1 U6231 ( .B1(n4994), .B2(n4993), .A(n4992), .ZN(n6598) );
  OAI21_X1 U6232 ( .B1(n5950), .B2(n6575), .A(n6598), .ZN(n6571) );
  NOR2_X1 U6233 ( .A1(n4859), .A2(n4996), .ZN(n4997) );
  OR2_X1 U6234 ( .A1(n4995), .A2(n4997), .ZN(n5498) );
  NAND2_X1 U6235 ( .A1(n6586), .A2(REIP_REG_5__SCAN_IN), .ZN(n5744) );
  OAI21_X1 U6236 ( .B1(n5951), .B2(n5498), .A(n5744), .ZN(n4998) );
  AOI21_X1 U6237 ( .B1(n4999), .B2(n6571), .A(n4998), .ZN(n5000) );
  OAI21_X1 U6238 ( .B1(n5957), .B2(n5749), .A(n5000), .ZN(U3013) );
  NAND2_X1 U6239 ( .A1(n4857), .A2(n5001), .ZN(n5380) );
  XNOR2_X1 U6240 ( .A(n5346), .B(n5380), .ZN(n6518) );
  INV_X1 U6241 ( .A(n6518), .ZN(n5377) );
  OAI222_X1 U6242 ( .A1(n5560), .A2(n5003), .B1(n5561), .B2(n5377), .C1(n5002), 
        .C2(n5559), .ZN(U2885) );
  OAI21_X1 U6243 ( .B1(n5004), .B2(n3336), .A(n5005), .ZN(n5717) );
  OR2_X1 U6244 ( .A1(n5007), .A2(n5008), .ZN(n5009) );
  AOI22_X1 U6245 ( .A1(n6543), .A2(n6492), .B1(n5493), .B2(EBX_REG_10__SCAN_IN), .ZN(n5010) );
  OAI21_X1 U6246 ( .B1(n5717), .B2(n5490), .A(n5010), .ZN(U2849) );
  INV_X1 U6247 ( .A(n5566), .ZN(n5013) );
  XNOR2_X1 U6248 ( .A(n5014), .B(n5751), .ZN(n5758) );
  NAND2_X1 U6249 ( .A1(n5725), .A2(n5015), .ZN(n5016) );
  NAND2_X1 U6250 ( .A1(n6586), .A2(REIP_REG_30__SCAN_IN), .ZN(n5752) );
  OAI211_X1 U6251 ( .C1(n5017), .C2(n5722), .A(n5016), .B(n5752), .ZN(n5018)
         );
  AOI21_X1 U6252 ( .B1(n5020), .B2(n6536), .A(n5018), .ZN(n5019) );
  OAI21_X1 U6253 ( .B1(n5758), .B2(n5750), .A(n5019), .ZN(U2956) );
  AOI22_X1 U6254 ( .A1(n5535), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5542), .ZN(n5023) );
  AND2_X1 U6255 ( .A1(n4145), .A2(n3636), .ZN(n5021) );
  NAND2_X1 U6256 ( .A1(n5536), .A2(DATAI_14_), .ZN(n5022) );
  OAI211_X1 U6257 ( .C1(n5024), .C2(n5561), .A(n5023), .B(n5022), .ZN(U2861)
         );
  INV_X1 U6258 ( .A(n5025), .ZN(n5962) );
  AOI21_X1 U6259 ( .B1(n6784), .B2(n5962), .A(n5037), .ZN(n5040) );
  NOR2_X1 U6260 ( .A1(n7079), .A2(n7015), .ZN(n5048) );
  OAI22_X1 U6261 ( .A1(n5027), .A2(n5026), .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5047) );
  INV_X1 U6262 ( .A(n5047), .ZN(n5036) );
  NOR3_X1 U6263 ( .A1(n5979), .A2(n3112), .A3(n5962), .ZN(n5035) );
  NAND2_X1 U6264 ( .A1(n5028), .A2(n5063), .ZN(n5966) );
  XNOR2_X1 U6265 ( .A(n5025), .B(n3112), .ZN(n5033) );
  XNOR2_X1 U6266 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3112), .ZN(n5029)
         );
  OAI22_X1 U6267 ( .A1(n6412), .A2(n5029), .B1(n5969), .B2(n5033), .ZN(n5032)
         );
  NOR2_X1 U6268 ( .A1(n5030), .A2(n5959), .ZN(n5031) );
  AOI211_X1 U6269 ( .C1(n5966), .C2(n5033), .A(n5032), .B(n5031), .ZN(n6407)
         );
  INV_X1 U6270 ( .A(n6442), .ZN(n5980) );
  NOR2_X1 U6271 ( .A1(n6407), .A2(n5980), .ZN(n5034) );
  AOI211_X1 U6272 ( .C1(n5048), .C2(n5036), .A(n5035), .B(n5034), .ZN(n5038)
         );
  OAI22_X1 U6273 ( .A1(n5040), .A2(n5039), .B1(n5038), .B2(n5037), .ZN(U3459)
         );
  OAI22_X1 U6274 ( .A1(n5041), .A2(n5497), .B1(n5042), .B2(n6495), .ZN(U2828)
         );
  NOR3_X1 U6275 ( .A1(n5043), .A2(n5025), .A3(n4683), .ZN(n5045) );
  AOI22_X1 U6276 ( .A1(n6784), .A2(n5046), .B1(n5048), .B2(n5047), .ZN(n5049)
         );
  OAI21_X1 U6277 ( .B1(n6414), .B2(n5980), .A(n5049), .ZN(n5051) );
  AOI22_X1 U6278 ( .A1(n5981), .A2(n5051), .B1(n5050), .B2(n6784), .ZN(n5052)
         );
  OAI21_X1 U6279 ( .B1(n5981), .B2(n5053), .A(n5052), .ZN(U3460) );
  AND2_X1 U6280 ( .A1(n6691), .A2(n7079), .ZN(n6447) );
  OR2_X1 U6281 ( .A1(n6447), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6282 ( .A1(n5054), .A2(n4334), .ZN(n5055) );
  MUX2_X1 U6283 ( .A(n5056), .B(n5055), .S(n5059), .Z(U3474) );
  AOI211_X1 U6284 ( .C1(n3487), .C2(n7046), .A(n6956), .B(n5057), .ZN(n5058)
         );
  OAI21_X1 U6285 ( .B1(n5058), .B2(n7091), .A(n6791), .ZN(n5062) );
  AOI211_X1 U6286 ( .C1(n6443), .C2(n6502), .A(n5060), .B(n5059), .ZN(n5061)
         );
  MUX2_X1 U6287 ( .A(n5062), .B(REQUESTPENDING_REG_SCAN_IN), .S(n5061), .Z(
        U3472) );
  NAND3_X1 U6288 ( .A1(n5064), .A2(n5063), .A3(n6424), .ZN(n5066) );
  MUX2_X1 U6289 ( .A(n5067), .B(n5066), .S(n5065), .Z(n5068) );
  AOI21_X1 U6290 ( .B1(n4309), .B2(n5069), .A(n5068), .ZN(n6425) );
  INV_X1 U6291 ( .A(n6425), .ZN(n5071) );
  MUX2_X1 U6292 ( .A(n5071), .B(MORE_REG_SCAN_IN), .S(n5070), .Z(U3471) );
  NAND2_X1 U6293 ( .A1(n5072), .A2(n4375), .ZN(n5075) );
  INV_X1 U6294 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6295 ( .A1(n5075), .A2(n5074), .ZN(n5076) );
  OR2_X1 U6296 ( .A1(n4553), .A2(n5076), .ZN(n5077) );
  NAND2_X1 U6297 ( .A1(n5078), .A2(n5077), .ZN(n5769) );
  OAI21_X1 U6298 ( .B1(n5079), .B2(n5081), .A(n5080), .ZN(n5571) );
  INV_X1 U6299 ( .A(n5571), .ZN(n5082) );
  NAND2_X1 U6300 ( .A1(n5082), .A2(n6488), .ZN(n5089) );
  INV_X1 U6301 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5083) );
  OAI22_X1 U6302 ( .A1(n5414), .A2(n5564), .B1(n5083), .B2(n6478), .ZN(n5087)
         );
  INV_X1 U6303 ( .A(n5084), .ZN(n5085) );
  MUX2_X1 U6304 ( .A(n5085), .B(n5093), .S(REIP_REG_29__SCAN_IN), .Z(n5086) );
  AOI211_X1 U6305 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6480), .A(n5087), .B(n5086), 
        .ZN(n5088) );
  OAI211_X1 U6306 ( .C1(n5415), .C2(n5769), .A(n5089), .B(n5088), .ZN(U2798)
         );
  INV_X1 U6307 ( .A(n5578), .ZN(n5505) );
  INV_X1 U6308 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5092) );
  OAI22_X1 U6309 ( .A1(n5414), .A2(n5576), .B1(n5092), .B2(n6478), .ZN(n5096)
         );
  AND2_X1 U6310 ( .A1(n3134), .A2(REIP_REG_27__SCAN_IN), .ZN(n5094) );
  MUX2_X1 U6311 ( .A(n5094), .B(n5093), .S(REIP_REG_28__SCAN_IN), .Z(n5095) );
  AOI211_X1 U6312 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6480), .A(n5096), .B(n5095), 
        .ZN(n5099) );
  AOI21_X1 U6313 ( .B1(n5097), .B2(n3124), .A(n4553), .ZN(n5775) );
  NAND2_X1 U6314 ( .A1(n5775), .A2(n6473), .ZN(n5098) );
  OAI211_X1 U6315 ( .C1(n5505), .C2(n5385), .A(n5099), .B(n5098), .ZN(U2799)
         );
  OR2_X1 U6316 ( .A1(n5100), .A2(n5101), .ZN(n5102) );
  AOI22_X1 U6317 ( .A1(n6487), .A2(n5586), .B1(n5454), .B2(
        PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6318 ( .A1(n6480), .A2(EBX_REG_27__SCAN_IN), .ZN(n5103) );
  OAI211_X1 U6319 ( .C1(n5118), .C2(n5109), .A(n5104), .B(n5103), .ZN(n5108)
         );
  NAND2_X1 U6320 ( .A1(n3144), .A2(n5105), .ZN(n5106) );
  NAND2_X1 U6321 ( .A1(n3124), .A2(n5106), .ZN(n5779) );
  NOR2_X1 U6322 ( .A1(n5779), .A2(n5415), .ZN(n5107) );
  AOI211_X1 U6323 ( .C1(n3134), .C2(n5109), .A(n5108), .B(n5107), .ZN(n5110)
         );
  OAI21_X1 U6324 ( .B1(n5583), .B2(n5385), .A(n5110), .ZN(U2800) );
  OR2_X1 U6325 ( .A1(n5111), .A2(n5112), .ZN(n5113) );
  NAND2_X1 U6326 ( .A1(n3144), .A2(n5113), .ZN(n5788) );
  AOI21_X1 U6327 ( .B1(n5116), .B2(n5124), .A(n5100), .ZN(n5595) );
  NAND2_X1 U6328 ( .A1(n5595), .A2(n6488), .ZN(n5123) );
  INV_X1 U6329 ( .A(n5591), .ZN(n5117) );
  OAI22_X1 U6330 ( .A1(n5414), .A2(n5117), .B1(n5593), .B2(n6478), .ZN(n5121)
         );
  AOI21_X1 U6331 ( .B1(n5119), .B2(n7105), .A(n5118), .ZN(n5120) );
  AOI211_X1 U6332 ( .C1(n6480), .C2(EBX_REG_26__SCAN_IN), .A(n5121), .B(n5120), 
        .ZN(n5122) );
  OAI211_X1 U6333 ( .C1(n5415), .C2(n5788), .A(n5123), .B(n5122), .ZN(U2801)
         );
  AOI21_X1 U6334 ( .B1(n5125), .B2(n4521), .A(n5115), .ZN(n5603) );
  INV_X1 U6335 ( .A(n5603), .ZN(n5513) );
  AOI21_X1 U6336 ( .B1(n5126), .B2(n5138), .A(n5111), .ZN(n5801) );
  XNOR2_X1 U6337 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5132) );
  OAI22_X1 U6338 ( .A1(n5414), .A2(n5601), .B1(n5127), .B2(n6478), .ZN(n5128)
         );
  AOI21_X1 U6339 ( .B1(n6480), .B2(EBX_REG_25__SCAN_IN), .A(n5128), .ZN(n5131)
         );
  AND2_X1 U6340 ( .A1(n5459), .A2(n5129), .ZN(n5150) );
  NAND2_X1 U6341 ( .A1(n5150), .A2(REIP_REG_25__SCAN_IN), .ZN(n5130) );
  OAI211_X1 U6342 ( .C1(n5144), .C2(n5132), .A(n5131), .B(n5130), .ZN(n5133)
         );
  AOI21_X1 U6343 ( .B1(n5801), .B2(n6473), .A(n5133), .ZN(n5134) );
  OAI21_X1 U6344 ( .B1(n5513), .B2(n5385), .A(n5134), .ZN(U2802) );
  NAND2_X1 U6345 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  NAND2_X1 U6346 ( .A1(n5138), .A2(n5137), .ZN(n5468) );
  INV_X1 U6347 ( .A(n5468), .ZN(n5809) );
  OAI22_X1 U6348 ( .A1(n5414), .A2(n5140), .B1(n5139), .B2(n6478), .ZN(n5141)
         );
  AOI21_X1 U6349 ( .B1(n6480), .B2(EBX_REG_24__SCAN_IN), .A(n5141), .ZN(n5143)
         );
  NAND2_X1 U6350 ( .A1(n5150), .A2(REIP_REG_24__SCAN_IN), .ZN(n5142) );
  OAI211_X1 U6351 ( .C1(n5144), .C2(REIP_REG_24__SCAN_IN), .A(n5143), .B(n5142), .ZN(n5145) );
  AOI21_X1 U6352 ( .B1(n5809), .B2(n6473), .A(n5145), .ZN(n5146) );
  OAI21_X1 U6353 ( .B1(n5516), .B2(n5385), .A(n5146), .ZN(U2803) );
  OAI22_X1 U6354 ( .A1(n5414), .A2(n5148), .B1(n5147), .B2(n6478), .ZN(n5149)
         );
  AOI21_X1 U6355 ( .B1(n6480), .B2(EBX_REG_23__SCAN_IN), .A(n5149), .ZN(n5153)
         );
  OAI21_X1 U6356 ( .B1(n5151), .B2(REIP_REG_23__SCAN_IN), .A(n5150), .ZN(n5152) );
  OAI211_X1 U6357 ( .C1(n5469), .C2(n5415), .A(n5153), .B(n5152), .ZN(n5154)
         );
  INV_X1 U6358 ( .A(n5154), .ZN(n5155) );
  OAI21_X1 U6359 ( .B1(n5519), .B2(n5385), .A(n5155), .ZN(U2804) );
  OR2_X1 U6360 ( .A1(n5182), .A2(n5172), .ZN(n5170) );
  AND2_X1 U6361 ( .A1(n5170), .A2(n5156), .ZN(n5158) );
  INV_X1 U6362 ( .A(n5159), .ZN(n5161) );
  AOI21_X1 U6363 ( .B1(n3161), .B2(n5161), .A(n5160), .ZN(n5818) );
  XNOR2_X1 U6364 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .ZN(
        n5162) );
  NOR2_X1 U6365 ( .A1(n5174), .A2(n5162), .ZN(n5168) );
  INV_X1 U6366 ( .A(n5459), .ZN(n5164) );
  OR2_X1 U6367 ( .A1(n5164), .A2(n5163), .ZN(n5192) );
  AOI22_X1 U6368 ( .A1(n6487), .A2(n5615), .B1(n5454), .B2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6369 ( .A1(n6480), .A2(EBX_REG_22__SCAN_IN), .ZN(n5165) );
  OAI211_X1 U6370 ( .C1(n5192), .C2(n4672), .A(n5166), .B(n5165), .ZN(n5167)
         );
  AOI211_X1 U6371 ( .C1(n5818), .C2(n6473), .A(n5168), .B(n5167), .ZN(n5169)
         );
  OAI21_X1 U6372 ( .B1(n5612), .B2(n5385), .A(n5169), .ZN(U2805) );
  INV_X1 U6373 ( .A(n5170), .ZN(n5171) );
  AOI21_X1 U6374 ( .B1(n5172), .B2(n5182), .A(n5171), .ZN(n5623) );
  INV_X1 U6375 ( .A(n5623), .ZN(n5524) );
  AOI21_X1 U6376 ( .B1(n3152), .B2(n5173), .A(n5159), .ZN(n5826) );
  NOR2_X1 U6377 ( .A1(n5174), .A2(REIP_REG_21__SCAN_IN), .ZN(n5179) );
  AOI22_X1 U6378 ( .A1(n6487), .A2(n5619), .B1(n5454), .B2(
        PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6379 ( .A1(n6480), .A2(EBX_REG_21__SCAN_IN), .ZN(n5175) );
  OAI211_X1 U6380 ( .C1(n5192), .C2(n5177), .A(n5176), .B(n5175), .ZN(n5178)
         );
  AOI211_X1 U6381 ( .C1(n5826), .C2(n6473), .A(n5179), .B(n5178), .ZN(n5180)
         );
  OAI21_X1 U6382 ( .B1(n5524), .B2(n5385), .A(n5180), .ZN(U2806) );
  OAI21_X1 U6383 ( .B1(n5181), .B2(n5183), .A(n5182), .ZN(n5628) );
  MUX2_X1 U6384 ( .A(n5185), .B(n5184), .S(n5199), .Z(n5187) );
  XNOR2_X1 U6385 ( .A(n5187), .B(n5186), .ZN(n5841) );
  INV_X1 U6386 ( .A(n5222), .ZN(n5189) );
  AOI21_X1 U6387 ( .B1(n5189), .B2(n5188), .A(REIP_REG_20__SCAN_IN), .ZN(n5193) );
  AOI22_X1 U6388 ( .A1(n6487), .A2(n5631), .B1(n5454), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6389 ( .A1(n6480), .A2(EBX_REG_20__SCAN_IN), .ZN(n5190) );
  OAI211_X1 U6390 ( .C1(n5193), .C2(n5192), .A(n5191), .B(n5190), .ZN(n5194)
         );
  AOI21_X1 U6391 ( .B1(n5841), .B2(n6473), .A(n5194), .ZN(n5195) );
  OAI21_X1 U6392 ( .B1(n5628), .B2(n5385), .A(n5195), .ZN(U2807) );
  NOR2_X1 U6393 ( .A1(n5196), .A2(n5197), .ZN(n5198) );
  NAND2_X1 U6394 ( .A1(n5201), .A2(n5200), .ZN(n5217) );
  AOI21_X1 U6395 ( .B1(n5202), .B2(n5217), .A(n5203), .ZN(n5204) );
  AOI21_X1 U6396 ( .B1(n3301), .B2(n5217), .A(n5204), .ZN(n5850) );
  XNOR2_X1 U6397 ( .A(REIP_REG_19__SCAN_IN), .B(REIP_REG_18__SCAN_IN), .ZN(
        n5211) );
  NAND2_X1 U6398 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5205)
         );
  NAND2_X1 U6399 ( .A1(n5420), .A2(n6447), .ZN(n6477) );
  OAI211_X1 U6400 ( .C1(n5414), .C2(n5637), .A(n5205), .B(n6477), .ZN(n5206)
         );
  AOI21_X1 U6401 ( .B1(n6480), .B2(EBX_REG_19__SCAN_IN), .A(n5206), .ZN(n5210)
         );
  INV_X1 U6402 ( .A(n5207), .ZN(n5208) );
  AND2_X1 U6403 ( .A1(n5208), .A2(n5459), .ZN(n5235) );
  NAND2_X1 U6404 ( .A1(n5235), .A2(REIP_REG_19__SCAN_IN), .ZN(n5209) );
  OAI211_X1 U6405 ( .C1(n5211), .C2(n5222), .A(n5210), .B(n5209), .ZN(n5212)
         );
  AOI21_X1 U6406 ( .B1(n5850), .B2(n6473), .A(n5212), .ZN(n5213) );
  OAI21_X1 U6407 ( .B1(n5635), .B2(n5385), .A(n5213), .ZN(U2808) );
  AOI21_X1 U6408 ( .B1(n5216), .B2(n5215), .A(n5196), .ZN(n5651) );
  INV_X1 U6409 ( .A(n5651), .ZN(n5531) );
  XOR2_X1 U6410 ( .A(n5217), .B(n5202), .Z(n5859) );
  NAND2_X1 U6411 ( .A1(n6487), .A2(n5648), .ZN(n5218) );
  OAI211_X1 U6412 ( .C1(n6478), .C2(n3274), .A(n5218), .B(n6477), .ZN(n5219)
         );
  AOI21_X1 U6413 ( .B1(EBX_REG_18__SCAN_IN), .B2(n6480), .A(n5219), .ZN(n5221)
         );
  NAND2_X1 U6414 ( .A1(n5235), .A2(REIP_REG_18__SCAN_IN), .ZN(n5220) );
  OAI211_X1 U6415 ( .C1(n5222), .C2(REIP_REG_18__SCAN_IN), .A(n5221), .B(n5220), .ZN(n5223) );
  AOI21_X1 U6416 ( .B1(n5859), .B2(n6473), .A(n5223), .ZN(n5224) );
  OAI21_X1 U6417 ( .B1(n5531), .B2(n5385), .A(n5224), .ZN(U2809) );
  NOR2_X1 U6418 ( .A1(n5241), .A2(n5225), .ZN(n5226) );
  INV_X1 U6419 ( .A(n5215), .ZN(n5228) );
  AOI21_X1 U6420 ( .B1(n5229), .B2(n5227), .A(n5228), .ZN(n5659) );
  NAND2_X1 U6421 ( .A1(n5659), .A2(n6488), .ZN(n5238) );
  NAND2_X1 U6422 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5245) );
  OAI21_X1 U6423 ( .B1(n5259), .B2(n5245), .A(n5230), .ZN(n5236) );
  NAND2_X1 U6424 ( .A1(n6480), .A2(EBX_REG_17__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6425 ( .A1(n6487), .A2(n5655), .ZN(n5232) );
  NAND2_X1 U6426 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5231)
         );
  NAND4_X1 U6427 ( .A1(n5233), .A2(n6477), .A3(n5232), .A4(n5231), .ZN(n5234)
         );
  AOI21_X1 U6428 ( .B1(n5236), .B2(n5235), .A(n5234), .ZN(n5237) );
  OAI211_X1 U6429 ( .C1(n5864), .C2(n5415), .A(n5238), .B(n5237), .ZN(U2810)
         );
  OAI21_X1 U6430 ( .B1(n5239), .B2(n5240), .A(n5227), .ZN(n5667) );
  AOI21_X1 U6431 ( .B1(n5242), .B2(n5255), .A(n5241), .ZN(n5884) );
  NAND2_X1 U6432 ( .A1(n5459), .A2(n5243), .ZN(n5271) );
  NAND2_X1 U6433 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5244)
         );
  OAI211_X1 U6434 ( .C1(n5414), .C2(n5663), .A(n6477), .B(n5244), .ZN(n5248)
         );
  OAI21_X1 U6435 ( .B1(REIP_REG_15__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .A(
        n5245), .ZN(n5246) );
  NOR2_X1 U6436 ( .A1(n5259), .A2(n5246), .ZN(n5247) );
  AOI211_X1 U6437 ( .C1(n6480), .C2(EBX_REG_16__SCAN_IN), .A(n5248), .B(n5247), 
        .ZN(n5249) );
  OAI21_X1 U6438 ( .B1(n5662), .B2(n5271), .A(n5249), .ZN(n5250) );
  AOI21_X1 U6439 ( .B1(n5884), .B2(n6473), .A(n5250), .ZN(n5251) );
  OAI21_X1 U6440 ( .B1(n5667), .B2(n5385), .A(n5251), .ZN(U2811) );
  AOI21_X1 U6441 ( .B1(n5253), .B2(n5252), .A(n5239), .ZN(n5673) );
  INV_X1 U6442 ( .A(n5673), .ZN(n5541) );
  INV_X1 U6443 ( .A(n5255), .ZN(n5256) );
  AOI21_X1 U6444 ( .B1(n5257), .B2(n5254), .A(n5256), .ZN(n5890) );
  NAND2_X1 U6445 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5258)
         );
  OAI211_X1 U6446 ( .C1(n5414), .C2(n5671), .A(n6477), .B(n5258), .ZN(n5261)
         );
  NOR2_X1 U6447 ( .A1(n5259), .A2(REIP_REG_15__SCAN_IN), .ZN(n5260) );
  AOI211_X1 U6448 ( .C1(EBX_REG_15__SCAN_IN), .C2(n6480), .A(n5261), .B(n5260), 
        .ZN(n5262) );
  OAI21_X1 U6449 ( .B1(n6971), .B2(n5271), .A(n5262), .ZN(n5263) );
  AOI21_X1 U6450 ( .B1(n5890), .B2(n6473), .A(n5263), .ZN(n5264) );
  OAI21_X1 U6451 ( .B1(n5541), .B2(n5385), .A(n5264), .ZN(U2812) );
  INV_X1 U6452 ( .A(n5252), .ZN(n5266) );
  AOI21_X1 U6453 ( .B1(n5267), .B2(n5265), .A(n5266), .ZN(n5681) );
  INV_X1 U6454 ( .A(n5681), .ZN(n5545) );
  INV_X1 U6455 ( .A(n5254), .ZN(n5269) );
  AOI21_X1 U6456 ( .B1(n5270), .B2(n5268), .A(n5269), .ZN(n5909) );
  AOI21_X1 U6457 ( .B1(n3135), .B2(REIP_REG_13__SCAN_IN), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5272) );
  NOR2_X1 U6458 ( .A1(n5272), .A2(n5271), .ZN(n5278) );
  INV_X1 U6459 ( .A(n6480), .ZN(n5457) );
  INV_X1 U6460 ( .A(n5679), .ZN(n5273) );
  INV_X1 U6461 ( .A(n6477), .ZN(n5403) );
  AOI21_X1 U6462 ( .B1(n6487), .B2(n5273), .A(n5403), .ZN(n5275) );
  NAND2_X1 U6463 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5274)
         );
  OAI211_X1 U6464 ( .C1(n5457), .C2(n5276), .A(n5275), .B(n5274), .ZN(n5277)
         );
  AOI211_X1 U6465 ( .C1(n5909), .C2(n6473), .A(n5278), .B(n5277), .ZN(n5279)
         );
  OAI21_X1 U6466 ( .B1(n5545), .B2(n5385), .A(n5279), .ZN(U2813) );
  AOI21_X1 U6467 ( .B1(n5282), .B2(n5281), .A(n3285), .ZN(n5688) );
  INV_X1 U6468 ( .A(n5688), .ZN(n5548) );
  INV_X1 U6469 ( .A(n5420), .ZN(n5442) );
  INV_X1 U6470 ( .A(n5296), .ZN(n5283) );
  OAI21_X1 U6471 ( .B1(n5442), .B2(n5283), .A(n5459), .ZN(n5314) );
  OAI21_X1 U6472 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5429), .A(n5314), .ZN(n5290) );
  INV_X1 U6473 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6474 ( .A1(n3135), .A2(n6965), .ZN(n5284) );
  OAI211_X1 U6475 ( .C1(n5457), .C2(n5286), .A(n5285), .B(n5284), .ZN(n5289)
         );
  OAI21_X1 U6476 ( .B1(n5294), .B2(n5287), .A(n5268), .ZN(n5912) );
  NOR2_X1 U6477 ( .A1(n5912), .A2(n5415), .ZN(n5288) );
  AOI211_X1 U6478 ( .C1(REIP_REG_13__SCAN_IN), .C2(n5290), .A(n5289), .B(n5288), .ZN(n5291) );
  OAI21_X1 U6479 ( .B1(n5548), .B2(n5385), .A(n5291), .ZN(U2814) );
  OAI21_X1 U6480 ( .B1(n5292), .B2(n5293), .A(n5281), .ZN(n5694) );
  AOI21_X1 U6481 ( .B1(n5295), .B2(n5309), .A(n5294), .ZN(n5933) );
  OAI21_X1 U6482 ( .B1(n6478), .B2(n3277), .A(n6477), .ZN(n5300) );
  NAND3_X1 U6483 ( .A1(n5441), .A2(n5296), .A3(n5302), .ZN(n5297) );
  OAI21_X1 U6484 ( .B1(n5457), .B2(n5298), .A(n5297), .ZN(n5299) );
  AOI211_X1 U6485 ( .C1(n5697), .C2(n6487), .A(n5300), .B(n5299), .ZN(n5301)
         );
  OAI21_X1 U6486 ( .B1(n5302), .B2(n5314), .A(n5301), .ZN(n5303) );
  AOI21_X1 U6487 ( .B1(n6473), .B2(n5933), .A(n5303), .ZN(n5304) );
  OAI21_X1 U6488 ( .B1(n5694), .B2(n5385), .A(n5304), .ZN(U2815) );
  AND2_X1 U6489 ( .A1(n5005), .A2(n5305), .ZN(n5306) );
  NAND2_X1 U6490 ( .A1(n5006), .A2(n5307), .ZN(n5308) );
  NAND2_X1 U6491 ( .A1(n5309), .A2(n5308), .ZN(n5936) );
  INV_X1 U6492 ( .A(n5936), .ZN(n5318) );
  INV_X1 U6493 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5481) );
  INV_X1 U6494 ( .A(n5705), .ZN(n5310) );
  AOI21_X1 U6495 ( .B1(n6487), .B2(n5310), .A(n5403), .ZN(n5312) );
  NAND2_X1 U6496 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5311)
         );
  OAI211_X1 U6497 ( .C1(n5457), .C2(n5481), .A(n5312), .B(n5311), .ZN(n5317)
         );
  AOI21_X1 U6498 ( .B1(n5441), .B2(n5313), .A(REIP_REG_11__SCAN_IN), .ZN(n5315) );
  NOR2_X1 U6499 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  AOI211_X1 U6500 ( .C1(n5318), .C2(n6473), .A(n5317), .B(n5316), .ZN(n5319)
         );
  OAI21_X1 U6501 ( .B1(n5708), .B2(n5385), .A(n5319), .ZN(U2816) );
  INV_X1 U6502 ( .A(n5340), .ZN(n5320) );
  OAI21_X1 U6503 ( .B1(n5429), .B2(n5320), .A(n5420), .ZN(n6475) );
  NAND2_X1 U6504 ( .A1(n4667), .A2(n5320), .ZN(n5321) );
  NOR2_X1 U6505 ( .A1(n5429), .A2(n5321), .ZN(n6476) );
  OAI21_X1 U6506 ( .B1(n6475), .B2(n6476), .A(REIP_REG_10__SCAN_IN), .ZN(n5330) );
  INV_X1 U6507 ( .A(n5713), .ZN(n5324) );
  INV_X1 U6508 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5322) );
  OAI21_X1 U6509 ( .B1(n6478), .B2(n5322), .A(n6477), .ZN(n5323) );
  AOI21_X1 U6510 ( .B1(n5324), .B2(n6487), .A(n5323), .ZN(n5329) );
  NAND2_X1 U6511 ( .A1(n6480), .A2(EBX_REG_10__SCAN_IN), .ZN(n5328) );
  NAND3_X1 U6512 ( .A1(n5441), .A2(n5326), .A3(n5325), .ZN(n5327) );
  NAND4_X1 U6513 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n5332)
         );
  NOR2_X1 U6514 ( .A1(n5717), .A2(n5385), .ZN(n5331) );
  AOI211_X1 U6515 ( .C1(n6543), .C2(n6473), .A(n5332), .B(n5331), .ZN(n5333)
         );
  INV_X1 U6516 ( .A(n5333), .ZN(U2817) );
  INV_X1 U6517 ( .A(n5731), .ZN(n5335) );
  OAI21_X1 U6518 ( .B1(n6478), .B2(n3731), .A(n6477), .ZN(n5334) );
  AOI21_X1 U6519 ( .B1(n5335), .B2(n6487), .A(n5334), .ZN(n5344) );
  AND2_X1 U6520 ( .A1(n5336), .A2(n5337), .ZN(n5338) );
  OR2_X1 U6521 ( .A1(n5338), .A2(n3159), .ZN(n5492) );
  INV_X1 U6522 ( .A(n5492), .ZN(n6552) );
  NAND2_X1 U6523 ( .A1(n6473), .A2(n6552), .ZN(n5343) );
  NAND2_X1 U6524 ( .A1(n6480), .A2(EBX_REG_8__SCAN_IN), .ZN(n5342) );
  NAND3_X1 U6525 ( .A1(n5441), .A2(n5340), .A3(n5339), .ZN(n5341) );
  NAND4_X1 U6526 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n5352)
         );
  INV_X1 U6527 ( .A(n5345), .ZN(n5350) );
  INV_X1 U6528 ( .A(n5346), .ZN(n5347) );
  NOR2_X1 U6529 ( .A1(n5380), .A2(n5347), .ZN(n5354) );
  NAND2_X1 U6530 ( .A1(n5354), .A2(n5348), .ZN(n5349) );
  NOR2_X1 U6531 ( .A1(n5349), .A2(n5350), .ZN(n5484) );
  AOI21_X1 U6532 ( .B1(n5350), .B2(n5349), .A(n5484), .ZN(n5733) );
  INV_X1 U6533 ( .A(n5733), .ZN(n5556) );
  NOR2_X1 U6534 ( .A1(n5556), .A2(n5385), .ZN(n5351) );
  AOI211_X1 U6535 ( .C1(REIP_REG_8__SCAN_IN), .C2(n6475), .A(n5352), .B(n5351), 
        .ZN(n5353) );
  INV_X1 U6536 ( .A(n5353), .ZN(U2819) );
  XOR2_X1 U6537 ( .A(n5348), .B(n5354), .Z(n5741) );
  INV_X1 U6538 ( .A(n5741), .ZN(n5558) );
  NOR4_X1 U6539 ( .A1(n5429), .A2(n5362), .A3(REIP_REG_7__SCAN_IN), .A4(n6978), 
        .ZN(n5361) );
  AOI21_X1 U6540 ( .B1(n5454), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5403), 
        .ZN(n5359) );
  INV_X1 U6541 ( .A(n5336), .ZN(n5356) );
  AOI21_X1 U6542 ( .B1(n5357), .B2(n5355), .A(n5356), .ZN(n6562) );
  NAND2_X1 U6543 ( .A1(n6473), .A2(n6562), .ZN(n5358) );
  OAI211_X1 U6544 ( .C1(n5414), .C2(n5739), .A(n5359), .B(n5358), .ZN(n5360)
         );
  AOI211_X1 U6545 ( .C1(n6480), .C2(EBX_REG_7__SCAN_IN), .A(n5361), .B(n5360), 
        .ZN(n5367) );
  INV_X1 U6546 ( .A(n5362), .ZN(n5364) );
  NAND2_X1 U6547 ( .A1(n5420), .A2(n5364), .ZN(n5363) );
  NAND2_X1 U6548 ( .A1(n6978), .A2(n5364), .ZN(n5365) );
  NOR2_X1 U6549 ( .A1(n5429), .A2(n5365), .ZN(n5369) );
  OAI21_X1 U6550 ( .B1(n5379), .B2(n5369), .A(REIP_REG_7__SCAN_IN), .ZN(n5366)
         );
  OAI211_X1 U6551 ( .C1(n5558), .C2(n5385), .A(n5367), .B(n5366), .ZN(U2820)
         );
  OR2_X1 U6552 ( .A1(n4995), .A2(n3333), .ZN(n5368) );
  AND2_X1 U6553 ( .A1(n5355), .A2(n5368), .ZN(n6570) );
  AOI22_X1 U6554 ( .A1(n6473), .A2(n6570), .B1(n6480), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n5374) );
  INV_X1 U6555 ( .A(n5369), .ZN(n5373) );
  INV_X1 U6556 ( .A(n6521), .ZN(n5370) );
  AOI21_X1 U6557 ( .B1(n6487), .B2(n5370), .A(n5403), .ZN(n5372) );
  NAND2_X1 U6558 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5371)
         );
  NAND4_X1 U6559 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n5375)
         );
  AOI21_X1 U6560 ( .B1(n5379), .B2(REIP_REG_6__SCAN_IN), .A(n5375), .ZN(n5376)
         );
  OAI21_X1 U6561 ( .B1(n5377), .B2(n5385), .A(n5376), .ZN(U2821) );
  AOI21_X1 U6562 ( .B1(n5441), .B2(n5378), .A(REIP_REG_5__SCAN_IN), .ZN(n5394)
         );
  INV_X1 U6563 ( .A(n5379), .ZN(n5393) );
  INV_X1 U6564 ( .A(n5001), .ZN(n5383) );
  INV_X1 U6565 ( .A(n4857), .ZN(n5382) );
  INV_X1 U6566 ( .A(n5380), .ZN(n5381) );
  AOI21_X1 U6567 ( .B1(n5383), .B2(n5382), .A(n5381), .ZN(n5747) );
  NAND2_X1 U6568 ( .A1(n5400), .A2(n3181), .ZN(n5384) );
  NAND2_X1 U6569 ( .A1(n5385), .A2(n5384), .ZN(n5449) );
  NAND2_X1 U6570 ( .A1(n5747), .A2(n5449), .ZN(n5392) );
  NAND2_X1 U6571 ( .A1(n6480), .A2(EBX_REG_5__SCAN_IN), .ZN(n5386) );
  OAI21_X1 U6572 ( .B1(n5498), .B2(n5415), .A(n5386), .ZN(n5390) );
  INV_X1 U6573 ( .A(n5745), .ZN(n5387) );
  NAND2_X1 U6574 ( .A1(n6487), .A2(n5387), .ZN(n5388) );
  OAI211_X1 U6575 ( .C1(n6478), .C2(n7111), .A(n5388), .B(n6477), .ZN(n5389)
         );
  NOR2_X1 U6576 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  OAI211_X1 U6577 ( .C1(n5394), .C2(n5393), .A(n5392), .B(n5391), .ZN(U2822)
         );
  INV_X1 U6578 ( .A(n5395), .ZN(n6526) );
  INV_X1 U6579 ( .A(n5401), .ZN(n5396) );
  NAND2_X1 U6580 ( .A1(n5420), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U6581 ( .A1(n5459), .A2(n5397), .ZN(n5422) );
  NOR2_X1 U6582 ( .A1(n5422), .A2(n4670), .ZN(n5410) );
  INV_X1 U6583 ( .A(n5398), .ZN(n5399) );
  AND2_X1 U6584 ( .A1(n5400), .A2(n5399), .ZN(n5452) );
  AOI22_X1 U6585 ( .A1(n6473), .A2(n6581), .B1(n5452), .B2(n6423), .ZN(n5408)
         );
  NOR2_X1 U6586 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5401), .ZN(n5402) );
  AOI22_X1 U6587 ( .A1(n5441), .A2(n5402), .B1(n6480), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5407) );
  INV_X1 U6588 ( .A(n6529), .ZN(n5404) );
  AOI21_X1 U6589 ( .B1(n6487), .B2(n5404), .A(n5403), .ZN(n5406) );
  OR2_X1 U6590 ( .A1(n6478), .A2(n3685), .ZN(n5405) );
  NAND4_X1 U6591 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n5409)
         );
  AOI211_X1 U6592 ( .C1(n6526), .C2(n5449), .A(n5410), .B(n5409), .ZN(n5411)
         );
  INV_X1 U6593 ( .A(n5411), .ZN(U2823) );
  OAI22_X1 U6594 ( .A1(n5414), .A2(n5413), .B1(n5412), .B2(n6478), .ZN(n5419)
         );
  INV_X1 U6595 ( .A(n5452), .ZN(n5417) );
  INV_X1 U6596 ( .A(n6587), .ZN(n5416) );
  OAI22_X1 U6597 ( .A1(n5417), .A2(n6224), .B1(n5416), .B2(n5415), .ZN(n5418)
         );
  AOI211_X1 U6598 ( .C1(n6480), .C2(EBX_REG_3__SCAN_IN), .A(n5419), .B(n5418), 
        .ZN(n5425) );
  NAND2_X1 U6599 ( .A1(n5420), .A2(REIP_REG_1__SCAN_IN), .ZN(n5421) );
  AOI21_X1 U6600 ( .B1(n5459), .B2(n5421), .A(n5428), .ZN(n5427) );
  INV_X1 U6601 ( .A(n5422), .ZN(n5423) );
  OAI21_X1 U6602 ( .B1(n5427), .B2(REIP_REG_3__SCAN_IN), .A(n5423), .ZN(n5424)
         );
  OAI211_X1 U6603 ( .C1(n5426), .C2(n5462), .A(n5425), .B(n5424), .ZN(U2824)
         );
  INV_X1 U6604 ( .A(n5427), .ZN(n5438) );
  OAI21_X1 U6605 ( .B1(n5429), .B2(n6888), .A(n5428), .ZN(n5437) );
  INV_X1 U6606 ( .A(n6540), .ZN(n5430) );
  AOI22_X1 U6607 ( .A1(n6487), .A2(n5430), .B1(n5454), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6608 ( .A1(n6480), .A2(EBX_REG_2__SCAN_IN), .ZN(n5434) );
  INV_X1 U6609 ( .A(n5431), .ZN(n6596) );
  NAND2_X1 U6610 ( .A1(n6473), .A2(n6596), .ZN(n5433) );
  NAND2_X1 U6611 ( .A1(n5452), .A2(n4837), .ZN(n5432) );
  NAND4_X1 U6612 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n5436)
         );
  AOI21_X1 U6613 ( .B1(n5438), .B2(n5437), .A(n5436), .ZN(n5439) );
  OAI21_X1 U6614 ( .B1(n5440), .B2(n5462), .A(n5439), .ZN(U2825) );
  AOI22_X1 U6615 ( .A1(n6473), .A2(n4808), .B1(n5452), .B2(n3116), .ZN(n5447)
         );
  AOI22_X1 U6616 ( .A1(n5441), .A2(n6888), .B1(n6480), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5446) );
  AOI22_X1 U6617 ( .A1(n6487), .A2(n5443), .B1(REIP_REG_1__SCAN_IN), .B2(n5442), .ZN(n5445) );
  NAND2_X1 U6618 ( .A1(n5454), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5444)
         );
  NAND4_X1 U6619 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n5448)
         );
  AOI21_X1 U6620 ( .B1(n5450), .B2(n5449), .A(n5448), .ZN(n5451) );
  INV_X1 U6621 ( .A(n5451), .ZN(U2826) );
  AOI22_X1 U6622 ( .A1(n6473), .A2(n5453), .B1(n5452), .B2(n6695), .ZN(n5456)
         );
  OAI21_X1 U6623 ( .B1(n6487), .B2(n5454), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5455) );
  OAI211_X1 U6624 ( .C1(n4344), .C2(n5457), .A(n5456), .B(n5455), .ZN(n5458)
         );
  AOI21_X1 U6625 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5459), .A(n5458), .ZN(n5460)
         );
  OAI21_X1 U6626 ( .B1(n5462), .B2(n5461), .A(n5460), .ZN(U2827) );
  OAI222_X1 U6627 ( .A1(n5463), .A2(n6495), .B1(n5497), .B2(n5769), .C1(n5571), 
        .C2(n5490), .ZN(U2830) );
  AOI22_X1 U6628 ( .A1(n5775), .A2(n6492), .B1(n5493), .B2(EBX_REG_28__SCAN_IN), .ZN(n5464) );
  OAI21_X1 U6629 ( .B1(n5505), .B2(n5495), .A(n5464), .ZN(U2831) );
  INV_X1 U6630 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5465) );
  OAI222_X1 U6631 ( .A1(n5465), .A2(n6495), .B1(n5497), .B2(n5779), .C1(n5583), 
        .C2(n5495), .ZN(U2832) );
  INV_X1 U6632 ( .A(n5595), .ZN(n5510) );
  OAI222_X1 U6633 ( .A1(n5466), .A2(n6495), .B1(n5497), .B2(n5788), .C1(n5510), 
        .C2(n5495), .ZN(U2833) );
  AOI22_X1 U6634 ( .A1(n5801), .A2(n6492), .B1(n5493), .B2(EBX_REG_25__SCAN_IN), .ZN(n5467) );
  OAI21_X1 U6635 ( .B1(n5513), .B2(n5495), .A(n5467), .ZN(U2834) );
  INV_X1 U6636 ( .A(EBX_REG_24__SCAN_IN), .ZN(n7064) );
  OAI222_X1 U6637 ( .A1(n7064), .A2(n6495), .B1(n5497), .B2(n5468), .C1(n5516), 
        .C2(n5490), .ZN(U2835) );
  OAI222_X1 U6638 ( .A1(n5470), .A2(n6495), .B1(n5497), .B2(n5469), .C1(n5519), 
        .C2(n5490), .ZN(U2836) );
  INV_X1 U6639 ( .A(EBX_REG_22__SCAN_IN), .ZN(n7031) );
  INV_X1 U6640 ( .A(n5818), .ZN(n5471) );
  OAI222_X1 U6641 ( .A1(n7031), .A2(n6495), .B1(n5497), .B2(n5471), .C1(n5612), 
        .C2(n5490), .ZN(U2837) );
  INV_X1 U6642 ( .A(n5826), .ZN(n5472) );
  INV_X1 U6643 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6893) );
  OAI222_X1 U6644 ( .A1(n5472), .A2(n5497), .B1(n6893), .B2(n6495), .C1(n5524), 
        .C2(n5490), .ZN(U2838) );
  AOI22_X1 U6645 ( .A1(n5841), .A2(n6492), .B1(n5493), .B2(EBX_REG_20__SCAN_IN), .ZN(n5473) );
  OAI21_X1 U6646 ( .B1(n5628), .B2(n5495), .A(n5473), .ZN(U2839) );
  AOI22_X1 U6647 ( .A1(n5850), .A2(n6492), .B1(n5493), .B2(EBX_REG_19__SCAN_IN), .ZN(n5474) );
  OAI21_X1 U6648 ( .B1(n5635), .B2(n5495), .A(n5474), .ZN(U2840) );
  INV_X1 U6649 ( .A(n5859), .ZN(n5475) );
  INV_X1 U6650 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7127) );
  OAI222_X1 U6651 ( .A1(n5531), .A2(n5495), .B1(n5497), .B2(n5475), .C1(n7127), 
        .C2(n6495), .ZN(U2841) );
  INV_X1 U6652 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5476) );
  INV_X1 U6653 ( .A(n5659), .ZN(n5534) );
  OAI222_X1 U6654 ( .A1(n5864), .A2(n5497), .B1(n5476), .B2(n6495), .C1(n5534), 
        .C2(n5490), .ZN(U2842) );
  AOI22_X1 U6655 ( .A1(n5884), .A2(n6492), .B1(n5493), .B2(EBX_REG_16__SCAN_IN), .ZN(n5477) );
  OAI21_X1 U6656 ( .B1(n5667), .B2(n5495), .A(n5477), .ZN(U2843) );
  AOI22_X1 U6657 ( .A1(n5890), .A2(n6492), .B1(n5493), .B2(EBX_REG_15__SCAN_IN), .ZN(n5478) );
  OAI21_X1 U6658 ( .B1(n5541), .B2(n5490), .A(n5478), .ZN(U2844) );
  AOI22_X1 U6659 ( .A1(n5909), .A2(n6492), .B1(n5493), .B2(EBX_REG_14__SCAN_IN), .ZN(n5479) );
  OAI21_X1 U6660 ( .B1(n5545), .B2(n5490), .A(n5479), .ZN(U2845) );
  OAI222_X1 U6661 ( .A1(n5912), .A2(n5497), .B1(n6495), .B2(n5286), .C1(n5490), 
        .C2(n5548), .ZN(U2846) );
  AOI22_X1 U6662 ( .A1(n5933), .A2(n6492), .B1(n5493), .B2(EBX_REG_12__SCAN_IN), .ZN(n5480) );
  OAI21_X1 U6663 ( .B1(n5694), .B2(n5495), .A(n5480), .ZN(U2847) );
  OAI222_X1 U6664 ( .A1(n5936), .A2(n5497), .B1(n5481), .B2(n6495), .C1(n5708), 
        .C2(n5490), .ZN(U2848) );
  OAI21_X1 U6665 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n6485) );
  NOR2_X1 U6666 ( .A1(n3159), .A2(n5485), .ZN(n5486) );
  OR2_X1 U6667 ( .A1(n5007), .A2(n5486), .ZN(n6472) );
  OAI22_X1 U6668 ( .A1(n6472), .A2(n5497), .B1(n5487), .B2(n6495), .ZN(n5488)
         );
  INV_X1 U6669 ( .A(n5488), .ZN(n5489) );
  OAI21_X1 U6670 ( .B1(n6485), .B2(n5495), .A(n5489), .ZN(U2850) );
  INV_X1 U6671 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5491) );
  OAI222_X1 U6672 ( .A1(n5492), .A2(n5497), .B1(n5491), .B2(n6495), .C1(n5490), 
        .C2(n5556), .ZN(U2851) );
  AOI22_X1 U6673 ( .A1(n6562), .A2(n6492), .B1(n5493), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5494) );
  OAI21_X1 U6674 ( .B1(n5558), .B2(n5495), .A(n5494), .ZN(U2852) );
  OAI22_X1 U6675 ( .A1(n5498), .A2(n5497), .B1(n5496), .B2(n6495), .ZN(n5499)
         );
  AOI21_X1 U6676 ( .B1(n5747), .B2(n6493), .A(n5499), .ZN(n5500) );
  INV_X1 U6677 ( .A(n5500), .ZN(U2854) );
  AOI22_X1 U6678 ( .A1(n5535), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5542), .ZN(n5502) );
  NAND2_X1 U6679 ( .A1(n5536), .A2(DATAI_13_), .ZN(n5501) );
  OAI211_X1 U6680 ( .C1(n5571), .C2(n5561), .A(n5502), .B(n5501), .ZN(U2862)
         );
  AOI22_X1 U6681 ( .A1(n5535), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5542), .ZN(n5504) );
  NAND2_X1 U6682 ( .A1(n5536), .A2(DATAI_12_), .ZN(n5503) );
  OAI211_X1 U6683 ( .C1(n5505), .C2(n5561), .A(n5504), .B(n5503), .ZN(U2863)
         );
  AOI22_X1 U6684 ( .A1(n5535), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5542), .ZN(n5507) );
  NAND2_X1 U6685 ( .A1(n5536), .A2(DATAI_11_), .ZN(n5506) );
  OAI211_X1 U6686 ( .C1(n5583), .C2(n5561), .A(n5507), .B(n5506), .ZN(U2864)
         );
  AOI22_X1 U6687 ( .A1(n5535), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5542), .ZN(n5509) );
  NAND2_X1 U6688 ( .A1(n5536), .A2(DATAI_10_), .ZN(n5508) );
  OAI211_X1 U6689 ( .C1(n5510), .C2(n5561), .A(n5509), .B(n5508), .ZN(U2865)
         );
  AOI22_X1 U6690 ( .A1(n5535), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5542), .ZN(n5512) );
  NAND2_X1 U6691 ( .A1(n5536), .A2(DATAI_9_), .ZN(n5511) );
  OAI211_X1 U6692 ( .C1(n5513), .C2(n5561), .A(n5512), .B(n5511), .ZN(U2866)
         );
  AOI22_X1 U6693 ( .A1(n5535), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5542), .ZN(n5515) );
  NAND2_X1 U6694 ( .A1(n5536), .A2(DATAI_8_), .ZN(n5514) );
  OAI211_X1 U6695 ( .C1(n5516), .C2(n5561), .A(n5515), .B(n5514), .ZN(U2867)
         );
  AOI22_X1 U6696 ( .A1(n5535), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5542), .ZN(n5518) );
  NAND2_X1 U6697 ( .A1(n5536), .A2(DATAI_7_), .ZN(n5517) );
  OAI211_X1 U6698 ( .C1(n5519), .C2(n5561), .A(n5518), .B(n5517), .ZN(U2868)
         );
  AOI22_X1 U6699 ( .A1(n5535), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5542), .ZN(n5521) );
  NAND2_X1 U6700 ( .A1(n5536), .A2(DATAI_6_), .ZN(n5520) );
  OAI211_X1 U6701 ( .C1(n5612), .C2(n5561), .A(n5521), .B(n5520), .ZN(U2869)
         );
  AOI22_X1 U6702 ( .A1(n5535), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5542), .ZN(n5523) );
  NAND2_X1 U6703 ( .A1(n5536), .A2(DATAI_5_), .ZN(n5522) );
  OAI211_X1 U6704 ( .C1(n5524), .C2(n5561), .A(n5523), .B(n5522), .ZN(U2870)
         );
  AOI22_X1 U6705 ( .A1(n5535), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5542), .ZN(n5526) );
  NAND2_X1 U6706 ( .A1(n5536), .A2(DATAI_4_), .ZN(n5525) );
  OAI211_X1 U6707 ( .C1(n5628), .C2(n5561), .A(n5526), .B(n5525), .ZN(U2871)
         );
  AOI22_X1 U6708 ( .A1(n5535), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5542), .ZN(n5528) );
  NAND2_X1 U6709 ( .A1(n5536), .A2(DATAI_3_), .ZN(n5527) );
  OAI211_X1 U6710 ( .C1(n5635), .C2(n5561), .A(n5528), .B(n5527), .ZN(U2872)
         );
  AOI22_X1 U6711 ( .A1(n5535), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5542), .ZN(n5530) );
  NAND2_X1 U6712 ( .A1(n5536), .A2(DATAI_2_), .ZN(n5529) );
  OAI211_X1 U6713 ( .C1(n5531), .C2(n5561), .A(n5530), .B(n5529), .ZN(U2873)
         );
  AOI22_X1 U6714 ( .A1(n5535), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5542), .ZN(n5533) );
  NAND2_X1 U6715 ( .A1(n5536), .A2(DATAI_1_), .ZN(n5532) );
  OAI211_X1 U6716 ( .C1(n5534), .C2(n5561), .A(n5533), .B(n5532), .ZN(U2874)
         );
  AOI22_X1 U6717 ( .A1(n5535), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5542), .ZN(n5538) );
  NAND2_X1 U6718 ( .A1(n5536), .A2(DATAI_0_), .ZN(n5537) );
  OAI211_X1 U6719 ( .C1(n5667), .C2(n5561), .A(n5538), .B(n5537), .ZN(U2875)
         );
  OAI222_X1 U6720 ( .A1(n5541), .A2(n5561), .B1(n5559), .B2(n5540), .C1(n5539), 
        .C2(n5560), .ZN(U2876) );
  INV_X1 U6721 ( .A(n5560), .ZN(n5543) );
  AOI22_X1 U6722 ( .A1(n5543), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5542), .ZN(n5544) );
  OAI21_X1 U6723 ( .B1(n5545), .B2(n5561), .A(n5544), .ZN(U2877) );
  INV_X1 U6724 ( .A(DATAI_13_), .ZN(n5546) );
  OAI222_X1 U6725 ( .A1(n5548), .A2(n5561), .B1(n5559), .B2(n5547), .C1(n5546), 
        .C2(n5560), .ZN(U2878) );
  INV_X1 U6726 ( .A(DATAI_12_), .ZN(n5549) );
  OAI222_X1 U6727 ( .A1(n5694), .A2(n5561), .B1(n5559), .B2(n5550), .C1(n5549), 
        .C2(n5560), .ZN(U2879) );
  INV_X1 U6728 ( .A(DATAI_11_), .ZN(n5551) );
  OAI222_X1 U6729 ( .A1(n5708), .A2(n5561), .B1(n5559), .B2(n5552), .C1(n5551), 
        .C2(n5560), .ZN(U2880) );
  INV_X1 U6730 ( .A(DATAI_10_), .ZN(n5553) );
  OAI222_X1 U6731 ( .A1(n5717), .A2(n5561), .B1(n5559), .B2(n5554), .C1(n5553), 
        .C2(n5560), .ZN(U2881) );
  OAI222_X1 U6732 ( .A1(n6485), .A2(n5561), .B1(n5560), .B2(n5555), .C1(n5559), 
        .C2(n4701), .ZN(U2882) );
  INV_X1 U6733 ( .A(DATAI_8_), .ZN(n6905) );
  OAI222_X1 U6734 ( .A1(n5556), .A2(n5561), .B1(n5560), .B2(n6905), .C1(n5559), 
        .C2(n4723), .ZN(U2883) );
  OAI222_X1 U6735 ( .A1(n5561), .A2(n5558), .B1(n5560), .B2(n5557), .C1(n5559), 
        .C2(n4707), .ZN(U2884) );
  INV_X1 U6736 ( .A(n5747), .ZN(n5562) );
  OAI222_X1 U6737 ( .A1(n5562), .A2(n5561), .B1(n5560), .B2(n7066), .C1(n5559), 
        .C2(n4782), .ZN(U2886) );
  NOR2_X1 U6738 ( .A1(n6522), .A2(n5563), .ZN(n5764) );
  NOR2_X1 U6739 ( .A1(n6541), .A2(n5564), .ZN(n5565) );
  AOI211_X1 U6740 ( .C1(n6531), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5764), 
        .B(n5565), .ZN(n5570) );
  NAND2_X1 U6741 ( .A1(n5759), .A2(n6535), .ZN(n5569) );
  OAI211_X1 U6742 ( .C1(n5571), .C2(n5718), .A(n5569), .B(n5570), .ZN(U2957)
         );
  INV_X1 U6743 ( .A(n5598), .ZN(n5573) );
  NOR2_X1 U6744 ( .A1(n6522), .A2(n7018), .ZN(n5774) );
  AOI21_X1 U6745 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5774), 
        .ZN(n5575) );
  OAI21_X1 U6746 ( .B1(n5576), .B2(n6541), .A(n5575), .ZN(n5577) );
  AOI21_X1 U6747 ( .B1(n5578), .B2(n6536), .A(n5577), .ZN(n5579) );
  OAI21_X1 U6748 ( .B1(n5750), .B2(n5778), .A(n5579), .ZN(U2958) );
  NAND2_X1 U6749 ( .A1(n3137), .A2(n5580), .ZN(n5581) );
  XNOR2_X1 U6750 ( .A(n5581), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5787)
         );
  NAND2_X1 U6751 ( .A1(n6586), .A2(REIP_REG_27__SCAN_IN), .ZN(n5781) );
  OAI21_X1 U6752 ( .B1(n5722), .B2(n5582), .A(n5781), .ZN(n5585) );
  NOR2_X1 U6753 ( .A1(n5583), .A2(n5718), .ZN(n5584) );
  OAI21_X1 U6754 ( .B1(n5787), .B2(n5750), .A(n5587), .ZN(U2959) );
  NAND2_X1 U6755 ( .A1(n3222), .A2(n5589), .ZN(n5590) );
  XNOR2_X1 U6756 ( .A(n3098), .B(n5590), .ZN(n5795) );
  NAND2_X1 U6757 ( .A1(n5725), .A2(n5591), .ZN(n5592) );
  NAND2_X1 U6758 ( .A1(n6586), .A2(REIP_REG_26__SCAN_IN), .ZN(n5789) );
  OAI211_X1 U6759 ( .C1(n5722), .C2(n5593), .A(n5592), .B(n5789), .ZN(n5594)
         );
  AOI21_X1 U6760 ( .B1(n5595), .B2(n6536), .A(n5594), .ZN(n5596) );
  OAI21_X1 U6761 ( .B1(n5795), .B2(n5750), .A(n5596), .ZN(U2960) );
  AOI21_X1 U6762 ( .B1(n5599), .B2(n5598), .A(n5597), .ZN(n5803) );
  NAND2_X1 U6763 ( .A1(n6586), .A2(REIP_REG_25__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U6764 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5600)
         );
  OAI211_X1 U6765 ( .C1(n6541), .C2(n5601), .A(n5797), .B(n5600), .ZN(n5602)
         );
  AOI21_X1 U6766 ( .B1(n5603), .B2(n6536), .A(n5602), .ZN(n5604) );
  OAI21_X1 U6767 ( .B1(n5803), .B2(n5750), .A(n5604), .ZN(U2961) );
  AOI21_X1 U6768 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5641), .A(n5605), 
        .ZN(n5610) );
  INV_X1 U6769 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5606) );
  XOR2_X1 U6770 ( .A(n5610), .B(n5609), .Z(n5820) );
  NAND2_X1 U6771 ( .A1(n6586), .A2(REIP_REG_22__SCAN_IN), .ZN(n5814) );
  OAI21_X1 U6772 ( .B1(n5722), .B2(n5611), .A(n5814), .ZN(n5614) );
  NOR2_X1 U6773 ( .A1(n5612), .A2(n5718), .ZN(n5613) );
  AOI211_X1 U6774 ( .C1(n5725), .C2(n5615), .A(n5614), .B(n5613), .ZN(n5616)
         );
  OAI21_X1 U6775 ( .B1(n5820), .B2(n5750), .A(n5616), .ZN(U2964) );
  AOI21_X1 U6776 ( .B1(n5618), .B2(n5617), .A(n5608), .ZN(n5828) );
  NAND2_X1 U6777 ( .A1(n5725), .A2(n5619), .ZN(n5620) );
  NAND2_X1 U6778 ( .A1(n6586), .A2(REIP_REG_21__SCAN_IN), .ZN(n5822) );
  OAI211_X1 U6779 ( .C1(n5722), .C2(n5621), .A(n5620), .B(n5822), .ZN(n5622)
         );
  AOI21_X1 U6780 ( .B1(n5623), .B2(n6536), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6781 ( .B1(n5828), .B2(n5750), .A(n5624), .ZN(U2965) );
  OAI21_X1 U6782 ( .B1(n5627), .B2(n5626), .A(n5625), .ZN(n5844) );
  NAND2_X1 U6783 ( .A1(n6586), .A2(REIP_REG_20__SCAN_IN), .ZN(n5835) );
  OAI21_X1 U6784 ( .B1(n5722), .B2(n3275), .A(n5835), .ZN(n5630) );
  NOR2_X1 U6785 ( .A1(n5628), .A2(n5718), .ZN(n5629) );
  AOI211_X1 U6786 ( .C1(n5725), .C2(n5631), .A(n5630), .B(n5629), .ZN(n5632)
         );
  OAI21_X1 U6787 ( .B1(n5750), .B2(n5844), .A(n5632), .ZN(U2966) );
  XOR2_X1 U6788 ( .A(n5634), .B(n5633), .Z(n5852) );
  INV_X1 U6789 ( .A(n5635), .ZN(n5639) );
  NAND2_X1 U6790 ( .A1(n6586), .A2(REIP_REG_19__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U6791 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5636)
         );
  OAI211_X1 U6792 ( .C1(n6541), .C2(n5637), .A(n5846), .B(n5636), .ZN(n5638)
         );
  AOI21_X1 U6793 ( .B1(n5639), .B2(n6536), .A(n5638), .ZN(n5640) );
  OAI21_X1 U6794 ( .B1(n5852), .B2(n5750), .A(n5640), .ZN(U2967) );
  NAND3_X1 U6795 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5646) );
  BUF_X1 U6796 ( .A(n5642), .Z(n5643) );
  NAND4_X1 U6797 ( .A1(n5643), .A2(n5644), .A3(n5829), .A4(n5878), .ZN(n5645)
         );
  OAI21_X1 U6798 ( .B1(n5646), .B2(n5643), .A(n5645), .ZN(n5647) );
  XNOR2_X1 U6799 ( .A(n5647), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5861)
         );
  NAND2_X1 U6800 ( .A1(n5725), .A2(n5648), .ZN(n5649) );
  NAND2_X1 U6801 ( .A1(n6586), .A2(REIP_REG_18__SCAN_IN), .ZN(n5855) );
  OAI211_X1 U6802 ( .C1(n5722), .C2(n3274), .A(n5649), .B(n5855), .ZN(n5650)
         );
  AOI21_X1 U6803 ( .B1(n5651), .B2(n6536), .A(n5650), .ZN(n5652) );
  OAI21_X1 U6804 ( .B1(n5861), .B2(n5750), .A(n5652), .ZN(U2968) );
  MUX2_X1 U6805 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n5699), .S(n5643), 
        .Z(n5653) );
  OAI21_X1 U6806 ( .B1(n5878), .B2(n5720), .A(n5653), .ZN(n5654) );
  XNOR2_X1 U6807 ( .A(n5654), .B(n5829), .ZN(n5869) );
  NAND2_X1 U6808 ( .A1(n5725), .A2(n5655), .ZN(n5656) );
  NAND2_X1 U6809 ( .A1(n6586), .A2(REIP_REG_17__SCAN_IN), .ZN(n5862) );
  OAI211_X1 U6810 ( .C1(n5722), .C2(n5657), .A(n5656), .B(n5862), .ZN(n5658)
         );
  AOI21_X1 U6811 ( .B1(n5659), .B2(n6536), .A(n5658), .ZN(n5660) );
  OAI21_X1 U6812 ( .B1(n5869), .B2(n5750), .A(n5660), .ZN(U2969) );
  XNOR2_X1 U6813 ( .A(n5720), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5661)
         );
  XNOR2_X1 U6814 ( .A(n5643), .B(n5661), .ZN(n5870) );
  NAND2_X1 U6815 ( .A1(n5870), .A2(n6535), .ZN(n5666) );
  NOR2_X1 U6816 ( .A1(n6522), .A2(n5662), .ZN(n5877) );
  NOR2_X1 U6817 ( .A1(n6541), .A2(n5663), .ZN(n5664) );
  AOI211_X1 U6818 ( .C1(n6531), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5877), 
        .B(n5664), .ZN(n5665) );
  OAI211_X1 U6819 ( .C1(n5718), .C2(n5667), .A(n5666), .B(n5665), .ZN(U2970)
         );
  AOI21_X1 U6820 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5699), .A(n3142), 
        .ZN(n5669) );
  XNOR2_X1 U6821 ( .A(n5720), .B(n5875), .ZN(n5668) );
  XNOR2_X1 U6822 ( .A(n5669), .B(n5668), .ZN(n5893) );
  NOR2_X1 U6823 ( .A1(n6522), .A2(n6971), .ZN(n5887) );
  AOI21_X1 U6824 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5887), 
        .ZN(n5670) );
  OAI21_X1 U6825 ( .B1(n5671), .B2(n6541), .A(n5670), .ZN(n5672) );
  AOI21_X1 U6826 ( .B1(n5673), .B2(n6536), .A(n5672), .ZN(n5674) );
  OAI21_X1 U6827 ( .B1(n5893), .B2(n5750), .A(n5674), .ZN(U2971) );
  OAI21_X1 U6828 ( .B1(n5699), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5675), 
        .ZN(n5677) );
  INV_X1 U6829 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5907) );
  XNOR2_X1 U6830 ( .A(n5720), .B(n5907), .ZN(n5676) );
  XNOR2_X1 U6831 ( .A(n5677), .B(n5676), .ZN(n5911) );
  NAND2_X1 U6832 ( .A1(n6586), .A2(REIP_REG_14__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U6833 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5678)
         );
  OAI211_X1 U6834 ( .C1(n6541), .C2(n5679), .A(n5906), .B(n5678), .ZN(n5680)
         );
  AOI21_X1 U6835 ( .B1(n5681), .B2(n6536), .A(n5680), .ZN(n5682) );
  OAI21_X1 U6836 ( .B1(n5911), .B2(n5750), .A(n5682), .ZN(U2972) );
  XOR2_X1 U6837 ( .A(n5683), .B(n5684), .Z(n5925) );
  NAND2_X1 U6838 ( .A1(n6586), .A2(REIP_REG_13__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U6839 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5685)
         );
  OAI211_X1 U6840 ( .C1(n6541), .C2(n5686), .A(n5918), .B(n5685), .ZN(n5687)
         );
  AOI21_X1 U6841 ( .B1(n5688), .B2(n6536), .A(n5687), .ZN(n5689) );
  OAI21_X1 U6842 ( .B1(n5925), .B2(n5750), .A(n5689), .ZN(U2973) );
  NAND2_X1 U6843 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  XNOR2_X1 U6844 ( .A(n3113), .B(n5693), .ZN(n5935) );
  NAND2_X1 U6845 ( .A1(n6586), .A2(REIP_REG_12__SCAN_IN), .ZN(n5930) );
  OAI21_X1 U6846 ( .B1(n5722), .B2(n3277), .A(n5930), .ZN(n5696) );
  NOR2_X1 U6847 ( .A1(n5694), .A2(n5718), .ZN(n5695) );
  AOI211_X1 U6848 ( .C1(n5725), .C2(n5697), .A(n5696), .B(n5695), .ZN(n5698)
         );
  OAI21_X1 U6849 ( .B1(n5935), .B2(n5750), .A(n5698), .ZN(U2974) );
  AOI21_X1 U6850 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5699), .A(n3141), 
        .ZN(n5712) );
  INV_X1 U6851 ( .A(n5712), .ZN(n5702) );
  AOI21_X1 U6852 ( .B1(n5712), .B2(n5700), .A(n5641), .ZN(n5701) );
  AOI21_X1 U6853 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5702), .A(n5701), 
        .ZN(n5704) );
  XNOR2_X1 U6854 ( .A(n5720), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5703)
         );
  XNOR2_X1 U6855 ( .A(n5704), .B(n5703), .ZN(n5944) );
  NOR2_X1 U6856 ( .A1(n6522), .A2(n4662), .ZN(n5937) );
  AOI21_X1 U6857 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5937), 
        .ZN(n5707) );
  OR2_X1 U6858 ( .A1(n6541), .A2(n5705), .ZN(n5706) );
  OAI211_X1 U6859 ( .C1(n5708), .C2(n5718), .A(n5707), .B(n5706), .ZN(n5709)
         );
  AOI21_X1 U6860 ( .B1(n5944), .B2(n6535), .A(n5709), .ZN(n5710) );
  INV_X1 U6861 ( .A(n5710), .ZN(U2975) );
  XNOR2_X1 U6862 ( .A(n5720), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5711)
         );
  XNOR2_X1 U6863 ( .A(n5712), .B(n5711), .ZN(n6545) );
  NAND2_X1 U6864 ( .A1(n6545), .A2(n6535), .ZN(n5716) );
  NOR2_X1 U6865 ( .A1(n6522), .A2(n5326), .ZN(n6542) );
  NOR2_X1 U6866 ( .A1(n6541), .A2(n5713), .ZN(n5714) );
  AOI211_X1 U6867 ( .C1(n6531), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6542), 
        .B(n5714), .ZN(n5715) );
  OAI211_X1 U6868 ( .C1(n5718), .C2(n5717), .A(n5716), .B(n5715), .ZN(U2976)
         );
  XNOR2_X1 U6869 ( .A(n5720), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5721)
         );
  XNOR2_X1 U6870 ( .A(n5719), .B(n5721), .ZN(n5958) );
  NAND2_X1 U6871 ( .A1(n6586), .A2(REIP_REG_9__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U6872 ( .B1(n5722), .B2(n7041), .A(n5953), .ZN(n5724) );
  NOR2_X1 U6873 ( .A1(n6485), .A2(n5718), .ZN(n5723) );
  AOI211_X1 U6874 ( .C1(n5725), .C2(n6486), .A(n5724), .B(n5723), .ZN(n5726)
         );
  OAI21_X1 U6875 ( .B1(n5958), .B2(n5750), .A(n5726), .ZN(U2977) );
  OAI21_X1 U6876 ( .B1(n5727), .B2(n5729), .A(n5728), .ZN(n6553) );
  NAND2_X1 U6877 ( .A1(n6586), .A2(REIP_REG_8__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U6878 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5730)
         );
  OAI211_X1 U6879 ( .C1(n6541), .C2(n5731), .A(n6550), .B(n5730), .ZN(n5732)
         );
  AOI21_X1 U6880 ( .B1(n5733), .B2(n6536), .A(n5732), .ZN(n5734) );
  OAI21_X1 U6881 ( .B1(n5750), .B2(n6553), .A(n5734), .ZN(U2978) );
  OAI21_X1 U6882 ( .B1(n5735), .B2(n5737), .A(n5736), .ZN(n6563) );
  NAND2_X1 U6883 ( .A1(n6586), .A2(REIP_REG_7__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U6884 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5738)
         );
  OAI211_X1 U6885 ( .C1(n6541), .C2(n5739), .A(n6560), .B(n5738), .ZN(n5740)
         );
  AOI21_X1 U6886 ( .B1(n5741), .B2(n6536), .A(n5740), .ZN(n5742) );
  OAI21_X1 U6887 ( .B1(n5750), .B2(n6563), .A(n5742), .ZN(U2979) );
  NAND2_X1 U6888 ( .A1(n6531), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5743)
         );
  OAI211_X1 U6889 ( .C1(n6541), .C2(n5745), .A(n5744), .B(n5743), .ZN(n5746)
         );
  AOI21_X1 U6890 ( .B1(n5747), .B2(n6536), .A(n5746), .ZN(n5748) );
  OAI21_X1 U6891 ( .B1(n5750), .B2(n5749), .A(n5748), .ZN(U2981) );
  AOI211_X1 U6892 ( .C1(n5762), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5751), .B(n5761), .ZN(n5755) );
  NAND2_X1 U6893 ( .A1(n5751), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5753) );
  OAI21_X1 U6894 ( .B1(n5760), .B2(n5753), .A(n5752), .ZN(n5754) );
  OAI21_X1 U6895 ( .B1(n5758), .B2(n5957), .A(n5757), .ZN(U2988) );
  NAND2_X1 U6896 ( .A1(n5759), .A2(n6602), .ZN(n5768) );
  INV_X1 U6897 ( .A(n5760), .ZN(n5766) );
  INV_X1 U6898 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5765) );
  NOR3_X1 U6899 ( .A1(n5762), .A2(n5761), .A3(n5765), .ZN(n5763) );
  AOI211_X1 U6900 ( .C1(n5766), .C2(n5765), .A(n5764), .B(n5763), .ZN(n5767)
         );
  OAI211_X1 U6901 ( .C1(n5951), .C2(n5769), .A(n5768), .B(n5767), .ZN(U2989)
         );
  INV_X1 U6902 ( .A(n5770), .ZN(n5783) );
  NOR3_X1 U6903 ( .A1(n5783), .A2(n5772), .A3(n5771), .ZN(n5773) );
  AOI211_X1 U6904 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5780), .A(n5774), .B(n5773), .ZN(n5777) );
  NAND2_X1 U6905 ( .A1(n5775), .A2(n6597), .ZN(n5776) );
  INV_X1 U6906 ( .A(n5779), .ZN(n5785) );
  NAND2_X1 U6907 ( .A1(n5780), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5782) );
  OAI211_X1 U6908 ( .C1(n5783), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5782), .B(n5781), .ZN(n5784) );
  AOI21_X1 U6909 ( .B1(n5785), .B2(n6597), .A(n5784), .ZN(n5786) );
  OAI21_X1 U6910 ( .B1(n5787), .B2(n5957), .A(n5786), .ZN(U2991) );
  INV_X1 U6911 ( .A(n5788), .ZN(n5793) );
  XNOR2_X1 U6912 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U6913 ( .A1(n5796), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5790) );
  OAI211_X1 U6914 ( .C1(n5791), .C2(n5799), .A(n5790), .B(n5789), .ZN(n5792)
         );
  AOI21_X1 U6915 ( .B1(n5793), .B2(n6597), .A(n5792), .ZN(n5794) );
  OAI21_X1 U6916 ( .B1(n5795), .B2(n5957), .A(n5794), .ZN(U2992) );
  NAND2_X1 U6917 ( .A1(n5796), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5798) );
  OAI211_X1 U6918 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5799), .A(n5798), .B(n5797), .ZN(n5800) );
  AOI21_X1 U6919 ( .B1(n5801), .B2(n6597), .A(n5800), .ZN(n5802) );
  OAI21_X1 U6920 ( .B1(n5803), .B2(n5957), .A(n5802), .ZN(U2993) );
  AOI211_X1 U6921 ( .C1(n7060), .C2(n5806), .A(n5805), .B(n5804), .ZN(n5807)
         );
  AOI211_X1 U6922 ( .C1(n5809), .C2(n6597), .A(n5808), .B(n5807), .ZN(n5810)
         );
  OAI21_X1 U6923 ( .B1(n5811), .B2(n5957), .A(n5810), .ZN(U2994) );
  NOR3_X1 U6924 ( .A1(n5824), .A2(n5813), .A3(n5812), .ZN(n5817) );
  INV_X1 U6925 ( .A(n5821), .ZN(n5815) );
  OAI21_X1 U6926 ( .B1(n5815), .B2(n7077), .A(n5814), .ZN(n5816) );
  AOI211_X1 U6927 ( .C1(n5818), .C2(n6597), .A(n5817), .B(n5816), .ZN(n5819)
         );
  OAI21_X1 U6928 ( .B1(n5820), .B2(n5957), .A(n5819), .ZN(U2996) );
  NAND2_X1 U6929 ( .A1(n5821), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5823) );
  OAI211_X1 U6930 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5824), .A(n5823), .B(n5822), .ZN(n5825) );
  AOI21_X1 U6931 ( .B1(n5826), .B2(n6597), .A(n5825), .ZN(n5827) );
  OAI21_X1 U6932 ( .B1(n5828), .B2(n5957), .A(n5827), .ZN(U2997) );
  NOR2_X1 U6933 ( .A1(n5830), .A2(n5829), .ZN(n5832) );
  OAI21_X1 U6934 ( .B1(n5832), .B2(n6599), .A(n5831), .ZN(n5867) );
  NOR2_X1 U6935 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5833), .ZN(n5834)
         );
  NOR2_X1 U6936 ( .A1(n5867), .A2(n5834), .ZN(n5857) );
  OAI21_X1 U6937 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5950), .A(n5857), 
        .ZN(n5845) );
  INV_X1 U6938 ( .A(n5835), .ZN(n5840) );
  INV_X1 U6939 ( .A(n5836), .ZN(n5848) );
  NOR3_X1 U6940 ( .A1(n5848), .A2(n5838), .A3(n5837), .ZN(n5839) );
  AOI211_X1 U6941 ( .C1(n5845), .C2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5840), .B(n5839), .ZN(n5843) );
  NAND2_X1 U6942 ( .A1(n5841), .A2(n6597), .ZN(n5842) );
  OAI211_X1 U6943 ( .C1(n5844), .C2(n5957), .A(n5843), .B(n5842), .ZN(U2998)
         );
  NAND2_X1 U6944 ( .A1(n5845), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5847) );
  OAI211_X1 U6945 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5848), .A(n5847), .B(n5846), .ZN(n5849) );
  AOI21_X1 U6946 ( .B1(n5850), .B2(n6597), .A(n5849), .ZN(n5851) );
  OAI21_X1 U6947 ( .B1(n5852), .B2(n5957), .A(n5851), .ZN(U2999) );
  INV_X1 U6948 ( .A(n5863), .ZN(n5853) );
  NAND3_X1 U6949 ( .A1(n5853), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5856), .ZN(n5854) );
  OAI211_X1 U6950 ( .C1(n5857), .C2(n5856), .A(n5855), .B(n5854), .ZN(n5858)
         );
  AOI21_X1 U6951 ( .B1(n5859), .B2(n6597), .A(n5858), .ZN(n5860) );
  OAI21_X1 U6952 ( .B1(n5861), .B2(n5957), .A(n5860), .ZN(U3000) );
  OAI21_X1 U6953 ( .B1(n5863), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5862), 
        .ZN(n5866) );
  NOR2_X1 U6954 ( .A1(n5864), .A2(n5951), .ZN(n5865) );
  AOI211_X1 U6955 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5867), .A(n5866), .B(n5865), .ZN(n5868) );
  OAI21_X1 U6956 ( .B1(n5869), .B2(n5957), .A(n5868), .ZN(U3001) );
  INV_X1 U6957 ( .A(n5870), .ZN(n5886) );
  INV_X1 U6958 ( .A(n5871), .ZN(n5872) );
  NOR2_X1 U6959 ( .A1(n6599), .A2(n5872), .ZN(n5873) );
  NOR2_X1 U6960 ( .A1(n5874), .A2(n5873), .ZN(n5941) );
  OAI21_X1 U6961 ( .B1(n5950), .B2(n5879), .A(n5941), .ZN(n5889) );
  AND2_X1 U6962 ( .A1(n5879), .A2(n5875), .ZN(n5876) );
  AND2_X1 U6963 ( .A1(n5938), .A2(n5876), .ZN(n5888) );
  OAI21_X1 U6964 ( .B1(n5889), .B2(n5888), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5882) );
  INV_X1 U6965 ( .A(n5877), .ZN(n5881) );
  NAND4_X1 U6966 ( .A1(n5938), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5879), .A4(n5878), .ZN(n5880) );
  NAND3_X1 U6967 ( .A1(n5882), .A2(n5881), .A3(n5880), .ZN(n5883) );
  AOI21_X1 U6968 ( .B1(n5884), .B2(n6597), .A(n5883), .ZN(n5885) );
  OAI21_X1 U6969 ( .B1(n5886), .B2(n5957), .A(n5885), .ZN(U3002) );
  AOI211_X1 U6970 ( .C1(n5889), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5888), .B(n5887), .ZN(n5892) );
  NAND2_X1 U6971 ( .A1(n5890), .A2(n6597), .ZN(n5891) );
  OAI211_X1 U6972 ( .C1(n5893), .C2(n5957), .A(n5892), .B(n5891), .ZN(U3003)
         );
  INV_X1 U6973 ( .A(n5941), .ZN(n5927) );
  NAND3_X1 U6974 ( .A1(n5894), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5916), 
        .ZN(n5897) );
  INV_X1 U6975 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5895) );
  NOR2_X1 U6976 ( .A1(n5940), .A2(n5928), .ZN(n5898) );
  NAND2_X1 U6977 ( .A1(n5895), .A2(n5898), .ZN(n5914) );
  AOI21_X1 U6978 ( .B1(n5897), .B2(n5896), .A(n5914), .ZN(n5913) );
  INV_X1 U6979 ( .A(n5898), .ZN(n5899) );
  NAND2_X1 U6980 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  OAI21_X1 U6981 ( .B1(n5904), .B2(n5902), .A(n5901), .ZN(n5903) );
  NOR3_X1 U6982 ( .A1(n5927), .A2(n5913), .A3(n5903), .ZN(n5921) );
  NAND3_X1 U6983 ( .A1(n5938), .A2(n5904), .A3(n5907), .ZN(n5905) );
  OAI211_X1 U6984 ( .C1(n5921), .C2(n5907), .A(n5906), .B(n5905), .ZN(n5908)
         );
  AOI21_X1 U6985 ( .B1(n5909), .B2(n6597), .A(n5908), .ZN(n5910) );
  OAI21_X1 U6986 ( .B1(n5911), .B2(n5957), .A(n5910), .ZN(U3004) );
  INV_X1 U6987 ( .A(n5912), .ZN(n5923) );
  NOR2_X1 U6988 ( .A1(n5913), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5920)
         );
  INV_X1 U6989 ( .A(n5914), .ZN(n5915) );
  NAND3_X1 U6990 ( .A1(n5917), .A2(n5916), .A3(n5915), .ZN(n5919) );
  OAI211_X1 U6991 ( .C1(n5921), .C2(n5920), .A(n5919), .B(n5918), .ZN(n5922)
         );
  AOI21_X1 U6992 ( .B1(n6597), .B2(n5923), .A(n5922), .ZN(n5924) );
  OAI21_X1 U6993 ( .B1(n5925), .B2(n5957), .A(n5924), .ZN(U3005) );
  NAND2_X1 U6994 ( .A1(n5950), .A2(n5926), .ZN(n5949) );
  OAI211_X1 U6995 ( .C1(n5927), .C2(n5940), .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(n5949), .ZN(n5931) );
  NAND3_X1 U6996 ( .A1(n5938), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n5928), .ZN(n5929) );
  NAND3_X1 U6997 ( .A1(n5931), .A2(n5930), .A3(n5929), .ZN(n5932) );
  AOI21_X1 U6998 ( .B1(n6597), .B2(n5933), .A(n5932), .ZN(n5934) );
  OAI21_X1 U6999 ( .B1(n5935), .B2(n5957), .A(n5934), .ZN(U3006) );
  NOR2_X1 U7000 ( .A1(n5936), .A2(n5951), .ZN(n5943) );
  AOI21_X1 U7001 ( .B1(n5938), .B2(n5940), .A(n5937), .ZN(n5939) );
  OAI21_X1 U7002 ( .B1(n5941), .B2(n5940), .A(n5939), .ZN(n5942) );
  AOI211_X1 U7003 ( .C1(n5944), .C2(n6602), .A(n5943), .B(n5942), .ZN(n5945)
         );
  INV_X1 U7004 ( .A(n5945), .ZN(U3007) );
  INV_X1 U7005 ( .A(n5946), .ZN(n5952) );
  NAND2_X1 U7006 ( .A1(n5948), .A2(n5947), .ZN(n6594) );
  NAND2_X1 U7007 ( .A1(n6598), .A2(n6594), .ZN(n6590) );
  OAI21_X1 U7008 ( .B1(n5952), .B2(n6590), .A(n5949), .ZN(n6568) );
  OAI21_X1 U7009 ( .B1(n5950), .B2(n6554), .A(n6568), .ZN(n6544) );
  NOR2_X1 U7010 ( .A1(n6472), .A2(n5951), .ZN(n5955) );
  NOR2_X1 U7011 ( .A1(n5952), .A2(n6593), .ZN(n6564) );
  NAND2_X1 U7012 ( .A1(n6554), .A2(n6564), .ZN(n6549) );
  OAI21_X1 U7013 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6549), .A(n5953), 
        .ZN(n5954) );
  AOI211_X1 U7014 ( .C1(n6544), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5955), 
        .B(n5954), .ZN(n5956) );
  OAI21_X1 U7015 ( .B1(n5958), .B2(n5957), .A(n5956), .ZN(U3009) );
  AOI21_X1 U7016 ( .B1(n5960), .B2(n5962), .A(n5961), .ZN(n5964) );
  NAND2_X1 U7017 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  NAND2_X1 U7018 ( .A1(n5966), .A2(n5965), .ZN(n5975) );
  NAND2_X1 U7019 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n3112), .ZN(n5967) );
  INV_X1 U7020 ( .A(n5967), .ZN(n5968) );
  MUX2_X1 U7021 ( .A(n5968), .B(n5967), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n5972) );
  INV_X1 U7022 ( .A(n5969), .ZN(n5971) );
  AOI21_X1 U7023 ( .B1(n3524), .B2(n3339), .A(n5970), .ZN(n5977) );
  AOI22_X1 U7024 ( .A1(n5973), .A2(n5972), .B1(n5971), .B2(n5977), .ZN(n5974)
         );
  NAND2_X1 U7025 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  AOI21_X1 U7026 ( .B1(n4889), .B2(n3199), .A(n5976), .ZN(n6409) );
  INV_X1 U7027 ( .A(n5977), .ZN(n5978) );
  OAI22_X1 U7028 ( .A1(n6409), .A2(n5980), .B1(n5979), .B2(n5978), .ZN(n5982)
         );
  MUX2_X1 U7029 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5982), .S(n5981), 
        .Z(U3456) );
  AND2_X1 U7030 ( .A1(n6022), .A2(n6140), .ZN(n6056) );
  NAND3_X1 U7031 ( .A1(n6982), .A2(n6421), .A3(n6417), .ZN(n6024) );
  OR2_X1 U7032 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6024), .ZN(n6013)
         );
  NOR2_X1 U7033 ( .A1(n6372), .A2(n6218), .ZN(n6104) );
  OAI21_X1 U7034 ( .B1(n6104), .B2(n6956), .A(n6063), .ZN(n6101) );
  AOI211_X1 U7035 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6013), .A(n6347), .B(
        n6101), .ZN(n5986) );
  OAI21_X1 U7036 ( .B1(n6056), .B2(n6016), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5984) );
  NAND2_X1 U7037 ( .A1(n6224), .A2(n3130), .ZN(n6020) );
  NAND3_X1 U7038 ( .A1(n5984), .A2(n6691), .A3(n6020), .ZN(n5985) );
  NAND2_X1 U7039 ( .A1(n6012), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5993) );
  INV_X1 U7040 ( .A(n6020), .ZN(n5987) );
  NAND2_X1 U7041 ( .A1(n5987), .A2(n6691), .ZN(n5990) );
  NAND2_X1 U7042 ( .A1(n6104), .A2(n6297), .ZN(n5989) );
  OAI22_X1 U7043 ( .A1(n6014), .A2(n6644), .B1(n6013), .B2(n6688), .ZN(n5991)
         );
  AOI21_X1 U7044 ( .B1(n6016), .B2(n6634), .A(n5991), .ZN(n5992) );
  OAI211_X1 U7045 ( .C1(n6019), .C2(n6707), .A(n5993), .B(n5992), .ZN(U3020)
         );
  NAND2_X1 U7046 ( .A1(n6012), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5996) );
  OAI22_X1 U7047 ( .A1(n6014), .A2(n6649), .B1(n6013), .B2(n6708), .ZN(n5994)
         );
  AOI21_X1 U7048 ( .B1(n6016), .B2(n6646), .A(n5994), .ZN(n5995) );
  OAI211_X1 U7049 ( .C1(n6019), .C2(n6709), .A(n5996), .B(n5995), .ZN(U3021)
         );
  NAND2_X1 U7050 ( .A1(n6012), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5999) );
  OAI22_X1 U7051 ( .A1(n6014), .A2(n6655), .B1(n6013), .B2(n6715), .ZN(n5997)
         );
  AOI21_X1 U7052 ( .B1(n6016), .B2(n6651), .A(n5997), .ZN(n5998) );
  OAI211_X1 U7053 ( .C1(n6019), .C2(n6716), .A(n5999), .B(n5998), .ZN(U3022)
         );
  NAND2_X1 U7054 ( .A1(n6012), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6002) );
  OAI22_X1 U7055 ( .A1(n6014), .A2(n6661), .B1(n6013), .B2(n6722), .ZN(n6000)
         );
  AOI21_X1 U7056 ( .B1(n6016), .B2(n6657), .A(n6000), .ZN(n6001) );
  OAI211_X1 U7057 ( .C1(n6019), .C2(n6723), .A(n6002), .B(n6001), .ZN(U3023)
         );
  NAND2_X1 U7058 ( .A1(n6012), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6005) );
  OAI22_X1 U7059 ( .A1(n6014), .A2(n6665), .B1(n6013), .B2(n6729), .ZN(n6003)
         );
  AOI21_X1 U7060 ( .B1(n6016), .B2(n6662), .A(n6003), .ZN(n6004) );
  OAI211_X1 U7061 ( .C1(n6019), .C2(n6733), .A(n6005), .B(n6004), .ZN(U3024)
         );
  NAND2_X1 U7062 ( .A1(n6012), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6008) );
  OAI22_X1 U7063 ( .A1(n6014), .A2(n6671), .B1(n6013), .B2(n6734), .ZN(n6006)
         );
  AOI21_X1 U7064 ( .B1(n6016), .B2(n6667), .A(n6006), .ZN(n6007) );
  OAI211_X1 U7065 ( .C1(n6019), .C2(n6735), .A(n6008), .B(n6007), .ZN(U3025)
         );
  NAND2_X1 U7066 ( .A1(n6012), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6011) );
  OAI22_X1 U7067 ( .A1(n6014), .A2(n6676), .B1(n6013), .B2(n6739), .ZN(n6009)
         );
  AOI21_X1 U7068 ( .B1(n6016), .B2(n6673), .A(n6009), .ZN(n6010) );
  OAI211_X1 U7069 ( .C1(n6019), .C2(n6740), .A(n6011), .B(n6010), .ZN(U3026)
         );
  NAND2_X1 U7070 ( .A1(n6012), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6018) );
  OAI22_X1 U7071 ( .A1(n6014), .A2(n6685), .B1(n6013), .B2(n6745), .ZN(n6015)
         );
  AOI21_X1 U7072 ( .B1(n6016), .B2(n6681), .A(n6015), .ZN(n6017) );
  OAI211_X1 U7073 ( .C1(n6019), .C2(n6752), .A(n6018), .B(n6017), .ZN(U3027)
         );
  OAI21_X1 U7074 ( .B1(n6022), .B2(n6698), .A(n6338), .ZN(n6025) );
  NOR2_X1 U7075 ( .A1(n6907), .A2(n6024), .ZN(n6053) );
  INV_X1 U7076 ( .A(n6053), .ZN(n6030) );
  OAI21_X1 U7077 ( .B1(n6020), .B2(n6135), .A(n6030), .ZN(n6023) );
  INV_X1 U7078 ( .A(n6024), .ZN(n6021) );
  INV_X1 U7079 ( .A(n6096), .ZN(n6060) );
  INV_X1 U7080 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6029) );
  INV_X1 U7081 ( .A(n6023), .ZN(n6026) );
  AOI22_X1 U7082 ( .A1(n6026), .A2(n6025), .B1(n6024), .B2(n6698), .ZN(n6027)
         );
  NAND2_X1 U7083 ( .A1(n6638), .A2(n6027), .ZN(n6052) );
  INV_X1 U7084 ( .A(n6052), .ZN(n6028) );
  OAI22_X1 U7085 ( .A1(n6688), .A2(n6030), .B1(n6029), .B2(n6028), .ZN(n6031)
         );
  AOI21_X1 U7086 ( .B1(n6060), .B2(n6641), .A(n6031), .ZN(n6033) );
  NAND2_X1 U7087 ( .A1(n6056), .A2(n6634), .ZN(n6032) );
  OAI211_X1 U7088 ( .C1(n6058), .C2(n6644), .A(n6033), .B(n6032), .ZN(U3028)
         );
  AOI22_X1 U7089 ( .A1(n6611), .A2(n6053), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n6052), .ZN(n6034) );
  OAI21_X1 U7090 ( .B1(n6096), .B2(n6709), .A(n6034), .ZN(n6035) );
  AOI21_X1 U7091 ( .B1(n6646), .B2(n6056), .A(n6035), .ZN(n6036) );
  OAI21_X1 U7092 ( .B1(n6058), .B2(n6649), .A(n6036), .ZN(U3029) );
  AOI22_X1 U7093 ( .A1(n6650), .A2(n6053), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n6052), .ZN(n6037) );
  OAI21_X1 U7094 ( .B1(n6096), .B2(n6716), .A(n6037), .ZN(n6038) );
  AOI21_X1 U7095 ( .B1(n6651), .B2(n6056), .A(n6038), .ZN(n6039) );
  OAI21_X1 U7096 ( .B1(n6058), .B2(n6655), .A(n6039), .ZN(U3030) );
  AOI22_X1 U7097 ( .A1(n6656), .A2(n6053), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n6052), .ZN(n6040) );
  OAI21_X1 U7098 ( .B1(n6096), .B2(n6723), .A(n6040), .ZN(n6041) );
  AOI21_X1 U7099 ( .B1(n6657), .B2(n6056), .A(n6041), .ZN(n6042) );
  OAI21_X1 U7100 ( .B1(n6058), .B2(n6661), .A(n6042), .ZN(U3031) );
  AOI22_X1 U7101 ( .A1(n6754), .A2(n6053), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n6052), .ZN(n6043) );
  OAI21_X1 U7102 ( .B1(n6096), .B2(n6733), .A(n6043), .ZN(n6044) );
  AOI21_X1 U7103 ( .B1(n6662), .B2(n6056), .A(n6044), .ZN(n6045) );
  OAI21_X1 U7104 ( .B1(n6058), .B2(n6665), .A(n6045), .ZN(U3032) );
  AOI22_X1 U7105 ( .A1(n6760), .A2(n6053), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n6052), .ZN(n6046) );
  OAI21_X1 U7106 ( .B1(n6096), .B2(n6735), .A(n6046), .ZN(n6047) );
  AOI21_X1 U7107 ( .B1(n6667), .B2(n6056), .A(n6047), .ZN(n6048) );
  OAI21_X1 U7108 ( .B1(n6058), .B2(n6671), .A(n6048), .ZN(U3033) );
  AOI22_X1 U7109 ( .A1(n6766), .A2(n6053), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n6052), .ZN(n6049) );
  OAI21_X1 U7110 ( .B1(n6096), .B2(n6740), .A(n6049), .ZN(n6050) );
  AOI21_X1 U7111 ( .B1(n6673), .B2(n6056), .A(n6050), .ZN(n6051) );
  OAI21_X1 U7112 ( .B1(n6058), .B2(n6676), .A(n6051), .ZN(U3034) );
  AOI22_X1 U7113 ( .A1(n6772), .A2(n6053), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n6052), .ZN(n6054) );
  OAI21_X1 U7114 ( .B1(n6096), .B2(n6752), .A(n6054), .ZN(n6055) );
  AOI21_X1 U7115 ( .B1(n6681), .B2(n6056), .A(n6055), .ZN(n6057) );
  OAI21_X1 U7116 ( .B1(n6058), .B2(n6685), .A(n6057), .ZN(U3035) );
  NOR2_X1 U7117 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6059), .ZN(n6067)
         );
  OAI21_X1 U7118 ( .B1(n6060), .B2(n6093), .A(n6338), .ZN(n6062) );
  INV_X1 U7119 ( .A(n6066), .ZN(n6061) );
  NAND2_X1 U7120 ( .A1(n6062), .A2(n6061), .ZN(n6064) );
  OAI21_X1 U7121 ( .B1(n6372), .B2(n6956), .A(n6063), .ZN(n6183) );
  NOR2_X1 U7122 ( .A1(n6347), .A2(n6183), .ZN(n6304) );
  NAND2_X1 U7123 ( .A1(n6089), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6070) );
  INV_X1 U7124 ( .A(n6297), .ZN(n6341) );
  NOR2_X1 U7125 ( .A1(n6341), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6065)
         );
  AOI22_X1 U7126 ( .A1(n6066), .A2(n6691), .B1(n6372), .B2(n6065), .ZN(n6091)
         );
  INV_X1 U7127 ( .A(n6067), .ZN(n6090) );
  OAI22_X1 U7128 ( .A1(n6091), .A2(n6644), .B1(n6090), .B2(n6688), .ZN(n6068)
         );
  AOI21_X1 U7129 ( .B1(n6093), .B2(n6641), .A(n6068), .ZN(n6069) );
  OAI211_X1 U7130 ( .C1(n6096), .C2(n6689), .A(n6070), .B(n6069), .ZN(U3036)
         );
  NAND2_X1 U7131 ( .A1(n6089), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6073) );
  OAI22_X1 U7132 ( .A1(n6091), .A2(n6649), .B1(n6090), .B2(n6708), .ZN(n6071)
         );
  AOI21_X1 U7133 ( .B1(n6093), .B2(n6612), .A(n6071), .ZN(n6072) );
  OAI211_X1 U7134 ( .C1(n6714), .C2(n6096), .A(n6073), .B(n6072), .ZN(U3037)
         );
  NAND2_X1 U7135 ( .A1(n6089), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6076) );
  OAI22_X1 U7136 ( .A1(n6091), .A2(n6655), .B1(n6090), .B2(n6715), .ZN(n6074)
         );
  AOI21_X1 U7137 ( .B1(n6093), .B2(n6652), .A(n6074), .ZN(n6075) );
  OAI211_X1 U7138 ( .C1(n6096), .C2(n6721), .A(n6076), .B(n6075), .ZN(U3038)
         );
  NAND2_X1 U7139 ( .A1(n6089), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6079) );
  OAI22_X1 U7140 ( .A1(n6091), .A2(n6661), .B1(n6090), .B2(n6722), .ZN(n6077)
         );
  AOI21_X1 U7141 ( .B1(n6093), .B2(n6658), .A(n6077), .ZN(n6078) );
  OAI211_X1 U7142 ( .C1(n6096), .C2(n6728), .A(n6079), .B(n6078), .ZN(U3039)
         );
  NAND2_X1 U7143 ( .A1(n6089), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6082) );
  OAI22_X1 U7144 ( .A1(n6091), .A2(n6665), .B1(n6090), .B2(n6729), .ZN(n6080)
         );
  AOI21_X1 U7145 ( .B1(n6093), .B2(n6756), .A(n6080), .ZN(n6081) );
  OAI211_X1 U7146 ( .C1(n6096), .C2(n6759), .A(n6082), .B(n6081), .ZN(U3040)
         );
  NAND2_X1 U7147 ( .A1(n6089), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6085) );
  OAI22_X1 U7148 ( .A1(n6091), .A2(n6671), .B1(n6090), .B2(n6734), .ZN(n6083)
         );
  AOI21_X1 U7149 ( .B1(n6093), .B2(n6762), .A(n6083), .ZN(n6084) );
  OAI211_X1 U7150 ( .C1(n6096), .C2(n6765), .A(n6085), .B(n6084), .ZN(U3041)
         );
  NAND2_X1 U7151 ( .A1(n6089), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6088) );
  OAI22_X1 U7152 ( .A1(n6091), .A2(n6676), .B1(n6090), .B2(n6739), .ZN(n6086)
         );
  AOI21_X1 U7153 ( .B1(n6093), .B2(n6768), .A(n6086), .ZN(n6087) );
  OAI211_X1 U7154 ( .C1(n6096), .C2(n6771), .A(n6088), .B(n6087), .ZN(U3042)
         );
  NAND2_X1 U7155 ( .A1(n6089), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6095) );
  OAI22_X1 U7156 ( .A1(n6091), .A2(n6685), .B1(n6090), .B2(n6745), .ZN(n6092)
         );
  AOI21_X1 U7157 ( .B1(n6093), .B2(n6777), .A(n6092), .ZN(n6094) );
  OAI211_X1 U7158 ( .C1(n6096), .C2(n6782), .A(n6095), .B(n6094), .ZN(U3043)
         );
  OR2_X1 U7159 ( .A1(n6099), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6143)
         );
  NOR2_X1 U7160 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6143), .ZN(n6105)
         );
  OAI21_X1 U7161 ( .B1(n6172), .B2(n6624), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6100) );
  NAND2_X1 U7162 ( .A1(n6348), .A2(n6178), .ZN(n6136) );
  AND2_X1 U7163 ( .A1(n6100), .A2(n6136), .ZN(n6102) );
  AOI211_X1 U7164 ( .C1(n6691), .C2(n6102), .A(n6297), .B(n6101), .ZN(n6103)
         );
  NAND2_X1 U7165 ( .A1(n6127), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6108) );
  NOR2_X1 U7166 ( .A1(n4889), .A2(n6698), .ZN(n6177) );
  AOI22_X1 U7167 ( .A1(n6177), .A2(n6348), .B1(n6347), .B2(n6104), .ZN(n6129)
         );
  INV_X1 U7168 ( .A(n6105), .ZN(n6128) );
  OAI22_X1 U7169 ( .A1(n6129), .A2(n6644), .B1(n6128), .B2(n6688), .ZN(n6106)
         );
  AOI21_X1 U7170 ( .B1(n6624), .B2(n6634), .A(n6106), .ZN(n6107) );
  OAI211_X1 U7171 ( .C1(n6707), .C2(n6133), .A(n6108), .B(n6107), .ZN(U3052)
         );
  NAND2_X1 U7172 ( .A1(n6127), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6111) );
  OAI22_X1 U7173 ( .A1(n6129), .A2(n6649), .B1(n6128), .B2(n6708), .ZN(n6109)
         );
  AOI21_X1 U7174 ( .B1(n6624), .B2(n6646), .A(n6109), .ZN(n6110) );
  OAI211_X1 U7175 ( .C1(n6133), .C2(n6709), .A(n6111), .B(n6110), .ZN(U3053)
         );
  NAND2_X1 U7176 ( .A1(n6127), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6114) );
  OAI22_X1 U7177 ( .A1(n6129), .A2(n6655), .B1(n6128), .B2(n6715), .ZN(n6112)
         );
  AOI21_X1 U7178 ( .B1(n6624), .B2(n6651), .A(n6112), .ZN(n6113) );
  OAI211_X1 U7179 ( .C1(n6133), .C2(n6716), .A(n6114), .B(n6113), .ZN(U3054)
         );
  NAND2_X1 U7180 ( .A1(n6127), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6117) );
  OAI22_X1 U7181 ( .A1(n6129), .A2(n6661), .B1(n6128), .B2(n6722), .ZN(n6115)
         );
  AOI21_X1 U7182 ( .B1(n6624), .B2(n6657), .A(n6115), .ZN(n6116) );
  OAI211_X1 U7183 ( .C1(n6133), .C2(n6723), .A(n6117), .B(n6116), .ZN(U3055)
         );
  NAND2_X1 U7184 ( .A1(n6127), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6120) );
  OAI22_X1 U7185 ( .A1(n6129), .A2(n6665), .B1(n6128), .B2(n6729), .ZN(n6118)
         );
  AOI21_X1 U7186 ( .B1(n6624), .B2(n6662), .A(n6118), .ZN(n6119) );
  OAI211_X1 U7187 ( .C1(n6133), .C2(n6733), .A(n6120), .B(n6119), .ZN(U3056)
         );
  NAND2_X1 U7188 ( .A1(n6127), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6123) );
  OAI22_X1 U7189 ( .A1(n6129), .A2(n6671), .B1(n6128), .B2(n6734), .ZN(n6121)
         );
  AOI21_X1 U7190 ( .B1(n6624), .B2(n6667), .A(n6121), .ZN(n6122) );
  OAI211_X1 U7191 ( .C1(n6133), .C2(n6735), .A(n6123), .B(n6122), .ZN(U3057)
         );
  NAND2_X1 U7192 ( .A1(n6127), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6126) );
  OAI22_X1 U7193 ( .A1(n6129), .A2(n6676), .B1(n6128), .B2(n6739), .ZN(n6124)
         );
  AOI21_X1 U7194 ( .B1(n6624), .B2(n6673), .A(n6124), .ZN(n6125) );
  OAI211_X1 U7195 ( .C1(n6133), .C2(n6740), .A(n6126), .B(n6125), .ZN(U3058)
         );
  NAND2_X1 U7196 ( .A1(n6127), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6132) );
  OAI22_X1 U7197 ( .A1(n6129), .A2(n6685), .B1(n6128), .B2(n6745), .ZN(n6130)
         );
  AOI21_X1 U7198 ( .B1(n6624), .B2(n6681), .A(n6130), .ZN(n6131) );
  OAI211_X1 U7199 ( .C1(n6133), .C2(n6752), .A(n6132), .B(n6131), .ZN(U3059)
         );
  OAI21_X1 U7200 ( .B1(n6134), .B2(n6698), .A(n6338), .ZN(n6144) );
  INV_X1 U7201 ( .A(n6169), .ZN(n6137) );
  NAND2_X1 U7202 ( .A1(n6138), .A2(n6137), .ZN(n6142) );
  INV_X1 U7203 ( .A(n6143), .ZN(n6139) );
  OR2_X1 U7204 ( .A1(n4221), .A2(n6140), .ZN(n6262) );
  INV_X1 U7205 ( .A(n6262), .ZN(n6141) );
  INV_X1 U7206 ( .A(n6142), .ZN(n6145) );
  AOI22_X1 U7207 ( .A1(n6145), .A2(n6144), .B1(n6143), .B2(n6698), .ZN(n6146)
         );
  NAND2_X1 U7208 ( .A1(n6638), .A2(n6146), .ZN(n6168) );
  AOI22_X1 U7209 ( .A1(n6633), .A2(n6169), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n6168), .ZN(n6147) );
  OAI21_X1 U7210 ( .B1(n6179), .B2(n6707), .A(n6147), .ZN(n6148) );
  AOI21_X1 U7211 ( .B1(n6172), .B2(n6634), .A(n6148), .ZN(n6149) );
  OAI21_X1 U7212 ( .B1(n6174), .B2(n6644), .A(n6149), .ZN(U3060) );
  AOI22_X1 U7213 ( .A1(n6611), .A2(n6169), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n6168), .ZN(n6150) );
  OAI21_X1 U7214 ( .B1(n6179), .B2(n6709), .A(n6150), .ZN(n6151) );
  AOI21_X1 U7215 ( .B1(n6172), .B2(n6646), .A(n6151), .ZN(n6152) );
  OAI21_X1 U7216 ( .B1(n6174), .B2(n6649), .A(n6152), .ZN(U3061) );
  AOI22_X1 U7217 ( .A1(n6650), .A2(n6169), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n6168), .ZN(n6153) );
  OAI21_X1 U7218 ( .B1(n6179), .B2(n6716), .A(n6153), .ZN(n6154) );
  AOI21_X1 U7219 ( .B1(n6172), .B2(n6651), .A(n6154), .ZN(n6155) );
  OAI21_X1 U7220 ( .B1(n6174), .B2(n6655), .A(n6155), .ZN(U3062) );
  AOI22_X1 U7221 ( .A1(n6656), .A2(n6169), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n6168), .ZN(n6156) );
  OAI21_X1 U7222 ( .B1(n6179), .B2(n6723), .A(n6156), .ZN(n6157) );
  AOI21_X1 U7223 ( .B1(n6172), .B2(n6657), .A(n6157), .ZN(n6158) );
  OAI21_X1 U7224 ( .B1(n6174), .B2(n6661), .A(n6158), .ZN(U3063) );
  AOI22_X1 U7225 ( .A1(n6754), .A2(n6169), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n6168), .ZN(n6159) );
  OAI21_X1 U7226 ( .B1(n6179), .B2(n6733), .A(n6159), .ZN(n6160) );
  AOI21_X1 U7227 ( .B1(n6172), .B2(n6662), .A(n6160), .ZN(n6161) );
  OAI21_X1 U7228 ( .B1(n6174), .B2(n6665), .A(n6161), .ZN(U3064) );
  AOI22_X1 U7229 ( .A1(n6760), .A2(n6169), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n6168), .ZN(n6162) );
  OAI21_X1 U7230 ( .B1(n6179), .B2(n6735), .A(n6162), .ZN(n6163) );
  AOI21_X1 U7231 ( .B1(n6172), .B2(n6667), .A(n6163), .ZN(n6164) );
  OAI21_X1 U7232 ( .B1(n6174), .B2(n6671), .A(n6164), .ZN(U3065) );
  AOI22_X1 U7233 ( .A1(n6766), .A2(n6169), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n6168), .ZN(n6165) );
  OAI21_X1 U7234 ( .B1(n6179), .B2(n6740), .A(n6165), .ZN(n6166) );
  AOI21_X1 U7235 ( .B1(n6172), .B2(n6673), .A(n6166), .ZN(n6167) );
  OAI21_X1 U7236 ( .B1(n6174), .B2(n6676), .A(n6167), .ZN(U3066) );
  AOI22_X1 U7237 ( .A1(n6772), .A2(n6169), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n6168), .ZN(n6170) );
  OAI21_X1 U7238 ( .B1(n6179), .B2(n6752), .A(n6170), .ZN(n6171) );
  AOI21_X1 U7239 ( .B1(n6172), .B2(n6681), .A(n6171), .ZN(n6173) );
  OAI21_X1 U7240 ( .B1(n6174), .B2(n6685), .A(n6173), .ZN(U3067) );
  INV_X1 U7241 ( .A(n6636), .ZN(n6175) );
  INV_X1 U7242 ( .A(n6347), .ZN(n6370) );
  NOR2_X1 U7243 ( .A1(n6370), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6176)
         );
  AOI22_X1 U7244 ( .A1(n6177), .A2(n6373), .B1(n6372), .B2(n6176), .ZN(n6209)
         );
  NAND2_X1 U7245 ( .A1(n6907), .A2(n6640), .ZN(n6182) );
  INV_X1 U7246 ( .A(n6182), .ZN(n6207) );
  NAND2_X1 U7247 ( .A1(n6373), .A2(n6178), .ZN(n6630) );
  NAND2_X1 U7248 ( .A1(n6691), .A2(n6179), .ZN(n6180) );
  OAI21_X1 U7249 ( .B1(n6680), .B2(n6180), .A(n6338), .ZN(n6181) );
  AOI22_X1 U7250 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6182), .B1(n6630), .B2(
        n6181), .ZN(n6184) );
  NOR2_X1 U7251 ( .A1(n6297), .A2(n6183), .ZN(n6368) );
  NAND3_X1 U7252 ( .A1(n6982), .A2(n6184), .A3(n6368), .ZN(n6206) );
  AOI22_X1 U7253 ( .A1(n6633), .A2(n6207), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n6206), .ZN(n6185) );
  OAI21_X1 U7254 ( .B1(n6209), .B2(n6644), .A(n6185), .ZN(n6186) );
  AOI21_X1 U7255 ( .B1(n6211), .B2(n6634), .A(n6186), .ZN(n6187) );
  OAI21_X1 U7256 ( .B1(n6213), .B2(n6707), .A(n6187), .ZN(U3068) );
  AOI22_X1 U7257 ( .A1(n6611), .A2(n6207), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n6206), .ZN(n6188) );
  OAI21_X1 U7258 ( .B1(n6209), .B2(n6649), .A(n6188), .ZN(n6189) );
  AOI21_X1 U7259 ( .B1(n6211), .B2(n6646), .A(n6189), .ZN(n6190) );
  OAI21_X1 U7260 ( .B1(n6213), .B2(n6709), .A(n6190), .ZN(U3069) );
  AOI22_X1 U7261 ( .A1(n6650), .A2(n6207), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n6206), .ZN(n6191) );
  OAI21_X1 U7262 ( .B1(n6209), .B2(n6655), .A(n6191), .ZN(n6192) );
  AOI21_X1 U7263 ( .B1(n6211), .B2(n6651), .A(n6192), .ZN(n6193) );
  OAI21_X1 U7264 ( .B1(n6213), .B2(n6716), .A(n6193), .ZN(U3070) );
  AOI22_X1 U7265 ( .A1(n6656), .A2(n6207), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n6206), .ZN(n6194) );
  OAI21_X1 U7266 ( .B1(n6209), .B2(n6661), .A(n6194), .ZN(n6195) );
  AOI21_X1 U7267 ( .B1(n6211), .B2(n6657), .A(n6195), .ZN(n6196) );
  OAI21_X1 U7268 ( .B1(n6213), .B2(n6723), .A(n6196), .ZN(U3071) );
  AOI22_X1 U7269 ( .A1(n6754), .A2(n6207), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n6206), .ZN(n6197) );
  OAI21_X1 U7270 ( .B1(n6209), .B2(n6665), .A(n6197), .ZN(n6198) );
  AOI21_X1 U7271 ( .B1(n6211), .B2(n6662), .A(n6198), .ZN(n6199) );
  OAI21_X1 U7272 ( .B1(n6213), .B2(n6733), .A(n6199), .ZN(U3072) );
  AOI22_X1 U7273 ( .A1(n6760), .A2(n6207), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n6206), .ZN(n6200) );
  OAI21_X1 U7274 ( .B1(n6209), .B2(n6671), .A(n6200), .ZN(n6201) );
  AOI21_X1 U7275 ( .B1(n6211), .B2(n6667), .A(n6201), .ZN(n6202) );
  OAI21_X1 U7276 ( .B1(n6213), .B2(n6735), .A(n6202), .ZN(U3073) );
  AOI22_X1 U7277 ( .A1(n6766), .A2(n6207), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n6206), .ZN(n6203) );
  OAI21_X1 U7278 ( .B1(n6209), .B2(n6676), .A(n6203), .ZN(n6204) );
  AOI21_X1 U7279 ( .B1(n6211), .B2(n6673), .A(n6204), .ZN(n6205) );
  OAI21_X1 U7280 ( .B1(n6213), .B2(n6740), .A(n6205), .ZN(U3074) );
  AOI22_X1 U7281 ( .A1(n6772), .A2(n6207), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n6206), .ZN(n6208) );
  OAI21_X1 U7282 ( .B1(n6209), .B2(n6685), .A(n6208), .ZN(n6210) );
  AOI21_X1 U7283 ( .B1(n6211), .B2(n6681), .A(n6210), .ZN(n6212) );
  OAI21_X1 U7284 ( .B1(n6213), .B2(n6752), .A(n6212), .ZN(U3075) );
  OR2_X1 U7285 ( .A1(n4221), .A2(n6214), .ZN(n6215) );
  INV_X1 U7286 ( .A(n6335), .ZN(n6216) );
  NAND2_X1 U7287 ( .A1(n6636), .A2(n6216), .ZN(n6678) );
  AOI21_X1 U7288 ( .B1(n6291), .B2(n6678), .A(n7046), .ZN(n6217) );
  AOI211_X1 U7289 ( .C1(n3130), .C2(n4889), .A(n6698), .B(n6217), .ZN(n6223)
         );
  NAND3_X1 U7290 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6421), .A3(n6417), .ZN(n6259) );
  NOR2_X1 U7291 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6259), .ZN(n6226)
         );
  OAI21_X1 U7292 ( .B1(n6343), .B2(n6226), .A(n6370), .ZN(n6222) );
  INV_X1 U7293 ( .A(n6218), .ZN(n6219) );
  OR2_X1 U7294 ( .A1(n6219), .A2(n6372), .ZN(n6225) );
  AOI21_X1 U7295 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6225), .A(n6220), .ZN(
        n6342) );
  INV_X1 U7296 ( .A(n6342), .ZN(n6221) );
  NAND2_X1 U7297 ( .A1(n6248), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6229) );
  NOR2_X1 U7298 ( .A1(n6224), .A2(n6698), .ZN(n6374) );
  INV_X1 U7299 ( .A(n6225), .ZN(n6346) );
  AOI22_X1 U7300 ( .A1(n6374), .A2(n3130), .B1(n6297), .B2(n6346), .ZN(n6250)
         );
  INV_X1 U7301 ( .A(n6226), .ZN(n6249) );
  OAI22_X1 U7302 ( .A1(n6250), .A2(n6644), .B1(n6249), .B2(n6688), .ZN(n6227)
         );
  AOI21_X1 U7303 ( .B1(n6668), .B2(n6634), .A(n6227), .ZN(n6228) );
  OAI211_X1 U7304 ( .C1(n6291), .C2(n6707), .A(n6229), .B(n6228), .ZN(U3084)
         );
  NAND2_X1 U7305 ( .A1(n6248), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6232) );
  OAI22_X1 U7306 ( .A1(n6250), .A2(n6649), .B1(n6249), .B2(n6708), .ZN(n6230)
         );
  AOI21_X1 U7307 ( .B1(n6668), .B2(n6646), .A(n6230), .ZN(n6231) );
  OAI211_X1 U7308 ( .C1(n6291), .C2(n6709), .A(n6232), .B(n6231), .ZN(U3085)
         );
  NAND2_X1 U7309 ( .A1(n6248), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6235) );
  OAI22_X1 U7310 ( .A1(n6250), .A2(n6655), .B1(n6249), .B2(n6715), .ZN(n6233)
         );
  AOI21_X1 U7311 ( .B1(n6668), .B2(n6651), .A(n6233), .ZN(n6234) );
  OAI211_X1 U7312 ( .C1(n6291), .C2(n6716), .A(n6235), .B(n6234), .ZN(U3086)
         );
  NAND2_X1 U7313 ( .A1(n6248), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6238) );
  OAI22_X1 U7314 ( .A1(n6250), .A2(n6661), .B1(n6249), .B2(n6722), .ZN(n6236)
         );
  AOI21_X1 U7315 ( .B1(n6668), .B2(n6657), .A(n6236), .ZN(n6237) );
  OAI211_X1 U7316 ( .C1(n6291), .C2(n6723), .A(n6238), .B(n6237), .ZN(U3087)
         );
  NAND2_X1 U7317 ( .A1(n6248), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6241) );
  OAI22_X1 U7318 ( .A1(n6250), .A2(n6665), .B1(n6249), .B2(n6729), .ZN(n6239)
         );
  AOI21_X1 U7319 ( .B1(n6668), .B2(n6662), .A(n6239), .ZN(n6240) );
  OAI211_X1 U7320 ( .C1(n6291), .C2(n6733), .A(n6241), .B(n6240), .ZN(U3088)
         );
  NAND2_X1 U7321 ( .A1(n6248), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6244) );
  OAI22_X1 U7322 ( .A1(n6250), .A2(n6671), .B1(n6249), .B2(n6734), .ZN(n6242)
         );
  AOI21_X1 U7323 ( .B1(n6668), .B2(n6667), .A(n6242), .ZN(n6243) );
  OAI211_X1 U7324 ( .C1(n6291), .C2(n6735), .A(n6244), .B(n6243), .ZN(U3089)
         );
  NAND2_X1 U7325 ( .A1(n6248), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6247) );
  OAI22_X1 U7326 ( .A1(n6250), .A2(n6676), .B1(n6249), .B2(n6739), .ZN(n6245)
         );
  AOI21_X1 U7327 ( .B1(n6668), .B2(n6673), .A(n6245), .ZN(n6246) );
  OAI211_X1 U7328 ( .C1(n6291), .C2(n6740), .A(n6247), .B(n6246), .ZN(U3090)
         );
  NAND2_X1 U7329 ( .A1(n6248), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6253) );
  OAI22_X1 U7330 ( .A1(n6250), .A2(n6685), .B1(n6249), .B2(n6745), .ZN(n6251)
         );
  AOI21_X1 U7331 ( .B1(n6668), .B2(n6681), .A(n6251), .ZN(n6252) );
  OAI211_X1 U7332 ( .C1(n6291), .C2(n6752), .A(n6253), .B(n6252), .ZN(U3091)
         );
  NOR2_X1 U7333 ( .A1(n6907), .A2(n6259), .ZN(n6263) );
  AOI21_X1 U7334 ( .B1(n6254), .B2(n3130), .A(n6263), .ZN(n6261) );
  OR2_X1 U7335 ( .A1(n4221), .A2(n7046), .ZN(n6255) );
  OR2_X1 U7336 ( .A1(n6693), .A2(n6255), .ZN(n6256) );
  AND2_X1 U7337 ( .A1(n6256), .A2(n6691), .ZN(n6258) );
  AOI22_X1 U7338 ( .A1(n6261), .A2(n6258), .B1(n6698), .B2(n6259), .ZN(n6257)
         );
  NAND2_X1 U7339 ( .A1(n6638), .A2(n6257), .ZN(n6286) );
  INV_X1 U7340 ( .A(n6258), .ZN(n6260) );
  OAI22_X1 U7341 ( .A1(n6261), .A2(n6260), .B1(n6956), .B2(n6259), .ZN(n6285)
         );
  AOI22_X1 U7342 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6286), .B1(n6704), 
        .B2(n6285), .ZN(n6266) );
  OAI22_X1 U7343 ( .A1(n6329), .A2(n6707), .B1(n6688), .B2(n6287), .ZN(n6264)
         );
  INV_X1 U7344 ( .A(n6264), .ZN(n6265) );
  OAI211_X1 U7345 ( .C1(n6689), .C2(n6291), .A(n6266), .B(n6265), .ZN(U3092)
         );
  AOI22_X1 U7346 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6286), .B1(n6711), 
        .B2(n6285), .ZN(n6269) );
  OAI22_X1 U7347 ( .A1(n6329), .A2(n6709), .B1(n6708), .B2(n6287), .ZN(n6267)
         );
  INV_X1 U7348 ( .A(n6267), .ZN(n6268) );
  OAI211_X1 U7349 ( .C1(n6714), .C2(n6291), .A(n6269), .B(n6268), .ZN(U3093)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6286), .B1(n6718), 
        .B2(n6285), .ZN(n6272) );
  OAI22_X1 U7351 ( .A1(n6329), .A2(n6716), .B1(n6715), .B2(n6287), .ZN(n6270)
         );
  INV_X1 U7352 ( .A(n6270), .ZN(n6271) );
  OAI211_X1 U7353 ( .C1(n6721), .C2(n6291), .A(n6272), .B(n6271), .ZN(U3094)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6286), .B1(n6725), 
        .B2(n6285), .ZN(n6275) );
  OAI22_X1 U7355 ( .A1(n6329), .A2(n6723), .B1(n6722), .B2(n6287), .ZN(n6273)
         );
  INV_X1 U7356 ( .A(n6273), .ZN(n6274) );
  OAI211_X1 U7357 ( .C1(n6728), .C2(n6291), .A(n6275), .B(n6274), .ZN(U3095)
         );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6286), .B1(n6755), 
        .B2(n6285), .ZN(n6278) );
  OAI22_X1 U7359 ( .A1(n6329), .A2(n6733), .B1(n6729), .B2(n6287), .ZN(n6276)
         );
  INV_X1 U7360 ( .A(n6276), .ZN(n6277) );
  OAI211_X1 U7361 ( .C1(n6759), .C2(n6291), .A(n6278), .B(n6277), .ZN(U3096)
         );
  AOI22_X1 U7362 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6286), .B1(n6761), 
        .B2(n6285), .ZN(n6281) );
  OAI22_X1 U7363 ( .A1(n6329), .A2(n6735), .B1(n6734), .B2(n6287), .ZN(n6279)
         );
  INV_X1 U7364 ( .A(n6279), .ZN(n6280) );
  OAI211_X1 U7365 ( .C1(n6765), .C2(n6291), .A(n6281), .B(n6280), .ZN(U3097)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6286), .B1(n6767), 
        .B2(n6285), .ZN(n6284) );
  OAI22_X1 U7367 ( .A1(n6329), .A2(n6740), .B1(n6739), .B2(n6287), .ZN(n6282)
         );
  INV_X1 U7368 ( .A(n6282), .ZN(n6283) );
  OAI211_X1 U7369 ( .C1(n6771), .C2(n6291), .A(n6284), .B(n6283), .ZN(U3098)
         );
  AOI22_X1 U7370 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6286), .B1(n6774), 
        .B2(n6285), .ZN(n6290) );
  OAI22_X1 U7371 ( .A1(n6329), .A2(n6752), .B1(n6745), .B2(n6287), .ZN(n6288)
         );
  INV_X1 U7372 ( .A(n6288), .ZN(n6289) );
  OAI211_X1 U7373 ( .C1(n6782), .C2(n6291), .A(n6290), .B(n6289), .ZN(U3099)
         );
  NAND2_X1 U7374 ( .A1(n6746), .A2(n6329), .ZN(n6293) );
  NAND2_X1 U7375 ( .A1(n6293), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7376 ( .A1(n6294), .A2(n6691), .ZN(n6301) );
  INV_X1 U7377 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U7378 ( .A1(n6296), .A2(n4889), .ZN(n6300) );
  NAND3_X1 U7379 ( .A1(n6297), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6372), .ZN(n6298) );
  INV_X1 U7380 ( .A(n6300), .ZN(n6696) );
  NAND3_X1 U7381 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6421), .ZN(n6701) );
  NOR2_X1 U7382 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6701), .ZN(n6305)
         );
  OAI22_X1 U7383 ( .A1(n6301), .A2(n6696), .B1(n6305), .B2(n6343), .ZN(n6302)
         );
  INV_X1 U7384 ( .A(n6302), .ZN(n6303) );
  NAND2_X1 U7385 ( .A1(n6327), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6308)
         );
  INV_X1 U7386 ( .A(n6305), .ZN(n6328) );
  OAI22_X1 U7387 ( .A1(n6329), .A2(n6689), .B1(n6688), .B2(n6328), .ZN(n6306)
         );
  AOI21_X1 U7388 ( .B1(n6331), .B2(n6641), .A(n6306), .ZN(n6307) );
  OAI211_X1 U7389 ( .C1(n6644), .C2(n6334), .A(n6308), .B(n6307), .ZN(U3100)
         );
  NAND2_X1 U7390 ( .A1(n6327), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6311)
         );
  OAI22_X1 U7391 ( .A1(n6329), .A2(n6714), .B1(n6328), .B2(n6708), .ZN(n6309)
         );
  AOI21_X1 U7392 ( .B1(n6331), .B2(n6612), .A(n6309), .ZN(n6310) );
  OAI211_X1 U7393 ( .C1(n6334), .C2(n6649), .A(n6311), .B(n6310), .ZN(U3101)
         );
  NAND2_X1 U7394 ( .A1(n6327), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6314)
         );
  OAI22_X1 U7395 ( .A1(n6329), .A2(n6721), .B1(n6328), .B2(n6715), .ZN(n6312)
         );
  AOI21_X1 U7396 ( .B1(n6331), .B2(n6652), .A(n6312), .ZN(n6313) );
  OAI211_X1 U7397 ( .C1(n6334), .C2(n6655), .A(n6314), .B(n6313), .ZN(U3102)
         );
  NAND2_X1 U7398 ( .A1(n6327), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6317)
         );
  OAI22_X1 U7399 ( .A1(n6329), .A2(n6728), .B1(n6328), .B2(n6722), .ZN(n6315)
         );
  AOI21_X1 U7400 ( .B1(n6331), .B2(n6658), .A(n6315), .ZN(n6316) );
  OAI211_X1 U7401 ( .C1(n6334), .C2(n6661), .A(n6317), .B(n6316), .ZN(U3103)
         );
  NAND2_X1 U7402 ( .A1(n6327), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6320)
         );
  OAI22_X1 U7403 ( .A1(n6329), .A2(n6759), .B1(n6328), .B2(n6729), .ZN(n6318)
         );
  AOI21_X1 U7404 ( .B1(n6331), .B2(n6756), .A(n6318), .ZN(n6319) );
  OAI211_X1 U7405 ( .C1(n6334), .C2(n6665), .A(n6320), .B(n6319), .ZN(U3104)
         );
  NAND2_X1 U7406 ( .A1(n6327), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6323)
         );
  OAI22_X1 U7407 ( .A1(n6329), .A2(n6765), .B1(n6328), .B2(n6734), .ZN(n6321)
         );
  AOI21_X1 U7408 ( .B1(n6331), .B2(n6762), .A(n6321), .ZN(n6322) );
  OAI211_X1 U7409 ( .C1(n6334), .C2(n6671), .A(n6323), .B(n6322), .ZN(U3105)
         );
  NAND2_X1 U7410 ( .A1(n6327), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6326)
         );
  OAI22_X1 U7411 ( .A1(n6329), .A2(n6771), .B1(n6328), .B2(n6739), .ZN(n6324)
         );
  AOI21_X1 U7412 ( .B1(n6331), .B2(n6768), .A(n6324), .ZN(n6325) );
  OAI211_X1 U7413 ( .C1(n6334), .C2(n6676), .A(n6326), .B(n6325), .ZN(U3106)
         );
  NAND2_X1 U7414 ( .A1(n6327), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6333)
         );
  OAI22_X1 U7415 ( .A1(n6329), .A2(n6782), .B1(n6328), .B2(n6745), .ZN(n6330)
         );
  AOI21_X1 U7416 ( .B1(n6331), .B2(n6777), .A(n6330), .ZN(n6332) );
  OAI211_X1 U7417 ( .C1(n6334), .C2(n6685), .A(n6333), .B(n6332), .ZN(U3107)
         );
  INV_X1 U7418 ( .A(n6776), .ZN(n6336) );
  NAND3_X1 U7419 ( .A1(n6336), .A2(n6781), .A3(n6691), .ZN(n6339) );
  AOI22_X1 U7420 ( .A1(n6339), .A2(n6338), .B1(n6348), .B2(n6337), .ZN(n6345)
         );
  NOR2_X1 U7421 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6340), .ZN(n6773)
         );
  OAI211_X1 U7422 ( .C1(n6773), .C2(n6343), .A(n6342), .B(n6341), .ZN(n6344)
         );
  NAND2_X1 U7423 ( .A1(n6778), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6351)
         );
  AOI22_X1 U7424 ( .A1(n6374), .A2(n6348), .B1(n6347), .B2(n6346), .ZN(n6753)
         );
  INV_X1 U7425 ( .A(n6773), .ZN(n6358) );
  OAI22_X1 U7426 ( .A1(n6753), .A2(n6644), .B1(n6358), .B2(n6688), .ZN(n6349)
         );
  AOI21_X1 U7427 ( .B1(n6776), .B2(n6641), .A(n6349), .ZN(n6350) );
  OAI211_X1 U7428 ( .C1(n6781), .C2(n6689), .A(n6351), .B(n6350), .ZN(U3116)
         );
  NAND2_X1 U7429 ( .A1(n6778), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6354)
         );
  OAI22_X1 U7430 ( .A1(n6753), .A2(n6649), .B1(n6358), .B2(n6708), .ZN(n6352)
         );
  AOI21_X1 U7431 ( .B1(n6776), .B2(n6612), .A(n6352), .ZN(n6353) );
  OAI211_X1 U7432 ( .C1(n6781), .C2(n6714), .A(n6354), .B(n6353), .ZN(U3117)
         );
  NAND2_X1 U7433 ( .A1(n6778), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6357)
         );
  OAI22_X1 U7434 ( .A1(n6753), .A2(n6655), .B1(n6358), .B2(n6715), .ZN(n6355)
         );
  AOI21_X1 U7435 ( .B1(n6776), .B2(n6652), .A(n6355), .ZN(n6356) );
  OAI211_X1 U7436 ( .C1(n6781), .C2(n6721), .A(n6357), .B(n6356), .ZN(U3118)
         );
  NAND2_X1 U7437 ( .A1(n6778), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6361)
         );
  OAI22_X1 U7438 ( .A1(n6753), .A2(n6661), .B1(n6358), .B2(n6722), .ZN(n6359)
         );
  AOI21_X1 U7439 ( .B1(n6776), .B2(n6658), .A(n6359), .ZN(n6360) );
  OAI211_X1 U7440 ( .C1(n6781), .C2(n6728), .A(n6361), .B(n6360), .ZN(U3119)
         );
  INV_X1 U7441 ( .A(n6403), .ZN(n6363) );
  NOR3_X1 U7442 ( .A1(n6400), .A2(n6363), .A3(n6698), .ZN(n6365) );
  INV_X1 U7443 ( .A(n6373), .ZN(n6364) );
  OAI21_X1 U7444 ( .B1(n6365), .B2(n6809), .A(n6364), .ZN(n6369) );
  OR2_X1 U7445 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6366), .ZN(n6397)
         );
  AOI21_X1 U7446 ( .B1(n6397), .B2(STATE2_REG_3__SCAN_IN), .A(n6982), .ZN(
        n6367) );
  NAND3_X1 U7447 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n6396) );
  NAND2_X1 U7448 ( .A1(n6396), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6377)
         );
  NOR2_X1 U7449 ( .A1(n6370), .A2(n6982), .ZN(n6371) );
  AOI22_X1 U7450 ( .A1(n6374), .A2(n6373), .B1(n6372), .B2(n6371), .ZN(n6398)
         );
  OAI22_X1 U7451 ( .A1(n6398), .A2(n6644), .B1(n6397), .B2(n6688), .ZN(n6375)
         );
  AOI21_X1 U7452 ( .B1(n6400), .B2(n6634), .A(n6375), .ZN(n6376) );
  OAI211_X1 U7453 ( .C1(n6403), .C2(n6707), .A(n6377), .B(n6376), .ZN(U3132)
         );
  NAND2_X1 U7454 ( .A1(n6396), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6380)
         );
  OAI22_X1 U7455 ( .A1(n6398), .A2(n6649), .B1(n6397), .B2(n6708), .ZN(n6378)
         );
  AOI21_X1 U7456 ( .B1(n6400), .B2(n6646), .A(n6378), .ZN(n6379) );
  OAI211_X1 U7457 ( .C1(n6403), .C2(n6709), .A(n6380), .B(n6379), .ZN(U3133)
         );
  NAND2_X1 U7458 ( .A1(n6396), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6383)
         );
  OAI22_X1 U7459 ( .A1(n6398), .A2(n6655), .B1(n6397), .B2(n6715), .ZN(n6381)
         );
  AOI21_X1 U7460 ( .B1(n6400), .B2(n6651), .A(n6381), .ZN(n6382) );
  OAI211_X1 U7461 ( .C1(n6403), .C2(n6716), .A(n6383), .B(n6382), .ZN(U3134)
         );
  NAND2_X1 U7462 ( .A1(n6396), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6386)
         );
  OAI22_X1 U7463 ( .A1(n6398), .A2(n6661), .B1(n6397), .B2(n6722), .ZN(n6384)
         );
  AOI21_X1 U7464 ( .B1(n6400), .B2(n6657), .A(n6384), .ZN(n6385) );
  OAI211_X1 U7465 ( .C1(n6403), .C2(n6723), .A(n6386), .B(n6385), .ZN(U3135)
         );
  NAND2_X1 U7466 ( .A1(n6396), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6389)
         );
  OAI22_X1 U7467 ( .A1(n6398), .A2(n6665), .B1(n6397), .B2(n6729), .ZN(n6387)
         );
  AOI21_X1 U7468 ( .B1(n6400), .B2(n6662), .A(n6387), .ZN(n6388) );
  OAI211_X1 U7469 ( .C1(n6403), .C2(n6733), .A(n6389), .B(n6388), .ZN(U3136)
         );
  NAND2_X1 U7470 ( .A1(n6396), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6392)
         );
  OAI22_X1 U7471 ( .A1(n6398), .A2(n6671), .B1(n6397), .B2(n6734), .ZN(n6390)
         );
  AOI21_X1 U7472 ( .B1(n6400), .B2(n6667), .A(n6390), .ZN(n6391) );
  OAI211_X1 U7473 ( .C1(n6403), .C2(n6735), .A(n6392), .B(n6391), .ZN(U3137)
         );
  NAND2_X1 U7474 ( .A1(n6396), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6395)
         );
  OAI22_X1 U7475 ( .A1(n6398), .A2(n6676), .B1(n6397), .B2(n6739), .ZN(n6393)
         );
  AOI21_X1 U7476 ( .B1(n6400), .B2(n6673), .A(n6393), .ZN(n6394) );
  OAI211_X1 U7477 ( .C1(n6403), .C2(n6740), .A(n6395), .B(n6394), .ZN(U3138)
         );
  NAND2_X1 U7478 ( .A1(n6396), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6402)
         );
  OAI22_X1 U7479 ( .A1(n6398), .A2(n6685), .B1(n6397), .B2(n6745), .ZN(n6399)
         );
  AOI21_X1 U7480 ( .B1(n6400), .B2(n6681), .A(n6399), .ZN(n6401) );
  OAI211_X1 U7481 ( .C1(n6403), .C2(n6752), .A(n6402), .B(n6401), .ZN(U3139)
         );
  INV_X1 U7482 ( .A(n6404), .ZN(n6439) );
  INV_X1 U7483 ( .A(n6405), .ZN(n6438) );
  INV_X1 U7484 ( .A(n6415), .ZN(n6429) );
  NAND2_X1 U7485 ( .A1(n6429), .A2(n3112), .ZN(n6406) );
  OAI21_X1 U7486 ( .B1(n6407), .B2(n6429), .A(n6406), .ZN(n6436) );
  NOR2_X1 U7487 ( .A1(n6415), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6408)
         );
  AOI21_X1 U7488 ( .B1(n6409), .B2(n6415), .A(n6408), .ZN(n6435) );
  INV_X1 U7489 ( .A(n6410), .ZN(n6411) );
  OAI211_X1 U7490 ( .C1(n6413), .C2(n6412), .A(n6411), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6418) );
  OAI211_X1 U7491 ( .C1(n6417), .C2(n6418), .A(n6416), .B(n6415), .ZN(n6420)
         );
  NAND2_X1 U7492 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  INV_X1 U7493 ( .A(n6435), .ZN(n6422) );
  INV_X1 U7494 ( .A(n6423), .ZN(n6431) );
  NOR2_X1 U7495 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6427) );
  OAI211_X1 U7496 ( .C1(n6427), .C2(n6426), .A(n6425), .B(n6424), .ZN(n6428)
         );
  AOI21_X1 U7497 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6429), .A(n6428), 
        .ZN(n6430) );
  OAI21_X1 U7498 ( .B1(n6432), .B2(n6431), .A(n6430), .ZN(n6433) );
  AOI211_X1 U7499 ( .C1(n6436), .C2(n6435), .A(n6434), .B(n6433), .ZN(n6789)
         );
  AOI22_X1 U7500 ( .A1(n6789), .A2(n6440), .B1(n6502), .B2(READY_N), .ZN(n6437) );
  AOI21_X1 U7501 ( .B1(n6439), .B2(n6438), .A(n6437), .ZN(n6804) );
  NOR2_X1 U7502 ( .A1(n7091), .A2(READY_N), .ZN(n6441) );
  AOI21_X1 U7503 ( .B1(n6442), .B2(n6441), .A(n6440), .ZN(n6446) );
  NOR2_X1 U7504 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6443), .ZN(n6795) );
  NAND2_X1 U7505 ( .A1(n7091), .A2(n6956), .ZN(n6792) );
  OAI211_X1 U7506 ( .C1(n6804), .C2(n6795), .A(STATE2_REG_1__SCAN_IN), .B(
        n6792), .ZN(n6445) );
  OAI211_X1 U7507 ( .C1(n6804), .C2(n6446), .A(n6445), .B(n6444), .ZN(U3149)
         );
  AND2_X1 U7508 ( .A1(n6506), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7509 ( .A(n6447), .ZN(n6454) );
  AOI21_X1 U7510 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n6449), .A(n6448), .ZN(
        n6450) );
  NAND2_X1 U7511 ( .A1(n6454), .A2(n6450), .ZN(U2788) );
  INV_X1 U7512 ( .A(n6451), .ZN(n6452) );
  OAI21_X1 U7513 ( .B1(n6452), .B2(n6788), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6453) );
  OAI21_X1 U7514 ( .B1(n6454), .B2(n7091), .A(n6453), .ZN(U2790) );
  NOR2_X1 U7515 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6456) );
  OAI21_X1 U7516 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6456), .A(n6824), .ZN(n6455)
         );
  OAI21_X1 U7517 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6824), .A(n6455), .ZN(
        U2791) );
  OAI21_X1 U7518 ( .B1(n6456), .B2(BS16_N), .A(n6801), .ZN(n6799) );
  OAI21_X1 U7519 ( .B1(n6801), .B2(n7046), .A(n6799), .ZN(U2792) );
  NOR4_X1 U7520 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6460) );
  NOR4_X1 U7521 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6459) );
  NOR4_X1 U7522 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6458) );
  NOR4_X1 U7523 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6457) );
  NAND4_X1 U7524 ( .A1(n6460), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n6466)
         );
  NOR4_X1 U7525 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6464) );
  AOI211_X1 U7526 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_27__SCAN_IN), .B(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6463) );
  NOR4_X1 U7527 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n6462) );
  NOR4_X1 U7528 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n6461) );
  NAND4_X1 U7529 ( .A1(n6464), .A2(n6463), .A3(n6462), .A4(n6461), .ZN(n6465)
         );
  INV_X1 U7530 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6468) );
  NOR3_X1 U7531 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6469) );
  OAI21_X1 U7532 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6469), .A(n6818), .ZN(n6467)
         );
  OAI21_X1 U7533 ( .B1(n6818), .B2(n6468), .A(n6467), .ZN(U2794) );
  INV_X1 U7534 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6800) );
  AOI21_X1 U7535 ( .B1(n6888), .B2(n6800), .A(n6469), .ZN(n6471) );
  INV_X1 U7536 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6470) );
  INV_X1 U7537 ( .A(n6818), .ZN(n6821) );
  AOI22_X1 U7538 ( .A1(n6818), .A2(n6471), .B1(n6470), .B2(n6821), .ZN(U2795)
         );
  INV_X1 U7539 ( .A(n6472), .ZN(n6474) );
  NAND2_X1 U7540 ( .A1(n6474), .A2(n6473), .ZN(n6484) );
  NAND2_X1 U7541 ( .A1(n6475), .A2(REIP_REG_9__SCAN_IN), .ZN(n6483) );
  INV_X1 U7542 ( .A(n6476), .ZN(n6482) );
  OAI21_X1 U7543 ( .B1(n6478), .B2(n7041), .A(n6477), .ZN(n6479) );
  AOI21_X1 U7544 ( .B1(n6480), .B2(EBX_REG_9__SCAN_IN), .A(n6479), .ZN(n6481)
         );
  AND4_X1 U7545 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n6491)
         );
  INV_X1 U7546 ( .A(n6485), .ZN(n6489) );
  AOI22_X1 U7547 ( .A1(n6489), .A2(n6488), .B1(n6487), .B2(n6486), .ZN(n6490)
         );
  NAND2_X1 U7548 ( .A1(n6491), .A2(n6490), .ZN(U2818) );
  INV_X1 U7549 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6902) );
  AOI22_X1 U7550 ( .A1(n6518), .A2(n6493), .B1(n6492), .B2(n6570), .ZN(n6494)
         );
  OAI21_X1 U7551 ( .B1(n6902), .B2(n6495), .A(n6494), .ZN(U2853) );
  AOI22_X1 U7552 ( .A1(n6498), .A2(EAX_REG_30__SCAN_IN), .B1(n6506), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n6496) );
  OAI21_X1 U7553 ( .B1(n6508), .B2(n7019), .A(n6496), .ZN(U2893) );
  AOI22_X1 U7554 ( .A1(n6498), .A2(EAX_REG_28__SCAN_IN), .B1(n6506), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6497) );
  OAI21_X1 U7555 ( .B1(n6508), .B2(n6904), .A(n6497), .ZN(U2895) );
  INV_X1 U7556 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7557 ( .A1(n6498), .A2(EAX_REG_23__SCAN_IN), .B1(n6502), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n6499) );
  OAI21_X1 U7558 ( .B1(n6942), .B2(n6504), .A(n6499), .ZN(U2900) );
  AOI22_X1 U7559 ( .A1(n6506), .A2(DATAO_REG_15__SCAN_IN), .B1(n6505), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n6500) );
  OAI21_X1 U7560 ( .B1(n6508), .B2(n6944), .A(n6500), .ZN(U2908) );
  AOI22_X1 U7561 ( .A1(n6506), .A2(DATAO_REG_13__SCAN_IN), .B1(n6505), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6501) );
  OAI21_X1 U7562 ( .B1(n6508), .B2(n7013), .A(n6501), .ZN(U2910) );
  INV_X1 U7563 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U7564 ( .A1(n6505), .A2(EAX_REG_12__SCAN_IN), .B1(n6502), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6503) );
  OAI21_X1 U7565 ( .B1(n6997), .B2(n6504), .A(n6503), .ZN(U2911) );
  AOI22_X1 U7566 ( .A1(n6506), .A2(DATAO_REG_5__SCAN_IN), .B1(n6505), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6507) );
  OAI21_X1 U7567 ( .B1(n6508), .B2(n4781), .A(n6507), .ZN(U2918) );
  AOI22_X1 U7568 ( .A1(n6825), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6509), .ZN(n6511) );
  NAND2_X1 U7569 ( .A1(n6511), .A2(n6510), .ZN(U2951) );
  NOR2_X1 U7570 ( .A1(n6522), .A2(n6978), .ZN(n6569) );
  AOI21_X1 U7571 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6569), 
        .ZN(n6520) );
  INV_X1 U7572 ( .A(n6512), .ZN(n6514) );
  NAND3_X1 U7573 ( .A1(n6515), .A2(n6514), .A3(n6513), .ZN(n6516) );
  AND2_X1 U7574 ( .A1(n3114), .A2(n6516), .ZN(n6572) );
  AOI22_X1 U7575 ( .A1(n6572), .A2(n6535), .B1(n6536), .B2(n6518), .ZN(n6519)
         );
  OAI211_X1 U7576 ( .C1(n6541), .C2(n6521), .A(n6520), .B(n6519), .ZN(U2980)
         );
  NOR2_X1 U7577 ( .A1(n6522), .A2(n4670), .ZN(n6580) );
  AOI21_X1 U7578 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6580), 
        .ZN(n6528) );
  OAI21_X1 U7579 ( .B1(n6523), .B2(n6524), .A(n4984), .ZN(n6525) );
  INV_X1 U7580 ( .A(n6525), .ZN(n6582) );
  AOI22_X1 U7581 ( .A1(n6582), .A2(n6535), .B1(n6536), .B2(n6526), .ZN(n6527)
         );
  OAI211_X1 U7582 ( .C1(n6541), .C2(n6529), .A(n6528), .B(n6527), .ZN(U2982)
         );
  NAND2_X1 U7583 ( .A1(n6586), .A2(REIP_REG_2__SCAN_IN), .ZN(n6607) );
  INV_X1 U7584 ( .A(n6607), .ZN(n6530) );
  AOI21_X1 U7585 ( .B1(n6531), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6530), 
        .ZN(n6539) );
  XNOR2_X1 U7586 ( .A(n6533), .B(n6604), .ZN(n6534) );
  XNOR2_X1 U7587 ( .A(n3104), .B(n6534), .ZN(n6601) );
  AOI22_X1 U7588 ( .A1(n6537), .A2(n6536), .B1(n6535), .B2(n6601), .ZN(n6538)
         );
  OAI211_X1 U7589 ( .C1(n6541), .C2(n6540), .A(n6539), .B(n6538), .ZN(U2984)
         );
  AOI22_X1 U7590 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5700), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n4373), .ZN(n6548) );
  AOI21_X1 U7591 ( .B1(n6543), .B2(n6597), .A(n6542), .ZN(n6547) );
  AOI22_X1 U7592 ( .A1(n6545), .A2(n6602), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6544), .ZN(n6546) );
  OAI211_X1 U7593 ( .C1(n6549), .C2(n6548), .A(n6547), .B(n6546), .ZN(U3008)
         );
  INV_X1 U7594 ( .A(n6550), .ZN(n6551) );
  AOI21_X1 U7595 ( .B1(n6552), .B2(n6597), .A(n6551), .ZN(n6558) );
  INV_X1 U7596 ( .A(n6553), .ZN(n6556) );
  AOI21_X1 U7597 ( .B1(n7012), .B2(n6559), .A(n6554), .ZN(n6555) );
  AOI22_X1 U7598 ( .A1(n6556), .A2(n6602), .B1(n6564), .B2(n6555), .ZN(n6557)
         );
  OAI211_X1 U7599 ( .C1(n6559), .C2(n6568), .A(n6558), .B(n6557), .ZN(U3010)
         );
  INV_X1 U7600 ( .A(n6560), .ZN(n6561) );
  AOI21_X1 U7601 ( .B1(n6562), .B2(n6597), .A(n6561), .ZN(n6567) );
  INV_X1 U7602 ( .A(n6563), .ZN(n6565) );
  AOI22_X1 U7603 ( .A1(n6565), .A2(n6602), .B1(n6564), .B2(n7012), .ZN(n6566)
         );
  OAI211_X1 U7604 ( .C1(n7012), .C2(n6568), .A(n6567), .B(n6566), .ZN(U3011)
         );
  AOI21_X1 U7605 ( .B1(n6597), .B2(n6570), .A(n6569), .ZN(n6578) );
  AOI22_X1 U7606 ( .A1(n6572), .A2(n6602), .B1(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .B2(n6571), .ZN(n6577) );
  NAND3_X1 U7607 ( .A1(n6575), .A2(n6574), .A3(n6573), .ZN(n6576) );
  NAND3_X1 U7608 ( .A1(n6578), .A2(n6577), .A3(n6576), .ZN(U3012) );
  OAI21_X1 U7609 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6579), .ZN(n6585) );
  AOI21_X1 U7610 ( .B1(n6597), .B2(n6581), .A(n6580), .ZN(n6584) );
  AOI22_X1 U7611 ( .A1(n6582), .A2(n6602), .B1(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .B2(n6590), .ZN(n6583) );
  OAI211_X1 U7612 ( .C1(n6593), .C2(n6585), .A(n6584), .B(n6583), .ZN(U3014)
         );
  AOI22_X1 U7613 ( .A1(n6597), .A2(n6587), .B1(n6586), .B2(REIP_REG_3__SCAN_IN), .ZN(n6592) );
  INV_X1 U7614 ( .A(n6588), .ZN(n6589) );
  AOI22_X1 U7615 ( .A1(n6590), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6589), 
        .B2(n6602), .ZN(n6591) );
  OAI211_X1 U7616 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6593), .A(n6592), 
        .B(n6591), .ZN(U3015) );
  INV_X1 U7617 ( .A(n6594), .ZN(n6595) );
  AOI21_X1 U7618 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(n6609) );
  OAI21_X1 U7619 ( .B1(n6600), .B2(n6599), .A(n6598), .ZN(n6603) );
  AOI22_X1 U7620 ( .A1(n6603), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6602), 
        .B2(n6601), .ZN(n6608) );
  NAND3_X1 U7621 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6605), .A3(n6604), 
        .ZN(n6606) );
  NAND4_X1 U7622 ( .A1(n6609), .A2(n6608), .A3(n6607), .A4(n6606), .ZN(U3016)
         );
  INV_X1 U7623 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U7624 ( .A1(n6610), .A2(n6812), .ZN(U3019) );
  AOI22_X1 U7625 ( .A1(n6624), .A2(n6612), .B1(n6611), .B2(n6623), .ZN(n6614)
         );
  AOI22_X1 U7626 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6626), .B1(n6711), 
        .B2(n6625), .ZN(n6613) );
  OAI211_X1 U7627 ( .C1(n6629), .C2(n6714), .A(n6614), .B(n6613), .ZN(U3045)
         );
  AOI22_X1 U7628 ( .A1(n6624), .A2(n6652), .B1(n6650), .B2(n6623), .ZN(n6616)
         );
  AOI22_X1 U7629 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6626), .B1(n6718), 
        .B2(n6625), .ZN(n6615) );
  OAI211_X1 U7630 ( .C1(n6629), .C2(n6721), .A(n6616), .B(n6615), .ZN(U3046)
         );
  AOI22_X1 U7631 ( .A1(n6624), .A2(n6658), .B1(n6656), .B2(n6623), .ZN(n6618)
         );
  AOI22_X1 U7632 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6626), .B1(n6725), 
        .B2(n6625), .ZN(n6617) );
  OAI211_X1 U7633 ( .C1(n6629), .C2(n6728), .A(n6618), .B(n6617), .ZN(U3047)
         );
  AOI22_X1 U7634 ( .A1(n6624), .A2(n6756), .B1(n6754), .B2(n6623), .ZN(n6620)
         );
  AOI22_X1 U7635 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6626), .B1(n6755), 
        .B2(n6625), .ZN(n6619) );
  OAI211_X1 U7636 ( .C1(n6629), .C2(n6759), .A(n6620), .B(n6619), .ZN(U3048)
         );
  AOI22_X1 U7637 ( .A1(n6624), .A2(n6768), .B1(n6766), .B2(n6623), .ZN(n6622)
         );
  AOI22_X1 U7638 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6626), .B1(n6767), 
        .B2(n6625), .ZN(n6621) );
  OAI211_X1 U7639 ( .C1(n6629), .C2(n6771), .A(n6622), .B(n6621), .ZN(U3050)
         );
  AOI22_X1 U7640 ( .A1(n6624), .A2(n6777), .B1(n6772), .B2(n6623), .ZN(n6628)
         );
  AOI22_X1 U7641 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6626), .B1(n6774), 
        .B2(n6625), .ZN(n6627) );
  OAI211_X1 U7642 ( .C1(n6629), .C2(n6782), .A(n6628), .B(n6627), .ZN(U3051)
         );
  INV_X1 U7643 ( .A(n6630), .ZN(n6631) );
  AOI21_X1 U7644 ( .B1(n6631), .B2(n6695), .A(n6666), .ZN(n6637) );
  NOR2_X1 U7645 ( .A1(n6637), .A2(n6698), .ZN(n6632) );
  AOI21_X1 U7646 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6640), .A(n6632), .ZN(
        n6686) );
  AOI22_X1 U7647 ( .A1(n6680), .A2(n6634), .B1(n6666), .B2(n6633), .ZN(n6643)
         );
  NAND2_X1 U7648 ( .A1(n6636), .A2(n6635), .ZN(n6807) );
  NAND3_X1 U7649 ( .A1(n6807), .A2(n6691), .A3(n6637), .ZN(n6639) );
  OAI211_X1 U7650 ( .C1(n6640), .C2(n6691), .A(n6639), .B(n6638), .ZN(n6682)
         );
  AOI22_X1 U7651 ( .A1(n6682), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n6641), 
        .B2(n6668), .ZN(n6642) );
  OAI211_X1 U7652 ( .C1(n6686), .C2(n6644), .A(n6643), .B(n6642), .ZN(U3076)
         );
  OAI22_X1 U7653 ( .A1(n6678), .A2(n6709), .B1(n6677), .B2(n6708), .ZN(n6645)
         );
  INV_X1 U7654 ( .A(n6645), .ZN(n6648) );
  AOI22_X1 U7655 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6682), .B1(n6646), 
        .B2(n6680), .ZN(n6647) );
  OAI211_X1 U7656 ( .C1(n6686), .C2(n6649), .A(n6648), .B(n6647), .ZN(U3077)
         );
  AOI22_X1 U7657 ( .A1(n6680), .A2(n6651), .B1(n6666), .B2(n6650), .ZN(n6654)
         );
  AOI22_X1 U7658 ( .A1(n6682), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6652), 
        .B2(n6668), .ZN(n6653) );
  OAI211_X1 U7659 ( .C1(n6686), .C2(n6655), .A(n6654), .B(n6653), .ZN(U3078)
         );
  AOI22_X1 U7660 ( .A1(n6680), .A2(n6657), .B1(n6666), .B2(n6656), .ZN(n6660)
         );
  AOI22_X1 U7661 ( .A1(n6682), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n6658), 
        .B2(n6668), .ZN(n6659) );
  OAI211_X1 U7662 ( .C1(n6686), .C2(n6661), .A(n6660), .B(n6659), .ZN(U3079)
         );
  AOI22_X1 U7663 ( .A1(n6680), .A2(n6662), .B1(n6666), .B2(n6754), .ZN(n6664)
         );
  AOI22_X1 U7664 ( .A1(n6682), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6756), 
        .B2(n6668), .ZN(n6663) );
  OAI211_X1 U7665 ( .C1(n6686), .C2(n6665), .A(n6664), .B(n6663), .ZN(U3080)
         );
  AOI22_X1 U7666 ( .A1(n6680), .A2(n6667), .B1(n6666), .B2(n6760), .ZN(n6670)
         );
  AOI22_X1 U7667 ( .A1(n6682), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6762), 
        .B2(n6668), .ZN(n6669) );
  OAI211_X1 U7668 ( .C1(n6686), .C2(n6671), .A(n6670), .B(n6669), .ZN(U3081)
         );
  OAI22_X1 U7669 ( .A1(n6678), .A2(n6740), .B1(n6677), .B2(n6739), .ZN(n6672)
         );
  INV_X1 U7670 ( .A(n6672), .ZN(n6675) );
  AOI22_X1 U7671 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6682), .B1(n6673), 
        .B2(n6680), .ZN(n6674) );
  OAI211_X1 U7672 ( .C1(n6686), .C2(n6676), .A(n6675), .B(n6674), .ZN(U3082)
         );
  OAI22_X1 U7673 ( .A1(n6678), .A2(n6752), .B1(n6677), .B2(n6745), .ZN(n6679)
         );
  INV_X1 U7674 ( .A(n6679), .ZN(n6684) );
  AOI22_X1 U7675 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6682), .B1(n6681), 
        .B2(n6680), .ZN(n6683) );
  OAI211_X1 U7676 ( .C1(n6686), .C2(n6685), .A(n6684), .B(n6683), .ZN(U3083)
         );
  NOR2_X1 U7677 ( .A1(n6687), .A2(n6982), .ZN(n6694) );
  INV_X1 U7678 ( .A(n6694), .ZN(n6744) );
  OAI22_X1 U7679 ( .A1(n6746), .A2(n6689), .B1(n6688), .B2(n6744), .ZN(n6690)
         );
  INV_X1 U7680 ( .A(n6690), .ZN(n6706) );
  OAI21_X1 U7681 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6703) );
  AOI21_X1 U7682 ( .B1(n6696), .B2(n6695), .A(n6694), .ZN(n6702) );
  INV_X1 U7683 ( .A(n6702), .ZN(n6700) );
  AOI21_X1 U7684 ( .B1(n6698), .B2(n6701), .A(n6697), .ZN(n6699) );
  OAI22_X1 U7685 ( .A1(n6703), .A2(n6702), .B1(n6701), .B2(n6956), .ZN(n6748)
         );
  AOI22_X1 U7686 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6749), .B1(n6704), 
        .B2(n6748), .ZN(n6705) );
  OAI211_X1 U7687 ( .C1(n6707), .C2(n6781), .A(n6706), .B(n6705), .ZN(U3108)
         );
  OAI22_X1 U7688 ( .A1(n6781), .A2(n6709), .B1(n6708), .B2(n6744), .ZN(n6710)
         );
  INV_X1 U7689 ( .A(n6710), .ZN(n6713) );
  AOI22_X1 U7690 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6749), .B1(n6711), 
        .B2(n6748), .ZN(n6712) );
  OAI211_X1 U7691 ( .C1(n6714), .C2(n6746), .A(n6713), .B(n6712), .ZN(U3109)
         );
  OAI22_X1 U7692 ( .A1(n6781), .A2(n6716), .B1(n6715), .B2(n6744), .ZN(n6717)
         );
  INV_X1 U7693 ( .A(n6717), .ZN(n6720) );
  AOI22_X1 U7694 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6749), .B1(n6718), 
        .B2(n6748), .ZN(n6719) );
  OAI211_X1 U7695 ( .C1(n6721), .C2(n6746), .A(n6720), .B(n6719), .ZN(U3110)
         );
  OAI22_X1 U7696 ( .A1(n6781), .A2(n6723), .B1(n6722), .B2(n6744), .ZN(n6724)
         );
  INV_X1 U7697 ( .A(n6724), .ZN(n6727) );
  AOI22_X1 U7698 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6749), .B1(n6725), 
        .B2(n6748), .ZN(n6726) );
  OAI211_X1 U7699 ( .C1(n6728), .C2(n6746), .A(n6727), .B(n6726), .ZN(U3111)
         );
  OAI22_X1 U7700 ( .A1(n6746), .A2(n6759), .B1(n6729), .B2(n6744), .ZN(n6730)
         );
  INV_X1 U7701 ( .A(n6730), .ZN(n6732) );
  AOI22_X1 U7702 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6749), .B1(n6755), 
        .B2(n6748), .ZN(n6731) );
  OAI211_X1 U7703 ( .C1(n6733), .C2(n6781), .A(n6732), .B(n6731), .ZN(U3112)
         );
  OAI22_X1 U7704 ( .A1(n6781), .A2(n6735), .B1(n6734), .B2(n6744), .ZN(n6736)
         );
  INV_X1 U7705 ( .A(n6736), .ZN(n6738) );
  AOI22_X1 U7706 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6749), .B1(n6761), 
        .B2(n6748), .ZN(n6737) );
  OAI211_X1 U7707 ( .C1(n6765), .C2(n6746), .A(n6738), .B(n6737), .ZN(U3113)
         );
  OAI22_X1 U7708 ( .A1(n6781), .A2(n6740), .B1(n6739), .B2(n6744), .ZN(n6741)
         );
  INV_X1 U7709 ( .A(n6741), .ZN(n6743) );
  AOI22_X1 U7710 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6749), .B1(n6767), 
        .B2(n6748), .ZN(n6742) );
  OAI211_X1 U7711 ( .C1(n6771), .C2(n6746), .A(n6743), .B(n6742), .ZN(U3114)
         );
  OAI22_X1 U7712 ( .A1(n6746), .A2(n6782), .B1(n6745), .B2(n6744), .ZN(n6747)
         );
  INV_X1 U7713 ( .A(n6747), .ZN(n6751) );
  AOI22_X1 U7714 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6749), .B1(n6774), 
        .B2(n6748), .ZN(n6750) );
  OAI211_X1 U7715 ( .C1(n6752), .C2(n6781), .A(n6751), .B(n6750), .ZN(U3115)
         );
  INV_X1 U7716 ( .A(n6753), .ZN(n6775) );
  AOI22_X1 U7717 ( .A1(n6775), .A2(n6755), .B1(n6773), .B2(n6754), .ZN(n6758)
         );
  AOI22_X1 U7718 ( .A1(n6778), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6756), 
        .B2(n6776), .ZN(n6757) );
  OAI211_X1 U7719 ( .C1(n6759), .C2(n6781), .A(n6758), .B(n6757), .ZN(U3120)
         );
  AOI22_X1 U7720 ( .A1(n6775), .A2(n6761), .B1(n6773), .B2(n6760), .ZN(n6764)
         );
  AOI22_X1 U7721 ( .A1(n6778), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6762), 
        .B2(n6776), .ZN(n6763) );
  OAI211_X1 U7722 ( .C1(n6765), .C2(n6781), .A(n6764), .B(n6763), .ZN(U3121)
         );
  AOI22_X1 U7723 ( .A1(n6775), .A2(n6767), .B1(n6773), .B2(n6766), .ZN(n6770)
         );
  AOI22_X1 U7724 ( .A1(n6778), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6768), 
        .B2(n6776), .ZN(n6769) );
  OAI211_X1 U7725 ( .C1(n6771), .C2(n6781), .A(n6770), .B(n6769), .ZN(U3122)
         );
  AOI22_X1 U7726 ( .A1(n6775), .A2(n6774), .B1(n6773), .B2(n6772), .ZN(n6780)
         );
  AOI22_X1 U7727 ( .A1(n6778), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6777), 
        .B2(n6776), .ZN(n6779) );
  OAI211_X1 U7728 ( .C1(n6782), .C2(n6781), .A(n6780), .B(n6779), .ZN(U3123)
         );
  OR2_X1 U7729 ( .A1(n6795), .A2(n6804), .ZN(n6786) );
  INV_X1 U7730 ( .A(n6791), .ZN(n6785) );
  NAND3_X1 U7731 ( .A1(n6792), .A2(n6791), .A3(n6790), .ZN(n6794) );
  OAI21_X1 U7732 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(U3150) );
  INV_X1 U7733 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U7734 ( .A1(n6801), .A2(n6926), .ZN(U3151) );
  AND2_X1 U7735 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6796), .ZN(U3152) );
  INV_X1 U7736 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6919) );
  NOR2_X1 U7737 ( .A1(n6801), .A2(n6919), .ZN(U3153) );
  AND2_X1 U7738 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6796), .ZN(U3154) );
  INV_X1 U7739 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U7740 ( .A1(n6801), .A2(n7029), .ZN(U3155) );
  AND2_X1 U7741 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6796), .ZN(U3156) );
  AND2_X1 U7742 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6796), .ZN(U3157) );
  AND2_X1 U7743 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6796), .ZN(U3158) );
  AND2_X1 U7744 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6796), .ZN(U3159) );
  AND2_X1 U7745 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6796), .ZN(U3160) );
  AND2_X1 U7746 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6796), .ZN(U3161) );
  INV_X1 U7747 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6916) );
  NOR2_X1 U7748 ( .A1(n6801), .A2(n6916), .ZN(U3162) );
  AND2_X1 U7749 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6796), .ZN(U3163) );
  AND2_X1 U7750 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6796), .ZN(U3164) );
  AND2_X1 U7751 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6796), .ZN(U3165) );
  INV_X1 U7752 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6970) );
  NOR2_X1 U7753 ( .A1(n6801), .A2(n6970), .ZN(U3166) );
  AND2_X1 U7754 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6796), .ZN(U3167) );
  AND2_X1 U7755 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6796), .ZN(U3168) );
  INV_X1 U7756 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7106) );
  NOR2_X1 U7757 ( .A1(n6801), .A2(n7106), .ZN(U3169) );
  AND2_X1 U7758 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6796), .ZN(U3170) );
  AND2_X1 U7759 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6796), .ZN(U3171) );
  AND2_X1 U7760 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6796), .ZN(U3172) );
  AND2_X1 U7761 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6796), .ZN(U3173) );
  AND2_X1 U7762 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6796), .ZN(U3174) );
  AND2_X1 U7763 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6796), .ZN(U3175) );
  AND2_X1 U7764 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6796), .ZN(U3176) );
  AND2_X1 U7765 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6796), .ZN(U3177) );
  AND2_X1 U7766 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6796), .ZN(U3178) );
  AND2_X1 U7767 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6796), .ZN(U3179) );
  AND2_X1 U7768 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6796), .ZN(U3180) );
  MUX2_X1 U7769 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6824), .Z(U3445) );
  INV_X1 U7770 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6816) );
  INV_X1 U7771 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6879) );
  AOI22_X1 U7772 ( .A1(n6797), .A2(n6816), .B1(n6879), .B2(n6824), .ZN(U3446)
         );
  MUX2_X1 U7773 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6824), .Z(U3447) );
  INV_X1 U7774 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6822) );
  INV_X1 U7775 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U7776 ( .A1(n6797), .A2(n6822), .B1(n6917), .B2(n6824), .ZN(U3448)
         );
  OAI21_X1 U7777 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6801), .A(n6799), .ZN(
        n6798) );
  INV_X1 U7778 ( .A(n6798), .ZN(U3451) );
  OAI21_X1 U7779 ( .B1(n6801), .B2(n6800), .A(n6799), .ZN(U3452) );
  AOI211_X1 U7780 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6804), .A(n6803), .B(
        n6802), .ZN(n6805) );
  INV_X1 U7781 ( .A(n6805), .ZN(U3453) );
  INV_X1 U7782 ( .A(n6806), .ZN(n6808) );
  NAND2_X1 U7783 ( .A1(n6808), .A2(n6807), .ZN(n6811) );
  AOI222_X1 U7784 ( .A1(n6811), .A2(n6691), .B1(n4889), .B2(n6810), .C1(n3115), 
        .C2(n6809), .ZN(n6813) );
  AOI22_X1 U7785 ( .A1(n6814), .A2(n6982), .B1(n6813), .B2(n6812), .ZN(U3462)
         );
  AOI21_X1 U7786 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7787 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6815), .B2(n6888), .ZN(n6817) );
  AOI22_X1 U7788 ( .A1(n6818), .A2(n6817), .B1(n6816), .B2(n6821), .ZN(U3468)
         );
  NOR2_X1 U7789 ( .A1(n6821), .A2(REIP_REG_1__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7790 ( .A1(n6822), .A2(n6821), .B1(n6820), .B2(n6819), .ZN(U3469)
         );
  NAND2_X1 U7791 ( .A1(n6824), .A2(W_R_N_REG_SCAN_IN), .ZN(n6823) );
  OAI21_X1 U7792 ( .B1(n6824), .B2(READREQUEST_REG_SCAN_IN), .A(n6823), .ZN(
        U3470) );
  MUX2_X1 U7793 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6824), .Z(U3473) );
  NAND2_X1 U7794 ( .A1(n6825), .A2(LWORD_REG_2__SCAN_IN), .ZN(n6827) );
  OAI211_X1 U7795 ( .C1(n3668), .C2(n6828), .A(n6827), .B(n6826), .ZN(n7129)
         );
  OR4_X1 U7796 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(
        INSTQUEUE_REG_12__0__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6839) );
  NOR4_X1 U7797 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n7025), .A4(n6907), .ZN(n6832)
         );
  INV_X1 U7798 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n7048) );
  NOR4_X1 U7799 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        INSTQUEUE_REG_9__0__SCAN_IN), .A3(INSTQUEUE_REG_6__1__SCAN_IN), .A4(
        n7048), .ZN(n6831) );
  INV_X1 U7800 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6954) );
  INV_X1 U7801 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n7113) );
  NOR4_X1 U7802 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(
        INSTQUEUE_REG_0__4__SCAN_IN), .A3(n6954), .A4(n7113), .ZN(n6830) );
  INV_X1 U7803 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n7005) );
  NOR4_X1 U7804 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(
        INSTQUEUE_REG_3__4__SCAN_IN), .A3(INSTQUEUE_REG_7__4__SCAN_IN), .A4(
        n7005), .ZN(n6829) );
  NAND4_X1 U7805 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6838)
         );
  INV_X1 U7806 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6834) );
  INV_X1 U7807 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6833) );
  NOR4_X1 U7808 ( .A1(n6834), .A2(n6833), .A3(INSTQUEUE_REG_6__7__SCAN_IN), 
        .A4(STATE_REG_2__SCAN_IN), .ZN(n6835) );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n7044) );
  NAND4_X1 U7810 ( .A1(n6835), .A2(n6983), .A3(REQUESTPENDING_REG_SCAN_IN), 
        .A4(n7044), .ZN(n6837) );
  INV_X1 U7811 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6968) );
  NAND4_X1 U7812 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(
        INSTQUEUE_REG_2__6__SCAN_IN), .A3(INSTQUEUE_REG_1__6__SCAN_IN), .A4(
        n6968), .ZN(n6836) );
  NOR4_X1 U7813 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6873)
         );
  NOR4_X1 U7814 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(EAX_REG_17__SCAN_IN), 
        .A3(ADDRESS_REG_27__SCAN_IN), .A4(n7105), .ZN(n6840) );
  NAND3_X1 U7815 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(n6840), .ZN(n6850) );
  NAND4_X1 U7816 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(DATAI_30_), .A3(
        DATAO_REG_16__SCAN_IN), .A4(ADDRESS_REG_2__SCAN_IN), .ZN(n6841) );
  NOR3_X1 U7817 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n7066), .A3(n6841), .ZN(n6848) );
  INV_X1 U7818 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n7016) );
  NAND4_X1 U7819 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(
        INSTQUEUE_REG_9__2__SCAN_IN), .A3(INSTQUEUE_REG_1__2__SCAN_IN), .A4(
        n7016), .ZN(n6846) );
  NAND4_X1 U7820 ( .A1(EBX_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A3(REIP_REG_28__SCAN_IN), .A4(n5127), 
        .ZN(n6845) );
  NAND4_X1 U7821 ( .A1(ADDRESS_REG_8__SCAN_IN), .A2(D_C_N_REG_SCAN_IN), .A3(
        ADDRESS_REG_24__SCAN_IN), .A4(LWORD_REG_13__SCAN_IN), .ZN(n6844) );
  INV_X1 U7822 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6842) );
  INV_X1 U7823 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6896) );
  NAND4_X1 U7824 ( .A1(n6842), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .A3(
        INSTQUEUE_REG_13__3__SCAN_IN), .A4(n6896), .ZN(n6843) );
  NOR4_X1 U7825 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6847)
         );
  NAND4_X1 U7826 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6848), .A3(n6847), 
        .A4(n7060), .ZN(n6849) );
  NOR4_X1 U7827 ( .A1(EBX_REG_24__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        n6850), .A4(n6849), .ZN(n6872) );
  NAND4_X1 U7828 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(DATAO_REG_8__SCAN_IN), 
        .A3(n7031), .A4(n7028), .ZN(n6851) );
  NOR3_X1 U7829 ( .A1(DATAI_15_), .A2(BE_N_REG_2__SCAN_IN), .A3(n6851), .ZN(
        n6852) );
  NAND3_X1 U7830 ( .A1(n6852), .A2(n4344), .A3(n7041), .ZN(n6860) );
  NAND4_X1 U7831 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n5700), .A3(n6910), .A4(
        n6909), .ZN(n6859) );
  NAND4_X1 U7832 ( .A1(EBX_REG_6__SCAN_IN), .A2(DATAI_8_), .A3(
        LWORD_REG_5__SCAN_IN), .A4(ADDRESS_REG_15__SCAN_IN), .ZN(n6858) );
  NOR4_X1 U7833 ( .A1(STATEBS16_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .A3(
        UWORD_REG_10__SCAN_IN), .A4(n7002), .ZN(n6856) );
  NOR4_X1 U7834 ( .A1(DATAI_26_), .A2(DATAO_REG_12__SCAN_IN), .A3(n7015), .A4(
        n6995), .ZN(n6855) );
  NOR4_X1 U7835 ( .A1(DATAO_REG_1__SCAN_IN), .A2(ADDRESS_REG_25__SCAN_IN), 
        .A3(ADDRESS_REG_29__SCAN_IN), .A4(n6893), .ZN(n6854) );
  NOR4_X1 U7836 ( .A1(n6882), .A2(n6890), .A3(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .A4(REIP_REG_1__SCAN_IN), .ZN(n6853) );
  NAND4_X1 U7837 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6857)
         );
  NOR4_X1 U7838 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n6871)
         );
  NAND4_X1 U7839 ( .A1(n6502), .A2(UWORD_REG_14__SCAN_IN), .A3(
        DATAO_REG_25__SCAN_IN), .A4(n6978), .ZN(n6869) );
  NAND4_X1 U7840 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(DATAO_REG_26__SCAN_IN), 
        .A3(ADDRESS_REG_21__SCAN_IN), .A4(n6917), .ZN(n6861) );
  NOR3_X1 U7841 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6920), .A3(n6861), .ZN(
        n6867) );
  NAND4_X1 U7842 ( .A1(DATAI_19_), .A2(REIP_REG_17__SCAN_IN), .A3(
        DATAWIDTH_REG_0__SCAN_IN), .A4(n6957), .ZN(n6865) );
  NAND4_X1 U7843 ( .A1(UWORD_REG_0__SCAN_IN), .A2(ADDRESS_REG_6__SCAN_IN), 
        .A3(n6942), .A4(n6944), .ZN(n6864) );
  NAND4_X1 U7844 ( .A1(EAX_REG_24__SCAN_IN), .A2(EAX_REG_9__SCAN_IN), .A3(
        UWORD_REG_11__SCAN_IN), .A4(n4658), .ZN(n6863) );
  NAND4_X1 U7845 ( .A1(REIP_REG_15__SCAN_IN), .A2(DATAO_REG_9__SCAN_IN), .A3(
        DATAWIDTH_REG_16__SCAN_IN), .A4(n6965), .ZN(n6862) );
  NOR4_X1 U7846 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6866)
         );
  NAND4_X1 U7847 ( .A1(EBX_REG_30__SCAN_IN), .A2(EBX_REG_10__SCAN_IN), .A3(
        n6867), .A4(n6866), .ZN(n6868) );
  NOR4_X1 U7848 ( .A1(STATE_REG_1__SCAN_IN), .A2(EBX_REG_8__SCAN_IN), .A3(
        n6869), .A4(n6868), .ZN(n6870) );
  NAND4_X1 U7849 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n7126)
         );
  AOI22_X1 U7850 ( .A1(n4748), .A2(keyinput60), .B1(n6875), .B2(keyinput96), 
        .ZN(n6874) );
  OAI221_X1 U7851 ( .B1(n4748), .B2(keyinput60), .C1(n6875), .C2(keyinput96), 
        .A(n6874), .ZN(n6886) );
  INV_X1 U7852 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6877) );
  AOI22_X1 U7853 ( .A1(n5539), .A2(keyinput42), .B1(n6877), .B2(keyinput83), 
        .ZN(n6876) );
  OAI221_X1 U7854 ( .B1(n5539), .B2(keyinput42), .C1(n6877), .C2(keyinput83), 
        .A(n6876), .ZN(n6885) );
  AOI22_X1 U7855 ( .A1(n6879), .A2(keyinput110), .B1(n3278), .B2(keyinput78), 
        .ZN(n6878) );
  OAI221_X1 U7856 ( .B1(n6879), .B2(keyinput110), .C1(n3278), .C2(keyinput78), 
        .A(n6878), .ZN(n6884) );
  AOI22_X1 U7857 ( .A1(n6882), .A2(keyinput75), .B1(keyinput98), .B2(n6881), 
        .ZN(n6880) );
  OAI221_X1 U7858 ( .B1(n6882), .B2(keyinput75), .C1(n6881), .C2(keyinput98), 
        .A(n6880), .ZN(n6883) );
  NOR4_X1 U7859 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n6934)
         );
  AOI22_X1 U7860 ( .A1(n4750), .A2(keyinput41), .B1(n6888), .B2(keyinput70), 
        .ZN(n6887) );
  OAI221_X1 U7861 ( .B1(n4750), .B2(keyinput41), .C1(n6888), .C2(keyinput70), 
        .A(n6887), .ZN(n6900) );
  AOI22_X1 U7862 ( .A1(n6891), .A2(keyinput113), .B1(keyinput65), .B2(n6890), 
        .ZN(n6889) );
  OAI221_X1 U7863 ( .B1(n6891), .B2(keyinput113), .C1(n6890), .C2(keyinput65), 
        .A(n6889), .ZN(n6899) );
  AOI22_X1 U7864 ( .A1(n6894), .A2(keyinput79), .B1(n6893), .B2(keyinput7), 
        .ZN(n6892) );
  OAI221_X1 U7865 ( .B1(n6894), .B2(keyinput79), .C1(n6893), .C2(keyinput7), 
        .A(n6892), .ZN(n6898) );
  AOI22_X1 U7866 ( .A1(n4781), .A2(keyinput88), .B1(n6896), .B2(keyinput16), 
        .ZN(n6895) );
  OAI221_X1 U7867 ( .B1(n4781), .B2(keyinput88), .C1(n6896), .C2(keyinput16), 
        .A(n6895), .ZN(n6897) );
  NOR4_X1 U7868 ( .A1(n6900), .A2(n6899), .A3(n6898), .A4(n6897), .ZN(n6933)
         );
  AOI22_X1 U7869 ( .A1(n4671), .A2(keyinput86), .B1(n6902), .B2(keyinput109), 
        .ZN(n6901) );
  OAI221_X1 U7870 ( .B1(n4671), .B2(keyinput86), .C1(n6902), .C2(keyinput109), 
        .A(n6901), .ZN(n6914) );
  AOI22_X1 U7871 ( .A1(n6905), .A2(keyinput49), .B1(keyinput85), .B2(n6904), 
        .ZN(n6903) );
  OAI221_X1 U7872 ( .B1(n6905), .B2(keyinput49), .C1(n6904), .C2(keyinput85), 
        .A(n6903), .ZN(n6913) );
  AOI22_X1 U7873 ( .A1(n5700), .A2(keyinput100), .B1(n6907), .B2(keyinput55), 
        .ZN(n6906) );
  OAI221_X1 U7874 ( .B1(n5700), .B2(keyinput100), .C1(n6907), .C2(keyinput55), 
        .A(n6906), .ZN(n6912) );
  AOI22_X1 U7875 ( .A1(n6910), .A2(keyinput111), .B1(keyinput119), .B2(n6909), 
        .ZN(n6908) );
  OAI221_X1 U7876 ( .B1(n6910), .B2(keyinput111), .C1(n6909), .C2(keyinput119), 
        .A(n6908), .ZN(n6911) );
  NOR4_X1 U7877 ( .A1(n6914), .A2(n6913), .A3(n6912), .A4(n6911), .ZN(n6932)
         );
  AOI22_X1 U7878 ( .A1(n6917), .A2(keyinput120), .B1(keyinput9), .B2(n6916), 
        .ZN(n6915) );
  OAI221_X1 U7879 ( .B1(n6917), .B2(keyinput120), .C1(n6916), .C2(keyinput9), 
        .A(n6915), .ZN(n6930) );
  AOI22_X1 U7880 ( .A1(n6920), .A2(keyinput17), .B1(keyinput69), .B2(n6919), 
        .ZN(n6918) );
  OAI221_X1 U7881 ( .B1(n6920), .B2(keyinput17), .C1(n6919), .C2(keyinput69), 
        .A(n6918), .ZN(n6929) );
  AOI22_X1 U7882 ( .A1(n6923), .A2(keyinput114), .B1(keyinput102), .B2(n6922), 
        .ZN(n6921) );
  OAI221_X1 U7883 ( .B1(n6923), .B2(keyinput114), .C1(n6922), .C2(keyinput102), 
        .A(n6921), .ZN(n6928) );
  AOI22_X1 U7884 ( .A1(n6926), .A2(keyinput11), .B1(keyinput76), .B2(n6925), 
        .ZN(n6924) );
  OAI221_X1 U7885 ( .B1(n6926), .B2(keyinput11), .C1(n6925), .C2(keyinput76), 
        .A(n6924), .ZN(n6927) );
  NOR4_X1 U7886 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n6931)
         );
  NAND4_X1 U7887 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n7124)
         );
  INV_X1 U7888 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6937) );
  INV_X1 U7889 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7890 ( .A1(n6937), .A2(keyinput12), .B1(n6936), .B2(keyinput6), 
        .ZN(n6935) );
  OAI221_X1 U7891 ( .B1(n6937), .B2(keyinput12), .C1(n6936), .C2(keyinput6), 
        .A(n6935), .ZN(n6949) );
  AOI22_X1 U7892 ( .A1(n6939), .A2(keyinput51), .B1(keyinput22), .B2(n4784), 
        .ZN(n6938) );
  OAI221_X1 U7893 ( .B1(n6939), .B2(keyinput51), .C1(n4784), .C2(keyinput22), 
        .A(n6938), .ZN(n6948) );
  INV_X1 U7894 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6941) );
  AOI22_X1 U7895 ( .A1(n6942), .A2(keyinput58), .B1(n6941), .B2(keyinput56), 
        .ZN(n6940) );
  OAI221_X1 U7896 ( .B1(n6942), .B2(keyinput58), .C1(n6941), .C2(keyinput56), 
        .A(n6940), .ZN(n6947) );
  AOI22_X1 U7897 ( .A1(n6945), .A2(keyinput33), .B1(keyinput37), .B2(n6944), 
        .ZN(n6943) );
  OAI221_X1 U7898 ( .B1(n6945), .B2(keyinput33), .C1(n6944), .C2(keyinput37), 
        .A(n6943), .ZN(n6946) );
  NOR4_X1 U7899 ( .A1(n6949), .A2(n6948), .A3(n6947), .A4(n6946), .ZN(n6993)
         );
  INV_X1 U7900 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6951) );
  AOI22_X1 U7901 ( .A1(n6951), .A2(keyinput118), .B1(keyinput13), .B2(n4940), 
        .ZN(n6950) );
  OAI221_X1 U7902 ( .B1(n6951), .B2(keyinput118), .C1(n4940), .C2(keyinput13), 
        .A(n6950), .ZN(n6963) );
  INV_X1 U7903 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6953) );
  AOI22_X1 U7904 ( .A1(n6954), .A2(keyinput63), .B1(keyinput40), .B2(n6953), 
        .ZN(n6952) );
  OAI221_X1 U7905 ( .B1(n6954), .B2(keyinput63), .C1(n6953), .C2(keyinput40), 
        .A(n6952), .ZN(n6962) );
  AOI22_X1 U7906 ( .A1(n6957), .A2(keyinput15), .B1(n6956), .B2(keyinput61), 
        .ZN(n6955) );
  OAI221_X1 U7907 ( .B1(n6957), .B2(keyinput15), .C1(n6956), .C2(keyinput61), 
        .A(n6955), .ZN(n6961) );
  XNOR2_X1 U7908 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .B(keyinput91), .ZN(n6959)
         );
  XNOR2_X1 U7909 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput26), .ZN(n6958) );
  NAND2_X1 U7910 ( .A1(n6959), .A2(n6958), .ZN(n6960) );
  NOR4_X1 U7911 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6992)
         );
  INV_X1 U7912 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6966) );
  AOI22_X1 U7913 ( .A1(n6966), .A2(keyinput32), .B1(keyinput1), .B2(n6965), 
        .ZN(n6964) );
  OAI221_X1 U7914 ( .B1(n6966), .B2(keyinput32), .C1(n6965), .C2(keyinput1), 
        .A(n6964), .ZN(n6976) );
  AOI22_X1 U7915 ( .A1(n6968), .A2(keyinput67), .B1(keyinput50), .B2(n4746), 
        .ZN(n6967) );
  OAI221_X1 U7916 ( .B1(n6968), .B2(keyinput67), .C1(n4746), .C2(keyinput50), 
        .A(n6967), .ZN(n6975) );
  AOI22_X1 U7917 ( .A1(n6971), .A2(keyinput92), .B1(keyinput94), .B2(n6970), 
        .ZN(n6969) );
  OAI221_X1 U7918 ( .B1(n6971), .B2(keyinput92), .C1(n6970), .C2(keyinput94), 
        .A(n6969), .ZN(n6974) );
  AOI22_X1 U7919 ( .A1(n4701), .A2(keyinput81), .B1(keyinput80), .B2(n4658), 
        .ZN(n6972) );
  OAI221_X1 U7920 ( .B1(n4701), .B2(keyinput81), .C1(n4658), .C2(keyinput80), 
        .A(n6972), .ZN(n6973) );
  NOR4_X1 U7921 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n6973), .ZN(n6991)
         );
  AOI22_X1 U7922 ( .A1(n6978), .A2(keyinput108), .B1(keyinput73), .B2(n4844), 
        .ZN(n6977) );
  OAI221_X1 U7923 ( .B1(n6978), .B2(keyinput108), .C1(n4844), .C2(keyinput73), 
        .A(n6977), .ZN(n6989) );
  INV_X1 U7924 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U7925 ( .A1(n6980), .A2(keyinput107), .B1(n4712), .B2(keyinput28), 
        .ZN(n6979) );
  OAI221_X1 U7926 ( .B1(n6980), .B2(keyinput107), .C1(n4712), .C2(keyinput28), 
        .A(n6979), .ZN(n6988) );
  AOI22_X1 U7927 ( .A1(n6983), .A2(keyinput101), .B1(n6982), .B2(keyinput18), 
        .ZN(n6981) );
  OAI221_X1 U7928 ( .B1(n6983), .B2(keyinput101), .C1(n6982), .C2(keyinput18), 
        .A(n6981), .ZN(n6987) );
  XOR2_X1 U7929 ( .A(n5491), .B(keyinput4), .Z(n6985) );
  XNOR2_X1 U7930 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput89), .ZN(n6984) );
  NAND2_X1 U7931 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  NOR4_X1 U7932 ( .A1(n6989), .A2(n6988), .A3(n6987), .A4(n6986), .ZN(n6990)
         );
  NAND4_X1 U7933 ( .A1(n6993), .A2(n6992), .A3(n6991), .A4(n6990), .ZN(n7123)
         );
  INV_X1 U7934 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U7935 ( .A1(n6996), .A2(keyinput59), .B1(keyinput30), .B2(n6995), 
        .ZN(n6994) );
  OAI221_X1 U7936 ( .B1(n6996), .B2(keyinput59), .C1(n6995), .C2(keyinput30), 
        .A(n6994), .ZN(n7000) );
  XNOR2_X1 U7937 ( .A(n6997), .B(keyinput5), .ZN(n6999) );
  XOR2_X1 U7938 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .B(keyinput93), .Z(n6998)
         );
  OR3_X1 U7939 ( .A1(n7000), .A2(n6999), .A3(n6998), .ZN(n7009) );
  INV_X1 U7940 ( .A(DATAI_26_), .ZN(n7003) );
  AOI22_X1 U7941 ( .A1(n7003), .A2(keyinput10), .B1(n7002), .B2(keyinput0), 
        .ZN(n7001) );
  OAI221_X1 U7942 ( .B1(n7003), .B2(keyinput10), .C1(n7002), .C2(keyinput0), 
        .A(n7001), .ZN(n7008) );
  INV_X1 U7943 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n7006) );
  AOI22_X1 U7944 ( .A1(n7006), .A2(keyinput125), .B1(n7005), .B2(keyinput47), 
        .ZN(n7004) );
  OAI221_X1 U7945 ( .B1(n7006), .B2(keyinput125), .C1(n7005), .C2(keyinput47), 
        .A(n7004), .ZN(n7007) );
  NOR3_X1 U7946 ( .A1(n7009), .A2(n7008), .A3(n7007), .ZN(n7058) );
  AOI22_X1 U7947 ( .A1(n5286), .A2(keyinput52), .B1(keyinput106), .B2(n5127), 
        .ZN(n7010) );
  OAI221_X1 U7948 ( .B1(n5286), .B2(keyinput52), .C1(n5127), .C2(keyinput106), 
        .A(n7010), .ZN(n7023) );
  AOI22_X1 U7949 ( .A1(n7013), .A2(keyinput35), .B1(n7012), .B2(keyinput72), 
        .ZN(n7011) );
  OAI221_X1 U7950 ( .B1(n7013), .B2(keyinput35), .C1(n7012), .C2(keyinput72), 
        .A(n7011), .ZN(n7022) );
  AOI22_X1 U7951 ( .A1(n7016), .A2(keyinput90), .B1(keyinput36), .B2(n7015), 
        .ZN(n7014) );
  OAI221_X1 U7952 ( .B1(n7016), .B2(keyinput90), .C1(n7015), .C2(keyinput36), 
        .A(n7014), .ZN(n7021) );
  AOI22_X1 U7953 ( .A1(n7019), .A2(keyinput84), .B1(n7018), .B2(keyinput122), 
        .ZN(n7017) );
  OAI221_X1 U7954 ( .B1(n7019), .B2(keyinput84), .C1(n7018), .C2(keyinput122), 
        .A(n7017), .ZN(n7020) );
  NOR4_X1 U7955 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n7057)
         );
  INV_X1 U7956 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n7026) );
  AOI22_X1 U7957 ( .A1(n7026), .A2(keyinput44), .B1(keyinput8), .B2(n7025), 
        .ZN(n7024) );
  OAI221_X1 U7958 ( .B1(n7026), .B2(keyinput44), .C1(n7025), .C2(keyinput8), 
        .A(n7024), .ZN(n7039) );
  AOI22_X1 U7959 ( .A1(n7029), .A2(keyinput99), .B1(keyinput71), .B2(n7028), 
        .ZN(n7027) );
  OAI221_X1 U7960 ( .B1(n7029), .B2(keyinput99), .C1(n7028), .C2(keyinput71), 
        .A(n7027), .ZN(n7038) );
  AOI22_X1 U7961 ( .A1(n7032), .A2(keyinput39), .B1(n7031), .B2(keyinput126), 
        .ZN(n7030) );
  OAI221_X1 U7962 ( .B1(n7032), .B2(keyinput39), .C1(n7031), .C2(keyinput126), 
        .A(n7030), .ZN(n7037) );
  XOR2_X1 U7963 ( .A(n7033), .B(keyinput19), .Z(n7035) );
  XNOR2_X1 U7964 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .B(keyinput3), .ZN(n7034)
         );
  NAND2_X1 U7965 ( .A1(n7035), .A2(n7034), .ZN(n7036) );
  NOR4_X1 U7966 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7056)
         );
  AOI22_X1 U7967 ( .A1(n4344), .A2(keyinput103), .B1(keyinput87), .B2(n7041), 
        .ZN(n7040) );
  OAI221_X1 U7968 ( .B1(n4344), .B2(keyinput103), .C1(n7041), .C2(keyinput87), 
        .A(n7040), .ZN(n7054) );
  AOI22_X1 U7969 ( .A1(n7044), .A2(keyinput64), .B1(keyinput21), .B2(n7043), 
        .ZN(n7042) );
  OAI221_X1 U7970 ( .B1(n7044), .B2(keyinput64), .C1(n7043), .C2(keyinput21), 
        .A(n7042), .ZN(n7053) );
  INV_X1 U7971 ( .A(MORE_REG_SCAN_IN), .ZN(n7047) );
  AOI22_X1 U7972 ( .A1(n7047), .A2(keyinput74), .B1(n7046), .B2(keyinput48), 
        .ZN(n7045) );
  OAI221_X1 U7973 ( .B1(n7047), .B2(keyinput74), .C1(n7046), .C2(keyinput48), 
        .A(n7045), .ZN(n7052) );
  XOR2_X1 U7974 ( .A(n7048), .B(keyinput124), .Z(n7050) );
  XNOR2_X1 U7975 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .B(keyinput82), .ZN(n7049)
         );
  NAND2_X1 U7976 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NOR4_X1 U7977 ( .A1(n7054), .A2(n7053), .A3(n7052), .A4(n7051), .ZN(n7055)
         );
  NAND4_X1 U7978 ( .A1(n7058), .A2(n7057), .A3(n7056), .A4(n7055), .ZN(n7122)
         );
  AOI22_X1 U7979 ( .A1(n7060), .A2(keyinput45), .B1(keyinput112), .B2(n5443), 
        .ZN(n7059) );
  OAI221_X1 U7980 ( .B1(n7060), .B2(keyinput45), .C1(n5443), .C2(keyinput112), 
        .A(n7059), .ZN(n7072) );
  INV_X1 U7981 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n7062) );
  AOI22_X1 U7982 ( .A1(n3731), .A2(keyinput38), .B1(n7062), .B2(keyinput34), 
        .ZN(n7061) );
  OAI221_X1 U7983 ( .B1(n3731), .B2(keyinput38), .C1(n7062), .C2(keyinput34), 
        .A(n7061), .ZN(n7071) );
  AOI22_X1 U7984 ( .A1(n7065), .A2(keyinput115), .B1(n7064), .B2(keyinput62), 
        .ZN(n7063) );
  OAI221_X1 U7985 ( .B1(n7065), .B2(keyinput115), .C1(n7064), .C2(keyinput62), 
        .A(n7063), .ZN(n7070) );
  XOR2_X1 U7986 ( .A(n7066), .B(keyinput14), .Z(n7068) );
  XNOR2_X1 U7987 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput121), .ZN(n7067) );
  NAND2_X1 U7988 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  NOR4_X1 U7989 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), .ZN(n7120)
         );
  AOI22_X1 U7990 ( .A1(keyinput68), .A2(n7074), .B1(keyinput105), .B2(n7127), 
        .ZN(n7073) );
  OAI21_X1 U7991 ( .B1(n7074), .B2(keyinput68), .A(n7073), .ZN(n7086) );
  AOI22_X1 U7992 ( .A1(n7077), .A2(keyinput43), .B1(keyinput116), .B2(n7076), 
        .ZN(n7075) );
  OAI221_X1 U7993 ( .B1(n7077), .B2(keyinput43), .C1(n7076), .C2(keyinput116), 
        .A(n7075), .ZN(n7085) );
  INV_X1 U7994 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n7080) );
  AOI22_X1 U7995 ( .A1(n7080), .A2(keyinput53), .B1(n7079), .B2(keyinput46), 
        .ZN(n7078) );
  OAI221_X1 U7996 ( .B1(n7080), .B2(keyinput53), .C1(n7079), .C2(keyinput46), 
        .A(n7078), .ZN(n7084) );
  AOI22_X1 U7997 ( .A1(n6833), .A2(keyinput24), .B1(keyinput25), .B2(n7082), 
        .ZN(n7081) );
  OAI221_X1 U7998 ( .B1(n6833), .B2(keyinput24), .C1(n7082), .C2(keyinput25), 
        .A(n7081), .ZN(n7083) );
  NOR4_X1 U7999 ( .A1(n7086), .A2(n7085), .A3(n7084), .A4(n7083), .ZN(n7119)
         );
  INV_X1 U8000 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7088) );
  AOI22_X1 U8001 ( .A1(n7089), .A2(keyinput77), .B1(keyinput2), .B2(n7088), 
        .ZN(n7087) );
  OAI221_X1 U8002 ( .B1(n7089), .B2(keyinput77), .C1(n7088), .C2(keyinput2), 
        .A(n7087), .ZN(n7102) );
  AOI22_X1 U8003 ( .A1(n7092), .A2(keyinput31), .B1(n7091), .B2(keyinput66), 
        .ZN(n7090) );
  OAI221_X1 U8004 ( .B1(n7092), .B2(keyinput31), .C1(n7091), .C2(keyinput66), 
        .A(n7090), .ZN(n7101) );
  INV_X1 U8005 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n7095) );
  INV_X1 U8006 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U8007 ( .A1(n7095), .A2(keyinput20), .B1(keyinput95), .B2(n7094), 
        .ZN(n7093) );
  OAI221_X1 U8008 ( .B1(n7095), .B2(keyinput20), .C1(n7094), .C2(keyinput95), 
        .A(n7093), .ZN(n7100) );
  AOI22_X1 U8009 ( .A1(n7098), .A2(keyinput29), .B1(keyinput57), .B2(n7097), 
        .ZN(n7096) );
  OAI221_X1 U8010 ( .B1(n7098), .B2(keyinput29), .C1(n7097), .C2(keyinput57), 
        .A(n7096), .ZN(n7099) );
  NOR4_X1 U8011 ( .A1(n7102), .A2(n7101), .A3(n7100), .A4(n7099), .ZN(n7118)
         );
  INV_X1 U8012 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n7104) );
  AOI22_X1 U8013 ( .A1(n7105), .A2(keyinput23), .B1(n7104), .B2(keyinput27), 
        .ZN(n7103) );
  OAI221_X1 U8014 ( .B1(n7105), .B2(keyinput23), .C1(n7104), .C2(keyinput27), 
        .A(n7103), .ZN(n7109) );
  XOR2_X1 U8015 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput97), .Z(n7108)
         );
  XNOR2_X1 U8016 ( .A(n7106), .B(keyinput54), .ZN(n7107) );
  OR3_X1 U8017 ( .A1(n7109), .A2(n7108), .A3(n7107), .ZN(n7116) );
  AOI22_X1 U8018 ( .A1(n7111), .A2(keyinput127), .B1(keyinput117), .B2(n3869), 
        .ZN(n7110) );
  OAI221_X1 U8019 ( .B1(n7111), .B2(keyinput127), .C1(n3869), .C2(keyinput117), 
        .A(n7110), .ZN(n7115) );
  AOI22_X1 U8020 ( .A1(n6029), .A2(keyinput104), .B1(keyinput123), .B2(n7113), 
        .ZN(n7112) );
  OAI221_X1 U8021 ( .B1(n6029), .B2(keyinput104), .C1(n7113), .C2(keyinput123), 
        .A(n7112), .ZN(n7114) );
  NOR3_X1 U8022 ( .A1(n7116), .A2(n7115), .A3(n7114), .ZN(n7117) );
  NAND4_X1 U8023 ( .A1(n7120), .A2(n7119), .A3(n7118), .A4(n7117), .ZN(n7121)
         );
  NOR4_X1 U8024 ( .A1(n7124), .A2(n7123), .A3(n7122), .A4(n7121), .ZN(n7125)
         );
  OAI221_X1 U8025 ( .B1(keyinput105), .B2(n7127), .C1(keyinput105), .C2(n7126), 
        .A(n7125), .ZN(n7128) );
  XNOR2_X1 U8026 ( .A(n7129), .B(n7128), .ZN(U2941) );
  AND2_X1 U3575 ( .A1(n3322), .A2(n3224), .ZN(n3223) );
  CLKBUF_X1 U3577 ( .A(n4343), .Z(n4429) );
  NAND2_X1 U3587 ( .A1(n4247), .A2(n4246), .ZN(n4248) );
  CLKBUF_X1 U3595 ( .A(n3457), .Z(n4812) );
  CLKBUF_X1 U3686 ( .A(n6517), .Z(n3114) );
  CLKBUF_X1 U3707 ( .A(n3434), .Z(n4449) );
  NAND2_X1 U3722 ( .A1(n5100), .A2(n5101), .ZN(n5090) );
endmodule

