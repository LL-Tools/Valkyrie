

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n1996, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741;

  INV_X2 U2238 ( .A(n2480), .ZN(n2817) );
  NOR2_X1 U2239 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2343)
         );
  AND3_X1 U2240 ( .A1(n2417), .A2(n2355), .A3(n2344), .ZN(n2050) );
  INV_X1 U2241 ( .A(n2817), .ZN(n2861) );
  INV_X1 U2242 ( .A(n2473), .ZN(n2538) );
  OR2_X1 U2243 ( .A1(n2980), .A2(n2140), .ZN(n2045) );
  INV_X1 U2244 ( .A(n3984), .ZN(n3496) );
  INV_X1 U2245 ( .A(n3990), .ZN(n3212) );
  INV_X1 U2246 ( .A(n3988), .ZN(n3384) );
  OR2_X1 U2247 ( .A1(n4185), .A2(n4189), .ZN(n4186) );
  XNOR2_X1 U2248 ( .A(n2423), .B(IR_REG_30__SCAN_IN), .ZN(n4480) );
  NAND4_X2 U2249 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .ZN(n3988)
         );
  OAI21_X1 U2250 ( .B1(n3190), .B2(n1996), .A(n2467), .ZN(n2468) );
  NOR2_X1 U2251 ( .A1(n3667), .A2(n3668), .ZN(n3666) );
  NAND2_X2 U2252 ( .A1(n3642), .A2(n2806), .ZN(n3697) );
  AND2_X1 U2253 ( .A1(n2432), .A2(n4480), .ZN(n2475) );
  NAND2_X1 U2254 ( .A1(n2471), .A2(n4557), .ZN(n1996) );
  NAND2_X1 U2255 ( .A1(n2471), .A2(n4557), .ZN(n2498) );
  NAND2_X2 U2256 ( .A1(n2413), .A2(IR_REG_31__SCAN_IN), .ZN(n2341) );
  AOI22_X2 U2257 ( .A1(n3111), .A2(REG1_REG_3__SCAN_IN), .B1(n4493), .B2(n2381), .ZN(n2382) );
  AND2_X1 U2258 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  NAND2_X2 U2259 ( .A1(n3006), .A2(n3913), .ZN(n3908) );
  INV_X2 U2260 ( .A(n2817), .ZN(n2912) );
  INV_X1 U2261 ( .A(n3987), .ZN(n3281) );
  INV_X2 U2262 ( .A(n3198), .ZN(n3272) );
  INV_X4 U2263 ( .A(n2850), .ZN(n2517) );
  AND2_X2 U2264 ( .A1(n2440), .A2(n2910), .ZN(n2850) );
  XNOR2_X1 U2265 ( .A(n2338), .B(n2337), .ZN(n3241) );
  OR2_X1 U2266 ( .A1(n2422), .A2(n2258), .ZN(n2423) );
  NOR2_X1 U2267 ( .A1(n2420), .A2(IR_REG_29__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U2268 ( .A1(n2047), .A2(n2046), .ZN(n2063) );
  AOI21_X1 U2269 ( .B1(n4076), .B2(n4318), .A(n4075), .ZN(n4348) );
  NAND2_X1 U2270 ( .A1(n2045), .A2(n2044), .ZN(n4125) );
  AND2_X1 U2271 ( .A1(n3056), .A2(n3055), .ZN(n3057) );
  AND2_X1 U2272 ( .A1(n3063), .A2(n3062), .ZN(n3064) );
  AOI21_X1 U2273 ( .B1(n2325), .B2(REG2_REG_16__SCAN_IN), .A(n2105), .ZN(n2104) );
  NAND2_X1 U2274 ( .A1(n2232), .A2(n2230), .ZN(n3403) );
  AND2_X1 U2275 ( .A1(n2304), .A2(n2635), .ZN(n2305) );
  AND2_X1 U2276 ( .A1(n2618), .A2(n3656), .ZN(n3657) );
  NOR2_X1 U2277 ( .A1(n2605), .A2(n2209), .ZN(n2208) );
  AND2_X1 U2278 ( .A1(n2617), .A2(n2616), .ZN(n3656) );
  OR2_X1 U2279 ( .A1(n3655), .A2(n2619), .ZN(n2605) );
  AND2_X1 U2280 ( .A1(n2950), .A2(n3908), .ZN(n2126) );
  NOR2_X1 U2281 ( .A1(n3373), .A2(n2251), .ZN(n2389) );
  AND2_X1 U2282 ( .A1(n3902), .A2(n3899), .ZN(n3853) );
  INV_X1 U2283 ( .A(n3343), .ZN(n3336) );
  NAND2_X1 U2284 ( .A1(n2449), .A2(n2448), .ZN(n3048) );
  NAND2_X1 U2285 ( .A1(n2446), .A2(n2445), .ZN(n3992) );
  NAND2_X1 U2286 ( .A1(n3828), .A2(DATAI_0_), .ZN(n2448) );
  OR2_X1 U2287 ( .A1(n3189), .A2(n4485), .ZN(n4557) );
  CLKBUF_X3 U2288 ( .A(n2475), .Z(n3823) );
  AND3_X1 U2289 ( .A1(n2097), .A2(n2094), .A3(n2016), .ZN(n2273) );
  XNOR2_X1 U2290 ( .A(n2292), .B(IR_REG_10__SCAN_IN), .ZN(n4490) );
  CLKBUF_X3 U2291 ( .A(n2474), .Z(n2855) );
  XNOR2_X1 U2292 ( .A(n2363), .B(IR_REG_24__SCAN_IN), .ZN(n2889) );
  XNOR2_X1 U2293 ( .A(n2370), .B(IR_REG_26__SCAN_IN), .ZN(n4482) );
  AND2_X1 U2294 ( .A1(n2368), .A2(n2369), .ZN(n4483) );
  NAND2_X1 U2295 ( .A1(n2362), .A2(IR_REG_31__SCAN_IN), .ZN(n2363) );
  AOI21_X1 U2296 ( .B1(n2412), .B2(n2411), .A(n2410), .ZN(n2414) );
  XNOR2_X1 U2297 ( .A(n2259), .B(n4493), .ZN(n3112) );
  XNOR2_X1 U2298 ( .A(n2347), .B(IR_REG_22__SCAN_IN), .ZN(n4484) );
  NOR2_X1 U2299 ( .A1(n3996), .A2(n2244), .ZN(n2259) );
  MUX2_X1 U2300 ( .A(IR_REG_31__SCAN_IN), .B(n2418), .S(IR_REG_29__SCAN_IN), 
        .Z(n2419) );
  CLKBUF_X1 U2301 ( .A(n2422), .Z(n3610) );
  NOR2_X1 U2302 ( .A1(n2346), .A2(n2356), .ZN(n2349) );
  NAND2_X1 U2303 ( .A1(n2353), .A2(n2352), .ZN(n2364) );
  OR2_X1 U2304 ( .A1(n2257), .A2(n2258), .ZN(n2255) );
  NOR2_X1 U2305 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2189)
         );
  NOR2_X1 U2306 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2188)
         );
  NOR2_X1 U2307 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2192)
         );
  NOR2_X1 U2308 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2187)
         );
  NOR2_X2 U2309 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2344)
         );
  INV_X1 U2310 ( .A(IR_REG_21__SCAN_IN), .ZN(n2342) );
  NOR2_X1 U2311 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2190)
         );
  NOR2_X1 U2312 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2354)
         );
  NAND4_X4 U2313 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n2938)
         );
  NAND4_X2 U2314 ( .A1(n2558), .A2(n2557), .A3(n2556), .A4(n2555), .ZN(n3986)
         );
  INV_X2 U2315 ( .A(n2938), .ZN(n3190) );
  AND2_X1 U2316 ( .A1(n4480), .A2(n2425), .ZN(n2474) );
  AOI21_X2 U2317 ( .B1(n4356), .B2(n4578), .A(n4355), .ZN(n4429) );
  NOR2_X2 U2318 ( .A1(n4371), .A2(n3053), .ZN(n4155) );
  NOR2_X2 U2319 ( .A1(n3666), .A2(n2753), .ZN(n3070) );
  OR2_X1 U2320 ( .A1(n1999), .A2(n2655), .ZN(n2206) );
  NOR2_X1 U2321 ( .A1(n2818), .A2(n4651), .ZN(n2807) );
  INV_X1 U2322 ( .A(n4106), .ZN(n2992) );
  AND2_X1 U2323 ( .A1(n2707), .A2(n3726), .ZN(n2709) );
  NAND2_X1 U2325 ( .A1(n2143), .A2(n2981), .ZN(n2140) );
  INV_X1 U2326 ( .A(n2138), .ZN(n2137) );
  OAI21_X1 U2327 ( .B1(n2976), .B2(n2139), .A(n2979), .ZN(n2138) );
  NOR2_X1 U2328 ( .A1(n2693), .A2(n3719), .ZN(n2043) );
  INV_X1 U2329 ( .A(n2364), .ZN(n2355) );
  INV_X1 U2330 ( .A(n2269), .ZN(n2306) );
  AOI21_X1 U2331 ( .B1(n2206), .B2(n2003), .A(n2201), .ZN(n2200) );
  NOR2_X1 U2332 ( .A1(n2204), .A2(n2646), .ZN(n2201) );
  INV_X1 U2333 ( .A(n2204), .ZN(n2203) );
  OR2_X1 U2334 ( .A1(n2790), .A2(n2789), .ZN(n2818) );
  NAND2_X1 U2335 ( .A1(n2359), .A2(n2358), .ZN(n2176) );
  OR2_X1 U2336 ( .A1(n2372), .A2(n2415), .ZN(n2359) );
  INV_X1 U2337 ( .A(n2538), .ZN(n3824) );
  INV_X1 U2338 ( .A(n2855), .ZN(n2921) );
  NOR2_X1 U2339 ( .A1(n3120), .A2(n2102), .ZN(n3119) );
  NAND2_X1 U2340 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2102) );
  XNOR2_X1 U2341 ( .A(n2379), .B(n3265), .ZN(n3994) );
  INV_X1 U2342 ( .A(n3371), .ZN(n2290) );
  INV_X1 U2343 ( .A(n4548), .ZN(n2675) );
  NOR2_X1 U2344 ( .A1(n2994), .A2(n2149), .ZN(n2148) );
  INV_X1 U2345 ( .A(n2993), .ZN(n2149) );
  OAI22_X1 U2346 ( .A1(n4125), .A2(n2991), .B1(n4154), .B2(n4136), .ZN(n4106)
         );
  OR2_X1 U2347 ( .A1(n2768), .A2(n4653), .ZN(n2790) );
  NAND2_X1 U2348 ( .A1(n2042), .A2(REG3_REG_19__SCAN_IN), .ZN(n2755) );
  INV_X1 U2349 ( .A(n2739), .ZN(n2042) );
  AND2_X1 U2350 ( .A1(n4132), .A2(n4151), .ZN(n2986) );
  NAND2_X1 U2351 ( .A1(n3683), .A2(n2205), .ZN(n2204) );
  INV_X1 U2352 ( .A(n3614), .ZN(n2205) );
  INV_X1 U2353 ( .A(n3069), .ZN(n2229) );
  INV_X1 U2354 ( .A(n3846), .ZN(n3033) );
  AND2_X1 U2355 ( .A1(n3948), .A2(n3032), .ZN(n3816) );
  INV_X1 U2356 ( .A(n2978), .ZN(n2139) );
  AND2_X1 U2357 ( .A1(n3022), .A2(n3937), .ZN(n2086) );
  INV_X1 U2358 ( .A(n3940), .ZN(n3022) );
  INV_X1 U2359 ( .A(n4284), .ZN(n2976) );
  NOR2_X1 U2360 ( .A1(n3859), .A2(n2133), .ZN(n2132) );
  INV_X1 U2361 ( .A(n2965), .ZN(n2133) );
  NAND2_X1 U2362 ( .A1(n2514), .A2(n2015), .ZN(n3903) );
  NAND2_X1 U2363 ( .A1(n3905), .A2(n3903), .ZN(n3337) );
  INV_X1 U2364 ( .A(n4178), .ZN(n3053) );
  AND2_X1 U2365 ( .A1(n3619), .A2(n3637), .ZN(n2182) );
  INV_X1 U2366 ( .A(n2128), .ZN(n2367) );
  INV_X1 U2367 ( .A(n2356), .ZN(n2129) );
  OR2_X1 U2368 ( .A1(n2275), .A2(IR_REG_6__SCAN_IN), .ZN(n2284) );
  NAND2_X1 U2369 ( .A1(n3380), .A2(n3381), .ZN(n2235) );
  OR2_X1 U2370 ( .A1(n3380), .A2(n3381), .ZN(n2234) );
  NAND2_X1 U2371 ( .A1(n2031), .A2(n2221), .ZN(n2220) );
  INV_X1 U2372 ( .A(n3783), .ZN(n2221) );
  XNOR2_X1 U2373 ( .A(n2502), .B(n2850), .ZN(n2505) );
  NAND2_X1 U2374 ( .A1(n2194), .A2(n2195), .ZN(n3769) );
  AOI21_X1 U2375 ( .B1(n2196), .B2(n2202), .A(n2023), .ZN(n2195) );
  INV_X1 U2376 ( .A(n2220), .ZN(n2219) );
  NOR2_X1 U2377 ( .A1(n2219), .A2(n2215), .ZN(n2214) );
  INV_X1 U2378 ( .A(n2250), .ZN(n2215) );
  AND2_X1 U2379 ( .A1(n2451), .A2(n2450), .ZN(n2457) );
  INV_X1 U2380 ( .A(n4191), .ZN(n3764) );
  NAND2_X1 U2381 ( .A1(n2207), .A2(n2020), .ZN(n2212) );
  XNOR2_X1 U2382 ( .A(n2483), .B(n2517), .ZN(n2488) );
  OR2_X1 U2383 ( .A1(n2834), .A2(n3700), .ZN(n2838) );
  NOR2_X1 U2384 ( .A1(n3119), .A2(n2013), .ZN(n3998) );
  AOI21_X1 U2385 ( .B1(n3994), .B2(n3993), .A(n2237), .ZN(n2380) );
  NOR2_X1 U2386 ( .A1(n2259), .A2(n3114), .ZN(n2260) );
  OR2_X1 U2387 ( .A1(n2267), .A2(n2266), .ZN(n2269) );
  INV_X1 U2388 ( .A(IR_REG_4__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U2389 ( .A1(n3143), .A2(REG2_REG_6__SCAN_IN), .ZN(n2093) );
  NAND2_X1 U2390 ( .A1(n2274), .A2(n3088), .ZN(n2092) );
  INV_X1 U2391 ( .A(n3155), .ZN(n2090) );
  AND2_X1 U2392 ( .A1(n4490), .A2(REG1_REG_10__SCAN_IN), .ZN(n2164) );
  NAND2_X1 U2393 ( .A1(n2117), .A2(n4490), .ZN(n2108) );
  AOI21_X1 U2394 ( .B1(n2115), .B2(REG2_REG_10__SCAN_IN), .A(n4490), .ZN(n2111) );
  NAND2_X1 U2395 ( .A1(n3451), .A2(n2301), .ZN(n2304) );
  NAND2_X1 U2396 ( .A1(n2300), .A2(REG2_REG_11__SCAN_IN), .ZN(n2301) );
  OAI21_X1 U2397 ( .B1(n4489), .B2(n3561), .A(n3453), .ZN(n2390) );
  NAND2_X1 U2398 ( .A1(n4009), .A2(n2236), .ZN(n2393) );
  NAND2_X1 U2399 ( .A1(n4035), .A2(n2395), .ZN(n2396) );
  NAND2_X1 U2400 ( .A1(n4033), .A2(REG1_REG_15__SCAN_IN), .ZN(n2395) );
  INV_X1 U2401 ( .A(n4505), .ZN(n2105) );
  AOI21_X1 U2402 ( .B1(n2172), .B2(n2171), .A(n2398), .ZN(n2170) );
  INV_X1 U2403 ( .A(n4508), .ZN(n2171) );
  AND2_X1 U2404 ( .A1(n2926), .A2(n2925), .ZN(n3831) );
  OAI21_X1 U2405 ( .B1(n4127), .B2(n2077), .A(n2074), .ZN(n4068) );
  INV_X1 U2406 ( .A(n2079), .ZN(n2077) );
  AND2_X1 U2407 ( .A1(n2078), .A2(n2075), .ZN(n2074) );
  NAND2_X1 U2408 ( .A1(n2079), .A2(n2076), .ZN(n2075) );
  NAND2_X1 U2409 ( .A1(n2992), .A2(n2242), .ZN(n2152) );
  INV_X1 U2410 ( .A(n4118), .ZN(n4112) );
  OR2_X1 U2411 ( .A1(n2990), .A2(n2005), .ZN(n2044) );
  INV_X1 U2412 ( .A(n4094), .ZN(n4135) );
  INV_X1 U2413 ( .A(n4113), .ZN(n4154) );
  NAND2_X1 U2414 ( .A1(n4204), .A2(n2981), .ZN(n4143) );
  NAND2_X1 U2415 ( .A1(n2754), .A2(REG3_REG_20__SCAN_IN), .ZN(n2768) );
  INV_X1 U2416 ( .A(n4193), .ZN(n4228) );
  NAND2_X1 U2417 ( .A1(n2977), .A2(n2976), .ZN(n4281) );
  INV_X1 U2418 ( .A(n2691), .ZN(n2668) );
  INV_X1 U2419 ( .A(n2043), .ZN(n2723) );
  INV_X1 U2420 ( .A(n4275), .ZN(n4312) );
  OR2_X1 U2421 ( .A1(n3036), .A2(n2915), .ZN(n3234) );
  OR2_X1 U2422 ( .A1(n3036), .A2(n4481), .ZN(n4315) );
  NOR2_X2 U2423 ( .A1(n3601), .A2(n3052), .ZN(n4298) );
  INV_X1 U2424 ( .A(IR_REG_26__SCAN_IN), .ZN(n4596) );
  AND2_X1 U2425 ( .A1(n2891), .A2(n4482), .ZN(n3097) );
  NAND4_X1 U2426 ( .A1(n2051), .A2(n2050), .A3(n2313), .A4(n1998), .ZN(n2420)
         );
  AND2_X1 U2427 ( .A1(n2052), .A2(n2053), .ZN(n2051) );
  AND2_X1 U2428 ( .A1(n2354), .A2(n2342), .ZN(n2053) );
  XNOR2_X1 U2429 ( .A(n2277), .B(IR_REG_7__SCAN_IN), .ZN(n3150) );
  AND2_X1 U2430 ( .A1(n3643), .A2(n3644), .ZN(n2806) );
  NAND2_X1 U2431 ( .A1(n3759), .A2(n3760), .ZN(n3642) );
  INV_X1 U2432 ( .A(n4252), .ZN(n4206) );
  AND2_X1 U2433 ( .A1(n2819), .A2(n2820), .ZN(n4158) );
  NAND2_X1 U2434 ( .A1(n2860), .A2(n2859), .ZN(n3325) );
  NAND2_X1 U2435 ( .A1(n2745), .A2(n2744), .ZN(n4273) );
  NAND2_X1 U2436 ( .A1(n2168), .A2(n2167), .ZN(n3373) );
  NAND2_X1 U2437 ( .A1(n2388), .A2(n2169), .ZN(n2167) );
  XNOR2_X1 U2438 ( .A(n2390), .B(n3526), .ZN(n3529) );
  NAND2_X1 U2439 ( .A1(n3529), .A2(REG1_REG_12__SCAN_IN), .ZN(n3528) );
  NAND2_X1 U2440 ( .A1(n4011), .A2(n4010), .ZN(n4009) );
  XNOR2_X1 U2441 ( .A(n2393), .B(n4019), .ZN(n4023) );
  NAND2_X1 U2442 ( .A1(n4023), .A2(REG1_REG_14__SCAN_IN), .ZN(n4022) );
  XNOR2_X1 U2443 ( .A(n2396), .B(n4486), .ZN(n4041) );
  INV_X1 U2444 ( .A(n2339), .ZN(n2119) );
  AOI21_X1 U2445 ( .B1(n2339), .B2(n2335), .A(n4014), .ZN(n2121) );
  INV_X1 U2446 ( .A(n4534), .ZN(n4329) );
  OR2_X1 U2447 ( .A1(n4083), .A2(n4418), .ZN(n3056) );
  INV_X1 U2448 ( .A(n4088), .ZN(n2046) );
  NAND2_X1 U2449 ( .A1(n4082), .A2(n4578), .ZN(n2047) );
  OR2_X1 U2450 ( .A1(n4083), .A2(n4478), .ZN(n3063) );
  NAND2_X1 U2451 ( .A1(n2056), .A2(n2059), .ZN(n2054) );
  INV_X1 U2452 ( .A(n2012), .ZN(n2081) );
  INV_X1 U2453 ( .A(n3926), .ZN(n2061) );
  NOR2_X1 U2454 ( .A1(n3906), .A2(n2072), .ZN(n2071) );
  INV_X1 U2455 ( .A(n3193), .ZN(n3860) );
  OR2_X1 U2456 ( .A1(n2715), .A2(n3724), .ZN(n2720) );
  NOR2_X1 U2457 ( .A1(n2636), .A2(n2430), .ZN(n2040) );
  AND2_X1 U2458 ( .A1(n2607), .A2(n2606), .ZN(n2619) );
  INV_X1 U2459 ( .A(n2249), .ZN(n2209) );
  INV_X1 U2460 ( .A(IR_REG_27__SCAN_IN), .ZN(n2415) );
  INV_X1 U2461 ( .A(IR_REG_28__SCAN_IN), .ZN(n2416) );
  NOR2_X1 U2462 ( .A1(n2113), .A2(n2110), .ZN(n2109) );
  NOR2_X1 U2463 ( .A1(n2011), .A2(n2114), .ZN(n2113) );
  NAND2_X1 U2464 ( .A1(n4490), .A2(n2116), .ZN(n2115) );
  INV_X1 U2465 ( .A(n2238), .ZN(n2174) );
  NOR2_X1 U2466 ( .A1(n2081), .A2(n2080), .ZN(n2079) );
  INV_X1 U2467 ( .A(n3951), .ZN(n2080) );
  OR2_X1 U2468 ( .A1(n2082), .A2(n2081), .ZN(n2078) );
  AND2_X1 U2469 ( .A1(n4093), .A2(n2084), .ZN(n2082) );
  NAND2_X1 U2470 ( .A1(n2142), .A2(n2981), .ZN(n2141) );
  INV_X1 U2471 ( .A(n3851), .ZN(n2142) );
  OR2_X1 U2472 ( .A1(n2247), .A2(n2988), .ZN(n2989) );
  NAND2_X1 U2473 ( .A1(n4309), .A2(n4310), .ZN(n2087) );
  INV_X1 U2475 ( .A(n2060), .ZN(n2059) );
  AOI21_X1 U2476 ( .B1(n2060), .B2(n2058), .A(n2057), .ZN(n2056) );
  INV_X1 U2477 ( .A(n3915), .ZN(n2058) );
  INV_X1 U2478 ( .A(n2028), .ZN(n2062) );
  AOI21_X1 U2479 ( .B1(n2071), .B2(n2069), .A(n2068), .ZN(n2067) );
  INV_X1 U2480 ( .A(n3903), .ZN(n2069) );
  INV_X1 U2481 ( .A(n2071), .ZN(n2070) );
  NAND2_X1 U2482 ( .A1(n2938), .A2(n3204), .ZN(n3894) );
  INV_X1 U2483 ( .A(IR_REG_0__SCAN_IN), .ZN(n2186) );
  AND2_X1 U2484 ( .A1(n2345), .A2(n2343), .ZN(n2052) );
  NAND2_X1 U2485 ( .A1(n2365), .A2(IR_REG_31__SCAN_IN), .ZN(n2350) );
  INV_X1 U2486 ( .A(IR_REG_3__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2487 ( .A1(n2040), .A2(REG3_REG_14__SCAN_IN), .ZN(n2691) );
  INV_X1 U2488 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2593) );
  INV_X1 U2489 ( .A(n2471), .ZN(n2878) );
  NAND2_X1 U2490 ( .A1(n3270), .A2(n3271), .ZN(n2223) );
  XNOR2_X1 U2491 ( .A(n2441), .B(n2850), .ZN(n3614) );
  INV_X1 U2492 ( .A(n2040), .ZN(n2657) );
  NAND2_X1 U2493 ( .A1(n2229), .A2(n2227), .ZN(n2224) );
  NAND2_X1 U2494 ( .A1(n2229), .A2(n2226), .ZN(n2225) );
  NAND2_X1 U2495 ( .A1(n2228), .A2(n3067), .ZN(n2227) );
  INV_X1 U2496 ( .A(n2498), .ZN(n2866) );
  AND3_X1 U2497 ( .A1(n2512), .A2(n2511), .A3(n2510), .ZN(n2514) );
  NOR2_X1 U2498 ( .A1(n3132), .A2(n2100), .ZN(n2099) );
  INV_X1 U2499 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2100) );
  NAND2_X1 U2500 ( .A1(n2101), .A2(n2098), .ZN(n2097) );
  NOR2_X1 U2501 ( .A1(n3132), .A2(n2156), .ZN(n2098) );
  NAND2_X1 U2502 ( .A1(n2306), .A2(n2270), .ZN(n2275) );
  NAND2_X1 U2503 ( .A1(n2383), .A2(n2155), .ZN(n2154) );
  NOR2_X1 U2504 ( .A1(n3134), .A2(n2156), .ZN(n2155) );
  NAND2_X1 U2505 ( .A1(n3161), .A2(n2157), .ZN(n2153) );
  NOR2_X1 U2506 ( .A1(n3134), .A2(n2159), .ZN(n2157) );
  NAND2_X1 U2507 ( .A1(n2089), .A2(n2088), .ZN(n2280) );
  NAND2_X1 U2508 ( .A1(n3155), .A2(n2008), .ZN(n2088) );
  NAND2_X1 U2509 ( .A1(n2093), .A2(n2018), .ZN(n2089) );
  AOI22_X1 U2510 ( .A1(n3151), .A2(n2385), .B1(n2384), .B2(n3154), .ZN(n2387)
         );
  AND2_X1 U2511 ( .A1(n3230), .A2(REG1_REG_8__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U2512 ( .A1(n2117), .A2(n3412), .ZN(n2116) );
  OAI21_X1 U2513 ( .B1(n2293), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2295) );
  INV_X1 U2514 ( .A(IR_REG_11__SCAN_IN), .ZN(n2294) );
  AOI21_X1 U2515 ( .B1(n4004), .B2(n2309), .A(n2308), .ZN(n2315) );
  INV_X1 U2516 ( .A(n3832), .ZN(n4071) );
  NOR2_X1 U2517 ( .A1(n2180), .A2(n2179), .ZN(n2178) );
  OR2_X1 U2518 ( .A1(n2995), .A2(n4112), .ZN(n2180) );
  OR2_X1 U2519 ( .A1(n4100), .A2(n4131), .ZN(n2179) );
  NAND2_X1 U2520 ( .A1(n4108), .A2(n3951), .ZN(n2085) );
  AND2_X1 U2521 ( .A1(n2877), .A2(n2876), .ZN(n4096) );
  OR2_X1 U2522 ( .A1(n4085), .A2(n2921), .ZN(n2877) );
  NAND2_X1 U2523 ( .A1(n2048), .A2(n3848), .ZN(n4148) );
  AOI21_X1 U2524 ( .B1(n2137), .B2(n2139), .A(n2032), .ZN(n2135) );
  INV_X1 U2525 ( .A(n4272), .ZN(n4278) );
  NAND2_X1 U2526 ( .A1(n2043), .A2(n2721), .ZN(n2739) );
  AND2_X1 U2527 ( .A1(n4248), .A2(n4249), .ZN(n4284) );
  AND2_X1 U2528 ( .A1(n3937), .A2(n3935), .ZN(n4310) );
  AOI21_X1 U2529 ( .B1(n2132), .B2(n2966), .A(n2022), .ZN(n2130) );
  NAND2_X1 U2530 ( .A1(n2134), .A2(n2965), .ZN(n3581) );
  OR2_X1 U2531 ( .A1(n3570), .A2(n2966), .ZN(n2134) );
  INV_X1 U2532 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2580) );
  OR2_X1 U2533 ( .A1(n2581), .A2(n2580), .ZN(n2594) );
  INV_X1 U2534 ( .A(n3985), .ZN(n3461) );
  INV_X1 U2535 ( .A(n4315), .ZN(n4292) );
  NAND2_X1 U2536 ( .A1(n2073), .A2(n3905), .ZN(n3357) );
  NAND2_X1 U2537 ( .A1(n3003), .A2(n3903), .ZN(n2073) );
  NAND2_X1 U2538 ( .A1(n3248), .A2(n3336), .ZN(n3363) );
  NAND2_X1 U2539 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2541) );
  INV_X1 U2540 ( .A(n4253), .ZN(n4311) );
  INV_X1 U2541 ( .A(n3989), .ZN(n3359) );
  CLKBUF_X1 U2542 ( .A(n3196), .Z(n3213) );
  NAND2_X1 U2543 ( .A1(n4063), .A2(n4057), .ZN(n4055) );
  OAI21_X1 U2544 ( .B1(n2992), .B2(n2147), .A(n2144), .ZN(n4342) );
  AOI21_X1 U2545 ( .B1(n2146), .B2(n2145), .A(n2004), .ZN(n2144) );
  INV_X1 U2546 ( .A(n2242), .ZN(n2145) );
  AND2_X1 U2547 ( .A1(n2182), .A2(n3800), .ZN(n2181) );
  NAND2_X1 U2548 ( .A1(n3550), .A2(n2182), .ZN(n3603) );
  AND2_X1 U2549 ( .A1(n3550), .A2(n3619), .ZN(n3590) );
  INV_X1 U2550 ( .A(n3481), .ZN(n3517) );
  AND2_X1 U2551 ( .A1(n2010), .A2(n3654), .ZN(n2183) );
  NAND2_X1 U2552 ( .A1(n3050), .A2(n2001), .ZN(n3465) );
  NAND2_X1 U2553 ( .A1(n3050), .A2(n3049), .ZN(n3425) );
  INV_X1 U2554 ( .A(n4557), .ZN(n4575) );
  NOR2_X2 U2555 ( .A1(n2006), .A2(n3219), .ZN(n3250) );
  NAND2_X1 U2556 ( .A1(n4530), .A2(n2997), .ZN(n4558) );
  NAND2_X1 U2557 ( .A1(n2367), .A2(n4596), .ZN(n2177) );
  INV_X1 U2558 ( .A(IR_REG_24__SCAN_IN), .ZN(n2353) );
  INV_X1 U2559 ( .A(IR_REG_17__SCAN_IN), .ZN(n2328) );
  OR2_X1 U2560 ( .A1(n2288), .A2(IR_REG_9__SCAN_IN), .ZN(n2293) );
  NOR2_X1 U2561 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2257)
         );
  NAND2_X1 U2562 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2252)
         );
  NAND2_X1 U2563 ( .A1(n2235), .A2(n2537), .ZN(n2231) );
  NAND2_X1 U2564 ( .A1(n2216), .A2(n2220), .ZN(n3628) );
  NAND2_X1 U2565 ( .A1(n2222), .A2(n2000), .ZN(n2216) );
  NAND2_X1 U2566 ( .A1(n3682), .A2(n2198), .ZN(n2197) );
  INV_X1 U2567 ( .A(n3498), .ZN(n3654) );
  XNOR2_X1 U2568 ( .A(n2503), .B(n2505), .ZN(n3271) );
  OAI21_X1 U2569 ( .B1(n2735), .B2(n3770), .A(n3771), .ZN(n2738) );
  AND2_X1 U2570 ( .A1(n2909), .A2(n3773), .ZN(n2900) );
  NAND2_X1 U2571 ( .A1(n2213), .A2(n2217), .ZN(n2906) );
  AND2_X1 U2572 ( .A1(n2218), .A2(n3627), .ZN(n2217) );
  OR2_X1 U2573 ( .A1(n2000), .A2(n2219), .ZN(n2218) );
  NOR2_X1 U2574 ( .A1(n3751), .A2(n3071), .ZN(n3074) );
  NAND2_X1 U2575 ( .A1(n2223), .A2(n2506), .ZN(n3331) );
  NOR2_X1 U2576 ( .A1(n3070), .A2(n3749), .ZN(n3751) );
  INV_X1 U2577 ( .A(n3010), .ZN(n3619) );
  NAND2_X1 U2578 ( .A1(n2199), .A2(n3683), .ZN(n3617) );
  NAND2_X1 U2579 ( .A1(n2647), .A2(n2646), .ZN(n2199) );
  INV_X1 U2580 ( .A(n3787), .ZN(n3796) );
  INV_X1 U2581 ( .A(n3776), .ZN(n3798) );
  INV_X1 U2582 ( .A(n3805), .ZN(n3773) );
  INV_X1 U2583 ( .A(n3763), .ZN(n3778) );
  NAND2_X1 U2584 ( .A1(n3278), .A2(n2537), .ZN(n3383) );
  AND2_X1 U2585 ( .A1(n2870), .A2(n2841), .ZN(n4120) );
  NAND2_X1 U2586 ( .A1(n2920), .A2(n3184), .ZN(n3802) );
  NAND2_X1 U2587 ( .A1(n2813), .A2(n2812), .ZN(n4113) );
  NAND2_X1 U2588 ( .A1(n2041), .A2(n2824), .ZN(n4132) );
  NAND2_X1 U2589 ( .A1(n4158), .A2(n2855), .ZN(n2041) );
  NAND2_X1 U2590 ( .A1(n2797), .A2(n2796), .ZN(n4191) );
  NAND2_X1 U2591 ( .A1(n2785), .A2(n2784), .ZN(n4208) );
  NAND2_X1 U2592 ( .A1(n2774), .A2(n2773), .ZN(n4193) );
  OR2_X1 U2593 ( .A1(n4217), .A2(n2921), .ZN(n2774) );
  NAND2_X1 U2594 ( .A1(n2761), .A2(n2760), .ZN(n4252) );
  NAND2_X1 U2595 ( .A1(n2674), .A2(n2673), .ZN(n3979) );
  OAI211_X1 U2596 ( .C1(n4330), .C2(n2921), .A(n2683), .B(n2682), .ZN(n4291)
         );
  OAI211_X1 U2597 ( .C1(n3605), .C2(n2921), .A(n2697), .B(n2696), .ZN(n4313)
         );
  NAND2_X1 U2598 ( .A1(n2514), .A2(n2513), .ZN(n3989) );
  NAND4_X2 U2599 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n3990)
         );
  NAND2_X1 U2600 ( .A1(n2473), .A2(REG0_REG_2__SCAN_IN), .ZN(n2478) );
  AND3_X1 U2601 ( .A1(n2444), .A2(n2443), .A3(n2442), .ZN(n2446) );
  XNOR2_X1 U2602 ( .A(n2382), .B(n3083), .ZN(n3161) );
  AND2_X1 U2603 ( .A1(n2096), .A2(n2095), .ZN(n3133) );
  NAND2_X1 U2604 ( .A1(n2101), .A2(n3083), .ZN(n2095) );
  NAND2_X1 U2605 ( .A1(n3162), .A2(REG2_REG_4__SCAN_IN), .ZN(n2096) );
  AND2_X1 U2606 ( .A1(n2158), .A2(n2162), .ZN(n3135) );
  NAND2_X1 U2607 ( .A1(n2383), .A2(n3083), .ZN(n2162) );
  NAND2_X1 U2608 ( .A1(n3161), .A2(REG1_REG_4__SCAN_IN), .ZN(n2158) );
  XNOR2_X1 U2609 ( .A(n2161), .B(n2160), .ZN(n3142) );
  AOI22_X1 U2610 ( .A1(n3142), .A2(REG1_REG_6__SCAN_IN), .B1(n3088), .B2(n2161), .ZN(n3151) );
  INV_X1 U2611 ( .A(n2091), .ZN(n3156) );
  NAND2_X1 U2612 ( .A1(n2093), .A2(n2092), .ZN(n2091) );
  XNOR2_X1 U2613 ( .A(n2387), .B(n2386), .ZN(n3230) );
  XNOR2_X1 U2614 ( .A(n2389), .B(n4490), .ZN(n3415) );
  NAND2_X1 U2615 ( .A1(n3415), .A2(REG1_REG_10__SCAN_IN), .ZN(n3414) );
  OAI21_X1 U2616 ( .B1(n2389), .B2(n2029), .A(n2163), .ZN(n3455) );
  NAND2_X1 U2617 ( .A1(n2389), .A2(n2164), .ZN(n2163) );
  OR2_X1 U2618 ( .A1(n4490), .A2(n2166), .ZN(n2165) );
  INV_X1 U2619 ( .A(n3447), .ZN(n2298) );
  XNOR2_X1 U2620 ( .A(n2304), .B(n3526), .ZN(n3524) );
  NAND2_X1 U2621 ( .A1(n3528), .A2(n2239), .ZN(n4011) );
  OR2_X1 U2622 ( .A1(n2391), .A2(n3526), .ZN(n2239) );
  NAND2_X1 U2623 ( .A1(n4022), .A2(n2240), .ZN(n4037) );
  OR2_X1 U2624 ( .A1(n2394), .A2(n4019), .ZN(n2240) );
  OR2_X1 U2625 ( .A1(n4497), .A2(n4495), .ZN(n4514) );
  OAI21_X1 U2626 ( .B1(n4041), .B2(REG1_REG_16__SCAN_IN), .A(n2397), .ZN(n4507) );
  INV_X1 U2627 ( .A(n4031), .ZN(n4517) );
  NAND2_X1 U2628 ( .A1(n2106), .A2(n2325), .ZN(n4504) );
  OR2_X1 U2629 ( .A1(n4042), .A2(REG2_REG_16__SCAN_IN), .ZN(n2106) );
  OR2_X1 U2630 ( .A1(n4497), .A2(n4481), .ZN(n4529) );
  AOI21_X1 U2631 ( .B1(n4516), .B2(n4515), .A(n4514), .ZN(n4522) );
  NAND2_X1 U2632 ( .A1(n4506), .A2(n2238), .ZN(n4516) );
  NAND2_X1 U2633 ( .A1(n2039), .A2(n2150), .ZN(n4061) );
  NAND2_X1 U2634 ( .A1(n2152), .A2(n2148), .ZN(n2039) );
  OAI21_X1 U2635 ( .B1(n3039), .B2(n4210), .A(n3038), .ZN(n4088) );
  XNOR2_X1 U2636 ( .A(n4068), .B(n2083), .ZN(n3039) );
  NAND2_X1 U2637 ( .A1(n2152), .A2(n2993), .ZN(n4091) );
  NAND2_X1 U2638 ( .A1(n4281), .A2(n2978), .ZN(n4261) );
  INV_X1 U2639 ( .A(n4285), .ZN(n4333) );
  INV_X2 U2640 ( .A(n4538), .ZN(n4540) );
  NAND2_X2 U2641 ( .A1(n3240), .A2(n4329), .ZN(n4538) );
  AND2_X1 U2642 ( .A1(n3041), .A2(n3235), .ZN(n4534) );
  INV_X1 U2643 ( .A(n4243), .ZN(n4536) );
  XOR2_X1 U2644 ( .A(n4052), .B(n4055), .Z(n4422) );
  OAI21_X1 U2645 ( .B1(n4063), .B2(n4057), .A(n4055), .ZN(n4426) );
  AND2_X1 U2646 ( .A1(n2896), .A2(n2895), .ZN(n3102) );
  NAND2_X1 U2647 ( .A1(n2369), .A2(IR_REG_31__SCAN_IN), .ZN(n2370) );
  INV_X1 U2648 ( .A(IR_REG_19__SCAN_IN), .ZN(n2337) );
  XNOR2_X1 U2649 ( .A(n2279), .B(IR_REG_8__SCAN_IN), .ZN(n4491) );
  XNOR2_X1 U2650 ( .A(n2261), .B(IR_REG_3__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U2652 ( .A1(n2121), .A2(n2038), .ZN(n2120) );
  NAND2_X1 U2653 ( .A1(n2063), .A2(n4592), .ZN(n3058) );
  NAND2_X1 U2654 ( .A1(n2063), .A2(n4586), .ZN(n3065) );
  AND4_X2 U2655 ( .A1(n2189), .A2(n2188), .A3(n2187), .A4(n2186), .ZN(n1998)
         );
  NAND2_X1 U2656 ( .A1(n2024), .A2(n2153), .ZN(n2161) );
  NOR2_X1 U2657 ( .A1(n2654), .A2(n3614), .ZN(n1999) );
  AND2_X1 U2658 ( .A1(n2839), .A2(n2031), .ZN(n2000) );
  AND2_X1 U2659 ( .A1(n2185), .A2(n3049), .ZN(n2001) );
  OR2_X1 U2660 ( .A1(n2470), .A2(n2469), .ZN(n2002) );
  OR2_X1 U2661 ( .A1(n1999), .A2(n3684), .ZN(n2003) );
  INV_X1 U2662 ( .A(n2202), .ZN(n2198) );
  NOR2_X1 U2663 ( .A1(n2206), .A2(n2203), .ZN(n2202) );
  AND2_X1 U2664 ( .A1(n2151), .A2(n4060), .ZN(n2004) );
  AND3_X1 U2665 ( .A1(n2983), .A2(n2141), .A3(n4142), .ZN(n2005) );
  OR2_X1 U2666 ( .A1(n3674), .A2(n3048), .ZN(n2006) );
  AOI21_X1 U2667 ( .B1(n3112), .B2(REG2_REG_3__SCAN_IN), .A(n2260), .ZN(n2264)
         );
  INV_X1 U2668 ( .A(IR_REG_31__SCAN_IN), .ZN(n2258) );
  NAND2_X1 U2669 ( .A1(n2131), .A2(n2130), .ZN(n3600) );
  AND2_X1 U2670 ( .A1(n2197), .A2(n2200), .ZN(n2007) );
  XNOR2_X1 U2671 ( .A(n2466), .B(n2850), .ZN(n2469) );
  NAND2_X1 U2672 ( .A1(n3150), .A2(REG2_REG_7__SCAN_IN), .ZN(n2008) );
  AND2_X1 U2673 ( .A1(n3711), .A2(n2709), .ZN(n2708) );
  INV_X1 U2674 ( .A(n4060), .ZN(n2083) );
  OR2_X1 U2675 ( .A1(n4117), .A2(n4112), .ZN(n2009) );
  INV_X1 U2676 ( .A(n3466), .ZN(n2184) );
  INV_X1 U2677 ( .A(n3426), .ZN(n2185) );
  AND2_X1 U2678 ( .A1(n2001), .A2(n2184), .ZN(n2010) );
  AND2_X1 U2679 ( .A1(n4490), .A2(n2291), .ZN(n2011) );
  NOR2_X1 U2680 ( .A1(n4064), .A2(n4071), .ZN(n4063) );
  INV_X1 U2681 ( .A(IR_REG_30__SCAN_IN), .ZN(n4594) );
  OR2_X1 U2682 ( .A1(n3325), .A2(n3630), .ZN(n2012) );
  AND2_X1 U2683 ( .A1(n3079), .A2(REG2_REG_1__SCAN_IN), .ZN(n2013) );
  NOR3_X1 U2684 ( .A1(n4117), .A2(n4100), .A3(n4112), .ZN(n2014) );
  AND2_X1 U2685 ( .A1(n3343), .A2(n2513), .ZN(n2015) );
  NAND2_X1 U2686 ( .A1(n4492), .A2(REG2_REG_5__SCAN_IN), .ZN(n2016) );
  NAND2_X1 U2687 ( .A1(n3900), .A2(n3896), .ZN(n3867) );
  NAND2_X1 U2688 ( .A1(n4492), .A2(REG1_REG_5__SCAN_IN), .ZN(n2017) );
  INV_X1 U2689 ( .A(n3843), .ZN(n2084) );
  AND2_X1 U2690 ( .A1(n2092), .A2(n2008), .ZN(n2018) );
  INV_X1 U2691 ( .A(n3950), .ZN(n2076) );
  AND2_X1 U2692 ( .A1(n2648), .A2(n2649), .ZN(n3684) );
  NAND2_X1 U2693 ( .A1(n4506), .A2(n2172), .ZN(n2019) );
  AND2_X1 U2694 ( .A1(n3807), .A2(n3808), .ZN(n3859) );
  OR2_X1 U2695 ( .A1(n2619), .A2(n3657), .ZN(n2020) );
  OR2_X1 U2696 ( .A1(n3212), .A2(n1996), .ZN(n2021) );
  AND2_X1 U2697 ( .A1(n2968), .A2(n3637), .ZN(n2022) );
  NAND2_X1 U2698 ( .A1(n2720), .A2(n3728), .ZN(n2023) );
  INV_X1 U2699 ( .A(n2147), .ZN(n2146) );
  NAND2_X1 U2700 ( .A1(n4060), .A2(n2148), .ZN(n2147) );
  NAND2_X1 U2701 ( .A1(n2087), .A2(n3937), .ZN(n4244) );
  AND2_X1 U2702 ( .A1(n2289), .A2(n2293), .ZN(n2587) );
  AND2_X1 U2703 ( .A1(n2154), .A2(n2017), .ZN(n2024) );
  INV_X1 U2704 ( .A(n2151), .ZN(n2150) );
  NOR2_X1 U2705 ( .A1(n4116), .A2(n3630), .ZN(n2151) );
  NAND2_X1 U2706 ( .A1(n2136), .A2(n2135), .ZN(n4222) );
  AND2_X1 U2707 ( .A1(n2085), .A2(n2084), .ZN(n4092) );
  AND2_X1 U2708 ( .A1(n3927), .A2(n2054), .ZN(n2025) );
  INV_X1 U2709 ( .A(n2990), .ZN(n2143) );
  AND2_X1 U2710 ( .A1(n2169), .A2(REG1_REG_8__SCAN_IN), .ZN(n2026) );
  AND2_X1 U2711 ( .A1(n2355), .A2(n2354), .ZN(n2027) );
  AND2_X1 U2712 ( .A1(n2708), .A2(n2200), .ZN(n2196) );
  NAND2_X1 U2713 ( .A1(n2567), .A2(n2249), .ZN(n3432) );
  NAND2_X1 U2714 ( .A1(n3550), .A2(n2181), .ZN(n3601) );
  INV_X1 U2715 ( .A(n3749), .ZN(n2226) );
  NAND2_X1 U2716 ( .A1(n4298), .A2(n4278), .ZN(n4262) );
  NAND2_X1 U2717 ( .A1(n2184), .A2(n3984), .ZN(n2028) );
  AOI21_X1 U2718 ( .B1(n3524), .B2(REG2_REG_12__SCAN_IN), .A(n2305), .ZN(n4004) );
  INV_X1 U2719 ( .A(n3919), .ZN(n2065) );
  INV_X1 U2720 ( .A(n3905), .ZN(n2072) );
  INV_X1 U2721 ( .A(n3918), .ZN(n2068) );
  INV_X1 U2722 ( .A(n3925), .ZN(n2057) );
  NAND2_X1 U2723 ( .A1(n3455), .A2(n3454), .ZN(n3453) );
  NOR2_X1 U2724 ( .A1(n3502), .A2(n3517), .ZN(n3516) );
  AND2_X1 U2725 ( .A1(n3412), .A2(n2165), .ZN(n2029) );
  AND2_X1 U2726 ( .A1(n2134), .A2(n2132), .ZN(n2030) );
  NAND2_X1 U2727 ( .A1(n2854), .A2(n2853), .ZN(n2031) );
  NOR2_X1 U2728 ( .A1(n4273), .A2(n4263), .ZN(n2032) );
  AND2_X1 U2729 ( .A1(n3516), .A2(n3051), .ZN(n3550) );
  INV_X1 U2730 ( .A(n3071), .ZN(n2228) );
  NAND2_X1 U2731 ( .A1(n2587), .A2(REG2_REG_9__SCAN_IN), .ZN(n2291) );
  INV_X1 U2732 ( .A(n2291), .ZN(n2117) );
  AND2_X1 U2733 ( .A1(n3050), .A2(n2010), .ZN(n2033) );
  NOR2_X1 U2734 ( .A1(n3363), .A2(n3364), .ZN(n3294) );
  AND2_X1 U2735 ( .A1(n3250), .A2(n3273), .ZN(n3248) );
  XNOR2_X1 U2736 ( .A(n2264), .B(n3083), .ZN(n3162) );
  XNOR2_X1 U2737 ( .A(n2280), .B(n4491), .ZN(n3225) );
  XNOR2_X1 U2738 ( .A(n2273), .B(n3088), .ZN(n3143) );
  AND3_X1 U2739 ( .A1(n2944), .A2(n2943), .A3(n2942), .ZN(n3251) );
  NOR2_X1 U2740 ( .A1(n3228), .A2(n2388), .ZN(n2034) );
  NAND2_X1 U2741 ( .A1(n2153), .A2(n2154), .ZN(n2035) );
  AND2_X1 U2742 ( .A1(n2121), .A2(n2119), .ZN(n2036) );
  AND2_X1 U2743 ( .A1(n2091), .A2(n2090), .ZN(n2037) );
  INV_X1 U2744 ( .A(n2173), .ZN(n2172) );
  OR2_X1 U2745 ( .A1(n4515), .A2(n2174), .ZN(n2173) );
  XNOR2_X1 U2746 ( .A(n2263), .B(IR_REG_4__SCAN_IN), .ZN(n3083) );
  INV_X1 U2747 ( .A(n3083), .ZN(n2156) );
  INV_X1 U2748 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2159) );
  XNOR2_X1 U2749 ( .A(n2272), .B(IR_REG_6__SCAN_IN), .ZN(n3088) );
  INV_X1 U2750 ( .A(n3088), .ZN(n2160) );
  INV_X1 U2751 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2110) );
  OR2_X1 U2752 ( .A1(n2339), .A2(n2335), .ZN(n2038) );
  INV_X1 U2753 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2166) );
  NAND4_X1 U2754 ( .A1(REG3_REG_6__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .A4(REG3_REG_3__SCAN_IN), .ZN(n2553) );
  INV_X1 U2755 ( .A(n4148), .ZN(n3034) );
  NAND2_X1 U2756 ( .A1(n2049), .A2(n3816), .ZN(n2048) );
  NAND2_X1 U2757 ( .A1(n4165), .A2(n3945), .ZN(n2049) );
  OAI21_X1 U2758 ( .B1(n3459), .B2(n2059), .A(n2056), .ZN(n3508) );
  NAND2_X1 U2759 ( .A1(n2055), .A2(n2025), .ZN(n3017) );
  NAND2_X1 U2760 ( .A1(n3459), .A2(n2056), .ZN(n2055) );
  OAI21_X1 U2761 ( .B1(n3459), .B2(n2062), .A(n3915), .ZN(n3495) );
  AOI21_X1 U2762 ( .B1(n2062), .B2(n3915), .A(n2061), .ZN(n2060) );
  OAI21_X1 U2763 ( .B1(n3003), .B2(n2070), .A(n2067), .ZN(n3287) );
  NAND2_X1 U2764 ( .A1(n2066), .A2(n2064), .ZN(n3005) );
  AOI21_X1 U2765 ( .B1(n2067), .B2(n2070), .A(n2065), .ZN(n2064) );
  NAND2_X1 U2766 ( .A1(n3003), .A2(n2067), .ZN(n2066) );
  NAND2_X1 U2767 ( .A1(n4127), .A2(n3950), .ZN(n4108) );
  NAND2_X1 U2768 ( .A1(n2087), .A2(n2086), .ZN(n4224) );
  NAND2_X1 U2769 ( .A1(n3162), .A2(n2099), .ZN(n2094) );
  NAND2_X1 U2770 ( .A1(n2097), .A2(n2094), .ZN(n3131) );
  INV_X1 U2771 ( .A(n2264), .ZN(n2101) );
  NOR2_X2 U2772 ( .A1(n3998), .A2(n3997), .ZN(n3996) );
  MUX2_X1 U2773 ( .A(n2253), .B(REG2_REG_1__SCAN_IN), .S(n3079), .Z(n3120) );
  NAND2_X1 U2774 ( .A1(n2104), .A2(n2103), .ZN(n4503) );
  NAND2_X1 U2775 ( .A1(n4042), .A2(n2325), .ZN(n2103) );
  NAND2_X1 U2776 ( .A1(n3369), .A2(n2109), .ZN(n2107) );
  OAI211_X1 U2777 ( .C1(n3369), .C2(n2111), .A(n2107), .B(n2108), .ZN(n2299)
         );
  OAI211_X1 U2778 ( .C1(n3369), .C2(n4490), .A(n2112), .B(n2116), .ZN(n3410)
         );
  NAND2_X1 U2779 ( .A1(n3369), .A2(n2011), .ZN(n2112) );
  INV_X1 U2780 ( .A(n2116), .ZN(n2114) );
  INV_X1 U2781 ( .A(n2299), .ZN(n3448) );
  NAND2_X1 U2782 ( .A1(n4523), .A2(n2036), .ZN(n2118) );
  OAI211_X1 U2783 ( .C1(n4523), .C2(n2120), .A(n2118), .B(n2122), .ZN(U3259)
         );
  AND2_X1 U2784 ( .A1(n2408), .A2(n2407), .ZN(n2122) );
  NAND3_X1 U2785 ( .A1(n2126), .A2(n2946), .A3(n3340), .ZN(n2125) );
  NAND2_X1 U2786 ( .A1(n2946), .A2(n3340), .ZN(n2127) );
  NAND3_X1 U2787 ( .A1(n2125), .A2(n2123), .A3(n2952), .ZN(n3423) );
  NAND2_X1 U2788 ( .A1(n2124), .A2(n2126), .ZN(n2123) );
  INV_X1 U2789 ( .A(n2948), .ZN(n2124) );
  NAND2_X1 U2790 ( .A1(n2127), .A2(n2948), .ZN(n3291) );
  NAND4_X1 U2791 ( .A1(n2344), .A2(n2345), .A3(n2343), .A4(n2342), .ZN(n2356)
         );
  AND2_X2 U2792 ( .A1(n1998), .A2(n2313), .ZN(n2357) );
  NAND4_X1 U2793 ( .A1(n2129), .A2(n2027), .A3(n1998), .A4(n2313), .ZN(n2128)
         );
  AND4_X2 U2794 ( .A1(n2193), .A2(n2192), .A3(n2190), .A4(n2191), .ZN(n2313)
         );
  NAND2_X1 U2795 ( .A1(n3570), .A2(n2132), .ZN(n2131) );
  NAND2_X1 U2796 ( .A1(n2977), .A2(n2137), .ZN(n2136) );
  NAND2_X1 U2797 ( .A1(n2980), .A2(n3851), .ZN(n4204) );
  NAND2_X1 U2798 ( .A1(n3230), .A2(n2026), .ZN(n2168) );
  INV_X1 U2799 ( .A(n3374), .ZN(n2169) );
  OAI21_X1 U2800 ( .B1(n4507), .B2(n2173), .A(n2170), .ZN(n2175) );
  NAND2_X1 U2801 ( .A1(n4507), .A2(n4508), .ZN(n4506) );
  INV_X1 U2802 ( .A(n2175), .ZN(n2400) );
  INV_X2 U2803 ( .A(n2634), .ZN(n3828) );
  NAND2_X1 U2804 ( .A1(n2634), .A2(IR_REG_0__SCAN_IN), .ZN(n2449) );
  AND2_X4 U2805 ( .A1(n2176), .A2(n2360), .ZN(n2634) );
  NAND2_X2 U2806 ( .A1(n2177), .A2(IR_REG_31__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U2807 ( .A1(n2245), .A2(n2178), .ZN(n4064) );
  NAND2_X1 U2808 ( .A1(n2245), .A2(n4136), .ZN(n4117) );
  NAND2_X1 U2809 ( .A1(n3050), .A2(n2183), .ZN(n3502) );
  NOR2_X2 U2810 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2191)
         );
  NOR2_X1 U2811 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2193)
         );
  NAND2_X1 U2812 ( .A1(n2647), .A2(n2196), .ZN(n2194) );
  NAND2_X1 U2813 ( .A1(n2567), .A2(n2208), .ZN(n2207) );
  INV_X1 U2814 ( .A(n2212), .ZN(n3478) );
  NAND2_X1 U2815 ( .A1(n2210), .A2(n3475), .ZN(n2633) );
  NAND2_X1 U2816 ( .A1(n2212), .A2(n2211), .ZN(n2210) );
  INV_X1 U2817 ( .A(n3476), .ZN(n2211) );
  NAND2_X1 U2818 ( .A1(n3697), .A2(n2250), .ZN(n2222) );
  NAND2_X1 U2819 ( .A1(n3697), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2820 ( .A1(n2222), .A2(n2839), .ZN(n3782) );
  NAND3_X1 U2821 ( .A1(n2521), .A2(n2506), .A3(n2223), .ZN(n3329) );
  OAI21_X1 U2822 ( .B1(n3070), .B2(n2225), .A(n2224), .ZN(n3759) );
  AND2_X1 U2823 ( .A1(n2234), .A2(n3279), .ZN(n2233) );
  NAND2_X1 U2824 ( .A1(n3280), .A2(n3279), .ZN(n3278) );
  NAND2_X1 U2825 ( .A1(n2234), .A2(n2231), .ZN(n2230) );
  NAND2_X1 U2826 ( .A1(n3280), .A2(n2233), .ZN(n2232) );
  OR2_X2 U2827 ( .A1(n3769), .A2(n2736), .ZN(n2737) );
  AND2_X1 U2828 ( .A1(n3969), .A2(n3962), .ZN(n4530) );
  OR2_X1 U2829 ( .A1(n3189), .A2(n3962), .ZN(n4253) );
  AND2_X2 U2830 ( .A1(n2424), .A2(n2432), .ZN(n2473) );
  NAND2_X1 U2831 ( .A1(n2473), .A2(REG0_REG_1__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U2832 ( .A1(n2454), .A2(n3962), .ZN(n2437) );
  NAND2_X1 U2833 ( .A1(n3190), .A2(n3674), .ZN(n3897) );
  NAND2_X1 U2834 ( .A1(n3992), .A2(n2480), .ZN(n2451) );
  OR2_X1 U2835 ( .A1(n2392), .A2(n4413), .ZN(n2236) );
  AND2_X2 U2836 ( .A1(n3060), .A2(n3239), .ZN(n4586) );
  AND2_X1 U2837 ( .A1(n2379), .A2(REG1_REG_2__SCAN_IN), .ZN(n2237) );
  OR2_X1 U2838 ( .A1(n2675), .A2(REG1_REG_17__SCAN_IN), .ZN(n2238) );
  NOR2_X1 U2839 ( .A1(n4132), .A2(n4151), .ZN(n2241) );
  NAND2_X1 U2840 ( .A1(n4094), .A2(n4112), .ZN(n2242) );
  NOR2_X1 U2841 ( .A1(n2971), .A2(n4322), .ZN(n2243) );
  AND2_X1 U2842 ( .A1(n2379), .A2(REG2_REG_2__SCAN_IN), .ZN(n2244) );
  INV_X1 U2843 ( .A(n4341), .ZN(n4069) );
  NAND2_X1 U2844 ( .A1(n2487), .A2(n2486), .ZN(n3180) );
  AND2_X2 U2845 ( .A1(n4155), .A2(n4157), .ZN(n2245) );
  INV_X1 U2846 ( .A(n3893), .ZN(n3000) );
  AND3_X1 U2847 ( .A1(n2909), .A2(n3773), .A3(n2908), .ZN(n2246) );
  INV_X1 U2848 ( .A(n3630), .ZN(n4100) );
  INV_X1 U2849 ( .A(n3753), .ZN(n4234) );
  NOR2_X1 U2850 ( .A1(n2986), .A2(n4145), .ZN(n2247) );
  AND2_X1 U2851 ( .A1(n2594), .A2(n2582), .ZN(n2248) );
  OR2_X1 U2852 ( .A1(n2566), .A2(n2565), .ZN(n2249) );
  AND2_X2 U2853 ( .A1(n3060), .A2(n3059), .ZN(n4592) );
  INV_X1 U2854 ( .A(n3549), .ZN(n3051) );
  AND2_X1 U2855 ( .A1(n3698), .A2(n2833), .ZN(n2250) );
  NAND2_X1 U2856 ( .A1(n2633), .A2(n2632), .ZN(n3682) );
  INV_X1 U2857 ( .A(n4491), .ZN(n2386) );
  AND2_X1 U2858 ( .A1(n2587), .A2(REG1_REG_9__SCAN_IN), .ZN(n2251) );
  NAND2_X1 U2859 ( .A1(n2302), .A2(n2296), .ZN(n4489) );
  INV_X1 U2860 ( .A(n4489), .ZN(n2300) );
  INV_X1 U2861 ( .A(n4014), .ZN(n2375) );
  INV_X1 U2862 ( .A(n3388), .ZN(n2949) );
  OR2_X1 U2863 ( .A1(n3023), .A2(n4245), .ZN(n3940) );
  AND2_X1 U2864 ( .A1(n4169), .A2(n4167), .ZN(n3945) );
  AND2_X1 U2865 ( .A1(n4223), .A2(n3028), .ZN(n3939) );
  AND2_X1 U2866 ( .A1(n3194), .A2(n2941), .ZN(n2939) );
  AND2_X1 U2867 ( .A1(n3887), .A2(n4126), .ZN(n3950) );
  INV_X1 U2868 ( .A(IR_REG_0__SCAN_IN), .ZN(n2447) );
  AND2_X1 U2869 ( .A1(n3844), .A2(n4107), .ZN(n3951) );
  INV_X1 U2870 ( .A(n2755), .ZN(n2754) );
  INV_X1 U2871 ( .A(n3982), .ZN(n3543) );
  INV_X1 U2872 ( .A(n2437), .ZN(n2996) );
  AOI21_X1 U2873 ( .B1(n3600), .B2(n2972), .A(n2243), .ZN(n4304) );
  AND3_X1 U2874 ( .A1(n4596), .A2(n2416), .A3(n2415), .ZN(n2417) );
  INV_X1 U2875 ( .A(n2553), .ZN(n2426) );
  INV_X1 U2876 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2568) );
  INV_X1 U2877 ( .A(n2623), .ZN(n2427) );
  AND2_X1 U2878 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  NAND2_X1 U2879 ( .A1(n2807), .A2(REG3_REG_25__SCAN_IN), .ZN(n2840) );
  INV_X1 U2880 ( .A(n3823), .ZN(n2874) );
  INV_X1 U2881 ( .A(n2331), .ZN(n2332) );
  INV_X1 U2882 ( .A(n4157), .ZN(n4151) );
  OR2_X1 U2883 ( .A1(n4208), .A2(n4199), .ZN(n4169) );
  NAND2_X1 U2884 ( .A1(n3272), .A2(n3219), .ZN(n3896) );
  OR2_X1 U2885 ( .A1(n4299), .A2(n4327), .ZN(n3052) );
  INV_X1 U2886 ( .A(n3311), .ZN(n3049) );
  INV_X1 U2887 ( .A(n4484), .ZN(n2997) );
  INV_X1 U2888 ( .A(IR_REG_5__SCAN_IN), .ZN(n2270) );
  NAND2_X1 U2889 ( .A1(n2426), .A2(REG3_REG_7__SCAN_IN), .ZN(n2569) );
  OR2_X1 U2890 ( .A1(n2594), .A2(n2593), .ZN(n2623) );
  OR2_X1 U2891 ( .A1(n2569), .A2(n2568), .ZN(n2581) );
  INV_X1 U2892 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U2893 ( .A1(n2427), .A2(REG3_REG_11__SCAN_IN), .ZN(n2636) );
  OR2_X1 U2894 ( .A1(n2840), .A2(n4668), .ZN(n2870) );
  OR2_X1 U2895 ( .A1(n4237), .A2(n2921), .ZN(n2761) );
  NAND2_X1 U2896 ( .A1(n2668), .A2(REG3_REG_15__SCAN_IN), .ZN(n2693) );
  AND2_X1 U2897 ( .A1(n2387), .A2(n4491), .ZN(n2388) );
  AND2_X1 U2898 ( .A1(n4169), .A2(n3031), .ZN(n4189) );
  OR2_X1 U2899 ( .A1(n3036), .A2(n3168), .ZN(n4275) );
  AND2_X1 U2900 ( .A1(n3967), .A2(n3035), .ZN(n4210) );
  INV_X1 U2901 ( .A(n2967), .ZN(n3637) );
  NAND2_X1 U2902 ( .A1(n3066), .A2(n3101), .ZN(n3040) );
  INV_X1 U2903 ( .A(n2933), .ZN(n2934) );
  NAND2_X1 U2904 ( .A1(n3329), .A2(n2524), .ZN(n3280) );
  INV_X1 U2905 ( .A(n3241), .ZN(n3969) );
  OR2_X1 U2906 ( .A1(n3703), .A2(n2921), .ZN(n2813) );
  XNOR2_X1 U2907 ( .A(n2380), .B(n4493), .ZN(n3111) );
  INV_X1 U2908 ( .A(n3368), .ZN(n3372) );
  INV_X1 U2909 ( .A(n4514), .ZN(n4510) );
  INV_X1 U2910 ( .A(n4210), .ZN(n4318) );
  INV_X1 U2911 ( .A(n3255), .ZN(n3273) );
  AND2_X1 U2912 ( .A1(n4288), .A2(n4575), .ZN(n4328) );
  AOI21_X1 U2913 ( .B1(n3097), .B2(n3103), .A(n3102), .ZN(n3059) );
  INV_X1 U2914 ( .A(n4578), .ZN(n4569) );
  NAND2_X1 U2915 ( .A1(n4232), .A2(n4558), .ZN(n4578) );
  AND3_X1 U2916 ( .A1(n3047), .A2(n3046), .A3(n3045), .ZN(n3060) );
  INV_X1 U2917 ( .A(n2889), .ZN(n2896) );
  INV_X1 U2918 ( .A(n3040), .ZN(n3235) );
  AND2_X1 U2919 ( .A1(n2319), .A2(n2321), .ZN(n4033) );
  OR2_X1 U2920 ( .A1(n2404), .A2(n2403), .ZN(n4031) );
  NOR2_X1 U2921 ( .A1(n2246), .A2(n2934), .ZN(n2935) );
  NAND2_X1 U2922 ( .A1(n2899), .A2(n2898), .ZN(n3805) );
  NAND2_X1 U2923 ( .A1(n2847), .A2(n2846), .ZN(n4094) );
  NAND2_X1 U2924 ( .A1(n2730), .A2(n2729), .ZN(n4293) );
  OR2_X1 U2925 ( .A1(n4497), .A2(n3971), .ZN(n4014) );
  AOI21_X1 U2926 ( .B1(n2019), .B2(n4522), .A(n4521), .ZN(n4528) );
  NAND2_X1 U2927 ( .A1(n4538), .A2(n3293), .ZN(n4285) );
  INV_X1 U2928 ( .A(n4328), .ZN(n4268) );
  NAND2_X1 U2929 ( .A1(n4592), .A2(n4575), .ZN(n4418) );
  INV_X1 U2930 ( .A(n4592), .ZN(n4590) );
  NAND2_X1 U2931 ( .A1(n4586), .A2(n4575), .ZN(n4478) );
  INV_X1 U2932 ( .A(n4586), .ZN(n4584) );
  INV_X1 U2933 ( .A(n4543), .ZN(n3101) );
  NAND2_X1 U2934 ( .A1(n3098), .A2(n3235), .ZN(n4593) );
  INV_X1 U2935 ( .A(n3991), .ZN(U4043) );
  INV_X2 U2936 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  XNOR2_X2 U2937 ( .A(n2252), .B(IR_REG_1__SCAN_IN), .ZN(n3079) );
  INV_X1 U2938 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2253) );
  INV_X1 U2939 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2254) );
  XNOR2_X2 U2940 ( .A(n2255), .B(IR_REG_2__SCAN_IN), .ZN(n2379) );
  MUX2_X1 U2941 ( .A(n3243), .B(REG2_REG_2__SCAN_IN), .S(n2379), .Z(n3997) );
  INV_X1 U2942 ( .A(IR_REG_2__SCAN_IN), .ZN(n2256) );
  NAND2_X1 U2943 ( .A1(n2257), .A2(n2256), .ZN(n2267) );
  NAND2_X1 U2944 ( .A1(n2267), .A2(IR_REG_31__SCAN_IN), .ZN(n2261) );
  NAND2_X1 U2945 ( .A1(n2261), .A2(n2265), .ZN(n2262) );
  NAND2_X1 U2946 ( .A1(n2262), .A2(IR_REG_31__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2947 ( .A1(n2265), .A2(n2312), .ZN(n2266) );
  NAND2_X1 U2948 ( .A1(n2269), .A2(IR_REG_31__SCAN_IN), .ZN(n2268) );
  MUX2_X1 U2949 ( .A(IR_REG_31__SCAN_IN), .B(n2268), .S(IR_REG_5__SCAN_IN), 
        .Z(n2271) );
  NAND2_X1 U2950 ( .A1(n2271), .A2(n2275), .ZN(n3137) );
  MUX2_X1 U2951 ( .A(REG2_REG_5__SCAN_IN), .B(n3362), .S(n3137), .Z(n3132) );
  INV_X1 U2952 ( .A(n3137), .ZN(n4492) );
  NAND2_X1 U2953 ( .A1(n2275), .A2(IR_REG_31__SCAN_IN), .ZN(n2272) );
  INV_X1 U2954 ( .A(n2273), .ZN(n2274) );
  INV_X1 U2955 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U2956 ( .A1(n2284), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  MUX2_X1 U2957 ( .A(n3315), .B(REG2_REG_7__SCAN_IN), .S(n3150), .Z(n3155) );
  INV_X1 U2958 ( .A(IR_REG_7__SCAN_IN), .ZN(n2276) );
  NAND2_X1 U2959 ( .A1(n2277), .A2(n2276), .ZN(n2278) );
  NAND2_X1 U2960 ( .A1(n2278), .A2(IR_REG_31__SCAN_IN), .ZN(n2279) );
  NAND2_X1 U2961 ( .A1(n3225), .A2(REG2_REG_8__SCAN_IN), .ZN(n2283) );
  INV_X1 U2962 ( .A(n2280), .ZN(n2281) );
  NAND2_X1 U2963 ( .A1(n2281), .A2(n4491), .ZN(n2282) );
  NAND2_X1 U2964 ( .A1(n2283), .A2(n2282), .ZN(n3368) );
  INV_X1 U2965 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4624) );
  INV_X1 U2966 ( .A(n2284), .ZN(n2286) );
  NOR2_X1 U2967 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2285)
         );
  NAND2_X1 U2968 ( .A1(n2286), .A2(n2285), .ZN(n2288) );
  NAND2_X1 U2969 ( .A1(n2288), .A2(IR_REG_31__SCAN_IN), .ZN(n2287) );
  MUX2_X1 U2970 ( .A(IR_REG_31__SCAN_IN), .B(n2287), .S(IR_REG_9__SCAN_IN), 
        .Z(n2289) );
  MUX2_X1 U2971 ( .A(n4624), .B(REG2_REG_9__SCAN_IN), .S(n2587), .Z(n3371) );
  NAND2_X1 U2972 ( .A1(n3368), .A2(n2290), .ZN(n3369) );
  INV_X1 U2973 ( .A(n2587), .ZN(n3376) );
  NAND2_X1 U2974 ( .A1(n2293), .A2(IR_REG_31__SCAN_IN), .ZN(n2292) );
  INV_X1 U2975 ( .A(n4490), .ZN(n3412) );
  INV_X1 U2976 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2297) );
  NAND2_X1 U2977 ( .A1(n2295), .A2(n2294), .ZN(n2302) );
  OR2_X1 U2978 ( .A1(n2295), .A2(n2294), .ZN(n2296) );
  MUX2_X1 U2979 ( .A(REG2_REG_11__SCAN_IN), .B(n2297), .S(n4489), .Z(n3447) );
  NAND2_X1 U2980 ( .A1(n2299), .A2(n2298), .ZN(n3451) );
  NAND2_X1 U2981 ( .A1(n2302), .A2(IR_REG_31__SCAN_IN), .ZN(n2303) );
  XNOR2_X1 U2982 ( .A(n2303), .B(IR_REG_12__SCAN_IN), .ZN(n2635) );
  INV_X1 U2983 ( .A(n2635), .ZN(n3526) );
  NAND2_X1 U2984 ( .A1(n2306), .A2(n2313), .ZN(n2310) );
  NAND2_X1 U2985 ( .A1(n2310), .A2(IR_REG_31__SCAN_IN), .ZN(n2307) );
  XNOR2_X1 U2986 ( .A(n2307), .B(IR_REG_13__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U2987 ( .A1(n4488), .A2(REG2_REG_13__SCAN_IN), .ZN(n2309) );
  NOR2_X1 U2988 ( .A1(n4488), .A2(REG2_REG_13__SCAN_IN), .ZN(n2308) );
  OAI21_X1 U2989 ( .B1(n2310), .B2(IR_REG_13__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2311) );
  MUX2_X1 U2990 ( .A(IR_REG_31__SCAN_IN), .B(n2311), .S(IR_REG_14__SCAN_IN), 
        .Z(n2314) );
  INV_X1 U2991 ( .A(n2357), .ZN(n2346) );
  AND2_X1 U2992 ( .A1(n2314), .A2(n2346), .ZN(n4487) );
  INV_X1 U2993 ( .A(n4487), .ZN(n4019) );
  XNOR2_X1 U2994 ( .A(n2315), .B(n4019), .ZN(n4017) );
  NAND2_X1 U2995 ( .A1(n4017), .A2(REG2_REG_14__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U2996 ( .A1(n2315), .A2(n4487), .ZN(n2316) );
  NAND2_X1 U2997 ( .A1(n4016), .A2(n2316), .ZN(n4029) );
  NAND2_X1 U2998 ( .A1(n2346), .A2(IR_REG_31__SCAN_IN), .ZN(n2318) );
  INV_X1 U2999 ( .A(n2318), .ZN(n2317) );
  NAND2_X1 U3000 ( .A1(n2317), .A2(IR_REG_15__SCAN_IN), .ZN(n2319) );
  INV_X1 U3001 ( .A(IR_REG_15__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U3002 ( .A1(n2318), .A2(n4604), .ZN(n2321) );
  XOR2_X1 U3003 ( .A(REG2_REG_15__SCAN_IN), .B(n4033), .Z(n4028) );
  NAND2_X1 U3004 ( .A1(n4029), .A2(n4028), .ZN(n4027) );
  NAND2_X1 U3005 ( .A1(n4033), .A2(REG2_REG_15__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U3006 ( .A1(n4027), .A2(n2320), .ZN(n2324) );
  NAND2_X1 U3007 ( .A1(n2321), .A2(IR_REG_31__SCAN_IN), .ZN(n2322) );
  XNOR2_X1 U3008 ( .A(n2322), .B(IR_REG_16__SCAN_IN), .ZN(n4486) );
  XNOR2_X1 U3009 ( .A(n2324), .B(n4486), .ZN(n4042) );
  INV_X1 U3010 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2323) );
  OR2_X1 U3011 ( .A1(n2324), .A2(n4486), .ZN(n2325) );
  NOR2_X2 U3012 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2345)
         );
  NAND2_X1 U3013 ( .A1(n2357), .A2(n2345), .ZN(n2327) );
  NAND2_X1 U3014 ( .A1(n2327), .A2(IR_REG_31__SCAN_IN), .ZN(n2326) );
  MUX2_X1 U3015 ( .A(IR_REG_31__SCAN_IN), .B(n2326), .S(IR_REG_17__SCAN_IN), 
        .Z(n2330) );
  INV_X1 U3016 ( .A(n2327), .ZN(n2329) );
  NAND2_X1 U3017 ( .A1(n2329), .A2(n2328), .ZN(n2336) );
  NAND2_X1 U3018 ( .A1(n2330), .A2(n2336), .ZN(n4548) );
  NOR2_X1 U3019 ( .A1(n2675), .A2(REG2_REG_17__SCAN_IN), .ZN(n2331) );
  AOI21_X1 U3020 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2675), .A(n2331), .ZN(n4505) );
  NAND2_X1 U3021 ( .A1(n4503), .A2(n2332), .ZN(n4524) );
  NAND2_X1 U3022 ( .A1(n2336), .A2(IR_REG_31__SCAN_IN), .ZN(n2333) );
  XNOR2_X1 U3023 ( .A(n2333), .B(IR_REG_18__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U3024 ( .A1(REG2_REG_18__SCAN_IN), .A2(n2731), .ZN(n2334) );
  OAI21_X1 U3025 ( .B1(REG2_REG_18__SCAN_IN), .B2(n2731), .A(n2334), .ZN(n4525) );
  NOR2_X2 U3026 ( .A1(n4524), .A2(n4525), .ZN(n4523) );
  AND2_X1 U3027 ( .A1(n2731), .A2(REG2_REG_18__SCAN_IN), .ZN(n2335) );
  INV_X1 U3028 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4627) );
  NOR2_X2 U3029 ( .A1(n2336), .A2(IR_REG_18__SCAN_IN), .ZN(n2340) );
  INV_X1 U3030 ( .A(n2340), .ZN(n2412) );
  NAND2_X1 U3031 ( .A1(n2412), .A2(IR_REG_31__SCAN_IN), .ZN(n2338) );
  MUX2_X1 U3032 ( .A(n4627), .B(REG2_REG_19__SCAN_IN), .S(n3241), .Z(n2339) );
  NAND2_X1 U3033 ( .A1(n2340), .A2(n2344), .ZN(n2413) );
  XNOR2_X2 U3034 ( .A(n2341), .B(IR_REG_21__SCAN_IN), .ZN(n2454) );
  OR2_X1 U3035 ( .A1(n2349), .A2(n2258), .ZN(n2347) );
  NAND2_X1 U3036 ( .A1(n2454), .A2(n4484), .ZN(n3036) );
  INV_X1 U3037 ( .A(IR_REG_22__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3038 ( .A1(n2349), .A2(n2348), .ZN(n2365) );
  INV_X2 U3039 ( .A(IR_REG_23__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3040 ( .A1(n2350), .A2(n2352), .ZN(n2362) );
  OR2_X1 U3041 ( .A1(n2350), .A2(n2352), .ZN(n2351) );
  NAND2_X1 U3042 ( .A1(n2362), .A2(n2351), .ZN(n2917) );
  INV_X1 U3043 ( .A(n2917), .ZN(n2371) );
  OR2_X1 U3044 ( .A1(n3036), .A2(n2371), .ZN(n2361) );
  NAND2_X1 U3045 ( .A1(n2372), .A2(n2416), .ZN(n2358) );
  NAND2_X1 U3046 ( .A1(n2416), .A2(IR_REG_27__SCAN_IN), .ZN(n2360) );
  INV_X2 U3047 ( .A(n2634), .ZN(n3821) );
  AND2_X1 U3048 ( .A1(n2361), .A2(n3821), .ZN(n2404) );
  OAI21_X1 U3049 ( .B1(n2365), .B2(n2364), .A(IR_REG_31__SCAN_IN), .ZN(n2366)
         );
  MUX2_X1 U3050 ( .A(IR_REG_31__SCAN_IN), .B(n2366), .S(IR_REG_25__SCAN_IN), 
        .Z(n2368) );
  INV_X1 U3051 ( .A(n2367), .ZN(n2369) );
  NAND3_X2 U3052 ( .A1(n2889), .A2(n4483), .A3(n4482), .ZN(n3066) );
  NAND2_X1 U3053 ( .A1(n2917), .A2(STATE_REG_SCAN_IN), .ZN(n4543) );
  NAND2_X1 U3054 ( .A1(n2371), .A2(STATE_REG_SCAN_IN), .ZN(n3975) );
  NAND2_X1 U3055 ( .A1(n3040), .A2(n3975), .ZN(n2402) );
  NAND2_X1 U3056 ( .A1(n2404), .A2(n2402), .ZN(n4497) );
  XNOR2_X1 U3057 ( .A(n2372), .B(IR_REG_27__SCAN_IN), .ZN(n4495) );
  INV_X1 U3058 ( .A(n4495), .ZN(n3167) );
  NAND2_X1 U3059 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3060 ( .A1(n2372), .A2(n2373), .ZN(n2374) );
  XNOR2_X1 U3061 ( .A(n2374), .B(IR_REG_28__SCAN_IN), .ZN(n3168) );
  OR2_X1 U3062 ( .A1(n3167), .A2(n3168), .ZN(n3971) );
  INV_X1 U3063 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3561) );
  INV_X1 U3064 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3265) );
  INV_X1 U3065 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2376) );
  XNOR2_X1 U3066 ( .A(n3079), .B(n2376), .ZN(n3123) );
  AND2_X1 U3067 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2377)
         );
  NAND2_X1 U3068 ( .A1(n3123), .A2(n2377), .ZN(n3122) );
  NAND2_X1 U3069 ( .A1(n3079), .A2(REG1_REG_1__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3070 ( .A1(n3122), .A2(n2378), .ZN(n3993) );
  INV_X1 U3071 ( .A(n2380), .ZN(n2381) );
  INV_X1 U3072 ( .A(n2382), .ZN(n2383) );
  INV_X1 U3073 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4722) );
  MUX2_X1 U3074 ( .A(REG1_REG_5__SCAN_IN), .B(n4722), .S(n3137), .Z(n3134) );
  NAND2_X1 U3075 ( .A1(n3150), .A2(REG1_REG_7__SCAN_IN), .ZN(n2385) );
  INV_X1 U3076 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2384) );
  INV_X1 U3077 ( .A(n3150), .ZN(n3154) );
  XNOR2_X1 U3078 ( .A(n2587), .B(REG1_REG_9__SCAN_IN), .ZN(n3374) );
  XNOR2_X1 U3079 ( .A(n4489), .B(REG1_REG_11__SCAN_IN), .ZN(n3454) );
  INV_X1 U3080 ( .A(n2390), .ZN(n2391) );
  XOR2_X1 U3081 ( .A(REG1_REG_13__SCAN_IN), .B(n4488), .Z(n4010) );
  INV_X1 U3082 ( .A(n4488), .ZN(n2392) );
  INV_X1 U3083 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4413) );
  INV_X1 U3084 ( .A(n2393), .ZN(n2394) );
  XOR2_X1 U3085 ( .A(REG1_REG_15__SCAN_IN), .B(n4033), .Z(n4036) );
  NAND2_X1 U3086 ( .A1(n4037), .A2(n4036), .ZN(n4035) );
  INV_X1 U3087 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4405) );
  OR2_X1 U3088 ( .A1(n2396), .A2(n4486), .ZN(n2397) );
  INV_X1 U3089 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2671) );
  AOI22_X1 U3090 ( .A1(n2675), .A2(REG1_REG_17__SCAN_IN), .B1(n2671), .B2(
        n4548), .ZN(n4508) );
  INV_X1 U3091 ( .A(n2731), .ZN(n4546) );
  INV_X1 U3092 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2727) );
  AOI22_X1 U3093 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4546), .B1(n2731), .B2(
        n2727), .ZN(n4515) );
  AND2_X1 U3094 ( .A1(n2731), .A2(REG1_REG_18__SCAN_IN), .ZN(n2398) );
  XNOR2_X1 U3095 ( .A(n3241), .B(REG1_REG_19__SCAN_IN), .ZN(n2399) );
  XNOR2_X1 U3096 ( .A(n2400), .B(n2399), .ZN(n2401) );
  NAND2_X1 U3097 ( .A1(n2401), .A2(n4510), .ZN(n2408) );
  INV_X1 U3098 ( .A(n3168), .ZN(n4481) );
  NAND2_X1 U3099 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3669) );
  INV_X1 U3100 ( .A(n2402), .ZN(n2403) );
  NAND2_X1 U3101 ( .A1(n4517), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2405) );
  OAI211_X1 U3102 ( .C1(n4529), .C2(n3241), .A(n3669), .B(n2405), .ZN(n2406)
         );
  INV_X1 U3103 ( .A(n2406), .ZN(n2407) );
  AND2_X1 U3104 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2411)
         );
  NAND2_X1 U3105 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2409) );
  AOI22_X1 U3106 ( .A1(IR_REG_20__SCAN_IN), .A2(n2258), .B1(n2409), .B2(
        IR_REG_31__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3107 ( .A1(n2414), .A2(n2413), .ZN(n3962) );
  AND2_X4 U3108 ( .A1(n2996), .A2(n3066), .ZN(n2480) );
  NAND2_X1 U3109 ( .A1(n2420), .A2(IR_REG_31__SCAN_IN), .ZN(n2418) );
  INV_X1 U3110 ( .A(n2419), .ZN(n2421) );
  NOR2_X2 U3111 ( .A1(n2421), .A2(n3610), .ZN(n2425) );
  INV_X1 U3112 ( .A(n4480), .ZN(n2424) );
  AND2_X2 U3113 ( .A1(n2425), .A2(n2424), .ZN(n2472) );
  INV_X2 U3114 ( .A(n2472), .ZN(n2493) );
  INV_X4 U3115 ( .A(n2493), .ZN(n3822) );
  NAND2_X1 U3116 ( .A1(n3822), .A2(REG1_REG_13__SCAN_IN), .ZN(n2436) );
  INV_X1 U3117 ( .A(n2425), .ZN(n2432) );
  NAND2_X1 U3118 ( .A1(n3824), .A2(REG0_REG_13__SCAN_IN), .ZN(n2435) );
  INV_X1 U3119 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2429) );
  INV_X1 U3120 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2428) );
  OAI21_X1 U3121 ( .B1(n2636), .B2(n2429), .A(n2428), .ZN(n2431) );
  NAND2_X1 U3122 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2430) );
  AND2_X1 U3123 ( .A1(n2431), .A2(n2657), .ZN(n3621) );
  NAND2_X1 U3124 ( .A1(n2855), .A2(n3621), .ZN(n2434) );
  NAND2_X1 U3125 ( .A1(n3823), .A2(REG2_REG_13__SCAN_IN), .ZN(n2433) );
  NAND4_X1 U3126 ( .A1(n2436), .A2(n2435), .A3(n2434), .A4(n2433), .ZN(n3980)
         );
  NAND2_X1 U3127 ( .A1(n2480), .A2(n3980), .ZN(n2439) );
  AND2_X4 U3128 ( .A1(n2440), .A2(n3066), .ZN(n2471) );
  MUX2_X1 U3129 ( .A(n4488), .B(DATAI_13_), .S(n3821), .Z(n3010) );
  NAND2_X1 U3130 ( .A1(n2471), .A2(n3010), .ZN(n2438) );
  NAND2_X1 U3131 ( .A1(n2439), .A2(n2438), .ZN(n2441) );
  NAND2_X1 U3132 ( .A1(n3241), .A2(n4484), .ZN(n2910) );
  NAND2_X1 U3133 ( .A1(n2473), .A2(REG0_REG_0__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3134 ( .A1(n2474), .A2(REG3_REG_0__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3135 ( .A1(n2475), .A2(REG2_REG_0__SCAN_IN), .ZN(n2442) );
  NAND2_X1 U3136 ( .A1(n2472), .A2(REG1_REG_0__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3137 ( .A1(n2471), .A2(n3048), .ZN(n2450) );
  INV_X1 U3138 ( .A(n3066), .ZN(n2452) );
  NAND2_X1 U3139 ( .A1(n2452), .A2(REG1_REG_0__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3140 ( .A1(n2457), .A2(n2453), .ZN(n3164) );
  INV_X1 U3141 ( .A(n3992), .ZN(n2999) );
  INV_X1 U3142 ( .A(n2454), .ZN(n3874) );
  NAND2_X1 U3143 ( .A1(n3874), .A2(n2997), .ZN(n3189) );
  INV_X1 U3144 ( .A(n3962), .ZN(n4485) );
  NOR2_X1 U3145 ( .A1(n3066), .A2(n2447), .ZN(n2455) );
  AOI21_X1 U3146 ( .B1(n2480), .B2(n3048), .A(n2455), .ZN(n2456) );
  OAI21_X1 U3147 ( .B1(n2999), .B2(n2498), .A(n2456), .ZN(n3165) );
  NAND2_X1 U31480 ( .A1(n3164), .A2(n3165), .ZN(n2459) );
  NAND2_X1 U31490 ( .A1(n2457), .A2(n2850), .ZN(n2458) );
  NAND2_X1 U3150 ( .A1(n2459), .A2(n2458), .ZN(n3677) );
  NAND2_X1 U3151 ( .A1(n2472), .A2(REG1_REG_1__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3152 ( .A1(n2475), .A2(REG2_REG_1__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3153 ( .A1(n2474), .A2(REG3_REG_1__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3154 ( .A1(n2480), .A2(n2938), .ZN(n2465) );
  MUX2_X1 U3155 ( .A(DATAI_1_), .B(n3079), .S(n2634), .Z(n3674) );
  NAND2_X1 U3156 ( .A1(n2471), .A2(n3674), .ZN(n2464) );
  NAND2_X1 U3157 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  NAND2_X1 U3158 ( .A1(n2480), .A2(n3674), .ZN(n2467) );
  XNOR2_X1 U3159 ( .A(n2469), .B(n2468), .ZN(n3676) );
  NAND2_X1 U3160 ( .A1(n3677), .A2(n3676), .ZN(n3678) );
  INV_X1 U3161 ( .A(n2468), .ZN(n2470) );
  NAND2_X1 U3162 ( .A1(n3678), .A2(n2002), .ZN(n3179) );
  INV_X1 U3163 ( .A(n3179), .ZN(n2487) );
  MUX2_X1 U3164 ( .A(DATAI_2_), .B(n2379), .S(n2634), .Z(n3219) );
  NAND2_X1 U3165 ( .A1(n2471), .A2(n3219), .ZN(n2482) );
  NAND2_X1 U3166 ( .A1(n2472), .A2(REG1_REG_2__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3167 ( .A1(n2474), .A2(REG3_REG_2__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3168 ( .A1(n2475), .A2(REG2_REG_2__SCAN_IN), .ZN(n2476) );
  NAND4_X2 U3169 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n3198)
         );
  NAND2_X1 U3170 ( .A1(n2480), .A2(n3198), .ZN(n2481) );
  NAND2_X1 U3171 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  OR2_X1 U3172 ( .A1(n3272), .A2(n2498), .ZN(n2485) );
  NAND2_X1 U3173 ( .A1(n2480), .A2(n3219), .ZN(n2484) );
  NAND2_X1 U3174 ( .A1(n2485), .A2(n2484), .ZN(n2489) );
  XNOR2_X1 U3175 ( .A(n2488), .B(n2489), .ZN(n3182) );
  INV_X1 U3176 ( .A(n3182), .ZN(n2486) );
  INV_X1 U3177 ( .A(n2488), .ZN(n2491) );
  INV_X1 U3178 ( .A(n2489), .ZN(n2490) );
  NAND2_X1 U3179 ( .A1(n2491), .A2(n2490), .ZN(n2492) );
  NAND2_X1 U3180 ( .A1(n3180), .A2(n2492), .ZN(n3270) );
  NAND2_X1 U3181 ( .A1(n3822), .A2(REG1_REG_3__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3182 ( .A1(n2621), .A2(REG0_REG_3__SCAN_IN), .ZN(n2496) );
  INV_X1 U3183 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3184 ( .A1(n2855), .A2(n2507), .ZN(n2495) );
  NAND2_X1 U3185 ( .A1(n3823), .A2(REG2_REG_3__SCAN_IN), .ZN(n2494) );
  MUX2_X1 U3186 ( .A(n4493), .B(DATAI_3_), .S(n3828), .Z(n3255) );
  NAND2_X1 U3187 ( .A1(n2480), .A2(n3255), .ZN(n2499) );
  NAND2_X1 U3188 ( .A1(n2021), .A2(n2499), .ZN(n2503) );
  NAND2_X1 U3189 ( .A1(n2480), .A2(n3990), .ZN(n2501) );
  NAND2_X1 U3190 ( .A1(n2471), .A2(n3255), .ZN(n2500) );
  NAND2_X1 U3191 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  INV_X1 U3192 ( .A(n2503), .ZN(n2504) );
  NAND2_X1 U3193 ( .A1(n2505), .A2(n2504), .ZN(n2506) );
  NAND2_X1 U3194 ( .A1(n3822), .A2(REG1_REG_4__SCAN_IN), .ZN(n2512) );
  INV_X1 U3195 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3196 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  AND2_X1 U3197 ( .A1(n2509), .A2(n2541), .ZN(n3350) );
  NAND2_X1 U3198 ( .A1(n2855), .A2(n3350), .ZN(n2511) );
  NAND2_X1 U3199 ( .A1(n2621), .A2(REG0_REG_4__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U3200 ( .A1(n3823), .A2(REG2_REG_4__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U3201 ( .A1(n2480), .A2(n3989), .ZN(n2516) );
  MUX2_X1 U3202 ( .A(n3083), .B(DATAI_4_), .S(n3821), .Z(n3343) );
  NAND2_X1 U3203 ( .A1(n2471), .A2(n3343), .ZN(n2515) );
  NAND2_X1 U3204 ( .A1(n2516), .A2(n2515), .ZN(n2518) );
  XNOR2_X1 U3205 ( .A(n2518), .B(n2517), .ZN(n2523) );
  OR2_X1 U3206 ( .A1(n3359), .A2(n2498), .ZN(n2520) );
  NAND2_X1 U3207 ( .A1(n2480), .A2(n3343), .ZN(n2519) );
  NAND2_X1 U3208 ( .A1(n2520), .A2(n2519), .ZN(n2522) );
  XNOR2_X1 U3209 ( .A(n2523), .B(n2522), .ZN(n3332) );
  INV_X1 U32100 ( .A(n3332), .ZN(n2521) );
  NAND2_X1 U32110 ( .A1(n2523), .A2(n2522), .ZN(n2524) );
  NAND2_X1 U32120 ( .A1(n2621), .A2(REG0_REG_5__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32130 ( .A1(n3822), .A2(REG1_REG_5__SCAN_IN), .ZN(n2527) );
  XNOR2_X1 U32140 ( .A(n2541), .B(REG3_REG_5__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U32150 ( .A1(n2855), .A2(n3365), .ZN(n2526) );
  NAND2_X1 U32160 ( .A1(n3823), .A2(REG2_REG_5__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32170 ( .A1(n2912), .A2(n3988), .ZN(n2530) );
  MUX2_X1 U32180 ( .A(n4492), .B(DATAI_5_), .S(n3828), .Z(n3364) );
  NAND2_X1 U32190 ( .A1(n2471), .A2(n3364), .ZN(n2529) );
  NAND2_X1 U32200 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  XNOR2_X1 U32210 ( .A(n2531), .B(n2850), .ZN(n2534) );
  OR2_X1 U32220 ( .A1(n3384), .A2(n1996), .ZN(n2533) );
  NAND2_X1 U32230 ( .A1(n2912), .A2(n3364), .ZN(n2532) );
  NAND2_X1 U32240 ( .A1(n2533), .A2(n2532), .ZN(n2535) );
  XNOR2_X1 U32250 ( .A(n2534), .B(n2535), .ZN(n3279) );
  INV_X1 U32260 ( .A(n2534), .ZN(n2536) );
  NAND2_X1 U32270 ( .A1(n2536), .A2(n2535), .ZN(n2537) );
  NAND2_X1 U32280 ( .A1(n3822), .A2(REG1_REG_6__SCAN_IN), .ZN(n2546) );
  INV_X2 U32290 ( .A(n2538), .ZN(n2621) );
  NAND2_X1 U32300 ( .A1(n2621), .A2(REG0_REG_6__SCAN_IN), .ZN(n2545) );
  INV_X1 U32310 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2540) );
  INV_X1 U32320 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2539) );
  OAI21_X1 U32330 ( .B1(n2541), .B2(n2540), .A(n2539), .ZN(n2542) );
  AND2_X1 U32340 ( .A1(n2553), .A2(n2542), .ZN(n3389) );
  NAND2_X1 U32350 ( .A1(n2855), .A2(n3389), .ZN(n2544) );
  NAND2_X1 U32360 ( .A1(n3823), .A2(REG2_REG_6__SCAN_IN), .ZN(n2543) );
  NAND4_X1 U32370 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(n3987)
         );
  OR2_X1 U32380 ( .A1(n3281), .A2(n2498), .ZN(n2548) );
  MUX2_X1 U32390 ( .A(n3088), .B(DATAI_6_), .S(n3828), .Z(n3388) );
  NAND2_X1 U32400 ( .A1(n2912), .A2(n3388), .ZN(n2547) );
  NAND2_X1 U32410 ( .A1(n2548), .A2(n2547), .ZN(n3381) );
  NAND2_X1 U32420 ( .A1(n2912), .A2(n3987), .ZN(n2550) );
  NAND2_X1 U32430 ( .A1(n2471), .A2(n3388), .ZN(n2549) );
  NAND2_X1 U32440 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  XNOR2_X1 U32450 ( .A(n2551), .B(n2517), .ZN(n3380) );
  NAND2_X1 U32460 ( .A1(n3822), .A2(REG1_REG_7__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U32470 ( .A1(n2621), .A2(REG0_REG_7__SCAN_IN), .ZN(n2557) );
  INV_X1 U32480 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32490 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  AND2_X1 U32500 ( .A1(n2569), .A2(n2554), .ZN(n3407) );
  NAND2_X1 U32510 ( .A1(n2855), .A2(n3407), .ZN(n2556) );
  NAND2_X1 U32520 ( .A1(n3823), .A2(REG2_REG_7__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32530 ( .A1(n2912), .A2(n3986), .ZN(n2560) );
  MUX2_X1 U32540 ( .A(n3150), .B(DATAI_7_), .S(n3828), .Z(n3311) );
  NAND2_X1 U32550 ( .A1(n2471), .A2(n3311), .ZN(n2559) );
  NAND2_X1 U32560 ( .A1(n2560), .A2(n2559), .ZN(n2561) );
  XNOR2_X1 U32570 ( .A(n2561), .B(n2850), .ZN(n2565) );
  INV_X1 U32580 ( .A(n3986), .ZN(n3385) );
  OR2_X1 U32590 ( .A1(n3385), .A2(n1996), .ZN(n2563) );
  NAND2_X1 U32600 ( .A1(n2912), .A2(n3311), .ZN(n2562) );
  NAND2_X1 U32610 ( .A1(n2563), .A2(n2562), .ZN(n2564) );
  XNOR2_X1 U32620 ( .A(n2565), .B(n2564), .ZN(n3402) );
  NAND2_X1 U32630 ( .A1(n3403), .A2(n3402), .ZN(n2567) );
  INV_X1 U32640 ( .A(n2564), .ZN(n2566) );
  NAND2_X1 U32650 ( .A1(n2621), .A2(REG0_REG_8__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U32660 ( .A1(n3822), .A2(REG1_REG_8__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32670 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  AND2_X1 U32680 ( .A1(n2581), .A2(n2570), .ZN(n3438) );
  NAND2_X1 U32690 ( .A1(n2855), .A2(n3438), .ZN(n2572) );
  NAND2_X1 U32700 ( .A1(n3823), .A2(REG2_REG_8__SCAN_IN), .ZN(n2571) );
  NAND4_X1 U32710 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(n3985)
         );
  NAND2_X1 U32720 ( .A1(n2912), .A2(n3985), .ZN(n2576) );
  MUX2_X1 U32730 ( .A(n4491), .B(DATAI_8_), .S(n3828), .Z(n3426) );
  NAND2_X1 U32740 ( .A1(n2471), .A2(n3426), .ZN(n2575) );
  NAND2_X1 U32750 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  XNOR2_X1 U32760 ( .A(n2577), .B(n2517), .ZN(n2608) );
  OR2_X1 U32770 ( .A1(n3461), .A2(n2498), .ZN(n2579) );
  NAND2_X1 U32780 ( .A1(n2912), .A2(n3426), .ZN(n2578) );
  NAND2_X1 U32790 ( .A1(n2579), .A2(n2578), .ZN(n2609) );
  AND2_X1 U32800 ( .A1(n2608), .A2(n2609), .ZN(n3485) );
  NAND2_X1 U32810 ( .A1(n3822), .A2(REG1_REG_9__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32820 ( .A1(n2621), .A2(REG0_REG_9__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32830 ( .A1(n2581), .A2(n2580), .ZN(n2582) );
  NAND2_X1 U32840 ( .A1(n2855), .A2(n2248), .ZN(n2584) );
  NAND2_X1 U32850 ( .A1(n3823), .A2(REG2_REG_9__SCAN_IN), .ZN(n2583) );
  NAND4_X1 U32860 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), .ZN(n3984)
         );
  NAND2_X1 U32870 ( .A1(n2480), .A2(n3984), .ZN(n2589) );
  MUX2_X1 U32880 ( .A(n2587), .B(DATAI_9_), .S(n3828), .Z(n3466) );
  NAND2_X1 U32890 ( .A1(n2471), .A2(n3466), .ZN(n2588) );
  NAND2_X1 U32900 ( .A1(n2589), .A2(n2588), .ZN(n2590) );
  XNOR2_X1 U32910 ( .A(n2590), .B(n2850), .ZN(n2615) );
  OR2_X1 U32920 ( .A1(n3496), .A2(n2498), .ZN(n2592) );
  NAND2_X1 U32930 ( .A1(n2480), .A2(n3466), .ZN(n2591) );
  NAND2_X1 U32940 ( .A1(n2592), .A2(n2591), .ZN(n2613) );
  XNOR2_X1 U32950 ( .A(n2615), .B(n2613), .ZN(n3489) );
  INV_X1 U32960 ( .A(n3489), .ZN(n2612) );
  OR2_X1 U32970 ( .A1(n3485), .A2(n2612), .ZN(n3655) );
  NAND2_X1 U32980 ( .A1(n2621), .A2(REG0_REG_10__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U32990 ( .A1(n3822), .A2(REG1_REG_10__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33000 ( .A1(n2594), .A2(n2593), .ZN(n2595) );
  AND2_X1 U33010 ( .A1(n2623), .A2(n2595), .ZN(n3664) );
  NAND2_X1 U33020 ( .A1(n2855), .A2(n3664), .ZN(n2597) );
  NAND2_X1 U33030 ( .A1(n3823), .A2(REG2_REG_10__SCAN_IN), .ZN(n2596) );
  NAND4_X1 U33040 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n3983)
         );
  NAND2_X1 U33050 ( .A1(n2480), .A2(n3983), .ZN(n2601) );
  MUX2_X1 U33060 ( .A(n4490), .B(DATAI_10_), .S(n3828), .Z(n3498) );
  NAND2_X1 U33070 ( .A1(n2471), .A2(n3498), .ZN(n2600) );
  NAND2_X1 U33080 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  XNOR2_X1 U33090 ( .A(n2602), .B(n2517), .ZN(n2607) );
  INV_X1 U33100 ( .A(n3983), .ZN(n3009) );
  OR2_X1 U33110 ( .A1(n3009), .A2(n1996), .ZN(n2604) );
  NAND2_X1 U33120 ( .A1(n2480), .A2(n3498), .ZN(n2603) );
  NAND2_X1 U33130 ( .A1(n2604), .A2(n2603), .ZN(n2606) );
  XNOR2_X1 U33140 ( .A(n2607), .B(n2606), .ZN(n3661) );
  INV_X1 U33150 ( .A(n3661), .ZN(n2618) );
  INV_X1 U33160 ( .A(n2608), .ZN(n2611) );
  INV_X1 U33170 ( .A(n2609), .ZN(n2610) );
  NAND2_X1 U33180 ( .A1(n2611), .A2(n2610), .ZN(n3486) );
  OR2_X1 U33190 ( .A1(n2612), .A2(n3486), .ZN(n2617) );
  INV_X1 U33200 ( .A(n2613), .ZN(n2614) );
  NAND2_X1 U33210 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  INV_X1 U33220 ( .A(DATAI_11_), .ZN(n2620) );
  MUX2_X1 U33230 ( .A(n4489), .B(n2620), .S(n3828), .Z(n3481) );
  NAND2_X1 U33240 ( .A1(n2621), .A2(REG0_REG_11__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U33250 ( .A1(n3822), .A2(REG1_REG_11__SCAN_IN), .ZN(n2627) );
  INV_X1 U33260 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U33270 ( .A1(n2623), .A2(n2622), .ZN(n2624) );
  AND2_X1 U33280 ( .A1(n2636), .A2(n2624), .ZN(n3519) );
  NAND2_X1 U33290 ( .A1(n2855), .A2(n3519), .ZN(n2626) );
  NAND2_X1 U33300 ( .A1(n3823), .A2(REG2_REG_11__SCAN_IN), .ZN(n2625) );
  NAND4_X1 U33310 ( .A1(n2628), .A2(n2627), .A3(n2626), .A4(n2625), .ZN(n3982)
         );
  OR2_X1 U33320 ( .A1(n3543), .A2(n1996), .ZN(n2629) );
  OAI21_X1 U33330 ( .B1(n2817), .B2(n3481), .A(n2629), .ZN(n3476) );
  NAND2_X1 U33340 ( .A1(n2480), .A2(n3982), .ZN(n2630) );
  OAI21_X1 U33350 ( .B1(n3481), .B2(n2878), .A(n2630), .ZN(n2631) );
  XNOR2_X1 U33360 ( .A(n2631), .B(n2517), .ZN(n3475) );
  NAND2_X1 U33370 ( .A1(n3478), .A2(n3476), .ZN(n2632) );
  INV_X1 U33380 ( .A(n3682), .ZN(n2647) );
  MUX2_X1 U33390 ( .A(DATAI_12_), .B(n2635), .S(n2634), .Z(n3549) );
  NAND2_X1 U33400 ( .A1(n3549), .A2(n2471), .ZN(n2642) );
  NAND2_X1 U33410 ( .A1(n3822), .A2(REG1_REG_12__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U33420 ( .A1(n3824), .A2(REG0_REG_12__SCAN_IN), .ZN(n2639) );
  XNOR2_X1 U33430 ( .A(n2636), .B(REG3_REG_12__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U33440 ( .A1(n2855), .A2(n3690), .ZN(n2638) );
  NAND2_X1 U33450 ( .A1(n3823), .A2(REG2_REG_12__SCAN_IN), .ZN(n2637) );
  NAND4_X1 U33460 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .ZN(n3981)
         );
  NAND2_X1 U33470 ( .A1(n2480), .A2(n3981), .ZN(n2641) );
  NAND2_X1 U33480 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  XNOR2_X1 U33490 ( .A(n2643), .B(n2517), .ZN(n2648) );
  NAND2_X1 U33500 ( .A1(n3549), .A2(n2861), .ZN(n2645) );
  NAND2_X1 U33510 ( .A1(n2866), .A2(n3981), .ZN(n2644) );
  NAND2_X1 U33520 ( .A1(n2645), .A2(n2644), .ZN(n2649) );
  INV_X1 U3353 ( .A(n3684), .ZN(n2646) );
  INV_X1 U33540 ( .A(n2648), .ZN(n2651) );
  INV_X1 U3355 ( .A(n2649), .ZN(n2650) );
  NAND2_X1 U3356 ( .A1(n2651), .A2(n2650), .ZN(n3683) );
  INV_X1 U3357 ( .A(n3980), .ZN(n3582) );
  OR2_X1 U3358 ( .A1(n3582), .A2(n2498), .ZN(n2653) );
  NAND2_X1 U3359 ( .A1(n2480), .A2(n3010), .ZN(n2652) );
  NAND2_X1 U3360 ( .A1(n2653), .A2(n2652), .ZN(n3615) );
  AND2_X1 U3361 ( .A1(n3683), .A2(n3615), .ZN(n2655) );
  INV_X1 U3362 ( .A(n3615), .ZN(n2654) );
  INV_X1 U3363 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3364 ( .A1(n2657), .A2(n2656), .ZN(n2658) );
  AND2_X1 U3365 ( .A1(n2691), .A2(n2658), .ZN(n3639) );
  NAND2_X1 U3366 ( .A1(n3639), .A2(n2855), .ZN(n2662) );
  NAND2_X1 U3367 ( .A1(n3824), .A2(REG0_REG_14__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3368 ( .A1(n3822), .A2(REG1_REG_14__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3369 ( .A1(n3823), .A2(REG2_REG_14__SCAN_IN), .ZN(n2659) );
  NAND4_X1 U3370 ( .A1(n2662), .A2(n2661), .A3(n2660), .A4(n2659), .ZN(n3797)
         );
  NAND2_X1 U3371 ( .A1(n2480), .A2(n3797), .ZN(n2664) );
  MUX2_X1 U3372 ( .A(n4487), .B(DATAI_14_), .S(n3821), .Z(n2967) );
  NAND2_X1 U3373 ( .A1(n2471), .A2(n2967), .ZN(n2663) );
  NAND2_X1 U3374 ( .A1(n2664), .A2(n2663), .ZN(n2665) );
  XNOR2_X1 U3375 ( .A(n2665), .B(n2517), .ZN(n2710) );
  NAND2_X1 U3376 ( .A1(n2866), .A2(n3797), .ZN(n2667) );
  NAND2_X1 U3377 ( .A1(n2861), .A2(n2967), .ZN(n2666) );
  NAND2_X1 U3378 ( .A1(n2667), .A2(n2666), .ZN(n2711) );
  NAND2_X1 U3379 ( .A1(n2710), .A2(n2711), .ZN(n3711) );
  XNOR2_X1 U3380 ( .A(n2723), .B(REG3_REG_17__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U3381 ( .A1(n4300), .A2(n2855), .ZN(n2674) );
  NAND2_X1 U3382 ( .A1(n3824), .A2(REG0_REG_17__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3383 ( .A1(n3823), .A2(REG2_REG_17__SCAN_IN), .ZN(n2669) );
  OAI211_X1 U3384 ( .C1(n2493), .C2(n2671), .A(n2670), .B(n2669), .ZN(n2672)
         );
  INV_X1 U3385 ( .A(n2672), .ZN(n2673) );
  NAND2_X1 U3386 ( .A1(n3979), .A2(n2861), .ZN(n2677) );
  MUX2_X1 U3387 ( .A(n2675), .B(DATAI_17_), .S(n3821), .Z(n4299) );
  NAND2_X1 U3388 ( .A1(n2471), .A2(n4299), .ZN(n2676) );
  NAND2_X1 U3389 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  XNOR2_X1 U3390 ( .A(n2678), .B(n2517), .ZN(n2716) );
  NAND2_X1 U3391 ( .A1(n3979), .A2(n2866), .ZN(n2680) );
  NAND2_X1 U3392 ( .A1(n2861), .A2(n4299), .ZN(n2679) );
  NAND2_X1 U3393 ( .A1(n2680), .A2(n2679), .ZN(n2717) );
  AND2_X1 U3394 ( .A1(n2716), .A2(n2717), .ZN(n3729) );
  INV_X1 U3395 ( .A(n3729), .ZN(n2707) );
  NAND2_X1 U3396 ( .A1(n2693), .A2(n3719), .ZN(n2681) );
  NAND2_X1 U3397 ( .A1(n2723), .A2(n2681), .ZN(n4330) );
  AOI22_X1 U3398 ( .A1(n3822), .A2(REG1_REG_16__SCAN_IN), .B1(n3824), .B2(
        REG0_REG_16__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3399 ( .A1(n3823), .A2(REG2_REG_16__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3400 ( .A1(n4291), .A2(n2861), .ZN(n2685) );
  MUX2_X1 U3401 ( .A(n4486), .B(DATAI_16_), .S(n3821), .Z(n4327) );
  NAND2_X1 U3402 ( .A1(n2471), .A2(n4327), .ZN(n2684) );
  NAND2_X1 U3403 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  XNOR2_X1 U3404 ( .A(n2686), .B(n2850), .ZN(n2705) );
  INV_X1 U3405 ( .A(n2705), .ZN(n2689) );
  INV_X1 U3406 ( .A(n4327), .ZN(n2970) );
  NOR2_X1 U3407 ( .A1(n2817), .A2(n2970), .ZN(n2687) );
  AOI21_X1 U3408 ( .B1(n4291), .B2(n2866), .A(n2687), .ZN(n2704) );
  INV_X1 U3409 ( .A(n2704), .ZN(n2688) );
  NAND2_X1 U3410 ( .A1(n2689), .A2(n2688), .ZN(n3709) );
  INV_X1 U3411 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3412 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U3413 ( .A1(n2693), .A2(n2692), .ZN(n3605) );
  NAND2_X1 U3414 ( .A1(n3822), .A2(REG1_REG_15__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U3415 ( .A1(n3824), .A2(REG0_REG_15__SCAN_IN), .ZN(n2694) );
  AND2_X1 U3416 ( .A1(n2695), .A2(n2694), .ZN(n2697) );
  NAND2_X1 U3417 ( .A1(n3823), .A2(REG2_REG_15__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3418 ( .A1(n4313), .A2(n2861), .ZN(n2699) );
  MUX2_X1 U3419 ( .A(n4033), .B(DATAI_15_), .S(n3821), .Z(n3602) );
  NAND2_X1 U3420 ( .A1(n2471), .A2(n3602), .ZN(n2698) );
  NAND2_X1 U3421 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  XNOR2_X1 U3422 ( .A(n2700), .B(n2517), .ZN(n3713) );
  NAND2_X1 U3423 ( .A1(n2866), .A2(n4313), .ZN(n2702) );
  NAND2_X1 U3424 ( .A1(n2861), .A2(n3602), .ZN(n2701) );
  NAND2_X1 U3425 ( .A1(n2702), .A2(n2701), .ZN(n3794) );
  NAND2_X1 U3426 ( .A1(n3713), .A2(n3794), .ZN(n2703) );
  NAND2_X1 U3427 ( .A1(n3709), .A2(n2703), .ZN(n2706) );
  NAND2_X1 U3428 ( .A1(n2705), .A2(n2704), .ZN(n3710) );
  NAND2_X1 U3429 ( .A1(n2706), .A2(n3710), .ZN(n3726) );
  INV_X1 U3430 ( .A(n2709), .ZN(n2715) );
  INV_X1 U3431 ( .A(n2710), .ZN(n2713) );
  INV_X1 U3432 ( .A(n2711), .ZN(n2712) );
  NAND2_X1 U3433 ( .A1(n2713), .A2(n2712), .ZN(n3712) );
  OAI211_X1 U3434 ( .C1(n3794), .C2(n3713), .A(n3710), .B(n3712), .ZN(n2714)
         );
  INV_X1 U3435 ( .A(n2714), .ZN(n3724) );
  INV_X1 U3436 ( .A(n2716), .ZN(n2719) );
  INV_X1 U3437 ( .A(n2717), .ZN(n2718) );
  NAND2_X1 U3438 ( .A1(n2719), .A2(n2718), .ZN(n3728) );
  INV_X1 U3439 ( .A(n3769), .ZN(n2735) );
  AND2_X1 U3440 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2721) );
  INV_X1 U3441 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3733) );
  INV_X1 U3442 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2722) );
  OAI21_X1 U3443 ( .B1(n2723), .B2(n3733), .A(n2722), .ZN(n2724) );
  NAND2_X1 U3444 ( .A1(n2739), .A2(n2724), .ZN(n4279) );
  OR2_X1 U3445 ( .A1(n4279), .A2(n2921), .ZN(n2730) );
  NAND2_X1 U3446 ( .A1(n3824), .A2(REG0_REG_18__SCAN_IN), .ZN(n2726) );
  NAND2_X1 U3447 ( .A1(n3823), .A2(REG2_REG_18__SCAN_IN), .ZN(n2725) );
  OAI211_X1 U3448 ( .C1(n2493), .C2(n2727), .A(n2726), .B(n2725), .ZN(n2728)
         );
  INV_X1 U3449 ( .A(n2728), .ZN(n2729) );
  NAND2_X1 U3450 ( .A1(n4293), .A2(n2866), .ZN(n2733) );
  MUX2_X1 U3451 ( .A(n2731), .B(DATAI_18_), .S(n3821), .Z(n4272) );
  NAND2_X1 U3452 ( .A1(n2912), .A2(n4272), .ZN(n2732) );
  NAND2_X1 U3453 ( .A1(n2733), .A2(n2732), .ZN(n3770) );
  AOI22_X1 U3454 ( .A1(n4293), .A2(n2861), .B1(n2471), .B2(n4272), .ZN(n2734)
         );
  XOR2_X1 U3455 ( .A(n2517), .B(n2734), .Z(n3771) );
  INV_X1 U3456 ( .A(n3770), .ZN(n2736) );
  NAND2_X1 U3457 ( .A1(n2738), .A2(n2737), .ZN(n3667) );
  INV_X1 U34580 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U34590 ( .A1(n2739), .A2(n4619), .ZN(n2740) );
  AND2_X1 U3460 ( .A1(n2755), .A2(n2740), .ZN(n4266) );
  NAND2_X1 U3461 ( .A1(n4266), .A2(n2855), .ZN(n2745) );
  NAND2_X1 U3462 ( .A1(n3822), .A2(REG1_REG_19__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U3463 ( .A1(n3824), .A2(REG0_REG_19__SCAN_IN), .ZN(n2741) );
  OAI211_X1 U3464 ( .C1(n4627), .C2(n2874), .A(n2742), .B(n2741), .ZN(n2743)
         );
  INV_X1 U3465 ( .A(n2743), .ZN(n2744) );
  NAND2_X1 U3466 ( .A1(n4273), .A2(n2861), .ZN(n2747) );
  MUX2_X1 U34670 ( .A(n3969), .B(DATAI_19_), .S(n3828), .Z(n4263) );
  NAND2_X1 U3468 ( .A1(n2471), .A2(n4263), .ZN(n2746) );
  NAND2_X1 U34690 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  XNOR2_X1 U3470 ( .A(n2748), .B(n2850), .ZN(n2751) );
  INV_X1 U34710 ( .A(n4263), .ZN(n4254) );
  NOR2_X1 U3472 ( .A1(n2817), .A2(n4254), .ZN(n2749) );
  AOI21_X1 U34730 ( .B1(n4273), .B2(n2866), .A(n2749), .ZN(n2750) );
  NAND2_X1 U3474 ( .A1(n2751), .A2(n2750), .ZN(n2752) );
  OAI21_X1 U34750 ( .B1(n2751), .B2(n2750), .A(n2752), .ZN(n3668) );
  INV_X1 U3476 ( .A(n2752), .ZN(n2753) );
  INV_X1 U34770 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3752) );
  NAND2_X1 U3478 ( .A1(n2755), .A2(n3752), .ZN(n2756) );
  NAND2_X1 U34790 ( .A1(n2768), .A2(n2756), .ZN(n4237) );
  INV_X1 U3480 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U34810 ( .A1(n3822), .A2(REG1_REG_20__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U3482 ( .A1(n3824), .A2(REG0_REG_20__SCAN_IN), .ZN(n2757) );
  OAI211_X1 U34830 ( .C1(n4238), .C2(n2874), .A(n2758), .B(n2757), .ZN(n2759)
         );
  INV_X1 U3484 ( .A(n2759), .ZN(n2760) );
  NAND2_X1 U34850 ( .A1(n4252), .A2(n2861), .ZN(n2763) );
  NAND2_X1 U3486 ( .A1(n3828), .A2(DATAI_20_), .ZN(n3753) );
  OR2_X1 U34870 ( .A1(n2878), .A2(n3753), .ZN(n2762) );
  NAND2_X1 U3488 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  XNOR2_X1 U34890 ( .A(n2764), .B(n2850), .ZN(n2767) );
  NOR2_X1 U3490 ( .A1(n2817), .A2(n3753), .ZN(n2765) );
  AOI21_X1 U34910 ( .B1(n4252), .B2(n2866), .A(n2765), .ZN(n2766) );
  NOR2_X1 U3492 ( .A1(n2767), .A2(n2766), .ZN(n3749) );
  AND2_X1 U34930 ( .A1(n2767), .A2(n2766), .ZN(n3071) );
  INV_X1 U3494 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U34950 ( .A1(n2768), .A2(n4653), .ZN(n2769) );
  NAND2_X1 U3496 ( .A1(n2790), .A2(n2769), .ZN(n4217) );
  INV_X1 U34970 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U3498 ( .A1(n3823), .A2(REG2_REG_21__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U34990 ( .A1(n3824), .A2(REG0_REG_21__SCAN_IN), .ZN(n2770) );
  OAI211_X1 U3500 ( .C1(n2493), .C2(n4696), .A(n2771), .B(n2770), .ZN(n2772)
         );
  INV_X1 U35010 ( .A(n2772), .ZN(n2773) );
  NAND2_X1 U3502 ( .A1(n4193), .A2(n2861), .ZN(n2776) );
  NAND2_X1 U35030 ( .A1(n3821), .A2(DATAI_21_), .ZN(n4215) );
  OR2_X1 U3504 ( .A1(n2878), .A2(n4215), .ZN(n2775) );
  NAND2_X1 U35050 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  XNOR2_X1 U35060 ( .A(n2777), .B(n2850), .ZN(n2780) );
  NOR2_X1 U35070 ( .A1(n2817), .A2(n4215), .ZN(n2778) );
  AOI21_X1 U35080 ( .B1(n4193), .B2(n2866), .A(n2778), .ZN(n2779) );
  NAND2_X1 U35090 ( .A1(n2780), .A2(n2779), .ZN(n3067) );
  NOR2_X1 U35100 ( .A1(n2780), .A2(n2779), .ZN(n3069) );
  XNOR2_X1 U35110 ( .A(n2790), .B(REG3_REG_22__SCAN_IN), .ZN(n4198) );
  NAND2_X1 U35120 ( .A1(n4198), .A2(n2855), .ZN(n2785) );
  INV_X1 U35130 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U35140 ( .A1(n3824), .A2(REG0_REG_22__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U35150 ( .A1(n3822), .A2(REG1_REG_22__SCAN_IN), .ZN(n2781) );
  OAI211_X1 U35160 ( .C1(n4613), .C2(n2874), .A(n2782), .B(n2781), .ZN(n2783)
         );
  INV_X1 U35170 ( .A(n2783), .ZN(n2784) );
  INV_X1 U35180 ( .A(n4208), .ZN(n3646) );
  NAND2_X1 U35190 ( .A1(n3821), .A2(DATAI_22_), .ZN(n4199) );
  OAI22_X1 U35200 ( .A1(n3646), .A2(n2498), .B1(n2817), .B2(n4199), .ZN(n2803)
         );
  NAND2_X1 U35210 ( .A1(n4208), .A2(n2861), .ZN(n2787) );
  OR2_X1 U35220 ( .A1(n2878), .A2(n4199), .ZN(n2786) );
  NAND2_X1 U35230 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  XNOR2_X1 U35240 ( .A(n2788), .B(n2517), .ZN(n2802) );
  XOR2_X1 U35250 ( .A(n2803), .B(n2802), .Z(n3760) );
  NAND2_X1 U35260 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2789) );
  INV_X1 U35270 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3762) );
  INV_X1 U35280 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3645) );
  OAI21_X1 U35290 ( .B1(n2790), .B2(n3762), .A(n3645), .ZN(n2791) );
  AND2_X1 U35300 ( .A1(n2818), .A2(n2791), .ZN(n4180) );
  NAND2_X1 U35310 ( .A1(n4180), .A2(n2855), .ZN(n2797) );
  INV_X1 U35320 ( .A(REG2_REG_23__SCAN_IN), .ZN(n2794) );
  NAND2_X1 U35330 ( .A1(n3822), .A2(REG1_REG_23__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U35340 ( .A1(n3824), .A2(REG0_REG_23__SCAN_IN), .ZN(n2792) );
  OAI211_X1 U35350 ( .C1(n2794), .C2(n2874), .A(n2793), .B(n2792), .ZN(n2795)
         );
  INV_X1 U35360 ( .A(n2795), .ZN(n2796) );
  NAND2_X1 U35370 ( .A1(n4191), .A2(n2861), .ZN(n2799) );
  NAND2_X1 U35380 ( .A1(n3828), .A2(DATAI_23_), .ZN(n4178) );
  OR2_X1 U35390 ( .A1(n2878), .A2(n4178), .ZN(n2798) );
  NAND2_X1 U35400 ( .A1(n2799), .A2(n2798), .ZN(n2800) );
  XNOR2_X1 U35410 ( .A(n2800), .B(n2517), .ZN(n2830) );
  NOR2_X1 U35420 ( .A1(n2817), .A2(n4178), .ZN(n2801) );
  AOI21_X1 U35430 ( .B1(n4191), .B2(n2866), .A(n2801), .ZN(n2828) );
  XNOR2_X1 U35440 ( .A(n2830), .B(n2828), .ZN(n3643) );
  INV_X1 U35450 ( .A(n2802), .ZN(n2805) );
  INV_X1 U35460 ( .A(n2803), .ZN(n2804) );
  NAND2_X1 U35470 ( .A1(n2805), .A2(n2804), .ZN(n3644) );
  INV_X1 U35480 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4651) );
  INV_X1 U35490 ( .A(n2807), .ZN(n2820) );
  INV_X1 U35500 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U35510 ( .A1(n2820), .A2(n3704), .ZN(n2808) );
  NAND2_X1 U35520 ( .A1(n2840), .A2(n2808), .ZN(n3703) );
  INV_X1 U35530 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U35540 ( .A1(n3822), .A2(REG1_REG_25__SCAN_IN), .ZN(n2810) );
  NAND2_X1 U35550 ( .A1(n3823), .A2(REG2_REG_25__SCAN_IN), .ZN(n2809) );
  OAI211_X1 U35560 ( .C1(n2538), .C2(n4667), .A(n2810), .B(n2809), .ZN(n2811)
         );
  INV_X1 U35570 ( .A(n2811), .ZN(n2812) );
  NAND2_X1 U35580 ( .A1(n4113), .A2(n2861), .ZN(n2815) );
  NAND2_X1 U35590 ( .A1(n3821), .A2(DATAI_25_), .ZN(n4136) );
  OR2_X1 U35600 ( .A1(n2878), .A2(n4136), .ZN(n2814) );
  NAND2_X1 U35610 ( .A1(n2815), .A2(n2814), .ZN(n2816) );
  XNOR2_X1 U35620 ( .A(n2816), .B(n2517), .ZN(n3700) );
  OAI22_X1 U35630 ( .A1(n4154), .A2(n2498), .B1(n2817), .B2(n4136), .ZN(n3699)
         );
  NAND2_X1 U35640 ( .A1(n3700), .A2(n3699), .ZN(n3698) );
  NAND2_X1 U35650 ( .A1(n2818), .A2(n4651), .ZN(n2819) );
  INV_X1 U35660 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U35670 ( .A1(n3822), .A2(REG1_REG_24__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U35680 ( .A1(n3823), .A2(REG2_REG_24__SCAN_IN), .ZN(n2821) );
  OAI211_X1 U35690 ( .C1(n2538), .C2(n4721), .A(n2822), .B(n2821), .ZN(n2823)
         );
  INV_X1 U35700 ( .A(n2823), .ZN(n2824) );
  NAND2_X1 U35710 ( .A1(n4132), .A2(n2861), .ZN(n2826) );
  NAND2_X1 U35720 ( .A1(n3821), .A2(DATAI_24_), .ZN(n4157) );
  OR2_X1 U35730 ( .A1(n2878), .A2(n4157), .ZN(n2825) );
  NAND2_X1 U35740 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
  XNOR2_X1 U35750 ( .A(n2827), .B(n2517), .ZN(n3743) );
  INV_X1 U35760 ( .A(n2828), .ZN(n2829) );
  NAND2_X1 U35770 ( .A1(n2830), .A2(n2829), .ZN(n3696) );
  INV_X1 U35780 ( .A(n3696), .ZN(n2832) );
  NOR2_X1 U35790 ( .A1(n2817), .A2(n4157), .ZN(n2831) );
  AOI21_X1 U35800 ( .B1(n4132), .B2(n2866), .A(n2831), .ZN(n3695) );
  NAND2_X1 U35810 ( .A1(n3696), .A2(n3695), .ZN(n3693) );
  OAI21_X1 U3582 ( .B1(n3743), .B2(n2832), .A(n3693), .ZN(n2833) );
  INV_X1 U3583 ( .A(n3743), .ZN(n2836) );
  INV_X1 U3584 ( .A(n3699), .ZN(n2835) );
  AOI21_X1 U3585 ( .B1(n2836), .B2(n3695), .A(n2835), .ZN(n2834) );
  NAND3_X1 U3586 ( .A1(n2836), .A2(n3695), .A3(n2835), .ZN(n2837) );
  INV_X1 U3587 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U3588 ( .A1(n2840), .A2(n4668), .ZN(n2841) );
  NAND2_X1 U3589 ( .A1(n4120), .A2(n2855), .ZN(n2847) );
  INV_X1 U3590 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2844) );
  NAND2_X1 U3591 ( .A1(n3822), .A2(REG1_REG_26__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3592 ( .A1(n3824), .A2(REG0_REG_26__SCAN_IN), .ZN(n2842) );
  OAI211_X1 U3593 ( .C1(n2844), .C2(n2874), .A(n2843), .B(n2842), .ZN(n2845)
         );
  INV_X1 U3594 ( .A(n2845), .ZN(n2846) );
  NAND2_X1 U3595 ( .A1(n4094), .A2(n2861), .ZN(n2849) );
  NAND2_X1 U3596 ( .A1(n3821), .A2(DATAI_26_), .ZN(n4118) );
  OR2_X1 U3597 ( .A1(n2878), .A2(n4118), .ZN(n2848) );
  NAND2_X1 U3598 ( .A1(n2849), .A2(n2848), .ZN(n2851) );
  XNOR2_X1 U3599 ( .A(n2851), .B(n2850), .ZN(n2854) );
  NOR2_X1 U3600 ( .A1(n2817), .A2(n4118), .ZN(n2852) );
  AOI21_X1 U3601 ( .B1(n4094), .B2(n2866), .A(n2852), .ZN(n2853) );
  OR2_X1 U3602 ( .A1(n2854), .A2(n2853), .ZN(n3783) );
  XNOR2_X1 U3603 ( .A(n2870), .B(REG3_REG_27__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U3604 ( .A1(n4099), .A2(n2855), .ZN(n2860) );
  INV_X1 U3605 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U3606 ( .A1(n3823), .A2(REG2_REG_27__SCAN_IN), .ZN(n2857) );
  NAND2_X1 U3607 ( .A1(n3822), .A2(REG1_REG_27__SCAN_IN), .ZN(n2856) );
  OAI211_X1 U3608 ( .C1(n2538), .C2(n4641), .A(n2857), .B(n2856), .ZN(n2858)
         );
  INV_X1 U3609 ( .A(n2858), .ZN(n2859) );
  NAND2_X1 U3610 ( .A1(n3325), .A2(n2861), .ZN(n2863) );
  NAND2_X1 U3611 ( .A1(n3821), .A2(DATAI_27_), .ZN(n3630) );
  OR2_X1 U3612 ( .A1(n2878), .A2(n3630), .ZN(n2862) );
  NAND2_X1 U3613 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  XNOR2_X1 U3614 ( .A(n2864), .B(n2517), .ZN(n2904) );
  NOR2_X1 U3615 ( .A1(n2817), .A2(n3630), .ZN(n2865) );
  AOI21_X1 U3616 ( .B1(n3325), .B2(n2866), .A(n2865), .ZN(n2902) );
  XNOR2_X1 U3617 ( .A(n2904), .B(n2902), .ZN(n3627) );
  INV_X1 U3618 ( .A(n2906), .ZN(n2901) );
  INV_X1 U3619 ( .A(n2870), .ZN(n2868) );
  AND2_X1 U3620 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2867) );
  NAND2_X1 U3621 ( .A1(n2868), .A2(n2867), .ZN(n4077) );
  INV_X1 U3622 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3629) );
  INV_X1 U3623 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2869) );
  OAI21_X1 U3624 ( .B1(n2870), .B2(n3629), .A(n2869), .ZN(n2871) );
  NAND2_X1 U3625 ( .A1(n4077), .A2(n2871), .ZN(n4085) );
  INV_X1 U3626 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4084) );
  NAND2_X1 U3627 ( .A1(n3822), .A2(REG1_REG_28__SCAN_IN), .ZN(n2873) );
  NAND2_X1 U3628 ( .A1(n3824), .A2(REG0_REG_28__SCAN_IN), .ZN(n2872) );
  OAI211_X1 U3629 ( .C1(n4084), .C2(n2874), .A(n2873), .B(n2872), .ZN(n2875)
         );
  INV_X1 U3630 ( .A(n2875), .ZN(n2876) );
  NAND2_X1 U3631 ( .A1(n3821), .A2(DATAI_28_), .ZN(n4062) );
  OAI22_X1 U3632 ( .A1(n4096), .A2(n2817), .B1(n2878), .B2(n4062), .ZN(n2879)
         );
  XNOR2_X1 U3633 ( .A(n2879), .B(n2517), .ZN(n2881) );
  OAI22_X1 U3634 ( .A1(n4096), .A2(n1996), .B1(n2817), .B2(n4062), .ZN(n2880)
         );
  XNOR2_X1 U3635 ( .A(n2881), .B(n2880), .ZN(n2909) );
  NOR4_X1 U3636 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2885) );
  NOR4_X1 U3637 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2884) );
  NOR4_X1 U3638 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2883) );
  NOR4_X1 U3639 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2882) );
  NAND4_X1 U3640 ( .A1(n2885), .A2(n2884), .A3(n2883), .A4(n2882), .ZN(n2893)
         );
  NOR4_X1 U3641 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n4603) );
  NOR2_X1 U3642 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .ZN(n2888)
         );
  NOR4_X1 U3643 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2887) );
  NOR4_X1 U3644 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2886) );
  NAND4_X1 U3645 ( .A1(n4603), .A2(n2888), .A3(n2887), .A4(n2886), .ZN(n2892)
         );
  INV_X1 U3646 ( .A(n4483), .ZN(n2894) );
  NAND2_X1 U3647 ( .A1(n2896), .A2(n2894), .ZN(n2890) );
  MUX2_X1 U3648 ( .A(n2896), .B(n2890), .S(B_REG_SCAN_IN), .Z(n2891) );
  OAI21_X1 U3649 ( .B1(n2893), .B2(n2892), .A(n3097), .ZN(n3045) );
  INV_X1 U3650 ( .A(n4482), .ZN(n2895) );
  NAND2_X1 U3651 ( .A1(n2894), .A2(n2895), .ZN(n3044) );
  AND2_X1 U3652 ( .A1(n3045), .A2(n3044), .ZN(n3238) );
  INV_X1 U3653 ( .A(D_REG_0__SCAN_IN), .ZN(n3103) );
  INV_X1 U3654 ( .A(D_REG_1__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U3655 ( .A1(n3097), .A2(n3100), .ZN(n3236) );
  NAND3_X1 U3656 ( .A1(n3238), .A2(n3059), .A3(n3236), .ZN(n2928) );
  INV_X1 U3657 ( .A(n2928), .ZN(n2899) );
  AND2_X1 U3658 ( .A1(n3241), .A2(n3962), .ZN(n2915) );
  OR2_X1 U3659 ( .A1(n3189), .A2(n2915), .ZN(n2897) );
  NAND2_X1 U3660 ( .A1(n2897), .A2(n3036), .ZN(n2913) );
  NOR2_X1 U3661 ( .A1(n2913), .A2(n3040), .ZN(n2898) );
  NAND2_X1 U3662 ( .A1(n2901), .A2(n2900), .ZN(n2937) );
  INV_X1 U3663 ( .A(n2909), .ZN(n2905) );
  INV_X1 U3664 ( .A(n2902), .ZN(n2903) );
  NAND2_X1 U3665 ( .A1(n2904), .A2(n2903), .ZN(n2907) );
  NAND4_X1 U3666 ( .A1(n2906), .A2(n3773), .A3(n2905), .A4(n2907), .ZN(n2936)
         );
  INV_X1 U3667 ( .A(n2907), .ZN(n2908) );
  NOR2_X1 U3668 ( .A1(n2910), .A2(n4543), .ZN(n2911) );
  NAND2_X1 U3669 ( .A1(n2912), .A2(n2911), .ZN(n3972) );
  NOR2_X1 U3670 ( .A1(n2928), .A2(n3972), .ZN(n2927) );
  NAND2_X1 U3671 ( .A1(n2927), .A2(n4481), .ZN(n3776) );
  NAND2_X1 U3672 ( .A1(n2913), .A2(n4253), .ZN(n2914) );
  NAND2_X1 U3673 ( .A1(n2928), .A2(n2914), .ZN(n2916) );
  NAND2_X1 U3674 ( .A1(n2916), .A2(n3234), .ZN(n3183) );
  NAND2_X1 U3675 ( .A1(n3066), .A2(n2917), .ZN(n2918) );
  OAI21_X1 U3676 ( .B1(n3183), .B2(n2918), .A(STATE_REG_SCAN_IN), .ZN(n2920)
         );
  INV_X1 U3677 ( .A(n3972), .ZN(n2919) );
  NAND2_X1 U3678 ( .A1(n2928), .A2(n2919), .ZN(n3184) );
  INV_X1 U3679 ( .A(n3802), .ZN(n3781) );
  NOR2_X1 U3680 ( .A1(n4085), .A2(n3781), .ZN(n2932) );
  OR2_X1 U3681 ( .A1(n4077), .A2(n2921), .ZN(n2926) );
  NAND2_X1 U3682 ( .A1(n3823), .A2(REG2_REG_29__SCAN_IN), .ZN(n2924) );
  NAND2_X1 U3683 ( .A1(n3822), .A2(REG1_REG_29__SCAN_IN), .ZN(n2923) );
  NAND2_X1 U3684 ( .A1(n3824), .A2(REG0_REG_29__SCAN_IN), .ZN(n2922) );
  AND3_X1 U3685 ( .A1(n2924), .A2(n2923), .A3(n2922), .ZN(n2925) );
  NAND2_X1 U3686 ( .A1(n2927), .A2(n3168), .ZN(n3787) );
  NOR3_X1 U3687 ( .A1(n2928), .A2(n3040), .A3(n4253), .ZN(n2929) );
  NOR2_X1 U3688 ( .A1(n4558), .A2(n2454), .ZN(n3041) );
  NOR2_X2 U3689 ( .A1(n2929), .A2(n4534), .ZN(n3763) );
  INV_X1 U3690 ( .A(n4062), .ZN(n2995) );
  AOI22_X1 U3691 ( .A1(n3778), .A2(n2995), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2930) );
  OAI21_X1 U3692 ( .B1(n3831), .B2(n3787), .A(n2930), .ZN(n2931) );
  AOI211_X1 U3693 ( .C1(n3798), .C2(n3325), .A(n2932), .B(n2931), .ZN(n2933)
         );
  NAND3_X1 U3694 ( .A1(n2937), .A2(n2936), .A3(n2935), .ZN(U3217) );
  AND2_X1 U3695 ( .A1(n3992), .A2(n3048), .ZN(n3194) );
  INV_X1 U3696 ( .A(n3219), .ZN(n2940) );
  NAND2_X1 U3697 ( .A1(n3272), .A2(n2940), .ZN(n2941) );
  INV_X1 U3698 ( .A(n3674), .ZN(n3204) );
  NAND2_X2 U3699 ( .A1(n3894), .A2(n3897), .ZN(n3193) );
  NAND2_X1 U3700 ( .A1(n2939), .A2(n3193), .ZN(n2944) );
  NAND2_X1 U3701 ( .A1(n2940), .A2(n3198), .ZN(n3900) );
  NAND2_X1 U3702 ( .A1(n3001), .A2(n2941), .ZN(n2943) );
  AND2_X1 U3703 ( .A1(n2938), .A2(n3674), .ZN(n3208) );
  NAND2_X1 U3704 ( .A1(n3208), .A2(n2941), .ZN(n2942) );
  NAND2_X1 U3705 ( .A1(n3990), .A2(n3255), .ZN(n2945) );
  NAND2_X1 U3706 ( .A1(n3251), .A2(n2945), .ZN(n3340) );
  NAND2_X1 U3707 ( .A1(n3336), .A2(n3989), .ZN(n3905) );
  INV_X1 U3708 ( .A(n3364), .ZN(n3004) );
  NAND2_X1 U3709 ( .A1(n3384), .A2(n3004), .ZN(n2947) );
  NAND2_X1 U3710 ( .A1(n3212), .A2(n3273), .ZN(n3339) );
  AND3_X1 U3711 ( .A1(n3337), .A2(n2947), .A3(n3339), .ZN(n2946) );
  AND2_X1 U3712 ( .A1(n3989), .A2(n3343), .ZN(n3353) );
  AOI22_X1 U3713 ( .A1(n2947), .A2(n3353), .B1(n3364), .B2(n3988), .ZN(n2948)
         );
  NAND2_X1 U3714 ( .A1(n3385), .A2(n3311), .ZN(n3006) );
  NAND2_X1 U3715 ( .A1(n3049), .A2(n3986), .ZN(n3913) );
  NAND2_X1 U3716 ( .A1(n3281), .A2(n2949), .ZN(n2950) );
  AND2_X1 U3717 ( .A1(n3987), .A2(n3388), .ZN(n2951) );
  AOI22_X1 U3718 ( .A1(n3908), .A2(n2951), .B1(n3311), .B2(n3986), .ZN(n2952)
         );
  NAND2_X1 U3719 ( .A1(n3461), .A2(n2185), .ZN(n2953) );
  NAND2_X1 U3720 ( .A1(n3423), .A2(n2953), .ZN(n2955) );
  NAND2_X1 U3721 ( .A1(n3985), .A2(n3426), .ZN(n2954) );
  NAND2_X1 U3722 ( .A1(n2955), .A2(n2954), .ZN(n3458) );
  AND2_X1 U3723 ( .A1(n3466), .A2(n3984), .ZN(n2956) );
  NAND2_X1 U3724 ( .A1(n3496), .A2(n2184), .ZN(n2957) );
  OAI21_X1 U3725 ( .B1(n3458), .B2(n2956), .A(n2957), .ZN(n2958) );
  INV_X1 U3726 ( .A(n2958), .ZN(n3501) );
  NAND2_X1 U3727 ( .A1(n3009), .A2(n3654), .ZN(n2960) );
  AND2_X1 U3728 ( .A1(n3983), .A2(n3498), .ZN(n2959) );
  AOI21_X1 U3729 ( .B1(n3501), .B2(n2960), .A(n2959), .ZN(n3510) );
  NAND2_X1 U3730 ( .A1(n3517), .A2(n3543), .ZN(n3540) );
  NAND2_X1 U3731 ( .A1(n3481), .A2(n3982), .ZN(n3542) );
  NAND2_X1 U3732 ( .A1(n3540), .A2(n3542), .ZN(n3852) );
  NAND2_X1 U3733 ( .A1(n3510), .A2(n3852), .ZN(n3509) );
  NAND2_X1 U3734 ( .A1(n3543), .A2(n3481), .ZN(n2961) );
  NAND2_X1 U3735 ( .A1(n3509), .A2(n2961), .ZN(n3547) );
  NAND2_X1 U3736 ( .A1(n3549), .A2(n3981), .ZN(n2962) );
  NAND2_X1 U3737 ( .A1(n3547), .A2(n2962), .ZN(n2964) );
  OR2_X1 U3738 ( .A1(n3549), .A2(n3981), .ZN(n2963) );
  NAND2_X1 U3739 ( .A1(n2964), .A2(n2963), .ZN(n3570) );
  NOR2_X1 U3740 ( .A1(n3980), .A2(n3010), .ZN(n2966) );
  NAND2_X1 U3741 ( .A1(n3980), .A2(n3010), .ZN(n2965) );
  INV_X1 U3742 ( .A(n3797), .ZN(n2968) );
  NAND2_X1 U3743 ( .A1(n2968), .A2(n2967), .ZN(n3807) );
  NAND2_X1 U3744 ( .A1(n3637), .A2(n3797), .ZN(n3808) );
  NAND2_X1 U3745 ( .A1(n4313), .A2(n3602), .ZN(n4320) );
  NAND2_X1 U3746 ( .A1(n4291), .A2(n4327), .ZN(n2969) );
  AND2_X1 U3747 ( .A1(n4320), .A2(n2969), .ZN(n2972) );
  INV_X1 U3748 ( .A(n2969), .ZN(n2971) );
  NAND2_X1 U3749 ( .A1(n4291), .A2(n2970), .ZN(n3937) );
  OR2_X1 U3750 ( .A1(n4291), .A2(n2970), .ZN(n3935) );
  INV_X1 U3751 ( .A(n4310), .ZN(n4325) );
  OR2_X1 U3752 ( .A1(n4313), .A2(n3602), .ZN(n4321) );
  AND2_X1 U3753 ( .A1(n4325), .A2(n4321), .ZN(n4322) );
  OR2_X1 U3754 ( .A1(n3979), .A2(n4299), .ZN(n2973) );
  NAND2_X1 U3755 ( .A1(n4304), .A2(n2973), .ZN(n2975) );
  NAND2_X1 U3756 ( .A1(n3979), .A2(n4299), .ZN(n2974) );
  NAND2_X1 U3757 ( .A1(n2975), .A2(n2974), .ZN(n4283) );
  INV_X1 U3758 ( .A(n4283), .ZN(n2977) );
  OR2_X1 U3759 ( .A1(n4293), .A2(n4278), .ZN(n4248) );
  NAND2_X1 U3760 ( .A1(n4293), .A2(n4278), .ZN(n4249) );
  OR2_X1 U3761 ( .A1(n4293), .A2(n4272), .ZN(n2978) );
  NAND2_X1 U3762 ( .A1(n4273), .A2(n4263), .ZN(n2979) );
  NAND2_X1 U3763 ( .A1(n4252), .A2(n4234), .ZN(n3850) );
  NAND2_X1 U3764 ( .A1(n4222), .A2(n3850), .ZN(n2980) );
  NAND2_X1 U3765 ( .A1(n4206), .A2(n3753), .ZN(n3851) );
  INV_X1 U3766 ( .A(n4215), .ZN(n3030) );
  NAND2_X1 U3767 ( .A1(n4193), .A2(n3030), .ZN(n2981) );
  NAND2_X1 U3768 ( .A1(n4208), .A2(n4199), .ZN(n3031) );
  NAND2_X1 U3769 ( .A1(n3764), .A2(n4178), .ZN(n4145) );
  OR2_X1 U3770 ( .A1(n4189), .A2(n2247), .ZN(n2982) );
  NOR2_X1 U3771 ( .A1(n2982), .A2(n2241), .ZN(n2983) );
  NAND2_X1 U3772 ( .A1(n4228), .A2(n4215), .ZN(n4142) );
  INV_X1 U3773 ( .A(n4199), .ZN(n2984) );
  NAND2_X1 U3774 ( .A1(n4208), .A2(n2984), .ZN(n4163) );
  NAND2_X1 U3775 ( .A1(n4191), .A2(n3053), .ZN(n2985) );
  AND2_X1 U3776 ( .A1(n4163), .A2(n2985), .ZN(n4144) );
  INV_X1 U3777 ( .A(n2986), .ZN(n2987) );
  AND2_X1 U3778 ( .A1(n4144), .A2(n2987), .ZN(n2988) );
  NOR2_X1 U3779 ( .A1(n2241), .A2(n2989), .ZN(n2990) );
  INV_X1 U3780 ( .A(n4136), .ZN(n4131) );
  NOR2_X1 U3781 ( .A1(n4113), .A2(n4131), .ZN(n2991) );
  NAND2_X1 U3782 ( .A1(n4135), .A2(n4118), .ZN(n2993) );
  NOR2_X1 U3783 ( .A1(n3325), .A2(n4100), .ZN(n2994) );
  INV_X1 U3784 ( .A(n3325), .ZN(n4116) );
  INV_X1 U3785 ( .A(n4096), .ZN(n3978) );
  NAND2_X1 U3786 ( .A1(n3978), .A2(n4062), .ZN(n4065) );
  NAND2_X1 U3787 ( .A1(n4096), .A2(n2995), .ZN(n4066) );
  NAND2_X1 U3788 ( .A1(n4065), .A2(n4066), .ZN(n4060) );
  XNOR2_X1 U3789 ( .A(n4061), .B(n2083), .ZN(n4082) );
  XNOR2_X1 U3790 ( .A(n2996), .B(n2997), .ZN(n2998) );
  NAND2_X1 U3791 ( .A1(n2998), .A2(n3241), .ZN(n4232) );
  NAND2_X1 U3792 ( .A1(n2999), .A2(n3048), .ZN(n3893) );
  NAND2_X1 U3793 ( .A1(n3860), .A2(n3000), .ZN(n3196) );
  NAND2_X1 U3794 ( .A1(n3196), .A2(n3897), .ZN(n3002) );
  INV_X1 U3795 ( .A(n3867), .ZN(n3001) );
  NAND2_X1 U3796 ( .A1(n3002), .A2(n3001), .ZN(n3215) );
  NAND2_X1 U3797 ( .A1(n3215), .A2(n3896), .ZN(n3253) );
  NAND2_X1 U3798 ( .A1(n3212), .A2(n3255), .ZN(n3902) );
  NAND2_X1 U3799 ( .A1(n3273), .A2(n3990), .ZN(n3899) );
  NAND2_X1 U3800 ( .A1(n3253), .A2(n3853), .ZN(n3252) );
  NAND2_X1 U3801 ( .A1(n3252), .A2(n3902), .ZN(n3338) );
  INV_X1 U3802 ( .A(n3338), .ZN(n3003) );
  AND2_X1 U3803 ( .A1(n3004), .A2(n3988), .ZN(n3906) );
  NAND2_X1 U3804 ( .A1(n3384), .A2(n3364), .ZN(n3918) );
  NAND2_X1 U3805 ( .A1(n2949), .A2(n3987), .ZN(n3919) );
  NAND2_X1 U3806 ( .A1(n3281), .A2(n3388), .ZN(n3907) );
  NAND2_X1 U3807 ( .A1(n3005), .A2(n3907), .ZN(n3306) );
  INV_X1 U3808 ( .A(n3006), .ZN(n3007) );
  OAI21_X2 U3809 ( .B1(n3306), .B2(n3007), .A(n3913), .ZN(n3419) );
  NAND2_X1 U3810 ( .A1(n3461), .A2(n3426), .ZN(n3914) );
  NAND2_X1 U3811 ( .A1(n3419), .A2(n3914), .ZN(n3008) );
  NAND2_X1 U3812 ( .A1(n2185), .A2(n3985), .ZN(n3912) );
  NAND2_X1 U3813 ( .A1(n3008), .A2(n3912), .ZN(n3459) );
  NAND2_X1 U3814 ( .A1(n3496), .A2(n3466), .ZN(n3915) );
  NAND2_X1 U3815 ( .A1(n3654), .A2(n3983), .ZN(n3926) );
  NAND2_X1 U3816 ( .A1(n3009), .A2(n3498), .ZN(n3925) );
  INV_X1 U3817 ( .A(n3981), .ZN(n3569) );
  OR2_X1 U3818 ( .A1(n3549), .A2(n3569), .ZN(n3564) );
  NAND2_X1 U3819 ( .A1(n3619), .A2(n3980), .ZN(n3011) );
  NAND2_X1 U3820 ( .A1(n3564), .A2(n3011), .ZN(n3013) );
  INV_X1 U3821 ( .A(n3542), .ZN(n3012) );
  NOR2_X1 U3822 ( .A1(n3013), .A2(n3012), .ZN(n3927) );
  INV_X1 U3823 ( .A(n3013), .ZN(n3016) );
  NAND2_X1 U3824 ( .A1(n3549), .A2(n3569), .ZN(n3566) );
  NAND2_X1 U3825 ( .A1(n3566), .A2(n3540), .ZN(n3015) );
  NOR2_X1 U3826 ( .A1(n3619), .A2(n3980), .ZN(n3014) );
  AOI21_X1 U3827 ( .B1(n3016), .B2(n3015), .A(n3014), .ZN(n3928) );
  NAND2_X1 U3828 ( .A1(n3017), .A2(n3928), .ZN(n3584) );
  NAND2_X1 U3829 ( .A1(n3584), .A2(n3859), .ZN(n3585) );
  INV_X1 U3830 ( .A(n3602), .ZN(n3800) );
  OR2_X1 U3831 ( .A1(n4313), .A2(n3800), .ZN(n3810) );
  NAND2_X1 U3832 ( .A1(n4313), .A2(n3800), .ZN(n3809) );
  NAND2_X1 U3833 ( .A1(n3810), .A2(n3809), .ZN(n3857) );
  INV_X1 U3834 ( .A(n3807), .ZN(n3018) );
  NOR2_X1 U3835 ( .A1(n3857), .A2(n3018), .ZN(n3019) );
  NAND2_X1 U3836 ( .A1(n3585), .A2(n3019), .ZN(n3020) );
  NAND2_X1 U3837 ( .A1(n3020), .A2(n3809), .ZN(n4309) );
  NAND2_X1 U3838 ( .A1(n4273), .A2(n4254), .ZN(n3021) );
  NAND2_X1 U3839 ( .A1(n3021), .A2(n4249), .ZN(n3023) );
  INV_X1 U3840 ( .A(n4299), .ZN(n3024) );
  AND2_X1 U3841 ( .A1(n3979), .A2(n3024), .ZN(n4245) );
  INV_X1 U3842 ( .A(n3023), .ZN(n3027) );
  OR2_X1 U3843 ( .A1(n3979), .A2(n3024), .ZN(n4246) );
  NAND2_X1 U3844 ( .A1(n4248), .A2(n4246), .ZN(n3026) );
  NOR2_X1 U3845 ( .A1(n4273), .A2(n4254), .ZN(n3025) );
  AOI21_X1 U3846 ( .B1(n3027), .B2(n3026), .A(n3025), .ZN(n4223) );
  NAND2_X1 U3847 ( .A1(n4206), .A2(n4234), .ZN(n3028) );
  NAND2_X1 U3848 ( .A1(n4224), .A2(n3939), .ZN(n3029) );
  NAND2_X1 U3849 ( .A1(n4252), .A2(n3753), .ZN(n3943) );
  NAND2_X1 U3850 ( .A1(n3029), .A2(n3943), .ZN(n4165) );
  NAND2_X1 U3851 ( .A1(n4228), .A2(n3030), .ZN(n4167) );
  NAND2_X1 U3852 ( .A1(n4191), .A2(n4178), .ZN(n3847) );
  AND2_X1 U3853 ( .A1(n3847), .A2(n3031), .ZN(n3948) );
  AND2_X1 U3854 ( .A1(n4193), .A2(n4215), .ZN(n4166) );
  NAND2_X1 U3855 ( .A1(n4169), .A2(n4166), .ZN(n3032) );
  NAND2_X1 U3856 ( .A1(n3764), .A2(n3053), .ZN(n3848) );
  NOR2_X1 U3857 ( .A1(n4132), .A2(n4157), .ZN(n3846) );
  NAND2_X1 U3858 ( .A1(n3034), .A2(n3033), .ZN(n4127) );
  NAND2_X1 U3859 ( .A1(n4113), .A2(n4136), .ZN(n3887) );
  NAND2_X1 U3860 ( .A1(n4132), .A2(n4157), .ZN(n4126) );
  NAND2_X1 U3861 ( .A1(n4135), .A2(n4112), .ZN(n3844) );
  NAND2_X1 U3862 ( .A1(n4154), .A2(n4131), .ZN(n4107) );
  AND2_X1 U3863 ( .A1(n4094), .A2(n4118), .ZN(n3843) );
  XNOR2_X1 U3864 ( .A(n3325), .B(n4100), .ZN(n4093) );
  NAND2_X1 U3865 ( .A1(n2454), .A2(n4485), .ZN(n3967) );
  NAND2_X1 U3866 ( .A1(n3969), .A2(n4484), .ZN(n3035) );
  OAI22_X1 U3867 ( .A1(n3831), .A2(n4315), .B1(n4253), .B2(n4062), .ZN(n3037)
         );
  AOI21_X1 U3868 ( .B1(n4312), .B2(n3325), .A(n3037), .ZN(n3038) );
  OR2_X1 U3869 ( .A1(n3041), .A2(n3040), .ZN(n3043) );
  INV_X1 U3870 ( .A(n3234), .ZN(n3042) );
  NOR2_X1 U3871 ( .A1(n3043), .A2(n3042), .ZN(n3047) );
  NAND2_X1 U3872 ( .A1(n3236), .A2(n3044), .ZN(n3046) );
  NAND2_X1 U3873 ( .A1(n3294), .A2(n2949), .ZN(n3312) );
  INV_X2 U3874 ( .A(n3312), .ZN(n3050) );
  NOR2_X2 U3875 ( .A1(n4262), .A2(n4263), .ZN(n4233) );
  AND2_X2 U3876 ( .A1(n4233), .A2(n3753), .ZN(n4212) );
  AND2_X2 U3877 ( .A1(n4212), .A2(n4215), .ZN(n4213) );
  NAND2_X2 U3878 ( .A1(n4213), .A2(n4199), .ZN(n4371) );
  OAI21_X1 U3879 ( .B1(n2014), .B2(n4062), .A(n4064), .ZN(n4083) );
  INV_X1 U3880 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3054) );
  OR2_X1 U3881 ( .A1(n4592), .A2(n3054), .ZN(n3055) );
  NAND2_X1 U3882 ( .A1(n3058), .A2(n3057), .ZN(U3546) );
  INV_X1 U3883 ( .A(n3059), .ZN(n3239) );
  INV_X1 U3884 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3061) );
  OR2_X1 U3885 ( .A1(n4586), .A2(n3061), .ZN(n3062) );
  NAND2_X1 U3886 ( .A1(n3065), .A2(n3064), .ZN(U3514) );
  OR2_X2 U3887 ( .A1(n3066), .A2(n4543), .ZN(n3991) );
  INV_X1 U3888 ( .A(n3067), .ZN(n3068) );
  NOR2_X1 U3889 ( .A1(n3069), .A2(n3068), .ZN(n3073) );
  AOI211_X1 U3890 ( .C1(n3070), .C2(n2228), .A(n3749), .B(n3073), .ZN(n3072)
         );
  AOI211_X1 U3891 ( .C1(n3074), .C2(n3073), .A(n3805), .B(n3072), .ZN(n3078)
         );
  NOR2_X1 U3892 ( .A1(n3781), .A2(n4217), .ZN(n3077) );
  OAI22_X1 U3893 ( .A1(n3763), .A2(n4215), .B1(STATE_REG_SCAN_IN), .B2(n4653), 
        .ZN(n3076) );
  OAI22_X1 U3894 ( .A1(n3646), .A2(n3787), .B1(n4206), .B2(n3776), .ZN(n3075)
         );
  OR4_X1 U3895 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(U3220) );
  INV_X1 U3896 ( .A(n3079), .ZN(n3130) );
  INV_X1 U3897 ( .A(DATAI_1_), .ZN(n3080) );
  MUX2_X1 U3898 ( .A(n3130), .B(n3080), .S(U3149), .Z(n3081) );
  INV_X1 U3899 ( .A(n3081), .ZN(U3351) );
  INV_X1 U3900 ( .A(DATAI_15_), .ZN(n4623) );
  NAND2_X1 U3901 ( .A1(n4033), .A2(STATE_REG_SCAN_IN), .ZN(n3082) );
  OAI21_X1 U3902 ( .B1(STATE_REG_SCAN_IN), .B2(n4623), .A(n3082), .ZN(U3337)
         );
  INV_X1 U3903 ( .A(DATAI_4_), .ZN(n3084) );
  MUX2_X1 U3904 ( .A(n3084), .B(n2156), .S(STATE_REG_SCAN_IN), .Z(n3085) );
  INV_X1 U3905 ( .A(n3085), .ZN(U3348) );
  INV_X1 U3906 ( .A(DATAI_29_), .ZN(n3087) );
  NAND2_X1 U3907 ( .A1(n2425), .A2(STATE_REG_SCAN_IN), .ZN(n3086) );
  OAI21_X1 U3908 ( .B1(STATE_REG_SCAN_IN), .B2(n3087), .A(n3086), .ZN(U3323)
         );
  INV_X1 U3909 ( .A(DATAI_6_), .ZN(n3089) );
  MUX2_X1 U3910 ( .A(n3089), .B(n2160), .S(STATE_REG_SCAN_IN), .Z(n3090) );
  INV_X1 U3911 ( .A(n3090), .ZN(U3346) );
  INV_X1 U3912 ( .A(DATAI_19_), .ZN(n3091) );
  MUX2_X1 U3913 ( .A(n3241), .B(n3091), .S(U3149), .Z(n3092) );
  INV_X1 U3914 ( .A(n3092), .ZN(U3333) );
  INV_X1 U3915 ( .A(DATAI_7_), .ZN(n3093) );
  MUX2_X1 U3916 ( .A(n3093), .B(n3154), .S(STATE_REG_SCAN_IN), .Z(n3094) );
  INV_X1 U3917 ( .A(n3094), .ZN(U3345) );
  INV_X1 U3918 ( .A(DATAI_9_), .ZN(n3095) );
  MUX2_X1 U3919 ( .A(n3376), .B(n3095), .S(U3149), .Z(n3096) );
  INV_X1 U3920 ( .A(n3096), .ZN(U3343) );
  INV_X1 U3921 ( .A(n3097), .ZN(n3098) );
  NOR3_X1 U3922 ( .A1(n4483), .A2(n4543), .A3(n4482), .ZN(n3099) );
  AOI21_X1 U3923 ( .B1(n4593), .B2(n3100), .A(n3099), .ZN(U3459) );
  AOI22_X1 U3924 ( .A1(n4593), .A2(n3103), .B1(n3102), .B2(n3101), .ZN(U3458)
         );
  INV_X1 U3925 ( .A(DATAI_12_), .ZN(n3104) );
  MUX2_X1 U3926 ( .A(n3104), .B(n3526), .S(STATE_REG_SCAN_IN), .Z(n3105) );
  INV_X1 U3927 ( .A(n3105), .ZN(U3340) );
  INV_X1 U3928 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U3929 ( .A1(n3822), .A2(REG1_REG_30__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U3930 ( .A1(n3823), .A2(REG2_REG_30__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3931 ( .A1(n3824), .A2(REG0_REG_30__SCAN_IN), .ZN(n3106) );
  NAND3_X1 U3932 ( .A1(n3108), .A2(n3107), .A3(n3106), .ZN(n4072) );
  NAND2_X1 U3933 ( .A1(n4072), .A2(U4043), .ZN(n3109) );
  OAI21_X1 U3934 ( .B1(U4043), .B2(n4723), .A(n3109), .ZN(U3580) );
  INV_X1 U3935 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U3936 ( .A1(n3797), .A2(U4043), .ZN(n3110) );
  OAI21_X1 U3937 ( .B1(U4043), .B2(n4631), .A(n3110), .ZN(U3564) );
  XNOR2_X1 U3938 ( .A(n3111), .B(REG1_REG_3__SCAN_IN), .ZN(n3118) );
  INV_X1 U3939 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3260) );
  XNOR2_X1 U3940 ( .A(n3112), .B(n3260), .ZN(n3116) );
  INV_X1 U3941 ( .A(n4493), .ZN(n3114) );
  AOI22_X1 U3942 ( .A1(n4517), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3113) );
  OAI21_X1 U3943 ( .B1(n3114), .B2(n4529), .A(n3113), .ZN(n3115) );
  AOI21_X1 U3944 ( .B1(n2375), .B2(n3116), .A(n3115), .ZN(n3117) );
  OAI21_X1 U3945 ( .B1(n3118), .B2(n4514), .A(n3117), .ZN(U3243) );
  NOR2_X1 U3946 ( .A1(n2447), .A2(n2254), .ZN(n3170) );
  INV_X1 U3947 ( .A(n3170), .ZN(n3121) );
  AOI211_X1 U3948 ( .C1(n3121), .C2(n3120), .A(n3119), .B(n4014), .ZN(n3127)
         );
  INV_X1 U3949 ( .A(n3122), .ZN(n3125) );
  AOI21_X1 U3950 ( .B1(REG1_REG_0__SCAN_IN), .B2(IR_REG_0__SCAN_IN), .A(n3123), 
        .ZN(n3124) );
  NOR3_X1 U3951 ( .A1(n4514), .A2(n3125), .A3(n3124), .ZN(n3126) );
  NOR2_X1 U3952 ( .A1(n3127), .A2(n3126), .ZN(n3129) );
  AOI22_X1 U3953 ( .A1(n4517), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3128) );
  OAI211_X1 U3954 ( .C1(n3130), .C2(n4529), .A(n3129), .B(n3128), .ZN(U3241)
         );
  AOI211_X1 U3955 ( .C1(n3133), .C2(n3132), .A(n4014), .B(n3131), .ZN(n3140)
         );
  AOI211_X1 U3956 ( .C1(n3135), .C2(n3134), .A(n4514), .B(n2035), .ZN(n3139)
         );
  AND2_X1 U3957 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3283) );
  AOI21_X1 U3958 ( .B1(n4517), .B2(ADDR_REG_5__SCAN_IN), .A(n3283), .ZN(n3136)
         );
  OAI21_X1 U3959 ( .B1(n3137), .B2(n4529), .A(n3136), .ZN(n3138) );
  OR3_X1 U3960 ( .A1(n3140), .A2(n3139), .A3(n3138), .ZN(U3245) );
  INV_X1 U3961 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U3962 ( .A1(n4252), .A2(U4043), .ZN(n3141) );
  OAI21_X1 U3963 ( .B1(U4043), .B2(n4683), .A(n3141), .ZN(U3570) );
  XNOR2_X1 U3964 ( .A(n3142), .B(REG1_REG_6__SCAN_IN), .ZN(n3148) );
  XOR2_X1 U3965 ( .A(n3143), .B(REG2_REG_6__SCAN_IN), .Z(n3146) );
  NOR2_X1 U3966 ( .A1(STATE_REG_SCAN_IN), .A2(n2539), .ZN(n3387) );
  AOI21_X1 U3967 ( .B1(n4517), .B2(ADDR_REG_6__SCAN_IN), .A(n3387), .ZN(n3144)
         );
  OAI21_X1 U3968 ( .B1(n2160), .B2(n4529), .A(n3144), .ZN(n3145) );
  AOI21_X1 U3969 ( .B1(n3146), .B2(n2375), .A(n3145), .ZN(n3147) );
  OAI21_X1 U3970 ( .B1(n3148), .B2(n4514), .A(n3147), .ZN(U3246) );
  INV_X1 U3971 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4639) );
  NAND2_X1 U3972 ( .A1(n4208), .A2(U4043), .ZN(n3149) );
  OAI21_X1 U3973 ( .B1(U4043), .B2(n4639), .A(n3149), .ZN(U3572) );
  MUX2_X1 U3974 ( .A(n2384), .B(REG1_REG_7__SCAN_IN), .S(n3150), .Z(n3152) );
  XOR2_X1 U3975 ( .A(n3152), .B(n3151), .Z(n3159) );
  NAND2_X1 U3976 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U3977 ( .A1(n4517), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3153) );
  OAI211_X1 U3978 ( .C1(n4529), .C2(n3154), .A(n3404), .B(n3153), .ZN(n3158)
         );
  AOI211_X1 U3979 ( .C1(n3156), .C2(n3155), .A(n4014), .B(n2037), .ZN(n3157)
         );
  AOI211_X1 U3980 ( .C1(n3159), .C2(n4510), .A(n3158), .B(n3157), .ZN(n3160)
         );
  INV_X1 U3981 ( .A(n3160), .ZN(U3247) );
  XNOR2_X1 U3982 ( .A(n3161), .B(REG1_REG_4__SCAN_IN), .ZN(n3178) );
  XOR2_X1 U3983 ( .A(n3162), .B(REG2_REG_4__SCAN_IN), .Z(n3176) );
  NAND2_X1 U3984 ( .A1(n4517), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U3985 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3327) );
  OAI211_X1 U3986 ( .C1(n2156), .C2(n4529), .A(n3163), .B(n3327), .ZN(n3175)
         );
  INV_X1 U3987 ( .A(n3165), .ZN(n3166) );
  XNOR2_X1 U3988 ( .A(n3164), .B(n3166), .ZN(n3624) );
  NAND2_X1 U3989 ( .A1(n4481), .A2(n3167), .ZN(n3173) );
  AOI21_X1 U3990 ( .B1(n4495), .B2(n2254), .A(n3168), .ZN(n4496) );
  INV_X1 U3991 ( .A(n4496), .ZN(n3171) );
  INV_X1 U3992 ( .A(n3971), .ZN(n3169) );
  AOI22_X1 U3993 ( .A1(n3171), .A2(n2447), .B1(n3170), .B2(n3169), .ZN(n3172)
         );
  OAI211_X1 U3994 ( .C1(n3624), .C2(n3173), .A(U4043), .B(n3172), .ZN(n4001)
         );
  INV_X1 U3995 ( .A(n4001), .ZN(n3174) );
  AOI211_X1 U3996 ( .C1(n3176), .C2(n2375), .A(n3175), .B(n3174), .ZN(n3177)
         );
  OAI21_X1 U3997 ( .B1(n3178), .B2(n4514), .A(n3177), .ZN(U3244) );
  INV_X1 U3998 ( .A(n3180), .ZN(n3181) );
  AOI21_X1 U3999 ( .B1(n3182), .B2(n3179), .A(n3181), .ZN(n3188) );
  AOI22_X1 U4000 ( .A1(n3778), .A2(n3219), .B1(n3798), .B2(n2938), .ZN(n3187)
         );
  INV_X1 U4001 ( .A(n3183), .ZN(n3185) );
  NAND3_X1 U4002 ( .A1(n3185), .A2(n3235), .A3(n3184), .ZN(n3675) );
  AOI22_X1 U4003 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3675), .B1(n3796), .B2(n3990), .ZN(n3186) );
  OAI211_X1 U4004 ( .C1(n3188), .C2(n3805), .A(n3187), .B(n3186), .ZN(U3234)
         );
  INV_X1 U4005 ( .A(n4558), .ZN(n4566) );
  INV_X1 U4006 ( .A(n3048), .ZN(n3205) );
  NAND2_X1 U4007 ( .A1(n3205), .A2(n3992), .ZN(n3895) );
  AND2_X1 U4008 ( .A1(n3893), .A2(n3895), .ZN(n3879) );
  INV_X1 U4009 ( .A(n3879), .ZN(n4535) );
  NOR2_X1 U4010 ( .A1(n3205), .A2(n3189), .ZN(n4533) );
  INV_X1 U4011 ( .A(n4232), .ZN(n3513) );
  NOR2_X1 U4012 ( .A1(n3513), .A2(n4318), .ZN(n3191) );
  OAI22_X1 U4013 ( .A1(n3191), .A2(n3879), .B1(n3190), .B2(n4315), .ZN(n4531)
         );
  AOI211_X1 U4014 ( .C1(n4566), .C2(n4535), .A(n4533), .B(n4531), .ZN(n4553)
         );
  NAND2_X1 U4015 ( .A1(n4590), .A2(REG1_REG_0__SCAN_IN), .ZN(n3192) );
  OAI21_X1 U4016 ( .B1(n4553), .B2(n4590), .A(n3192), .ZN(U3518) );
  AND2_X1 U4017 ( .A1(n3193), .A2(n3194), .ZN(n3209) );
  NOR2_X1 U4018 ( .A1(n3193), .A2(n3194), .ZN(n3195) );
  OR2_X1 U4019 ( .A1(n3209), .A2(n3195), .ZN(n3301) );
  NAND2_X1 U4020 ( .A1(n3193), .A2(n3893), .ZN(n3197) );
  NAND2_X1 U4021 ( .A1(n3213), .A2(n3197), .ZN(n3202) );
  NAND2_X1 U4022 ( .A1(n4312), .A2(n3992), .ZN(n3200) );
  NAND2_X1 U4023 ( .A1(n4292), .A2(n3198), .ZN(n3199) );
  OAI211_X1 U4024 ( .C1(n3204), .C2(n4253), .A(n3200), .B(n3199), .ZN(n3201)
         );
  AOI21_X1 U4025 ( .B1(n3202), .B2(n4318), .A(n3201), .ZN(n3203) );
  OAI21_X1 U4026 ( .B1(n3301), .B2(n4232), .A(n3203), .ZN(n3299) );
  OAI21_X1 U4027 ( .B1(n3205), .B2(n3204), .A(n2006), .ZN(n3305) );
  OAI22_X1 U4028 ( .A1(n3301), .A2(n4558), .B1(n4557), .B2(n3305), .ZN(n3206)
         );
  NOR2_X1 U4029 ( .A1(n3299), .A2(n3206), .ZN(n4555) );
  NAND2_X1 U4030 ( .A1(n4590), .A2(REG1_REG_1__SCAN_IN), .ZN(n3207) );
  OAI21_X1 U4031 ( .B1(n4555), .B2(n4590), .A(n3207), .ZN(U3519) );
  NOR2_X1 U4032 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  XNOR2_X1 U4033 ( .A(n3210), .B(n3867), .ZN(n3245) );
  INV_X1 U4034 ( .A(n3245), .ZN(n3218) );
  AOI22_X1 U4035 ( .A1(n3219), .A2(n4311), .B1(n4312), .B2(n2938), .ZN(n3211)
         );
  OAI21_X1 U4036 ( .B1(n3212), .B2(n4315), .A(n3211), .ZN(n3217) );
  NAND3_X1 U4037 ( .A1(n3213), .A2(n3897), .A3(n3867), .ZN(n3214) );
  AOI21_X1 U4038 ( .B1(n3215), .B2(n3214), .A(n4210), .ZN(n3216) );
  AOI211_X1 U4039 ( .C1(n3245), .C2(n3513), .A(n3217), .B(n3216), .ZN(n3242)
         );
  OAI21_X1 U4040 ( .B1(n4558), .B2(n3218), .A(n3242), .ZN(n3268) );
  INV_X1 U4041 ( .A(n3250), .ZN(n3221) );
  NAND2_X1 U4042 ( .A1(n2006), .A2(n3219), .ZN(n3220) );
  NAND2_X1 U40430 ( .A1(n3221), .A2(n3220), .ZN(n3266) );
  INV_X1 U4044 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3222) );
  OAI22_X1 U4045 ( .A1(n4478), .A2(n3266), .B1(n4586), .B2(n3222), .ZN(n3223)
         );
  AOI21_X1 U4046 ( .B1(n3268), .B2(n4586), .A(n3223), .ZN(n3224) );
  INV_X1 U4047 ( .A(n3224), .ZN(U3471) );
  XNOR2_X1 U4048 ( .A(n3225), .B(REG2_REG_8__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4049 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3435) );
  INV_X1 U4050 ( .A(n3435), .ZN(n3227) );
  NOR2_X1 U4051 ( .A1(n4529), .A2(n2386), .ZN(n3226) );
  AOI211_X1 U4052 ( .C1(n4517), .C2(ADDR_REG_8__SCAN_IN), .A(n3227), .B(n3226), 
        .ZN(n3232) );
  INV_X1 U4053 ( .A(n3228), .ZN(n3229) );
  OAI211_X1 U4054 ( .C1(REG1_REG_8__SCAN_IN), .C2(n3230), .A(n3229), .B(n4510), 
        .ZN(n3231) );
  OAI211_X1 U4055 ( .C1(n3233), .C2(n4014), .A(n3232), .B(n3231), .ZN(U3248)
         );
  AND3_X1 U4056 ( .A1(n3236), .A2(n3235), .A3(n3234), .ZN(n3237) );
  NAND3_X1 U4057 ( .A1(n3239), .A2(n3238), .A3(n3237), .ZN(n3240) );
  AND2_X1 U4058 ( .A1(n4538), .A2(n3241), .ZN(n4288) );
  INV_X1 U4059 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3243) );
  MUX2_X1 U4060 ( .A(n3243), .B(n3242), .S(n4538), .Z(n3247) );
  NAND2_X1 U4061 ( .A1(n2996), .A2(n3969), .ZN(n3292) );
  INV_X1 U4062 ( .A(n3292), .ZN(n3244) );
  NAND2_X1 U4063 ( .A1(n4538), .A2(n3244), .ZN(n4243) );
  AOI22_X1 U4064 ( .A1(n3245), .A2(n4536), .B1(REG3_REG_2__SCAN_IN), .B2(n4534), .ZN(n3246) );
  OAI211_X1 U4065 ( .C1(n4268), .C2(n3266), .A(n3247), .B(n3246), .ZN(U3288)
         );
  INV_X1 U4066 ( .A(n3248), .ZN(n3249) );
  OAI21_X1 U4067 ( .B1(n3250), .B2(n3273), .A(n3249), .ZN(n4556) );
  XNOR2_X1 U4068 ( .A(n3251), .B(n3853), .ZN(n4559) );
  OAI21_X1 U4069 ( .B1(n3853), .B2(n3253), .A(n3252), .ZN(n3254) );
  NAND2_X1 U4070 ( .A1(n3254), .A2(n4318), .ZN(n3257) );
  AOI22_X1 U4071 ( .A1(n4311), .A2(n3255), .B1(n4312), .B2(n3198), .ZN(n3256)
         );
  OAI211_X1 U4072 ( .C1(n3359), .C2(n4315), .A(n3257), .B(n3256), .ZN(n3258)
         );
  INV_X1 U4073 ( .A(n3258), .ZN(n3259) );
  OAI21_X1 U4074 ( .B1(n4232), .B2(n4559), .A(n3259), .ZN(n4561) );
  NAND2_X1 U4075 ( .A1(n4561), .A2(n4538), .ZN(n3264) );
  INV_X1 U4076 ( .A(n4559), .ZN(n3262) );
  OAI22_X1 U4077 ( .A1(n4538), .A2(n3260), .B1(REG3_REG_3__SCAN_IN), .B2(n4329), .ZN(n3261) );
  AOI21_X1 U4078 ( .B1(n3262), .B2(n4536), .A(n3261), .ZN(n3263) );
  OAI211_X1 U4079 ( .C1(n4268), .C2(n4556), .A(n3264), .B(n3263), .ZN(U3287)
         );
  OAI22_X1 U4080 ( .A1(n4418), .A2(n3266), .B1(n4592), .B2(n3265), .ZN(n3267)
         );
  AOI21_X1 U4081 ( .B1(n3268), .B2(n4592), .A(n3267), .ZN(n3269) );
  INV_X1 U4082 ( .A(n3269), .ZN(U3520) );
  XOR2_X1 U4083 ( .A(n3271), .B(n3270), .Z(n3277) );
  MUX2_X1 U4084 ( .A(n3802), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3275) );
  OAI22_X1 U4085 ( .A1(n3763), .A2(n3273), .B1(n3272), .B2(n3776), .ZN(n3274)
         );
  AOI211_X1 U4086 ( .C1(n3796), .C2(n3989), .A(n3275), .B(n3274), .ZN(n3276)
         );
  OAI21_X1 U4087 ( .B1(n3805), .B2(n3277), .A(n3276), .ZN(U3215) );
  INV_X1 U4088 ( .A(n3365), .ZN(n3286) );
  OAI211_X1 U4089 ( .C1(n3280), .C2(n3279), .A(n3278), .B(n3773), .ZN(n3285)
         );
  OAI22_X1 U4090 ( .A1(n3359), .A2(n3776), .B1(n3787), .B2(n3281), .ZN(n3282)
         );
  AOI211_X1 U4091 ( .C1(n3364), .C2(n3778), .A(n3283), .B(n3282), .ZN(n3284)
         );
  OAI211_X1 U4092 ( .C1(n3781), .C2(n3286), .A(n3285), .B(n3284), .ZN(U3224)
         );
  AND2_X1 U4093 ( .A1(n3907), .A2(n3919), .ZN(n3858) );
  XNOR2_X1 U4094 ( .A(n3287), .B(n3858), .ZN(n3288) );
  NAND2_X1 U4095 ( .A1(n3288), .A2(n4318), .ZN(n3290) );
  AOI22_X1 U4096 ( .A1(n3388), .A2(n4311), .B1(n4312), .B2(n3988), .ZN(n3289)
         );
  OAI211_X1 U4097 ( .C1(n3385), .C2(n4315), .A(n3290), .B(n3289), .ZN(n3393)
         );
  INV_X1 U4098 ( .A(n3393), .ZN(n3298) );
  XNOR2_X1 U4099 ( .A(n3291), .B(n3858), .ZN(n3394) );
  NAND2_X1 U4100 ( .A1(n4232), .A2(n3292), .ZN(n3293) );
  OAI21_X1 U4101 ( .B1(n3294), .B2(n2949), .A(n3312), .ZN(n3398) );
  AOI22_X1 U4102 ( .A1(n4540), .A2(REG2_REG_6__SCAN_IN), .B1(n3389), .B2(n4534), .ZN(n3295) );
  OAI21_X1 U4103 ( .B1(n4268), .B2(n3398), .A(n3295), .ZN(n3296) );
  AOI21_X1 U4104 ( .B1(n3394), .B2(n4333), .A(n3296), .ZN(n3297) );
  OAI21_X1 U4105 ( .B1(n3298), .B2(n4540), .A(n3297), .ZN(U3284) );
  MUX2_X1 U4106 ( .A(n3299), .B(REG2_REG_1__SCAN_IN), .S(n4540), .Z(n3300) );
  INV_X1 U4107 ( .A(n3300), .ZN(n3304) );
  INV_X1 U4108 ( .A(n3301), .ZN(n3302) );
  AOI22_X1 U4109 ( .A1(n4536), .A2(n3302), .B1(REG3_REG_1__SCAN_IN), .B2(n4534), .ZN(n3303) );
  OAI211_X1 U4110 ( .C1(n4268), .C2(n3305), .A(n3304), .B(n3303), .ZN(U3289)
         );
  INV_X1 U4111 ( .A(n3908), .ZN(n3854) );
  XNOR2_X1 U4112 ( .A(n3306), .B(n3854), .ZN(n3310) );
  NAND2_X1 U4113 ( .A1(n4292), .A2(n3985), .ZN(n3308) );
  NAND2_X1 U4114 ( .A1(n4312), .A2(n3987), .ZN(n3307) );
  OAI211_X1 U4115 ( .C1(n3049), .C2(n4253), .A(n3308), .B(n3307), .ZN(n3309)
         );
  AOI21_X1 U4116 ( .B1(n3310), .B2(n4318), .A(n3309), .ZN(n4583) );
  AOI21_X1 U4117 ( .B1(n3312), .B2(n3311), .A(n4557), .ZN(n3313) );
  NAND2_X1 U4118 ( .A1(n3313), .A2(n3425), .ZN(n4580) );
  INV_X1 U4119 ( .A(n4580), .ZN(n3317) );
  INV_X1 U4120 ( .A(n3407), .ZN(n3314) );
  OAI22_X1 U4121 ( .A1(n4538), .A2(n3315), .B1(n3314), .B2(n4329), .ZN(n3316)
         );
  AOI21_X1 U4122 ( .B1(n3317), .B2(n4288), .A(n3316), .ZN(n3324) );
  NAND2_X1 U4123 ( .A1(n3291), .A2(n3987), .ZN(n3318) );
  NAND2_X1 U4124 ( .A1(n3318), .A2(n2949), .ZN(n3320) );
  OR2_X1 U4125 ( .A1(n3291), .A2(n3987), .ZN(n3319) );
  AND2_X1 U4126 ( .A1(n3320), .A2(n3319), .ZN(n3321) );
  NAND2_X1 U4127 ( .A1(n3321), .A2(n3908), .ZN(n4579) );
  INV_X1 U4128 ( .A(n3321), .ZN(n3322) );
  NAND2_X1 U4129 ( .A1(n3322), .A2(n3854), .ZN(n4577) );
  NAND3_X1 U4130 ( .A1(n4579), .A2(n4333), .A3(n4577), .ZN(n3323) );
  OAI211_X1 U4131 ( .C1(n4583), .C2(n4540), .A(n3324), .B(n3323), .ZN(U3283)
         );
  INV_X1 U4132 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U4133 ( .A1(n3325), .A2(U4043), .ZN(n3326) );
  OAI21_X1 U4134 ( .B1(U4043), .B2(n4710), .A(n3326), .ZN(U3577) );
  AOI22_X1 U4135 ( .A1(n3796), .A2(n3988), .B1(n3798), .B2(n3990), .ZN(n3328)
         );
  OAI211_X1 U4136 ( .C1(n3763), .C2(n3336), .A(n3328), .B(n3327), .ZN(n3334)
         );
  INV_X1 U4137 ( .A(n3329), .ZN(n3330) );
  AOI211_X1 U4138 ( .C1(n3332), .C2(n3331), .A(n3805), .B(n3330), .ZN(n3333)
         );
  AOI211_X1 U4139 ( .C1(n3350), .C2(n3802), .A(n3334), .B(n3333), .ZN(n3335)
         );
  INV_X1 U4140 ( .A(n3335), .ZN(U3227) );
  OAI211_X1 U4141 ( .C1(n3248), .C2(n3336), .A(n4575), .B(n3363), .ZN(n4563)
         );
  NOR2_X1 U4142 ( .A1(n4563), .A2(n3969), .ZN(n3349) );
  INV_X1 U4143 ( .A(n3337), .ZN(n3855) );
  XNOR2_X1 U4144 ( .A(n3338), .B(n3855), .ZN(n3347) );
  NAND2_X1 U4145 ( .A1(n3340), .A2(n3339), .ZN(n3341) );
  NOR2_X1 U4146 ( .A1(n3341), .A2(n3855), .ZN(n3354) );
  AND2_X1 U4147 ( .A1(n3341), .A2(n3855), .ZN(n3342) );
  NOR2_X1 U4148 ( .A1(n3354), .A2(n3342), .ZN(n4567) );
  NAND2_X1 U4149 ( .A1(n4567), .A2(n3513), .ZN(n3345) );
  AOI22_X1 U4150 ( .A1(n3343), .A2(n4311), .B1(n4312), .B2(n3990), .ZN(n3344)
         );
  OAI211_X1 U4151 ( .C1(n3384), .C2(n4315), .A(n3345), .B(n3344), .ZN(n3346)
         );
  AOI21_X1 U4152 ( .B1(n3347), .B2(n4318), .A(n3346), .ZN(n3348) );
  INV_X1 U4153 ( .A(n3348), .ZN(n4564) );
  AOI211_X1 U4154 ( .C1(n4534), .C2(n3350), .A(n3349), .B(n4564), .ZN(n3352)
         );
  AOI22_X1 U4155 ( .A1(n4567), .A2(n4536), .B1(REG2_REG_4__SCAN_IN), .B2(n4540), .ZN(n3351) );
  OAI21_X1 U4156 ( .B1(n3352), .B2(n4540), .A(n3351), .ZN(U3286) );
  NOR2_X1 U4157 ( .A1(n3354), .A2(n3353), .ZN(n3356) );
  INV_X1 U4158 ( .A(n3906), .ZN(n3355) );
  AND2_X1 U4159 ( .A1(n3355), .A2(n3918), .ZN(n3866) );
  XNOR2_X1 U4160 ( .A(n3356), .B(n3866), .ZN(n4570) );
  XOR2_X1 U4161 ( .A(n3357), .B(n3866), .Z(n3361) );
  AOI22_X1 U4162 ( .A1(n4311), .A2(n3364), .B1(n4292), .B2(n3987), .ZN(n3358)
         );
  OAI21_X1 U4163 ( .B1(n3359), .B2(n4275), .A(n3358), .ZN(n3360) );
  AOI21_X1 U4164 ( .B1(n3361), .B2(n4318), .A(n3360), .ZN(n4571) );
  INV_X1 U4165 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3362) );
  MUX2_X1 U4166 ( .A(n4571), .B(n3362), .S(n4540), .Z(n3367) );
  AOI21_X1 U4167 ( .B1(n3364), .B2(n3363), .A(n3294), .ZN(n4574) );
  AOI22_X1 U4168 ( .A1(n4574), .A2(n4328), .B1(n3365), .B2(n4534), .ZN(n3366)
         );
  OAI211_X1 U4169 ( .C1(n4285), .C2(n4570), .A(n3367), .B(n3366), .ZN(U3285)
         );
  INV_X1 U4170 ( .A(n3369), .ZN(n3370) );
  AOI211_X1 U4171 ( .C1(n3372), .C2(n3371), .A(n4014), .B(n3370), .ZN(n3379)
         );
  AOI211_X1 U4172 ( .C1(n2034), .C2(n3374), .A(n4514), .B(n3373), .ZN(n3378)
         );
  NAND2_X1 U4173 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U4174 ( .A1(n4517), .A2(ADDR_REG_9__SCAN_IN), .ZN(n3375) );
  OAI211_X1 U4175 ( .C1(n4529), .C2(n3376), .A(n3490), .B(n3375), .ZN(n3377)
         );
  OR3_X1 U4176 ( .A1(n3379), .A2(n3378), .A3(n3377), .ZN(U3249) );
  XOR2_X1 U4177 ( .A(n3381), .B(n3380), .Z(n3382) );
  XNOR2_X1 U4178 ( .A(n3383), .B(n3382), .ZN(n3392) );
  OAI22_X1 U4179 ( .A1(n3385), .A2(n3787), .B1(n3776), .B2(n3384), .ZN(n3386)
         );
  AOI211_X1 U4180 ( .C1(n3388), .C2(n3778), .A(n3387), .B(n3386), .ZN(n3391)
         );
  NAND2_X1 U4181 ( .A1(n3802), .A2(n3389), .ZN(n3390) );
  OAI211_X1 U4182 ( .C1(n3392), .C2(n3805), .A(n3391), .B(n3390), .ZN(U3236)
         );
  AOI21_X1 U4183 ( .B1(n3394), .B2(n4578), .A(n3393), .ZN(n3401) );
  INV_X1 U4184 ( .A(n3398), .ZN(n3395) );
  INV_X1 U4185 ( .A(n4478), .ZN(n4459) );
  AOI22_X1 U4186 ( .A1(n3395), .A2(n4459), .B1(n4584), .B2(REG0_REG_6__SCAN_IN), .ZN(n3396) );
  OAI21_X1 U4187 ( .B1(n3401), .B2(n4584), .A(n3396), .ZN(U3479) );
  INV_X1 U4188 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3397) );
  OAI22_X1 U4189 ( .A1(n3398), .A2(n4418), .B1(n4592), .B2(n3397), .ZN(n3399)
         );
  INV_X1 U4190 ( .A(n3399), .ZN(n3400) );
  OAI21_X1 U4191 ( .B1(n3401), .B2(n4590), .A(n3400), .ZN(U3524) );
  XNOR2_X1 U4192 ( .A(n3403), .B(n3402), .ZN(n3409) );
  AOI22_X1 U4193 ( .A1(n3798), .A2(n3987), .B1(n3796), .B2(n3985), .ZN(n3405)
         );
  OAI211_X1 U4194 ( .C1(n3763), .C2(n3049), .A(n3405), .B(n3404), .ZN(n3406)
         );
  AOI21_X1 U4195 ( .B1(n3407), .B2(n3802), .A(n3406), .ZN(n3408) );
  OAI21_X1 U4196 ( .B1(n3409), .B2(n3805), .A(n3408), .ZN(U3210) );
  XNOR2_X1 U4197 ( .A(n3410), .B(REG2_REG_10__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4198 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4199 ( .A1(n4517), .A2(ADDR_REG_10__SCAN_IN), .ZN(n3411) );
  OAI211_X1 U4200 ( .C1(n4529), .C2(n3412), .A(n3652), .B(n3411), .ZN(n3413)
         );
  INV_X1 U4201 ( .A(n3413), .ZN(n3417) );
  OAI211_X1 U4202 ( .C1(n3415), .C2(REG1_REG_10__SCAN_IN), .A(n3414), .B(n4510), .ZN(n3416) );
  OAI211_X1 U4203 ( .C1(n3418), .C2(n4014), .A(n3417), .B(n3416), .ZN(U3250)
         );
  NAND2_X1 U4204 ( .A1(n3914), .A2(n3912), .ZN(n3877) );
  XNOR2_X1 U4205 ( .A(n3419), .B(n3877), .ZN(n3420) );
  NAND2_X1 U4206 ( .A1(n3420), .A2(n4318), .ZN(n3422) );
  AOI22_X1 U4207 ( .A1(n4292), .A2(n3984), .B1(n4312), .B2(n3986), .ZN(n3421)
         );
  OAI211_X1 U4208 ( .C1(n4253), .C2(n2185), .A(n3422), .B(n3421), .ZN(n3441)
         );
  INV_X1 U4209 ( .A(n3441), .ZN(n3431) );
  XOR2_X1 U4210 ( .A(n3423), .B(n3877), .Z(n3442) );
  INV_X1 U4211 ( .A(n3465), .ZN(n3424) );
  AOI21_X1 U4212 ( .B1(n3426), .B2(n3425), .A(n3424), .ZN(n3444) );
  INV_X1 U4213 ( .A(n3444), .ZN(n3428) );
  AOI22_X1 U4214 ( .A1(n4540), .A2(REG2_REG_8__SCAN_IN), .B1(n3438), .B2(n4534), .ZN(n3427) );
  OAI21_X1 U4215 ( .B1(n3428), .B2(n4268), .A(n3427), .ZN(n3429) );
  AOI21_X1 U4216 ( .B1(n3442), .B2(n4333), .A(n3429), .ZN(n3430) );
  OAI21_X1 U4217 ( .B1(n3431), .B2(n4540), .A(n3430), .ZN(U3282) );
  INV_X1 U4218 ( .A(n3486), .ZN(n3433) );
  NOR2_X1 U4219 ( .A1(n3433), .A2(n3485), .ZN(n3434) );
  XNOR2_X1 U4220 ( .A(n3432), .B(n3434), .ZN(n3440) );
  AOI22_X1 U4221 ( .A1(n3796), .A2(n3984), .B1(n3798), .B2(n3986), .ZN(n3436)
         );
  OAI211_X1 U4222 ( .C1(n3763), .C2(n2185), .A(n3436), .B(n3435), .ZN(n3437)
         );
  AOI21_X1 U4223 ( .B1(n3438), .B2(n3802), .A(n3437), .ZN(n3439) );
  OAI21_X1 U4224 ( .B1(n3440), .B2(n3805), .A(n3439), .ZN(U3218) );
  AOI21_X1 U4225 ( .B1(n3442), .B2(n4578), .A(n3441), .ZN(n3446) );
  INV_X1 U4226 ( .A(n4418), .ZN(n4396) );
  AOI22_X1 U4227 ( .A1(n3444), .A2(n4396), .B1(REG1_REG_8__SCAN_IN), .B2(n4590), .ZN(n3443) );
  OAI21_X1 U4228 ( .B1(n3446), .B2(n4590), .A(n3443), .ZN(U3526) );
  AOI22_X1 U4229 ( .A1(n3444), .A2(n4459), .B1(REG0_REG_8__SCAN_IN), .B2(n4584), .ZN(n3445) );
  OAI21_X1 U4230 ( .B1(n3446), .B2(n4584), .A(n3445), .ZN(U3483) );
  AOI21_X1 U4231 ( .B1(n3448), .B2(n3447), .A(n4014), .ZN(n3452) );
  NAND2_X1 U4232 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3479) );
  NAND2_X1 U4233 ( .A1(n4517), .A2(ADDR_REG_11__SCAN_IN), .ZN(n3449) );
  OAI211_X1 U4234 ( .C1(n4529), .C2(n4489), .A(n3479), .B(n3449), .ZN(n3450)
         );
  AOI21_X1 U4235 ( .B1(n3452), .B2(n3451), .A(n3450), .ZN(n3457) );
  OAI211_X1 U4236 ( .C1(n3455), .C2(n3454), .A(n3453), .B(n4510), .ZN(n3456)
         );
  NAND2_X1 U4237 ( .A1(n3457), .A2(n3456), .ZN(U3251) );
  NAND2_X1 U4238 ( .A1(n2028), .A2(n3915), .ZN(n3868) );
  XNOR2_X1 U4239 ( .A(n3458), .B(n3868), .ZN(n3474) );
  XNOR2_X1 U4240 ( .A(n3459), .B(n3868), .ZN(n3463) );
  AOI22_X1 U4241 ( .A1(n4311), .A2(n3466), .B1(n4292), .B2(n3983), .ZN(n3460)
         );
  OAI21_X1 U4242 ( .B1(n3461), .B2(n4275), .A(n3460), .ZN(n3462) );
  AOI21_X1 U4243 ( .B1(n3463), .B2(n4318), .A(n3462), .ZN(n3470) );
  OAI21_X1 U4244 ( .B1(n4569), .B2(n3474), .A(n3470), .ZN(n3464) );
  INV_X1 U4245 ( .A(n3464), .ZN(n3469) );
  AOI21_X1 U4246 ( .B1(n3466), .B2(n3465), .A(n2033), .ZN(n3471) );
  AOI22_X1 U4247 ( .A1(n3471), .A2(n4459), .B1(REG0_REG_9__SCAN_IN), .B2(n4584), .ZN(n3467) );
  OAI21_X1 U4248 ( .B1(n3469), .B2(n4584), .A(n3467), .ZN(U3485) );
  AOI22_X1 U4249 ( .A1(n3471), .A2(n4396), .B1(REG1_REG_9__SCAN_IN), .B2(n4590), .ZN(n3468) );
  OAI21_X1 U4250 ( .B1(n3469), .B2(n4590), .A(n3468), .ZN(U3527) );
  MUX2_X1 U4251 ( .A(n4624), .B(n3470), .S(n4538), .Z(n3473) );
  AOI22_X1 U4252 ( .A1(n3471), .A2(n4328), .B1(n2248), .B2(n4534), .ZN(n3472)
         );
  OAI211_X1 U4253 ( .C1(n4285), .C2(n3474), .A(n3473), .B(n3472), .ZN(U3281)
         );
  XOR2_X1 U4254 ( .A(n3476), .B(n3475), .Z(n3477) );
  XNOR2_X1 U4255 ( .A(n3478), .B(n3477), .ZN(n3484) );
  AOI22_X1 U4256 ( .A1(n3798), .A2(n3983), .B1(n3796), .B2(n3981), .ZN(n3480)
         );
  OAI211_X1 U4257 ( .C1(n3763), .C2(n3481), .A(n3480), .B(n3479), .ZN(n3482)
         );
  AOI21_X1 U4258 ( .B1(n3519), .B2(n3802), .A(n3482), .ZN(n3483) );
  OAI21_X1 U4259 ( .B1(n3484), .B2(n3805), .A(n3483), .ZN(U3233) );
  OR2_X1 U4260 ( .A1(n3432), .A2(n3485), .ZN(n3487) );
  NAND2_X1 U4261 ( .A1(n3487), .A2(n3486), .ZN(n3488) );
  XOR2_X1 U4262 ( .A(n3489), .B(n3488), .Z(n3494) );
  AOI22_X1 U4263 ( .A1(n3798), .A2(n3985), .B1(n3796), .B2(n3983), .ZN(n3491)
         );
  OAI211_X1 U4264 ( .C1(n3763), .C2(n2184), .A(n3491), .B(n3490), .ZN(n3492)
         );
  AOI21_X1 U4265 ( .B1(n2248), .B2(n3802), .A(n3492), .ZN(n3493) );
  OAI21_X1 U4266 ( .B1(n3494), .B2(n3805), .A(n3493), .ZN(U3228) );
  AND2_X1 U4267 ( .A1(n3925), .A2(n3926), .ZN(n3865) );
  XOR2_X1 U4268 ( .A(n3865), .B(n3495), .Z(n3500) );
  OAI22_X1 U4269 ( .A1(n3496), .A2(n4275), .B1(n3543), .B2(n4315), .ZN(n3497)
         );
  AOI21_X1 U4270 ( .B1(n3498), .B2(n4311), .A(n3497), .ZN(n3499) );
  OAI21_X1 U4271 ( .B1(n3500), .B2(n4210), .A(n3499), .ZN(n3533) );
  INV_X1 U4272 ( .A(n3533), .ZN(n3507) );
  XNOR2_X1 U4273 ( .A(n3501), .B(n3865), .ZN(n3534) );
  OR2_X1 U4274 ( .A1(n2033), .A2(n3654), .ZN(n3503) );
  NAND2_X1 U4275 ( .A1(n3502), .A2(n3503), .ZN(n3539) );
  AOI22_X1 U4276 ( .A1(n4540), .A2(REG2_REG_10__SCAN_IN), .B1(n3664), .B2(
        n4534), .ZN(n3504) );
  OAI21_X1 U4277 ( .B1(n3539), .B2(n4268), .A(n3504), .ZN(n3505) );
  AOI21_X1 U4278 ( .B1(n3534), .B2(n4333), .A(n3505), .ZN(n3506) );
  OAI21_X1 U4279 ( .B1(n3507), .B2(n4540), .A(n3506), .ZN(U3280) );
  XNOR2_X1 U4280 ( .A(n3508), .B(n3852), .ZN(n3515) );
  OAI21_X1 U4281 ( .B1(n3510), .B2(n3852), .A(n3509), .ZN(n3557) );
  AOI22_X1 U4282 ( .A1(n3517), .A2(n4311), .B1(n4312), .B2(n3983), .ZN(n3511)
         );
  OAI21_X1 U4283 ( .B1(n3569), .B2(n4315), .A(n3511), .ZN(n3512) );
  AOI21_X1 U4284 ( .B1(n3557), .B2(n3513), .A(n3512), .ZN(n3514) );
  OAI21_X1 U4285 ( .B1(n3515), .B2(n4210), .A(n3514), .ZN(n3556) );
  INV_X1 U4286 ( .A(n3556), .ZN(n3523) );
  INV_X1 U4287 ( .A(n3516), .ZN(n3548) );
  NAND2_X1 U4288 ( .A1(n3502), .A2(n3517), .ZN(n3518) );
  NAND2_X1 U4289 ( .A1(n3548), .A2(n3518), .ZN(n3563) );
  AOI22_X1 U4290 ( .A1(n4540), .A2(REG2_REG_11__SCAN_IN), .B1(n3519), .B2(
        n4534), .ZN(n3520) );
  OAI21_X1 U4291 ( .B1(n3563), .B2(n4268), .A(n3520), .ZN(n3521) );
  AOI21_X1 U4292 ( .B1(n3557), .B2(n4536), .A(n3521), .ZN(n3522) );
  OAI21_X1 U4293 ( .B1(n3523), .B2(n4540), .A(n3522), .ZN(U3279) );
  XNOR2_X1 U4294 ( .A(n3524), .B(REG2_REG_12__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U4295 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3687) );
  NAND2_X1 U4296 ( .A1(n4517), .A2(ADDR_REG_12__SCAN_IN), .ZN(n3525) );
  OAI211_X1 U4297 ( .C1(n4529), .C2(n3526), .A(n3687), .B(n3525), .ZN(n3527)
         );
  INV_X1 U4298 ( .A(n3527), .ZN(n3531) );
  OAI211_X1 U4299 ( .C1(n3529), .C2(REG1_REG_12__SCAN_IN), .A(n3528), .B(n4510), .ZN(n3530) );
  OAI211_X1 U4300 ( .C1(n3532), .C2(n4014), .A(n3531), .B(n3530), .ZN(U3252)
         );
  INV_X1 U4301 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3535) );
  AOI21_X1 U4302 ( .B1(n4578), .B2(n3534), .A(n3533), .ZN(n3537) );
  MUX2_X1 U4303 ( .A(n3535), .B(n3537), .S(n4586), .Z(n3536) );
  OAI21_X1 U4304 ( .B1(n3539), .B2(n4478), .A(n3536), .ZN(U3487) );
  MUX2_X1 U4305 ( .A(n2166), .B(n3537), .S(n4592), .Z(n3538) );
  OAI21_X1 U4306 ( .B1(n4418), .B2(n3539), .A(n3538), .ZN(U3528) );
  NAND2_X1 U4307 ( .A1(n3564), .A2(n3566), .ZN(n3849) );
  INV_X1 U4308 ( .A(n3540), .ZN(n3541) );
  AOI21_X1 U4309 ( .B1(n3508), .B2(n3542), .A(n3541), .ZN(n3567) );
  XOR2_X1 U4310 ( .A(n3849), .B(n3567), .Z(n3546) );
  OAI22_X1 U4311 ( .A1(n3543), .A2(n4275), .B1(n3582), .B2(n4315), .ZN(n3544)
         );
  AOI21_X1 U4312 ( .B1(n3549), .B2(n4311), .A(n3544), .ZN(n3545) );
  OAI21_X1 U4313 ( .B1(n3546), .B2(n4210), .A(n3545), .ZN(n4415) );
  INV_X1 U4314 ( .A(n4415), .ZN(n3555) );
  XNOR2_X1 U4315 ( .A(n3547), .B(n3849), .ZN(n4416) );
  INV_X1 U4316 ( .A(n3550), .ZN(n3551) );
  OAI21_X1 U4317 ( .B1(n3516), .B2(n3051), .A(n3551), .ZN(n4479) );
  AOI22_X1 U4318 ( .A1(n4540), .A2(REG2_REG_12__SCAN_IN), .B1(n3690), .B2(
        n4534), .ZN(n3552) );
  OAI21_X1 U4319 ( .B1(n4479), .B2(n4268), .A(n3552), .ZN(n3553) );
  AOI21_X1 U4320 ( .B1(n4416), .B2(n4333), .A(n3553), .ZN(n3554) );
  OAI21_X1 U4321 ( .B1(n3555), .B2(n4540), .A(n3554), .ZN(U3278) );
  INV_X1 U4322 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3558) );
  AOI21_X1 U4323 ( .B1(n4566), .B2(n3557), .A(n3556), .ZN(n3560) );
  MUX2_X1 U4324 ( .A(n3558), .B(n3560), .S(n4586), .Z(n3559) );
  OAI21_X1 U4325 ( .B1(n3563), .B2(n4478), .A(n3559), .ZN(U3489) );
  MUX2_X1 U4326 ( .A(n3561), .B(n3560), .S(n4592), .Z(n3562) );
  OAI21_X1 U4327 ( .B1(n4418), .B2(n3563), .A(n3562), .ZN(U3529) );
  INV_X1 U4328 ( .A(n3564), .ZN(n3565) );
  AOI21_X1 U4329 ( .B1(n3567), .B2(n3566), .A(n3565), .ZN(n3568) );
  XNOR2_X1 U4330 ( .A(n3619), .B(n3980), .ZN(n3881) );
  XNOR2_X1 U4331 ( .A(n3568), .B(n3881), .ZN(n3574) );
  OAI22_X1 U4332 ( .A1(n3569), .A2(n4275), .B1(n3619), .B2(n4253), .ZN(n3572)
         );
  XOR2_X1 U4333 ( .A(n3881), .B(n3570), .Z(n3575) );
  NOR2_X1 U4334 ( .A1(n3575), .A2(n4232), .ZN(n3571) );
  AOI211_X1 U4335 ( .C1(n4292), .C2(n3797), .A(n3572), .B(n3571), .ZN(n3573)
         );
  OAI21_X1 U4336 ( .B1(n4210), .B2(n3574), .A(n3573), .ZN(n4411) );
  INV_X1 U4337 ( .A(n4411), .ZN(n3580) );
  INV_X1 U4338 ( .A(n3575), .ZN(n4412) );
  NOR2_X1 U4339 ( .A1(n3550), .A2(n3619), .ZN(n3576) );
  OR2_X1 U4340 ( .A1(n3590), .A2(n3576), .ZN(n4474) );
  AOI22_X1 U4341 ( .A1(n4540), .A2(REG2_REG_13__SCAN_IN), .B1(n3621), .B2(
        n4534), .ZN(n3577) );
  OAI21_X1 U4342 ( .B1(n4474), .B2(n4268), .A(n3577), .ZN(n3578) );
  AOI21_X1 U4343 ( .B1(n4412), .B2(n4536), .A(n3578), .ZN(n3579) );
  OAI21_X1 U4344 ( .B1(n3580), .B2(n4540), .A(n3579), .ZN(U3277) );
  AOI21_X1 U4345 ( .B1(n3859), .B2(n3581), .A(n2030), .ZN(n3589) );
  OAI22_X1 U4346 ( .A1(n3582), .A2(n4275), .B1(n3637), .B2(n4253), .ZN(n3583)
         );
  AOI21_X1 U4347 ( .B1(n4292), .B2(n4313), .A(n3583), .ZN(n3588) );
  OAI21_X1 U4348 ( .B1(n3859), .B2(n3811), .A(n3585), .ZN(n3586) );
  NAND2_X1 U4349 ( .A1(n3586), .A2(n4318), .ZN(n3587) );
  OAI211_X1 U4350 ( .C1(n3589), .C2(n4232), .A(n3588), .B(n3587), .ZN(n4407)
         );
  INV_X1 U4351 ( .A(n4407), .ZN(n3595) );
  INV_X1 U4352 ( .A(n3589), .ZN(n4408) );
  OR2_X1 U4353 ( .A1(n3590), .A2(n3637), .ZN(n3591) );
  NAND2_X1 U4354 ( .A1(n3603), .A2(n3591), .ZN(n4470) );
  AOI22_X1 U4355 ( .A1(n4540), .A2(REG2_REG_14__SCAN_IN), .B1(n3639), .B2(
        n4534), .ZN(n3592) );
  OAI21_X1 U4356 ( .B1(n4470), .B2(n4268), .A(n3592), .ZN(n3593) );
  AOI21_X1 U4357 ( .B1(n4408), .B2(n4536), .A(n3593), .ZN(n3594) );
  OAI21_X1 U4358 ( .B1(n3595), .B2(n4540), .A(n3594), .ZN(U3276) );
  NAND2_X1 U4359 ( .A1(n3585), .A2(n3807), .ZN(n3596) );
  XNOR2_X1 U4360 ( .A(n3596), .B(n3857), .ZN(n3599) );
  INV_X1 U4361 ( .A(n4291), .ZN(n3734) );
  OAI22_X1 U4362 ( .A1(n3734), .A2(n4315), .B1(n4253), .B2(n3800), .ZN(n3597)
         );
  AOI21_X1 U4363 ( .B1(n4312), .B2(n3797), .A(n3597), .ZN(n3598) );
  OAI21_X1 U4364 ( .B1(n3599), .B2(n4210), .A(n3598), .ZN(n4403) );
  INV_X1 U4365 ( .A(n4403), .ZN(n3609) );
  XNOR2_X1 U4366 ( .A(n3600), .B(n3857), .ZN(n4404) );
  NAND2_X1 U4367 ( .A1(n3603), .A2(n3602), .ZN(n3604) );
  NAND2_X1 U4368 ( .A1(n3601), .A2(n3604), .ZN(n4466) );
  INV_X1 U4369 ( .A(n3605), .ZN(n3803) );
  AOI22_X1 U4370 ( .A1(n4540), .A2(REG2_REG_15__SCAN_IN), .B1(n3803), .B2(
        n4534), .ZN(n3606) );
  OAI21_X1 U4371 ( .B1(n4466), .B2(n4268), .A(n3606), .ZN(n3607) );
  AOI21_X1 U4372 ( .B1(n4404), .B2(n4333), .A(n3607), .ZN(n3608) );
  OAI21_X1 U4373 ( .B1(n3609), .B2(n4540), .A(n3608), .ZN(U3275) );
  AND2_X1 U4374 ( .A1(n4031), .A2(n3991), .ZN(U3148) );
  INV_X1 U4375 ( .A(n3610), .ZN(n3613) );
  NAND3_X1 U4376 ( .A1(n4594), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3612) );
  INV_X1 U4377 ( .A(DATAI_31_), .ZN(n3611) );
  OAI22_X1 U4378 ( .A1(n3613), .A2(n3612), .B1(STATE_REG_SCAN_IN), .B2(n3611), 
        .ZN(U3321) );
  XOR2_X1 U4379 ( .A(n3615), .B(n3614), .Z(n3616) );
  XNOR2_X1 U4380 ( .A(n3617), .B(n3616), .ZN(n3623) );
  AOI22_X1 U4381 ( .A1(n3798), .A2(n3981), .B1(n3796), .B2(n3797), .ZN(n3618)
         );
  NAND2_X1 U4382 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4006) );
  OAI211_X1 U4383 ( .C1(n3763), .C2(n3619), .A(n3618), .B(n4006), .ZN(n3620)
         );
  AOI21_X1 U4384 ( .B1(n3621), .B2(n3802), .A(n3620), .ZN(n3622) );
  OAI21_X1 U4385 ( .B1(n3623), .B2(n3805), .A(n3622), .ZN(U3231) );
  AOI22_X1 U4386 ( .A1(n3778), .A2(n3048), .B1(n3773), .B2(n3624), .ZN(n3626)
         );
  NAND2_X1 U4387 ( .A1(n3675), .A2(REG3_REG_0__SCAN_IN), .ZN(n3625) );
  OAI211_X1 U4388 ( .C1(n3190), .C2(n3787), .A(n3626), .B(n3625), .ZN(U3229)
         );
  XNOR2_X1 U4389 ( .A(n3628), .B(n3627), .ZN(n3634) );
  OAI22_X1 U4390 ( .A1(n3763), .A2(n3630), .B1(STATE_REG_SCAN_IN), .B2(n3629), 
        .ZN(n3632) );
  OAI22_X1 U4391 ( .A1(n4096), .A2(n3787), .B1(n4135), .B2(n3776), .ZN(n3631)
         );
  AOI211_X1 U4392 ( .C1(n4099), .C2(n3802), .A(n3632), .B(n3631), .ZN(n3633)
         );
  OAI21_X1 U4393 ( .B1(n3634), .B2(n3805), .A(n3633), .ZN(U3211) );
  NAND2_X1 U4394 ( .A1(n3712), .A2(n3711), .ZN(n3635) );
  XNOR2_X1 U4395 ( .A(n2007), .B(n3635), .ZN(n3641) );
  AOI22_X1 U4396 ( .A1(n3798), .A2(n3980), .B1(n3796), .B2(n4313), .ZN(n3636)
         );
  NAND2_X1 U4397 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4018) );
  OAI211_X1 U4398 ( .C1(n3763), .C2(n3637), .A(n3636), .B(n4018), .ZN(n3638)
         );
  AOI21_X1 U4399 ( .B1(n3639), .B2(n3802), .A(n3638), .ZN(n3640) );
  OAI21_X1 U4400 ( .B1(n3641), .B2(n3805), .A(n3640), .ZN(U3212) );
  NAND2_X1 U4401 ( .A1(n3697), .A2(n3773), .ZN(n3651) );
  AOI21_X1 U4402 ( .B1(n3642), .B2(n3644), .A(n3643), .ZN(n3650) );
  OAI22_X1 U4403 ( .A1(n3763), .A2(n4178), .B1(STATE_REG_SCAN_IN), .B2(n3645), 
        .ZN(n3648) );
  INV_X1 U4404 ( .A(n4132), .ZN(n4173) );
  OAI22_X1 U4405 ( .A1(n4173), .A2(n3787), .B1(n3646), .B2(n3776), .ZN(n3647)
         );
  AOI211_X1 U4406 ( .C1(n4180), .C2(n3802), .A(n3648), .B(n3647), .ZN(n3649)
         );
  OAI21_X1 U4407 ( .B1(n3651), .B2(n3650), .A(n3649), .ZN(U3213) );
  AOI22_X1 U4408 ( .A1(n3798), .A2(n3984), .B1(n3796), .B2(n3982), .ZN(n3653)
         );
  OAI211_X1 U4409 ( .C1(n3763), .C2(n3654), .A(n3653), .B(n3652), .ZN(n3663)
         );
  OR2_X1 U4410 ( .A1(n3432), .A2(n3655), .ZN(n3658) );
  NAND2_X1 U4411 ( .A1(n3658), .A2(n3656), .ZN(n3660) );
  AND2_X1 U4412 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  AOI211_X1 U4413 ( .C1(n3661), .C2(n3660), .A(n3805), .B(n3659), .ZN(n3662)
         );
  AOI211_X1 U4414 ( .C1(n3664), .C2(n3802), .A(n3663), .B(n3662), .ZN(n3665)
         );
  INV_X1 U4415 ( .A(n3665), .ZN(U3214) );
  AOI21_X1 U4416 ( .B1(n3668), .B2(n3667), .A(n3666), .ZN(n3673) );
  AOI22_X1 U4417 ( .A1(n3798), .A2(n4293), .B1(n3796), .B2(n4252), .ZN(n3670)
         );
  OAI211_X1 U4418 ( .C1(n3763), .C2(n4254), .A(n3670), .B(n3669), .ZN(n3671)
         );
  AOI21_X1 U4419 ( .B1(n4266), .B2(n3802), .A(n3671), .ZN(n3672) );
  OAI21_X1 U4420 ( .B1(n3673), .B2(n3805), .A(n3672), .ZN(U3216) );
  AOI22_X1 U4421 ( .A1(n3778), .A2(n3674), .B1(n3798), .B2(n3992), .ZN(n3681)
         );
  AOI22_X1 U4422 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3675), .B1(n3796), .B2(n3198), .ZN(n3680) );
  OAI211_X1 U4423 ( .C1(n3676), .C2(n3677), .A(n3678), .B(n3773), .ZN(n3679)
         );
  NAND3_X1 U4424 ( .A1(n3681), .A2(n3680), .A3(n3679), .ZN(U3219) );
  INV_X1 U4425 ( .A(n3683), .ZN(n3685) );
  NOR2_X1 U4426 ( .A1(n3685), .A2(n3684), .ZN(n3686) );
  XNOR2_X1 U4427 ( .A(n3682), .B(n3686), .ZN(n3692) );
  AOI22_X1 U4428 ( .A1(n3798), .A2(n3982), .B1(n3796), .B2(n3980), .ZN(n3688)
         );
  OAI211_X1 U4429 ( .C1(n3763), .C2(n3051), .A(n3688), .B(n3687), .ZN(n3689)
         );
  AOI21_X1 U4430 ( .B1(n3690), .B2(n3802), .A(n3689), .ZN(n3691) );
  OAI21_X1 U4431 ( .B1(n3692), .B2(n3805), .A(n3691), .ZN(U3221) );
  INV_X1 U4432 ( .A(n3693), .ZN(n3694) );
  NAND2_X1 U4433 ( .A1(n3697), .A2(n3694), .ZN(n3740) );
  AOI21_X1 U4434 ( .B1(n3697), .B2(n3696), .A(n3695), .ZN(n3742) );
  AOI21_X1 U4435 ( .B1(n3743), .B2(n3740), .A(n3742), .ZN(n3702) );
  OAI21_X1 U4436 ( .B1(n3700), .B2(n3699), .A(n3698), .ZN(n3701) );
  XNOR2_X1 U4437 ( .A(n3702), .B(n3701), .ZN(n3708) );
  INV_X1 U4438 ( .A(n3703), .ZN(n4137) );
  OAI22_X1 U4439 ( .A1(n3763), .A2(n4136), .B1(STATE_REG_SCAN_IN), .B2(n3704), 
        .ZN(n3706) );
  OAI22_X1 U4440 ( .A1(n4135), .A2(n3787), .B1(n4173), .B2(n3776), .ZN(n3705)
         );
  AOI211_X1 U4441 ( .C1(n4137), .C2(n3802), .A(n3706), .B(n3705), .ZN(n3707)
         );
  OAI21_X1 U4442 ( .B1(n3708), .B2(n3805), .A(n3707), .ZN(U3222) );
  NAND2_X1 U4443 ( .A1(n3710), .A2(n3709), .ZN(n3717) );
  NAND2_X1 U4444 ( .A1(n2007), .A2(n3711), .ZN(n3725) );
  NAND2_X1 U4445 ( .A1(n3725), .A2(n3712), .ZN(n3715) );
  INV_X1 U4446 ( .A(n3713), .ZN(n3714) );
  NOR2_X1 U4447 ( .A1(n3715), .A2(n3714), .ZN(n3793) );
  NAND2_X1 U4448 ( .A1(n3715), .A2(n3714), .ZN(n3791) );
  OAI21_X1 U4449 ( .B1(n3793), .B2(n3794), .A(n3791), .ZN(n3716) );
  XOR2_X1 U4450 ( .A(n3717), .B(n3716), .Z(n3718) );
  NAND2_X1 U4451 ( .A1(n3718), .A2(n3773), .ZN(n3723) );
  NOR2_X1 U4452 ( .A1(n3719), .A2(STATE_REG_SCAN_IN), .ZN(n4043) );
  INV_X1 U4453 ( .A(n4313), .ZN(n3720) );
  INV_X1 U4454 ( .A(n3979), .ZN(n4316) );
  OAI22_X1 U4455 ( .A1(n3720), .A2(n3776), .B1(n3787), .B2(n4316), .ZN(n3721)
         );
  AOI211_X1 U4456 ( .C1(n4327), .C2(n3778), .A(n4043), .B(n3721), .ZN(n3722)
         );
  OAI211_X1 U4457 ( .C1(n3781), .C2(n4330), .A(n3723), .B(n3722), .ZN(U3223)
         );
  NAND2_X1 U4458 ( .A1(n3725), .A2(n3724), .ZN(n3727) );
  NAND2_X1 U4459 ( .A1(n3727), .A2(n3726), .ZN(n3732) );
  INV_X1 U4460 ( .A(n3728), .ZN(n3730) );
  NOR2_X1 U4461 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  XNOR2_X1 U4462 ( .A(n3732), .B(n3731), .ZN(n3739) );
  NOR2_X1 U4463 ( .A1(n3733), .A2(STATE_REG_SCAN_IN), .ZN(n4502) );
  INV_X1 U4464 ( .A(n4293), .ZN(n3735) );
  OAI22_X1 U4465 ( .A1(n3735), .A2(n3787), .B1(n3776), .B2(n3734), .ZN(n3736)
         );
  AOI211_X1 U4466 ( .C1(n4299), .C2(n3778), .A(n4502), .B(n3736), .ZN(n3738)
         );
  NAND2_X1 U4467 ( .A1(n3802), .A2(n4300), .ZN(n3737) );
  OAI211_X1 U4468 ( .C1(n3739), .C2(n3805), .A(n3738), .B(n3737), .ZN(U3225)
         );
  INV_X1 U4469 ( .A(n3740), .ZN(n3741) );
  NOR2_X1 U4470 ( .A1(n3742), .A2(n3741), .ZN(n3744) );
  XNOR2_X1 U4471 ( .A(n3744), .B(n3743), .ZN(n3748) );
  OAI22_X1 U4472 ( .A1(n3763), .A2(n4157), .B1(STATE_REG_SCAN_IN), .B2(n4651), 
        .ZN(n3746) );
  OAI22_X1 U4473 ( .A1(n4154), .A2(n3787), .B1(n3764), .B2(n3776), .ZN(n3745)
         );
  AOI211_X1 U4474 ( .C1(n4158), .C2(n3802), .A(n3746), .B(n3745), .ZN(n3747)
         );
  OAI21_X1 U4475 ( .B1(n3748), .B2(n3805), .A(n3747), .ZN(U3226) );
  NAND2_X1 U4476 ( .A1(n2226), .A2(n2228), .ZN(n3750) );
  AOI22_X1 U4477 ( .A1(n3751), .A2(n2228), .B1(n3070), .B2(n3750), .ZN(n3758)
         );
  INV_X1 U4478 ( .A(n4237), .ZN(n3756) );
  INV_X1 U4479 ( .A(n4273), .ZN(n3775) );
  OAI22_X1 U4480 ( .A1(n4228), .A2(n3787), .B1(n3775), .B2(n3776), .ZN(n3755)
         );
  OAI22_X1 U4481 ( .A1(n3763), .A2(n3753), .B1(STATE_REG_SCAN_IN), .B2(n3752), 
        .ZN(n3754) );
  AOI211_X1 U4482 ( .C1(n3756), .C2(n3802), .A(n3755), .B(n3754), .ZN(n3757)
         );
  OAI21_X1 U4483 ( .B1(n3758), .B2(n3805), .A(n3757), .ZN(U3230) );
  OAI21_X1 U4484 ( .B1(n3760), .B2(n3759), .A(n3642), .ZN(n3761) );
  NAND2_X1 U4485 ( .A1(n3761), .A2(n3773), .ZN(n3768) );
  OAI22_X1 U4486 ( .A1(n3763), .A2(n4199), .B1(STATE_REG_SCAN_IN), .B2(n3762), 
        .ZN(n3766) );
  OAI22_X1 U4487 ( .A1(n3764), .A2(n3787), .B1(n4228), .B2(n3776), .ZN(n3765)
         );
  AOI211_X1 U4488 ( .C1(n4198), .C2(n3802), .A(n3766), .B(n3765), .ZN(n3767)
         );
  NAND2_X1 U4489 ( .A1(n3768), .A2(n3767), .ZN(U3232) );
  XNOR2_X1 U4490 ( .A(n3771), .B(n3770), .ZN(n3772) );
  XNOR2_X1 U4491 ( .A(n2735), .B(n3772), .ZN(n3774) );
  NAND2_X1 U4492 ( .A1(n3774), .A2(n3773), .ZN(n3780) );
  AND2_X1 U4493 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4518) );
  OAI22_X1 U4494 ( .A1(n4316), .A2(n3776), .B1(n3787), .B2(n3775), .ZN(n3777)
         );
  AOI211_X1 U4495 ( .C1(n4272), .C2(n3778), .A(n4518), .B(n3777), .ZN(n3779)
         );
  OAI211_X1 U4496 ( .C1(n3781), .C2(n4279), .A(n3780), .B(n3779), .ZN(U3235)
         );
  NAND2_X1 U4497 ( .A1(n2031), .A2(n3783), .ZN(n3784) );
  XNOR2_X1 U4498 ( .A(n3782), .B(n3784), .ZN(n3790) );
  OAI22_X1 U4499 ( .A1(n3763), .A2(n4118), .B1(STATE_REG_SCAN_IN), .B2(n4668), 
        .ZN(n3785) );
  AOI21_X1 U4500 ( .B1(n4113), .B2(n3798), .A(n3785), .ZN(n3786) );
  OAI21_X1 U4501 ( .B1(n4116), .B2(n3787), .A(n3786), .ZN(n3788) );
  AOI21_X1 U4502 ( .B1(n4120), .B2(n3802), .A(n3788), .ZN(n3789) );
  OAI21_X1 U4503 ( .B1(n3790), .B2(n3805), .A(n3789), .ZN(U3237) );
  INV_X1 U4504 ( .A(n3791), .ZN(n3792) );
  NOR2_X1 U4505 ( .A1(n3793), .A2(n3792), .ZN(n3795) );
  XNOR2_X1 U4506 ( .A(n3795), .B(n3794), .ZN(n3806) );
  AOI22_X1 U4507 ( .A1(n3798), .A2(n3797), .B1(n3796), .B2(n4291), .ZN(n3799)
         );
  NAND2_X1 U4508 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4030) );
  OAI211_X1 U4509 ( .C1(n3763), .C2(n3800), .A(n3799), .B(n4030), .ZN(n3801)
         );
  AOI21_X1 U4510 ( .B1(n3803), .B2(n3802), .A(n3801), .ZN(n3804) );
  OAI21_X1 U4511 ( .B1(n3806), .B2(n3805), .A(n3804), .ZN(U3238) );
  NAND2_X1 U4512 ( .A1(n3810), .A2(n3807), .ZN(n3930) );
  NAND2_X1 U4513 ( .A1(n3809), .A2(n3808), .ZN(n3917) );
  NAND2_X1 U4514 ( .A1(n3917), .A2(n3810), .ZN(n3929) );
  OAI21_X1 U4515 ( .B1(n3811), .B2(n3930), .A(n3929), .ZN(n3813) );
  INV_X1 U4516 ( .A(n3937), .ZN(n3812) );
  AOI211_X1 U4517 ( .C1(n3813), .C2(n3935), .A(n3812), .B(n3940), .ZN(n3815)
         );
  INV_X1 U4518 ( .A(n3939), .ZN(n3814) );
  OAI21_X1 U4519 ( .B1(n3815), .B2(n3814), .A(n3943), .ZN(n3818) );
  INV_X1 U4520 ( .A(n3816), .ZN(n3817) );
  AOI21_X1 U4521 ( .B1(n3818), .B2(n3945), .A(n3817), .ZN(n3820) );
  INV_X1 U4522 ( .A(n3848), .ZN(n3819) );
  OR2_X1 U4523 ( .A1(n3846), .A2(n3819), .ZN(n3947) );
  OAI21_X1 U4524 ( .B1(n3820), .B2(n3947), .A(n3950), .ZN(n3830) );
  AND2_X1 U4525 ( .A1(n2012), .A2(n4066), .ZN(n3835) );
  NAND2_X1 U4526 ( .A1(n3821), .A2(DATAI_29_), .ZN(n3832) );
  NAND2_X1 U4527 ( .A1(n3831), .A2(n4071), .ZN(n3841) );
  NAND2_X1 U4528 ( .A1(n3821), .A2(DATAI_30_), .ZN(n4057) );
  OR2_X1 U4529 ( .A1(n4072), .A2(n4057), .ZN(n3875) );
  NAND2_X1 U4530 ( .A1(n3822), .A2(REG1_REG_31__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4531 ( .A1(n3823), .A2(REG2_REG_31__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4532 ( .A1(n3824), .A2(REG0_REG_31__SCAN_IN), .ZN(n3825) );
  NAND3_X1 U4533 ( .A1(n3827), .A2(n3826), .A3(n3825), .ZN(n4051) );
  NAND2_X1 U4534 ( .A1(n3828), .A2(DATAI_31_), .ZN(n4052) );
  NAND2_X1 U4535 ( .A1(n4051), .A2(n4052), .ZN(n3959) );
  AND2_X1 U4536 ( .A1(n3875), .A2(n3959), .ZN(n3829) );
  AND2_X1 U4537 ( .A1(n3841), .A2(n3829), .ZN(n3833) );
  NAND4_X1 U4538 ( .A1(n3830), .A2(n3951), .A3(n3835), .A4(n3833), .ZN(n3840)
         );
  INV_X1 U4539 ( .A(n4052), .ZN(n3837) );
  AND2_X1 U4540 ( .A1(n4072), .A2(n4057), .ZN(n3864) );
  NOR2_X1 U4541 ( .A1(n4051), .A2(n4052), .ZN(n3873) );
  INV_X1 U4542 ( .A(n3831), .ZN(n3977) );
  NAND2_X1 U4543 ( .A1(n3977), .A2(n3832), .ZN(n3842) );
  NAND2_X1 U4544 ( .A1(n4065), .A2(n3842), .ZN(n3834) );
  NOR2_X1 U4545 ( .A1(n3834), .A2(n3843), .ZN(n3953) );
  OAI21_X1 U4546 ( .B1(n3835), .B2(n3834), .A(n3833), .ZN(n3955) );
  AOI21_X1 U4547 ( .B1(n4093), .B2(n3953), .A(n3955), .ZN(n3836) );
  AOI211_X1 U4548 ( .C1(n3837), .C2(n3864), .A(n3873), .B(n3836), .ZN(n3839)
         );
  INV_X1 U4549 ( .A(n4057), .ZN(n3838) );
  AOI22_X1 U4550 ( .A1(n3840), .A2(n3839), .B1(n3838), .B2(n4052), .ZN(n3968)
         );
  NAND2_X1 U4551 ( .A1(n3842), .A2(n3841), .ZN(n4341) );
  NAND2_X1 U4552 ( .A1(n2084), .A2(n3844), .ZN(n4110) );
  INV_X1 U4553 ( .A(n4110), .ZN(n3890) );
  INV_X1 U4554 ( .A(n4126), .ZN(n3845) );
  OR2_X1 U4555 ( .A1(n3846), .A2(n3845), .ZN(n4149) );
  NAND2_X1 U4556 ( .A1(n3848), .A2(n3847), .ZN(n4172) );
  INV_X1 U4557 ( .A(n4166), .ZN(n3942) );
  NAND2_X1 U4558 ( .A1(n3942), .A2(n4167), .ZN(n4205) );
  OR3_X1 U4559 ( .A1(n4172), .A2(n4205), .A3(n3849), .ZN(n3886) );
  NAND2_X1 U4560 ( .A1(n3851), .A2(n3850), .ZN(n4225) );
  INV_X1 U4561 ( .A(n3852), .ZN(n3856) );
  NAND4_X1 U4562 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3863)
         );
  INV_X1 U4563 ( .A(n3857), .ZN(n3861) );
  NAND4_X1 U4564 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3862)
         );
  NOR2_X1 U4565 ( .A1(n3863), .A2(n3862), .ZN(n3871) );
  INV_X1 U4566 ( .A(n3864), .ZN(n3956) );
  AND4_X1 U4567 ( .A1(n3866), .A2(n3865), .A3(n3959), .A4(n3956), .ZN(n3870)
         );
  NOR2_X1 U4568 ( .A1(n3868), .A2(n3867), .ZN(n3869) );
  NAND4_X1 U4569 ( .A1(n3871), .A2(n4284), .A3(n3870), .A4(n3869), .ZN(n3872)
         );
  XNOR2_X1 U4570 ( .A(n4273), .B(n4254), .ZN(n4260) );
  NOR2_X1 U4571 ( .A1(n3872), .A2(n4260), .ZN(n3884) );
  INV_X1 U4572 ( .A(n3873), .ZN(n3957) );
  NAND3_X1 U4573 ( .A1(n3957), .A2(n3875), .A3(n3874), .ZN(n3876) );
  NOR2_X1 U4574 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  AND3_X1 U4575 ( .A1(n4310), .A2(n3879), .A3(n3878), .ZN(n3883) );
  INV_X1 U4576 ( .A(n4245), .ZN(n3880) );
  NAND2_X1 U4577 ( .A1(n3880), .A2(n4246), .ZN(n4305) );
  NOR2_X1 U4578 ( .A1(n4305), .A2(n3881), .ZN(n3882) );
  NAND4_X1 U4579 ( .A1(n4225), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3885)
         );
  NOR3_X1 U4580 ( .A1(n4149), .A2(n3886), .A3(n3885), .ZN(n3889) );
  NAND2_X1 U4581 ( .A1(n4107), .A2(n3887), .ZN(n4128) );
  INV_X1 U4582 ( .A(n4189), .ZN(n4187) );
  NOR2_X1 U4583 ( .A1(n4128), .A2(n4187), .ZN(n3888) );
  NAND4_X1 U4584 ( .A1(n4069), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3892)
         );
  INV_X1 U4585 ( .A(n4093), .ZN(n3891) );
  NOR3_X1 U4586 ( .A1(n3892), .A2(n4060), .A3(n3891), .ZN(n3964) );
  OAI211_X1 U4587 ( .C1(n3000), .C2(n2454), .A(n3895), .B(n3894), .ZN(n3898)
         );
  NAND3_X1 U4588 ( .A1(n3898), .A2(n3897), .A3(n3896), .ZN(n3901) );
  NAND3_X1 U4589 ( .A1(n3901), .A2(n3900), .A3(n3899), .ZN(n3904) );
  NAND3_X1 U4590 ( .A1(n3904), .A2(n3903), .A3(n3902), .ZN(n3911) );
  NOR3_X1 U4591 ( .A1(n2065), .A2(n2072), .A3(n3906), .ZN(n3910) );
  INV_X1 U4592 ( .A(n3907), .ZN(n3909) );
  AOI211_X1 U4593 ( .C1(n3911), .C2(n3910), .A(n3909), .B(n3908), .ZN(n3916)
         );
  NAND2_X1 U4594 ( .A1(n3913), .A2(n3912), .ZN(n3920) );
  OAI211_X1 U4595 ( .C1(n3916), .C2(n3920), .A(n3915), .B(n3914), .ZN(n3924)
         );
  INV_X1 U4596 ( .A(n3917), .ZN(n3923) );
  NAND2_X1 U4597 ( .A1(n2068), .A2(n3919), .ZN(n3921) );
  OAI21_X1 U4598 ( .B1(n3921), .B2(n3920), .A(n3925), .ZN(n3922) );
  AOI22_X1 U4599 ( .A1(n3924), .A2(n3923), .B1(n3929), .B2(n3922), .ZN(n3934)
         );
  OAI211_X1 U4600 ( .C1(n2057), .C2(n2028), .A(n3927), .B(n3926), .ZN(n3933)
         );
  INV_X1 U4601 ( .A(n3928), .ZN(n3931) );
  OAI21_X1 U4602 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n3932) );
  OAI21_X1 U4603 ( .B1(n3934), .B2(n3933), .A(n3932), .ZN(n3938) );
  INV_X1 U4604 ( .A(n3935), .ZN(n3936) );
  AOI21_X1 U4605 ( .B1(n3938), .B2(n3937), .A(n3936), .ZN(n3941) );
  OAI21_X1 U4606 ( .B1(n3941), .B2(n3940), .A(n3939), .ZN(n3944) );
  NAND3_X1 U4607 ( .A1(n3944), .A2(n3943), .A3(n3942), .ZN(n3946) );
  NAND2_X1 U4608 ( .A1(n3946), .A2(n3945), .ZN(n3949) );
  AOI21_X1 U4609 ( .B1(n3949), .B2(n3948), .A(n3947), .ZN(n3952) );
  OAI21_X1 U4610 ( .B1(n3952), .B2(n2076), .A(n3951), .ZN(n3954) );
  OAI211_X1 U4611 ( .C1(n4116), .C2(n4100), .A(n3954), .B(n3953), .ZN(n3961)
         );
  INV_X1 U4612 ( .A(n3955), .ZN(n3960) );
  NAND2_X1 U4613 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  AOI22_X1 U4614 ( .A1(n3961), .A2(n3960), .B1(n3959), .B2(n3958), .ZN(n3963)
         );
  MUX2_X1 U4615 ( .A(n3964), .B(n3963), .S(n3962), .Z(n3965) );
  INV_X1 U4616 ( .A(n3965), .ZN(n3966) );
  OAI21_X1 U4617 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n3970) );
  XNOR2_X1 U4618 ( .A(n3970), .B(n3969), .ZN(n3976) );
  NOR2_X1 U4619 ( .A1(n3972), .A2(n3971), .ZN(n3974) );
  OAI21_X1 U4620 ( .B1(n3975), .B2(n4484), .A(B_REG_SCAN_IN), .ZN(n3973) );
  OAI22_X1 U4621 ( .A1(n3976), .A2(n3975), .B1(n3974), .B2(n3973), .ZN(U3239)
         );
  MUX2_X1 U4622 ( .A(n4051), .B(DATAO_REG_31__SCAN_IN), .S(n3991), .Z(U3581)
         );
  MUX2_X1 U4623 ( .A(n3977), .B(DATAO_REG_29__SCAN_IN), .S(n3991), .Z(U3579)
         );
  MUX2_X1 U4624 ( .A(n3978), .B(DATAO_REG_28__SCAN_IN), .S(n3991), .Z(U3578)
         );
  MUX2_X1 U4625 ( .A(n4094), .B(DATAO_REG_26__SCAN_IN), .S(n3991), .Z(U3576)
         );
  MUX2_X1 U4626 ( .A(n4113), .B(DATAO_REG_25__SCAN_IN), .S(n3991), .Z(U3575)
         );
  MUX2_X1 U4627 ( .A(n4132), .B(DATAO_REG_24__SCAN_IN), .S(n3991), .Z(U3574)
         );
  MUX2_X1 U4628 ( .A(n4191), .B(DATAO_REG_23__SCAN_IN), .S(n3991), .Z(U3573)
         );
  MUX2_X1 U4629 ( .A(n4193), .B(DATAO_REG_21__SCAN_IN), .S(n3991), .Z(U3571)
         );
  MUX2_X1 U4630 ( .A(n4273), .B(DATAO_REG_19__SCAN_IN), .S(n3991), .Z(U3569)
         );
  MUX2_X1 U4631 ( .A(n4293), .B(DATAO_REG_18__SCAN_IN), .S(n3991), .Z(U3568)
         );
  MUX2_X1 U4632 ( .A(n3979), .B(DATAO_REG_17__SCAN_IN), .S(n3991), .Z(U3567)
         );
  MUX2_X1 U4633 ( .A(n4291), .B(DATAO_REG_16__SCAN_IN), .S(n3991), .Z(U3566)
         );
  MUX2_X1 U4634 ( .A(n4313), .B(DATAO_REG_15__SCAN_IN), .S(n3991), .Z(U3565)
         );
  MUX2_X1 U4635 ( .A(n3980), .B(DATAO_REG_13__SCAN_IN), .S(n3991), .Z(U3563)
         );
  MUX2_X1 U4636 ( .A(n3981), .B(DATAO_REG_12__SCAN_IN), .S(n3991), .Z(U3562)
         );
  MUX2_X1 U4637 ( .A(n3982), .B(DATAO_REG_11__SCAN_IN), .S(n3991), .Z(U3561)
         );
  MUX2_X1 U4638 ( .A(n3983), .B(DATAO_REG_10__SCAN_IN), .S(n3991), .Z(U3560)
         );
  MUX2_X1 U4639 ( .A(n3984), .B(DATAO_REG_9__SCAN_IN), .S(n3991), .Z(U3559) );
  MUX2_X1 U4640 ( .A(n3985), .B(DATAO_REG_8__SCAN_IN), .S(n3991), .Z(U3558) );
  MUX2_X1 U4641 ( .A(n3986), .B(DATAO_REG_7__SCAN_IN), .S(n3991), .Z(U3557) );
  MUX2_X1 U4642 ( .A(n3987), .B(DATAO_REG_6__SCAN_IN), .S(n3991), .Z(U3556) );
  MUX2_X1 U4643 ( .A(n3988), .B(DATAO_REG_5__SCAN_IN), .S(n3991), .Z(U3555) );
  MUX2_X1 U4644 ( .A(n3989), .B(DATAO_REG_4__SCAN_IN), .S(n3991), .Z(U3554) );
  MUX2_X1 U4645 ( .A(n3990), .B(DATAO_REG_3__SCAN_IN), .S(n3991), .Z(U3553) );
  MUX2_X1 U4646 ( .A(n3198), .B(DATAO_REG_2__SCAN_IN), .S(n3991), .Z(U3552) );
  MUX2_X1 U4647 ( .A(n2938), .B(DATAO_REG_1__SCAN_IN), .S(n3991), .Z(U3551) );
  MUX2_X1 U4648 ( .A(n3992), .B(DATAO_REG_0__SCAN_IN), .S(n3991), .Z(U3550) );
  INV_X1 U4649 ( .A(n4529), .ZN(n4034) );
  XNOR2_X1 U4650 ( .A(n3994), .B(n3993), .ZN(n3995) );
  NOR2_X1 U4651 ( .A1(n4514), .A2(n3995), .ZN(n4000) );
  AOI211_X1 U4652 ( .C1(n3998), .C2(n3997), .A(n3996), .B(n4014), .ZN(n3999)
         );
  AOI211_X1 U4653 ( .C1(n4034), .C2(n2379), .A(n4000), .B(n3999), .ZN(n4003)
         );
  AOI22_X1 U4654 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4517), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4002) );
  NAND3_X1 U4655 ( .A1(n4003), .A2(n4002), .A3(n4001), .ZN(U3242) );
  XNOR2_X1 U4656 ( .A(n4488), .B(REG2_REG_13__SCAN_IN), .ZN(n4005) );
  XNOR2_X1 U4657 ( .A(n4004), .B(n4005), .ZN(n4015) );
  INV_X1 U4658 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4007) );
  OAI21_X1 U4659 ( .B1(n4031), .B2(n4007), .A(n4006), .ZN(n4008) );
  AOI21_X1 U4660 ( .B1(n4034), .B2(n4488), .A(n4008), .ZN(n4013) );
  OAI211_X1 U4661 ( .C1(n4011), .C2(n4010), .A(n4009), .B(n4510), .ZN(n4012)
         );
  OAI211_X1 U4662 ( .C1(n4015), .C2(n4014), .A(n4013), .B(n4012), .ZN(U3253)
         );
  OAI211_X1 U4663 ( .C1(n4017), .C2(REG2_REG_14__SCAN_IN), .A(n4016), .B(n2375), .ZN(n4026) );
  INV_X1 U4664 ( .A(n4018), .ZN(n4021) );
  NOR2_X1 U4665 ( .A1(n4529), .A2(n4019), .ZN(n4020) );
  AOI211_X1 U4666 ( .C1(n4517), .C2(ADDR_REG_14__SCAN_IN), .A(n4021), .B(n4020), .ZN(n4025) );
  OAI211_X1 U4667 ( .C1(n4023), .C2(REG1_REG_14__SCAN_IN), .A(n4022), .B(n4510), .ZN(n4024) );
  NAND3_X1 U4668 ( .A1(n4026), .A2(n4025), .A3(n4024), .ZN(U3254) );
  OAI211_X1 U4669 ( .C1(n4029), .C2(n4028), .A(n4027), .B(n2375), .ZN(n4040)
         );
  INV_X1 U4670 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U4671 ( .B1(n4031), .B2(n4662), .A(n4030), .ZN(n4032) );
  AOI21_X1 U4672 ( .B1(n4034), .B2(n4033), .A(n4032), .ZN(n4039) );
  OAI211_X1 U4673 ( .C1(n4037), .C2(n4036), .A(n4035), .B(n4510), .ZN(n4038)
         );
  NAND3_X1 U4674 ( .A1(n4040), .A2(n4039), .A3(n4038), .ZN(U3255) );
  XOR2_X1 U4675 ( .A(REG1_REG_16__SCAN_IN), .B(n4041), .Z(n4049) );
  XOR2_X1 U4676 ( .A(n2323), .B(n4042), .Z(n4047) );
  INV_X1 U4677 ( .A(n4486), .ZN(n4045) );
  AOI21_X1 U4678 ( .B1(n4517), .B2(ADDR_REG_16__SCAN_IN), .A(n4043), .ZN(n4044) );
  OAI21_X1 U4679 ( .B1(n4045), .B2(n4529), .A(n4044), .ZN(n4046) );
  AOI21_X1 U4680 ( .B1(n4047), .B2(n2375), .A(n4046), .ZN(n4048) );
  OAI21_X1 U4681 ( .B1(n4049), .B2(n4514), .A(n4048), .ZN(U3256) );
  AND2_X1 U4682 ( .A1(n4495), .A2(B_REG_SCAN_IN), .ZN(n4050) );
  NOR2_X1 U4683 ( .A1(n4315), .A2(n4050), .ZN(n4073) );
  NAND2_X1 U4684 ( .A1(n4073), .A2(n4051), .ZN(n4056) );
  OAI21_X1 U4685 ( .B1(n4052), .B2(n4253), .A(n4056), .ZN(n4419) );
  NAND2_X1 U4686 ( .A1(n4538), .A2(n4419), .ZN(n4054) );
  NAND2_X1 U4687 ( .A1(n4540), .A2(REG2_REG_31__SCAN_IN), .ZN(n4053) );
  OAI211_X1 U4688 ( .C1(n4422), .C2(n4268), .A(n4054), .B(n4053), .ZN(U3260)
         );
  OAI21_X1 U4689 ( .B1(n4057), .B2(n4253), .A(n4056), .ZN(n4423) );
  NAND2_X1 U4690 ( .A1(n4538), .A2(n4423), .ZN(n4059) );
  NAND2_X1 U4691 ( .A1(n4540), .A2(REG2_REG_30__SCAN_IN), .ZN(n4058) );
  OAI211_X1 U4692 ( .C1(n4426), .C2(n4268), .A(n4059), .B(n4058), .ZN(U3261)
         );
  NOR2_X1 U4693 ( .A1(n4096), .A2(n4062), .ZN(n4344) );
  NOR2_X1 U4694 ( .A1(n4342), .A2(n4344), .ZN(n4340) );
  XOR2_X1 U4695 ( .A(n4341), .B(n4340), .Z(n4081) );
  AOI21_X1 U4696 ( .B1(n4071), .B2(n4064), .A(n4063), .ZN(n4345) );
  AOI22_X1 U4697 ( .A1(n4345), .A2(n4328), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4540), .ZN(n4080) );
  INV_X1 U4698 ( .A(n4065), .ZN(n4067) );
  OAI21_X1 U4699 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n4070) );
  XNOR2_X1 U4700 ( .A(n4070), .B(n4069), .ZN(n4076) );
  AOI22_X1 U4701 ( .A1(n4073), .A2(n4072), .B1(n4311), .B2(n4071), .ZN(n4074)
         );
  OAI21_X1 U4702 ( .B1(n4096), .B2(n4275), .A(n4074), .ZN(n4075) );
  OAI21_X1 U4703 ( .B1(n4329), .B2(n4077), .A(n4348), .ZN(n4078) );
  NAND2_X1 U4704 ( .A1(n4078), .A2(n4538), .ZN(n4079) );
  OAI211_X1 U4705 ( .C1(n4081), .C2(n4285), .A(n4080), .B(n4079), .ZN(U3354)
         );
  INV_X1 U4706 ( .A(n4082), .ZN(n4090) );
  NOR2_X1 U4707 ( .A1(n4083), .A2(n4268), .ZN(n4087) );
  OAI22_X1 U4708 ( .A1(n4085), .A2(n4329), .B1(n4084), .B2(n4538), .ZN(n4086)
         );
  AOI211_X1 U4709 ( .C1(n4088), .C2(n4538), .A(n4087), .B(n4086), .ZN(n4089)
         );
  OAI21_X1 U4710 ( .B1(n4090), .B2(n4285), .A(n4089), .ZN(U3262) );
  XNOR2_X1 U4711 ( .A(n4091), .B(n4093), .ZN(n4354) );
  XNOR2_X1 U4712 ( .A(n4092), .B(n4093), .ZN(n4098) );
  AOI22_X1 U4713 ( .A1(n4094), .A2(n4312), .B1(n4100), .B2(n4311), .ZN(n4095)
         );
  OAI21_X1 U4714 ( .B1(n4096), .B2(n4315), .A(n4095), .ZN(n4097) );
  AOI21_X1 U4715 ( .B1(n4098), .B2(n4318), .A(n4097), .ZN(n4353) );
  AOI22_X1 U4716 ( .A1(n4099), .A2(n4534), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4540), .ZN(n4103) );
  AND2_X1 U4717 ( .A1(n2009), .A2(n4100), .ZN(n4101) );
  NOR2_X1 U4718 ( .A1(n2014), .A2(n4101), .ZN(n4351) );
  NAND2_X1 U4719 ( .A1(n4351), .A2(n4328), .ZN(n4102) );
  OAI211_X1 U4720 ( .C1(n4353), .C2(n4540), .A(n4103), .B(n4102), .ZN(n4104)
         );
  INV_X1 U4721 ( .A(n4104), .ZN(n4105) );
  OAI21_X1 U4722 ( .B1(n4354), .B2(n4285), .A(n4105), .ZN(U3263) );
  XOR2_X1 U4723 ( .A(n4110), .B(n4106), .Z(n4356) );
  INV_X1 U4724 ( .A(n4356), .ZN(n4124) );
  NAND2_X1 U4725 ( .A1(n4108), .A2(n4107), .ZN(n4109) );
  XOR2_X1 U4726 ( .A(n4110), .B(n4109), .Z(n4111) );
  NAND2_X1 U4727 ( .A1(n4111), .A2(n4318), .ZN(n4115) );
  AOI22_X1 U4728 ( .A1(n4113), .A2(n4312), .B1(n4112), .B2(n4311), .ZN(n4114)
         );
  OAI211_X1 U4729 ( .C1(n4116), .C2(n4315), .A(n4115), .B(n4114), .ZN(n4355)
         );
  INV_X1 U4730 ( .A(n4117), .ZN(n4119) );
  OAI21_X1 U4731 ( .B1(n4119), .B2(n4118), .A(n2009), .ZN(n4432) );
  AOI22_X1 U4732 ( .A1(n4120), .A2(n4534), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4540), .ZN(n4121) );
  OAI21_X1 U4733 ( .B1(n4432), .B2(n4268), .A(n4121), .ZN(n4122) );
  AOI21_X1 U4734 ( .B1(n4355), .B2(n4538), .A(n4122), .ZN(n4123) );
  OAI21_X1 U4735 ( .B1(n4124), .B2(n4285), .A(n4123), .ZN(U3264) );
  XNOR2_X1 U4736 ( .A(n4125), .B(n4128), .ZN(n4360) );
  INV_X1 U4737 ( .A(n4360), .ZN(n4141) );
  NAND2_X1 U4738 ( .A1(n4127), .A2(n4126), .ZN(n4129) );
  XNOR2_X1 U4739 ( .A(n4129), .B(n4128), .ZN(n4130) );
  NAND2_X1 U4740 ( .A1(n4130), .A2(n4318), .ZN(n4134) );
  AOI22_X1 U4741 ( .A1(n4132), .A2(n4312), .B1(n4311), .B2(n4131), .ZN(n4133)
         );
  OAI211_X1 U4742 ( .C1(n4135), .C2(n4315), .A(n4134), .B(n4133), .ZN(n4359)
         );
  OAI21_X1 U4743 ( .B1(n2245), .B2(n4136), .A(n4117), .ZN(n4435) );
  AOI22_X1 U4744 ( .A1(n4137), .A2(n4534), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4540), .ZN(n4138) );
  OAI21_X1 U4745 ( .B1(n4435), .B2(n4268), .A(n4138), .ZN(n4139) );
  AOI21_X1 U4746 ( .B1(n4359), .B2(n4538), .A(n4139), .ZN(n4140) );
  OAI21_X1 U4747 ( .B1(n4141), .B2(n4285), .A(n4140), .ZN(U3265) );
  NAND2_X1 U4748 ( .A1(n4143), .A2(n4142), .ZN(n4185) );
  NAND2_X1 U4749 ( .A1(n4186), .A2(n4144), .ZN(n4146) );
  XOR2_X1 U4750 ( .A(n4149), .B(n4147), .Z(n4364) );
  INV_X1 U4751 ( .A(n4364), .ZN(n4162) );
  XOR2_X1 U4752 ( .A(n4149), .B(n4148), .Z(n4150) );
  NAND2_X1 U4753 ( .A1(n4150), .A2(n4318), .ZN(n4153) );
  AOI22_X1 U4754 ( .A1(n4191), .A2(n4312), .B1(n4311), .B2(n4151), .ZN(n4152)
         );
  OAI211_X1 U4755 ( .C1(n4154), .C2(n4315), .A(n4153), .B(n4152), .ZN(n4363)
         );
  INV_X1 U4756 ( .A(n4155), .ZN(n4177) );
  INV_X1 U4757 ( .A(n2245), .ZN(n4156) );
  OAI21_X1 U4758 ( .B1(n4155), .B2(n4157), .A(n4156), .ZN(n4438) );
  AOI22_X1 U4759 ( .A1(n4158), .A2(n4534), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4540), .ZN(n4159) );
  OAI21_X1 U4760 ( .B1(n4438), .B2(n4268), .A(n4159), .ZN(n4160) );
  AOI21_X1 U4761 ( .B1(n4538), .B2(n4363), .A(n4160), .ZN(n4161) );
  OAI21_X1 U4762 ( .B1(n4162), .B2(n4285), .A(n4161), .ZN(U3266) );
  NAND2_X1 U4763 ( .A1(n4186), .A2(n4163), .ZN(n4164) );
  XOR2_X1 U4764 ( .A(n4172), .B(n4164), .Z(n4368) );
  INV_X1 U4765 ( .A(n4368), .ZN(n4184) );
  OR2_X1 U4766 ( .A1(n4165), .A2(n4166), .ZN(n4168) );
  NAND2_X1 U4767 ( .A1(n4168), .A2(n4167), .ZN(n4190) );
  INV_X1 U4768 ( .A(n4169), .ZN(n4170) );
  AOI21_X1 U4769 ( .B1(n4190), .B2(n4189), .A(n4170), .ZN(n4171) );
  XOR2_X1 U4770 ( .A(n4172), .B(n4171), .Z(n4176) );
  OAI22_X1 U4771 ( .A1(n4173), .A2(n4315), .B1(n4178), .B2(n4253), .ZN(n4174)
         );
  AOI21_X1 U4772 ( .B1(n4312), .B2(n4208), .A(n4174), .ZN(n4175) );
  OAI21_X1 U4773 ( .B1(n4176), .B2(n4210), .A(n4175), .ZN(n4367) );
  INV_X1 U4774 ( .A(n4371), .ZN(n4179) );
  OAI21_X1 U4775 ( .B1(n4179), .B2(n4178), .A(n4177), .ZN(n4442) );
  AOI22_X1 U4776 ( .A1(n4180), .A2(n4534), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4540), .ZN(n4181) );
  OAI21_X1 U4777 ( .B1(n4442), .B2(n4268), .A(n4181), .ZN(n4182) );
  AOI21_X1 U4778 ( .B1(n4367), .B2(n4538), .A(n4182), .ZN(n4183) );
  OAI21_X1 U4779 ( .B1(n4184), .B2(n4285), .A(n4183), .ZN(U3267) );
  INV_X1 U4780 ( .A(n4185), .ZN(n4188) );
  OAI21_X1 U4781 ( .B1(n4188), .B2(n4187), .A(n4186), .ZN(n4375) );
  XNOR2_X1 U4782 ( .A(n4190), .B(n4189), .ZN(n4197) );
  NAND2_X1 U4783 ( .A1(n4191), .A2(n4292), .ZN(n4195) );
  NOR2_X1 U4784 ( .A1(n4253), .A2(n4199), .ZN(n4192) );
  AOI21_X1 U4785 ( .B1(n4193), .B2(n4312), .A(n4192), .ZN(n4194) );
  NAND2_X1 U4786 ( .A1(n4195), .A2(n4194), .ZN(n4196) );
  AOI21_X1 U4787 ( .B1(n4197), .B2(n4318), .A(n4196), .ZN(n4374) );
  AOI22_X1 U4788 ( .A1(n4198), .A2(n4534), .B1(n4540), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4201) );
  OR2_X1 U4789 ( .A1(n4213), .A2(n4199), .ZN(n4372) );
  NAND3_X1 U4790 ( .A1(n4372), .A2(n4371), .A3(n4328), .ZN(n4200) );
  OAI211_X1 U4791 ( .C1(n4374), .C2(n4540), .A(n4201), .B(n4200), .ZN(n4202)
         );
  INV_X1 U4792 ( .A(n4202), .ZN(n4203) );
  OAI21_X1 U4793 ( .B1(n4375), .B2(n4285), .A(n4203), .ZN(U3268) );
  XNOR2_X1 U4794 ( .A(n4204), .B(n4205), .ZN(n4377) );
  INV_X1 U4795 ( .A(n4377), .ZN(n4221) );
  XOR2_X1 U4796 ( .A(n4205), .B(n4165), .Z(n4211) );
  OAI22_X1 U4797 ( .A1(n4206), .A2(n4275), .B1(n4215), .B2(n4253), .ZN(n4207)
         );
  AOI21_X1 U4798 ( .B1(n4292), .B2(n4208), .A(n4207), .ZN(n4209) );
  OAI21_X1 U4799 ( .B1(n4211), .B2(n4210), .A(n4209), .ZN(n4376) );
  INV_X1 U4800 ( .A(n4213), .ZN(n4214) );
  OAI21_X1 U4801 ( .B1(n4212), .B2(n4215), .A(n4214), .ZN(n4447) );
  NOR2_X1 U4802 ( .A1(n4447), .A2(n4268), .ZN(n4219) );
  INV_X1 U4803 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4216) );
  OAI22_X1 U4804 ( .A1(n4217), .A2(n4329), .B1(n4538), .B2(n4216), .ZN(n4218)
         );
  AOI211_X1 U4805 ( .C1(n4376), .C2(n4538), .A(n4219), .B(n4218), .ZN(n4220)
         );
  OAI21_X1 U4806 ( .B1(n4221), .B2(n4285), .A(n4220), .ZN(U3269) );
  XNOR2_X1 U4807 ( .A(n4222), .B(n4225), .ZN(n4379) );
  NAND2_X1 U4808 ( .A1(n4224), .A2(n4223), .ZN(n4226) );
  XNOR2_X1 U4809 ( .A(n4226), .B(n4225), .ZN(n4230) );
  AOI22_X1 U4810 ( .A1(n4273), .A2(n4312), .B1(n4234), .B2(n4311), .ZN(n4227)
         );
  OAI21_X1 U4811 ( .B1(n4228), .B2(n4315), .A(n4227), .ZN(n4229) );
  AOI21_X1 U4812 ( .B1(n4230), .B2(n4318), .A(n4229), .ZN(n4231) );
  OAI21_X1 U4813 ( .B1(n4379), .B2(n4232), .A(n4231), .ZN(n4380) );
  NAND2_X1 U4814 ( .A1(n4380), .A2(n4538), .ZN(n4242) );
  INV_X1 U4815 ( .A(n4212), .ZN(n4236) );
  INV_X1 U4816 ( .A(n4233), .ZN(n4265) );
  NAND2_X1 U4817 ( .A1(n4265), .A2(n4234), .ZN(n4235) );
  NAND2_X1 U4818 ( .A1(n4236), .A2(n4235), .ZN(n4451) );
  INV_X1 U4819 ( .A(n4451), .ZN(n4240) );
  OAI22_X1 U4820 ( .A1(n4538), .A2(n4238), .B1(n4237), .B2(n4329), .ZN(n4239)
         );
  AOI21_X1 U4821 ( .B1(n4240), .B2(n4328), .A(n4239), .ZN(n4241) );
  OAI211_X1 U4822 ( .C1(n4379), .C2(n4243), .A(n4242), .B(n4241), .ZN(U3270)
         );
  OR2_X1 U4823 ( .A1(n4244), .A2(n4245), .ZN(n4247) );
  NAND2_X1 U4824 ( .A1(n4247), .A2(n4246), .ZN(n4271) );
  INV_X1 U4825 ( .A(n4248), .ZN(n4250) );
  OAI21_X1 U4826 ( .B1(n4271), .B2(n4250), .A(n4249), .ZN(n4251) );
  XNOR2_X1 U4827 ( .A(n4251), .B(n4260), .ZN(n4259) );
  NAND2_X1 U4828 ( .A1(n4252), .A2(n4292), .ZN(n4257) );
  NOR2_X1 U4829 ( .A1(n4254), .A2(n4253), .ZN(n4255) );
  AOI21_X1 U4830 ( .B1(n4293), .B2(n4312), .A(n4255), .ZN(n4256) );
  NAND2_X1 U4831 ( .A1(n4257), .A2(n4256), .ZN(n4258) );
  AOI21_X1 U4832 ( .B1(n4259), .B2(n4318), .A(n4258), .ZN(n4386) );
  XNOR2_X1 U4833 ( .A(n4261), .B(n4260), .ZN(n4384) );
  NAND2_X1 U4834 ( .A1(n4262), .A2(n4263), .ZN(n4264) );
  NAND2_X1 U4835 ( .A1(n4265), .A2(n4264), .ZN(n4455) );
  AOI22_X1 U4836 ( .A1(n4540), .A2(REG2_REG_19__SCAN_IN), .B1(n4266), .B2(
        n4534), .ZN(n4267) );
  OAI21_X1 U4837 ( .B1(n4455), .B2(n4268), .A(n4267), .ZN(n4269) );
  AOI21_X1 U4838 ( .B1(n4384), .B2(n4333), .A(n4269), .ZN(n4270) );
  OAI21_X1 U4839 ( .B1(n4386), .B2(n4540), .A(n4270), .ZN(U3271) );
  XNOR2_X1 U4840 ( .A(n4271), .B(n4284), .ZN(n4277) );
  AOI22_X1 U4841 ( .A1(n4273), .A2(n4292), .B1(n4311), .B2(n4272), .ZN(n4274)
         );
  OAI21_X1 U4842 ( .B1(n4316), .B2(n4275), .A(n4274), .ZN(n4276) );
  AOI21_X1 U4843 ( .B1(n4277), .B2(n4318), .A(n4276), .ZN(n4390) );
  OAI211_X1 U4844 ( .C1(n4298), .C2(n4278), .A(n4262), .B(n4575), .ZN(n4389)
         );
  INV_X1 U4845 ( .A(n4389), .ZN(n4289) );
  INV_X1 U4846 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4280) );
  OAI22_X1 U4847 ( .A1(n4538), .A2(n4280), .B1(n4279), .B2(n4329), .ZN(n4287)
         );
  INV_X1 U4848 ( .A(n4281), .ZN(n4282) );
  AOI21_X1 U4849 ( .B1(n4284), .B2(n4283), .A(n4282), .ZN(n4391) );
  NOR2_X1 U4850 ( .A1(n4391), .A2(n4285), .ZN(n4286) );
  AOI211_X1 U4851 ( .C1(n4289), .C2(n4288), .A(n4287), .B(n4286), .ZN(n4290)
         );
  OAI21_X1 U4852 ( .B1(n4540), .B2(n4390), .A(n4290), .ZN(U3272) );
  XNOR2_X1 U4853 ( .A(n4244), .B(n4305), .ZN(n4297) );
  AOI22_X1 U4854 ( .A1(n4291), .A2(n4312), .B1(n4299), .B2(n4311), .ZN(n4295)
         );
  NAND2_X1 U4855 ( .A1(n4293), .A2(n4292), .ZN(n4294) );
  NAND2_X1 U4856 ( .A1(n4295), .A2(n4294), .ZN(n4296) );
  AOI21_X1 U4857 ( .B1(n4297), .B2(n4318), .A(n4296), .ZN(n4394) );
  OR2_X1 U4858 ( .A1(n3601), .A2(n4327), .ZN(n4399) );
  AOI21_X1 U4859 ( .B1(n4299), .B2(n4399), .A(n4298), .ZN(n4460) );
  INV_X1 U4860 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4302) );
  INV_X1 U4861 ( .A(n4300), .ZN(n4301) );
  OAI22_X1 U4862 ( .A1(n4538), .A2(n4302), .B1(n4301), .B2(n4329), .ZN(n4303)
         );
  AOI21_X1 U4863 ( .B1(n4460), .B2(n4328), .A(n4303), .ZN(n4308) );
  INV_X1 U4864 ( .A(n4305), .ZN(n4306) );
  XNOR2_X1 U4865 ( .A(n4304), .B(n4306), .ZN(n4392) );
  NAND2_X1 U4866 ( .A1(n4392), .A2(n4333), .ZN(n4307) );
  OAI211_X1 U4867 ( .C1(n4394), .C2(n4540), .A(n4308), .B(n4307), .ZN(U3273)
         );
  XOR2_X1 U4868 ( .A(n4309), .B(n4310), .Z(n4319) );
  AOI22_X1 U4869 ( .A1(n4313), .A2(n4312), .B1(n4327), .B2(n4311), .ZN(n4314)
         );
  OAI21_X1 U4870 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n4317) );
  AOI21_X1 U4871 ( .B1(n4319), .B2(n4318), .A(n4317), .ZN(n4401) );
  NAND2_X1 U4872 ( .A1(n3600), .A2(n4320), .ZN(n4323) );
  AND2_X1 U4873 ( .A1(n4323), .A2(n4321), .ZN(n4326) );
  NAND2_X1 U4874 ( .A1(n4323), .A2(n4322), .ZN(n4324) );
  OAI21_X1 U4875 ( .B1(n4326), .B2(n4325), .A(n4324), .ZN(n4402) );
  INV_X1 U4876 ( .A(n4402), .ZN(n4334) );
  NAND2_X1 U4877 ( .A1(n3601), .A2(n4327), .ZN(n4398) );
  AND3_X1 U4878 ( .A1(n4399), .A2(n4328), .A3(n4398), .ZN(n4332) );
  OAI22_X1 U4879 ( .A1(n4538), .A2(n2323), .B1(n4330), .B2(n4329), .ZN(n4331)
         );
  AOI211_X1 U4880 ( .C1(n4334), .C2(n4333), .A(n4332), .B(n4331), .ZN(n4335)
         );
  OAI21_X1 U4881 ( .B1(n4540), .B2(n4401), .A(n4335), .ZN(U3274) );
  NAND2_X1 U4882 ( .A1(n4592), .A2(n4419), .ZN(n4337) );
  NAND2_X1 U4883 ( .A1(n4590), .A2(REG1_REG_31__SCAN_IN), .ZN(n4336) );
  OAI211_X1 U4884 ( .C1(n4422), .C2(n4418), .A(n4337), .B(n4336), .ZN(U3549)
         );
  NAND2_X1 U4885 ( .A1(n4592), .A2(n4423), .ZN(n4339) );
  NAND2_X1 U4886 ( .A1(n4590), .A2(REG1_REG_30__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U4887 ( .C1(n4426), .C2(n4418), .A(n4339), .B(n4338), .ZN(U3548)
         );
  NAND3_X1 U4888 ( .A1(n4340), .A2(n4578), .A3(n4341), .ZN(n4350) );
  NOR2_X1 U4889 ( .A1(n4341), .A2(n4569), .ZN(n4343) );
  NAND2_X1 U4890 ( .A1(n4342), .A2(n4343), .ZN(n4347) );
  AOI22_X1 U4891 ( .A1(n4345), .A2(n4575), .B1(n4344), .B2(n4343), .ZN(n4346)
         );
  AND2_X1 U4892 ( .A1(n4347), .A2(n4346), .ZN(n4349) );
  NAND3_X1 U4893 ( .A1(n4350), .A2(n4349), .A3(n4348), .ZN(n4427) );
  MUX2_X1 U4894 ( .A(REG1_REG_29__SCAN_IN), .B(n4427), .S(n4592), .Z(U3547) );
  NAND2_X1 U4895 ( .A1(n4351), .A2(n4575), .ZN(n4352) );
  OAI211_X1 U4896 ( .C1(n4354), .C2(n4569), .A(n4353), .B(n4352), .ZN(n4428)
         );
  MUX2_X1 U4897 ( .A(REG1_REG_27__SCAN_IN), .B(n4428), .S(n4592), .Z(U3545) );
  INV_X1 U4898 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4357) );
  MUX2_X1 U4899 ( .A(n4357), .B(n4429), .S(n4592), .Z(n4358) );
  OAI21_X1 U4900 ( .B1(n4418), .B2(n4432), .A(n4358), .ZN(U3544) );
  AOI21_X1 U4901 ( .B1(n4360), .B2(n4578), .A(n4359), .ZN(n4433) );
  INV_X1 U4902 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4361) );
  MUX2_X1 U4903 ( .A(n4433), .B(n4361), .S(n4590), .Z(n4362) );
  OAI21_X1 U4904 ( .B1(n4418), .B2(n4435), .A(n4362), .ZN(U3543) );
  INV_X1 U4905 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4365) );
  AOI21_X1 U4906 ( .B1(n4364), .B2(n4578), .A(n4363), .ZN(n4436) );
  MUX2_X1 U4907 ( .A(n4365), .B(n4436), .S(n4592), .Z(n4366) );
  OAI21_X1 U4908 ( .B1(n4418), .B2(n4438), .A(n4366), .ZN(U3542) );
  AOI21_X1 U4909 ( .B1(n4368), .B2(n4578), .A(n4367), .ZN(n4440) );
  INV_X1 U4910 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4369) );
  MUX2_X1 U4911 ( .A(n4440), .B(n4369), .S(n4590), .Z(n4370) );
  OAI21_X1 U4912 ( .B1(n4418), .B2(n4442), .A(n4370), .ZN(U3541) );
  NAND3_X1 U4913 ( .A1(n4372), .A2(n4575), .A3(n4371), .ZN(n4373) );
  OAI211_X1 U4914 ( .C1(n4375), .C2(n4569), .A(n4374), .B(n4373), .ZN(n4443)
         );
  MUX2_X1 U4915 ( .A(REG1_REG_22__SCAN_IN), .B(n4443), .S(n4592), .Z(U3540) );
  AOI21_X1 U4916 ( .B1(n4377), .B2(n4578), .A(n4376), .ZN(n4444) );
  MUX2_X1 U4917 ( .A(n4696), .B(n4444), .S(n4592), .Z(n4378) );
  OAI21_X1 U4918 ( .B1(n4418), .B2(n4447), .A(n4378), .ZN(U3539) );
  INV_X1 U4919 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4382) );
  INV_X1 U4920 ( .A(n4379), .ZN(n4381) );
  AOI21_X1 U4921 ( .B1(n4566), .B2(n4381), .A(n4380), .ZN(n4448) );
  MUX2_X1 U4922 ( .A(n4382), .B(n4448), .S(n4592), .Z(n4383) );
  OAI21_X1 U4923 ( .B1(n4418), .B2(n4451), .A(n4383), .ZN(U3538) );
  NAND2_X1 U4924 ( .A1(n4384), .A2(n4578), .ZN(n4385) );
  NAND2_X1 U4925 ( .A1(n4386), .A2(n4385), .ZN(n4452) );
  MUX2_X1 U4926 ( .A(n4452), .B(REG1_REG_19__SCAN_IN), .S(n4590), .Z(n4387) );
  INV_X1 U4927 ( .A(n4387), .ZN(n4388) );
  OAI21_X1 U4928 ( .B1(n4418), .B2(n4455), .A(n4388), .ZN(U3537) );
  OAI211_X1 U4929 ( .C1(n4391), .C2(n4569), .A(n4390), .B(n4389), .ZN(n4456)
         );
  MUX2_X1 U4930 ( .A(REG1_REG_18__SCAN_IN), .B(n4456), .S(n4592), .Z(U3536) );
  NAND2_X1 U4931 ( .A1(n4392), .A2(n4578), .ZN(n4393) );
  NAND2_X1 U4932 ( .A1(n4394), .A2(n4393), .ZN(n4457) );
  MUX2_X1 U4933 ( .A(REG1_REG_17__SCAN_IN), .B(n4457), .S(n4592), .Z(n4395) );
  AOI21_X1 U4934 ( .B1(n4396), .B2(n4460), .A(n4395), .ZN(n4397) );
  INV_X1 U4935 ( .A(n4397), .ZN(U3535) );
  NAND3_X1 U4936 ( .A1(n4399), .A2(n4575), .A3(n4398), .ZN(n4400) );
  OAI211_X1 U4937 ( .C1(n4569), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4462)
         );
  MUX2_X1 U4938 ( .A(REG1_REG_16__SCAN_IN), .B(n4462), .S(n4592), .Z(U3534) );
  AOI21_X1 U4939 ( .B1(n4578), .B2(n4404), .A(n4403), .ZN(n4463) );
  MUX2_X1 U4940 ( .A(n4405), .B(n4463), .S(n4592), .Z(n4406) );
  OAI21_X1 U4941 ( .B1(n4418), .B2(n4466), .A(n4406), .ZN(U3533) );
  INV_X1 U4942 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4409) );
  AOI21_X1 U4943 ( .B1(n4566), .B2(n4408), .A(n4407), .ZN(n4467) );
  MUX2_X1 U4944 ( .A(n4409), .B(n4467), .S(n4592), .Z(n4410) );
  OAI21_X1 U4945 ( .B1(n4418), .B2(n4470), .A(n4410), .ZN(U3532) );
  AOI21_X1 U4946 ( .B1(n4566), .B2(n4412), .A(n4411), .ZN(n4471) );
  MUX2_X1 U4947 ( .A(n4413), .B(n4471), .S(n4592), .Z(n4414) );
  OAI21_X1 U4948 ( .B1(n4418), .B2(n4474), .A(n4414), .ZN(U3531) );
  INV_X1 U4949 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4680) );
  AOI21_X1 U4950 ( .B1(n4578), .B2(n4416), .A(n4415), .ZN(n4475) );
  MUX2_X1 U4951 ( .A(n4680), .B(n4475), .S(n4592), .Z(n4417) );
  OAI21_X1 U4952 ( .B1(n4418), .B2(n4479), .A(n4417), .ZN(U3530) );
  NAND2_X1 U4953 ( .A1(n4586), .A2(n4419), .ZN(n4421) );
  NAND2_X1 U4954 ( .A1(n4584), .A2(REG0_REG_31__SCAN_IN), .ZN(n4420) );
  OAI211_X1 U4955 ( .C1(n4422), .C2(n4478), .A(n4421), .B(n4420), .ZN(U3517)
         );
  NAND2_X1 U4956 ( .A1(n4586), .A2(n4423), .ZN(n4425) );
  NAND2_X1 U4957 ( .A1(n4584), .A2(REG0_REG_30__SCAN_IN), .ZN(n4424) );
  OAI211_X1 U4958 ( .C1(n4426), .C2(n4478), .A(n4425), .B(n4424), .ZN(U3516)
         );
  MUX2_X1 U4959 ( .A(REG0_REG_29__SCAN_IN), .B(n4427), .S(n4586), .Z(U3515) );
  MUX2_X1 U4960 ( .A(REG0_REG_27__SCAN_IN), .B(n4428), .S(n4586), .Z(U3513) );
  INV_X1 U4961 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4430) );
  MUX2_X1 U4962 ( .A(n4430), .B(n4429), .S(n4586), .Z(n4431) );
  OAI21_X1 U4963 ( .B1(n4432), .B2(n4478), .A(n4431), .ZN(U3512) );
  MUX2_X1 U4964 ( .A(n4433), .B(n4667), .S(n4584), .Z(n4434) );
  OAI21_X1 U4965 ( .B1(n4435), .B2(n4478), .A(n4434), .ZN(U3511) );
  MUX2_X1 U4966 ( .A(n4721), .B(n4436), .S(n4586), .Z(n4437) );
  OAI21_X1 U4967 ( .B1(n4438), .B2(n4478), .A(n4437), .ZN(U3510) );
  INV_X1 U4968 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4439) );
  MUX2_X1 U4969 ( .A(n4440), .B(n4439), .S(n4584), .Z(n4441) );
  OAI21_X1 U4970 ( .B1(n4442), .B2(n4478), .A(n4441), .ZN(U3509) );
  MUX2_X1 U4971 ( .A(REG0_REG_22__SCAN_IN), .B(n4443), .S(n4586), .Z(U3508) );
  INV_X1 U4972 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4445) );
  MUX2_X1 U4973 ( .A(n4445), .B(n4444), .S(n4586), .Z(n4446) );
  OAI21_X1 U4974 ( .B1(n4447), .B2(n4478), .A(n4446), .ZN(U3507) );
  INV_X1 U4975 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4449) );
  MUX2_X1 U4976 ( .A(n4449), .B(n4448), .S(n4586), .Z(n4450) );
  OAI21_X1 U4977 ( .B1(n4451), .B2(n4478), .A(n4450), .ZN(U3506) );
  MUX2_X1 U4978 ( .A(REG0_REG_19__SCAN_IN), .B(n4452), .S(n4586), .Z(n4453) );
  INV_X1 U4979 ( .A(n4453), .ZN(n4454) );
  OAI21_X1 U4980 ( .B1(n4455), .B2(n4478), .A(n4454), .ZN(U3505) );
  MUX2_X1 U4981 ( .A(REG0_REG_18__SCAN_IN), .B(n4456), .S(n4586), .Z(U3503) );
  MUX2_X1 U4982 ( .A(REG0_REG_17__SCAN_IN), .B(n4457), .S(n4586), .Z(n4458) );
  AOI21_X1 U4983 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n4461) );
  INV_X1 U4984 ( .A(n4461), .ZN(U3501) );
  MUX2_X1 U4985 ( .A(REG0_REG_16__SCAN_IN), .B(n4462), .S(n4586), .Z(U3499) );
  INV_X1 U4986 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4464) );
  MUX2_X1 U4987 ( .A(n4464), .B(n4463), .S(n4586), .Z(n4465) );
  OAI21_X1 U4988 ( .B1(n4466), .B2(n4478), .A(n4465), .ZN(U3497) );
  INV_X1 U4989 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4468) );
  MUX2_X1 U4990 ( .A(n4468), .B(n4467), .S(n4586), .Z(n4469) );
  OAI21_X1 U4991 ( .B1(n4470), .B2(n4478), .A(n4469), .ZN(U3495) );
  INV_X1 U4992 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4472) );
  MUX2_X1 U4993 ( .A(n4472), .B(n4471), .S(n4586), .Z(n4473) );
  OAI21_X1 U4994 ( .B1(n4474), .B2(n4478), .A(n4473), .ZN(U3493) );
  INV_X1 U4995 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4476) );
  MUX2_X1 U4996 ( .A(n4476), .B(n4475), .S(n4586), .Z(n4477) );
  OAI21_X1 U4997 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(U3491) );
  MUX2_X1 U4998 ( .A(DATAI_30_), .B(n4480), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4999 ( .A(DATAI_28_), .B(n4481), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5000 ( .A(n4495), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5001 ( .A(n4482), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5002 ( .A(n4483), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5003 ( .A(DATAI_24_), .B(n2889), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5004 ( .A(n4484), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5005 ( .A(n2454), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5006 ( .A(DATAI_20_), .B(n4485), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5007 ( .A(n4486), .B(DATAI_16_), .S(U3149), .Z(U3336) );
  MUX2_X1 U5008 ( .A(n4487), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5009 ( .A(n4488), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5010 ( .A(DATAI_11_), .B(n2300), .S(STATE_REG_SCAN_IN), .Z(U3341)
         );
  MUX2_X1 U5011 ( .A(n4490), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5012 ( .A(n4491), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U5013 ( .A(n4492), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5014 ( .A(DATAI_3_), .B(n4493), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5015 ( .A(n2379), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U5016 ( .A(n4497), .ZN(n4494) );
  OAI211_X1 U5017 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4495), .A(n4494), .B(n4496), 
        .ZN(n4501) );
  OAI22_X1 U5018 ( .A1(n4497), .A2(n4496), .B1(n4514), .B2(REG1_REG_0__SCAN_IN), .ZN(n4498) );
  INV_X1 U5019 ( .A(n4498), .ZN(n4500) );
  AOI22_X1 U5020 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4517), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4499) );
  OAI221_X1 U5021 ( .B1(IR_REG_0__SCAN_IN), .B2(n4501), .C1(n2447), .C2(n4500), 
        .A(n4499), .ZN(U3240) );
  AOI21_X1 U5022 ( .B1(n4517), .B2(ADDR_REG_17__SCAN_IN), .A(n4502), .ZN(n4513) );
  OAI21_X1 U5023 ( .B1(n4505), .B2(n4504), .A(n4503), .ZN(n4511) );
  OAI21_X1 U5024 ( .B1(n4508), .B2(n4507), .A(n4506), .ZN(n4509) );
  AOI22_X1 U5025 ( .A1(n2375), .A2(n4511), .B1(n4510), .B2(n4509), .ZN(n4512)
         );
  OAI211_X1 U5026 ( .C1(n4548), .C2(n4529), .A(n4513), .B(n4512), .ZN(U3257)
         );
  NAND2_X1 U5027 ( .A1(n4517), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4520) );
  INV_X1 U5028 ( .A(n4518), .ZN(n4519) );
  NAND2_X1 U5029 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  AOI21_X1 U5030 ( .B1(n4525), .B2(n4524), .A(n4523), .ZN(n4526) );
  NAND2_X1 U5031 ( .A1(n2375), .A2(n4526), .ZN(n4527) );
  OAI211_X1 U5032 ( .C1(n4529), .C2(n4546), .A(n4528), .B(n4527), .ZN(U3258)
         );
  INV_X1 U5033 ( .A(n4530), .ZN(n4532) );
  AOI21_X1 U5034 ( .B1(n4533), .B2(n4532), .A(n4531), .ZN(n4539) );
  AOI22_X1 U5035 ( .A1(n4536), .A2(n4535), .B1(REG3_REG_0__SCAN_IN), .B2(n4534), .ZN(n4537) );
  OAI221_X1 U5036 ( .B1(n4540), .B2(n4539), .C1(n4538), .C2(n2254), .A(n4537), 
        .ZN(U3290) );
  AND2_X1 U5037 ( .A1(D_REG_31__SCAN_IN), .A2(n4593), .ZN(U3291) );
  AND2_X1 U5038 ( .A1(D_REG_30__SCAN_IN), .A2(n4593), .ZN(U3292) );
  AND2_X1 U5039 ( .A1(D_REG_29__SCAN_IN), .A2(n4593), .ZN(U3293) );
  AND2_X1 U5040 ( .A1(D_REG_27__SCAN_IN), .A2(n4593), .ZN(U3295) );
  AND2_X1 U5041 ( .A1(D_REG_26__SCAN_IN), .A2(n4593), .ZN(U3296) );
  AND2_X1 U5042 ( .A1(D_REG_25__SCAN_IN), .A2(n4593), .ZN(U3297) );
  INV_X1 U5043 ( .A(n4593), .ZN(n4542) );
  INV_X1 U5044 ( .A(D_REG_24__SCAN_IN), .ZN(n4687) );
  NOR2_X1 U5045 ( .A1(n4542), .A2(n4687), .ZN(U3298) );
  INV_X1 U5046 ( .A(D_REG_23__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U5047 ( .A1(n4542), .A2(n4720), .ZN(U3299) );
  INV_X1 U5048 ( .A(D_REG_22__SCAN_IN), .ZN(n4686) );
  NOR2_X1 U5049 ( .A1(n4542), .A2(n4686), .ZN(U3300) );
  INV_X1 U5050 ( .A(D_REG_21__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5051 ( .A1(n4542), .A2(n4689), .ZN(U3301) );
  AND2_X1 U5052 ( .A1(D_REG_20__SCAN_IN), .A2(n4593), .ZN(U3302) );
  AND2_X1 U5053 ( .A1(D_REG_19__SCAN_IN), .A2(n4593), .ZN(U3303) );
  AND2_X1 U5054 ( .A1(D_REG_18__SCAN_IN), .A2(n4593), .ZN(U3304) );
  INV_X1 U5055 ( .A(D_REG_17__SCAN_IN), .ZN(n4708) );
  NOR2_X1 U5056 ( .A1(n4542), .A2(n4708), .ZN(U3305) );
  AND2_X1 U5057 ( .A1(D_REG_16__SCAN_IN), .A2(n4593), .ZN(U3306) );
  INV_X1 U5058 ( .A(D_REG_15__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U5059 ( .A1(n4542), .A2(n4663), .ZN(U3307) );
  AND2_X1 U5060 ( .A1(D_REG_14__SCAN_IN), .A2(n4593), .ZN(U3308) );
  AND2_X1 U5061 ( .A1(D_REG_13__SCAN_IN), .A2(n4593), .ZN(U3309) );
  AND2_X1 U5062 ( .A1(D_REG_12__SCAN_IN), .A2(n4593), .ZN(U3310) );
  AND2_X1 U5063 ( .A1(D_REG_11__SCAN_IN), .A2(n4593), .ZN(U3311) );
  AND2_X1 U5064 ( .A1(D_REG_10__SCAN_IN), .A2(n4593), .ZN(U3312) );
  AND2_X1 U5065 ( .A1(D_REG_9__SCAN_IN), .A2(n4593), .ZN(U3313) );
  AND2_X1 U5066 ( .A1(D_REG_8__SCAN_IN), .A2(n4593), .ZN(U3314) );
  AND2_X1 U5067 ( .A1(D_REG_7__SCAN_IN), .A2(n4593), .ZN(U3315) );
  INV_X1 U5068 ( .A(D_REG_6__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U5069 ( .A1(n4542), .A2(n4541), .ZN(U3316) );
  AND2_X1 U5070 ( .A1(D_REG_5__SCAN_IN), .A2(n4593), .ZN(U3317) );
  AND2_X1 U5071 ( .A1(D_REG_4__SCAN_IN), .A2(n4593), .ZN(U3318) );
  AND2_X1 U5072 ( .A1(D_REG_3__SCAN_IN), .A2(n4593), .ZN(U3319) );
  AND2_X1 U5073 ( .A1(D_REG_2__SCAN_IN), .A2(n4593), .ZN(U3320) );
  OAI21_X1 U5074 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4543), .ZN(
        n4544) );
  INV_X1 U5075 ( .A(n4544), .ZN(U3329) );
  INV_X1 U5076 ( .A(DATAI_18_), .ZN(n4545) );
  AOI22_X1 U5077 ( .A1(STATE_REG_SCAN_IN), .A2(n4546), .B1(n4545), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5078 ( .A(DATAI_17_), .ZN(n4547) );
  AOI22_X1 U5079 ( .A1(STATE_REG_SCAN_IN), .A2(n4548), .B1(n4547), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5080 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4551) );
  INV_X1 U5081 ( .A(n4551), .ZN(U3352) );
  INV_X1 U5082 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4552) );
  AOI22_X1 U5083 ( .A1(n4586), .A2(n4553), .B1(n4552), .B2(n4584), .ZN(U3467)
         );
  INV_X1 U5084 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5085 ( .A1(n4586), .A2(n4555), .B1(n4554), .B2(n4584), .ZN(U3469)
         );
  OAI22_X1 U5086 ( .A1(n4559), .A2(n4558), .B1(n4557), .B2(n4556), .ZN(n4560)
         );
  NOR2_X1 U5087 ( .A1(n4561), .A2(n4560), .ZN(n4587) );
  INV_X1 U5088 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5089 ( .A1(n4586), .A2(n4587), .B1(n4562), .B2(n4584), .ZN(U3473)
         );
  INV_X1 U5090 ( .A(n4563), .ZN(n4565) );
  AOI211_X1 U5091 ( .C1(n4567), .C2(n4566), .A(n4565), .B(n4564), .ZN(n4588)
         );
  INV_X1 U5092 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5093 ( .A1(n4586), .A2(n4588), .B1(n4568), .B2(n4584), .ZN(U3475)
         );
  NOR2_X1 U5094 ( .A1(n4570), .A2(n4569), .ZN(n4573) );
  INV_X1 U5095 ( .A(n4571), .ZN(n4572) );
  AOI211_X1 U5096 ( .C1(n4575), .C2(n4574), .A(n4573), .B(n4572), .ZN(n4589)
         );
  INV_X1 U5097 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5098 ( .A1(n4586), .A2(n4589), .B1(n4576), .B2(n4584), .ZN(U3477)
         );
  NAND3_X1 U5099 ( .A1(n4579), .A2(n4578), .A3(n4577), .ZN(n4581) );
  AND2_X1 U5100 ( .A1(n4581), .A2(n4580), .ZN(n4582) );
  AND2_X1 U5101 ( .A1(n4583), .A2(n4582), .ZN(n4591) );
  INV_X1 U5102 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5103 ( .A1(n4586), .A2(n4591), .B1(n4585), .B2(n4584), .ZN(U3481)
         );
  INV_X1 U5104 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5105 ( .A1(n4592), .A2(n4587), .B1(n4681), .B2(n4590), .ZN(U3521)
         );
  AOI22_X1 U5106 ( .A1(n4592), .A2(n4588), .B1(n2159), .B2(n4590), .ZN(U3522)
         );
  AOI22_X1 U5107 ( .A1(n4592), .A2(n4589), .B1(n4722), .B2(n4590), .ZN(U3523)
         );
  AOI22_X1 U5108 ( .A1(n4592), .A2(n4591), .B1(n2384), .B2(n4590), .ZN(U3525)
         );
  NAND2_X1 U5109 ( .A1(n4593), .A2(D_REG_28__SCAN_IN), .ZN(n4741) );
  INV_X1 U5110 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4711) );
  NAND4_X1 U5111 ( .A1(D_REG_17__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), .A3(
        n4711), .A4(n2539), .ZN(n4600) );
  INV_X1 U5112 ( .A(IR_REG_1__SCAN_IN), .ZN(n4595) );
  NAND4_X1 U5113 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(IR_REG_20__SCAN_IN), 
        .ZN(n4599) );
  NAND4_X1 U5114 ( .A1(D_REG_0__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(DATAO_REG_30__SCAN_IN), .ZN(n4598) );
  NAND4_X1 U5115 ( .A1(REG3_REG_9__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .A3(
        REG1_REG_5__SCAN_IN), .A4(REG0_REG_24__SCAN_IN), .ZN(n4597) );
  NOR4_X1 U5116 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4739)
         );
  NOR3_X1 U5117 ( .A1(DATAI_15_), .A2(REG2_REG_31__SCAN_IN), .A3(n4624), .ZN(
        n4602) );
  NOR4_X1 U5118 ( .A1(IR_REG_16__SCAN_IN), .A2(REG2_REG_19__SCAN_IN), .A3(
        DATAI_14_), .A4(DATAO_REG_14__SCAN_IN), .ZN(n4601) );
  NAND4_X1 U5119 ( .A1(n4603), .A2(REG3_REG_4__SCAN_IN), .A3(n4602), .A4(n4601), .ZN(n4618) );
  NOR4_X1 U5120 ( .A1(n4604), .A2(DATAI_25_), .A3(REG0_REG_9__SCAN_IN), .A4(
        DATAI_28_), .ZN(n4612) );
  NOR4_X1 U5121 ( .A1(REG0_REG_27__SCAN_IN), .A2(DATAI_16_), .A3(
        REG2_REG_10__SCAN_IN), .A4(REG1_REG_4__SCAN_IN), .ZN(n4606) );
  NOR4_X1 U5122 ( .A1(REG3_REG_26__SCAN_IN), .A2(REG3_REG_14__SCAN_IN), .A3(
        REG0_REG_25__SCAN_IN), .A4(n4662), .ZN(n4605) );
  NAND2_X1 U5123 ( .A1(n4606), .A2(n4605), .ZN(n4610) );
  NOR4_X1 U5124 ( .A1(REG1_REG_12__SCAN_IN), .A2(DATAI_3_), .A3(
        REG1_REG_3__SCAN_IN), .A4(n4683), .ZN(n4608) );
  INV_X1 U5125 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4649) );
  INV_X1 U5126 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4654) );
  NOR4_X1 U5127 ( .A1(REG3_REG_21__SCAN_IN), .A2(DATAI_11_), .A3(n4649), .A4(
        n4654), .ZN(n4607) );
  NAND3_X1 U5128 ( .A1(REG0_REG_6__SCAN_IN), .A2(n4608), .A3(n4607), .ZN(n4609) );
  NOR3_X1 U5129 ( .A1(IR_REG_6__SCAN_IN), .A2(n4610), .A3(n4609), .ZN(n4611)
         );
  NAND4_X1 U5130 ( .A1(n4612), .A2(IR_REG_24__SCAN_IN), .A3(IR_REG_28__SCAN_IN), .A4(n4611), .ZN(n4617) );
  NAND4_X1 U5131 ( .A1(n4613), .A2(n4696), .A3(REG2_REG_3__SCAN_IN), .A4(
        REG1_REG_25__SCAN_IN), .ZN(n4616) );
  INV_X1 U5132 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4614) );
  NAND4_X1 U5133 ( .A1(n4614), .A2(ADDR_REG_13__SCAN_IN), .A3(
        REG1_REG_30__SCAN_IN), .A4(DATAO_REG_22__SCAN_IN), .ZN(n4615) );
  NOR4_X1 U5134 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4621)
         );
  NOR4_X1 U5135 ( .A1(IR_REG_9__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .A3(n4619), .A4(n2794), .ZN(n4620) );
  AND2_X1 U5136 ( .A1(n4621), .A2(n4620), .ZN(n4738) );
  AOI22_X1 U5137 ( .A1(n4624), .A2(keyinput32), .B1(n4623), .B2(keyinput33), 
        .ZN(n4622) );
  OAI221_X1 U5138 ( .B1(n4624), .B2(keyinput32), .C1(n4623), .C2(keyinput33), 
        .A(n4622), .ZN(n4635) );
  INV_X1 U5139 ( .A(DATAI_14_), .ZN(n4626) );
  AOI22_X1 U5140 ( .A1(n4627), .A2(keyinput41), .B1(keyinput40), .B2(n4626), 
        .ZN(n4625) );
  OAI221_X1 U5141 ( .B1(n4627), .B2(keyinput41), .C1(n4626), .C2(keyinput40), 
        .A(n4625), .ZN(n4634) );
  XNOR2_X1 U5142 ( .A(IR_REG_16__SCAN_IN), .B(keyinput38), .ZN(n4630) );
  XNOR2_X1 U5143 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput37), .ZN(n4629) );
  XNOR2_X1 U5144 ( .A(REG2_REG_31__SCAN_IN), .B(keyinput34), .ZN(n4628) );
  NAND3_X1 U5145 ( .A1(n4630), .A2(n4629), .A3(n4628), .ZN(n4633) );
  XNOR2_X1 U5146 ( .A(n4631), .B(keyinput36), .ZN(n4632) );
  NOR4_X1 U5147 ( .A1(n4635), .A2(n4634), .A3(n4633), .A4(n4632), .ZN(n4678)
         );
  INV_X1 U5148 ( .A(DATAI_16_), .ZN(n4637) );
  AOI22_X1 U5149 ( .A1(n2159), .A2(keyinput26), .B1(n4637), .B2(keyinput29), 
        .ZN(n4636) );
  OAI221_X1 U5150 ( .B1(n2159), .B2(keyinput26), .C1(n4637), .C2(keyinput29), 
        .A(n4636), .ZN(n4647) );
  AOI22_X1 U5151 ( .A1(n3260), .A2(keyinput22), .B1(keyinput20), .B2(n4639), 
        .ZN(n4638) );
  OAI221_X1 U5152 ( .B1(n3260), .B2(keyinput22), .C1(n4639), .C2(keyinput20), 
        .A(n4638), .ZN(n4646) );
  AOI22_X1 U5153 ( .A1(n2110), .A2(keyinput30), .B1(n4641), .B2(keyinput28), 
        .ZN(n4640) );
  OAI221_X1 U5154 ( .B1(n2110), .B2(keyinput30), .C1(n4641), .C2(keyinput28), 
        .A(n4640), .ZN(n4645) );
  XOR2_X1 U5155 ( .A(n4007), .B(keyinput25), .Z(n4643) );
  XNOR2_X1 U5156 ( .A(IR_REG_6__SCAN_IN), .B(keyinput24), .ZN(n4642) );
  NAND2_X1 U5157 ( .A1(n4643), .A2(n4642), .ZN(n4644) );
  NOR4_X1 U5158 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4677)
         );
  AOI22_X1 U5159 ( .A1(n4649), .A2(keyinput57), .B1(keyinput56), .B2(n2620), 
        .ZN(n4648) );
  OAI221_X1 U5160 ( .B1(n4649), .B2(keyinput57), .C1(n2620), .C2(keyinput56), 
        .A(n4648), .ZN(n4660) );
  AOI22_X1 U5161 ( .A1(n4651), .A2(keyinput58), .B1(keyinput61), .B2(n2794), 
        .ZN(n4650) );
  OAI221_X1 U5162 ( .B1(n4651), .B2(keyinput58), .C1(n2794), .C2(keyinput61), 
        .A(n4650), .ZN(n4659) );
  AOI22_X1 U5163 ( .A1(n4654), .A2(keyinput52), .B1(n4653), .B2(keyinput54), 
        .ZN(n4652) );
  OAI221_X1 U5164 ( .B1(n4654), .B2(keyinput52), .C1(n4653), .C2(keyinput54), 
        .A(n4652), .ZN(n4658) );
  XNOR2_X1 U5165 ( .A(IR_REG_9__SCAN_IN), .B(keyinput62), .ZN(n4656) );
  XNOR2_X1 U5166 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput60), .ZN(n4655) );
  NAND2_X1 U5167 ( .A1(n4656), .A2(n4655), .ZN(n4657) );
  NOR4_X1 U5168 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4676)
         );
  AOI22_X1 U5169 ( .A1(n4663), .A2(keyinput49), .B1(keyinput48), .B2(n4662), 
        .ZN(n4661) );
  OAI221_X1 U5170 ( .B1(n4663), .B2(keyinput49), .C1(n4662), .C2(keyinput48), 
        .A(n4661), .ZN(n4674) );
  INV_X1 U5171 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4665) );
  AOI22_X1 U5172 ( .A1(n4665), .A2(keyinput45), .B1(keyinput42), .B2(n4614), 
        .ZN(n4664) );
  OAI221_X1 U5173 ( .B1(n4665), .B2(keyinput45), .C1(n4614), .C2(keyinput42), 
        .A(n4664), .ZN(n4673) );
  AOI22_X1 U5174 ( .A1(n4668), .A2(keyinput50), .B1(keyinput53), .B2(n4667), 
        .ZN(n4666) );
  OAI221_X1 U5175 ( .B1(n4668), .B2(keyinput50), .C1(n4667), .C2(keyinput53), 
        .A(n4666), .ZN(n4672) );
  XNOR2_X1 U5176 ( .A(REG1_REG_30__SCAN_IN), .B(keyinput44), .ZN(n4670) );
  XNOR2_X1 U5177 ( .A(IR_REG_28__SCAN_IN), .B(keyinput46), .ZN(n4669) );
  NAND2_X1 U5178 ( .A1(n4670), .A2(n4669), .ZN(n4671) );
  NOR4_X1 U5179 ( .A1(n4674), .A2(n4673), .A3(n4672), .A4(n4671), .ZN(n4675)
         );
  NAND4_X1 U5180 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4737)
         );
  AOI22_X1 U5181 ( .A1(n4681), .A2(keyinput15), .B1(n4680), .B2(keyinput31), 
        .ZN(n4679) );
  OAI221_X1 U5182 ( .B1(n4681), .B2(keyinput15), .C1(n4680), .C2(keyinput31), 
        .A(n4679), .ZN(n4694) );
  INV_X1 U5183 ( .A(DATAI_25_), .ZN(n4684) );
  AOI22_X1 U5184 ( .A1(n4684), .A2(keyinput3), .B1(keyinput7), .B2(n4683), 
        .ZN(n4682) );
  OAI221_X1 U5185 ( .B1(n4684), .B2(keyinput3), .C1(n4683), .C2(keyinput7), 
        .A(n4682), .ZN(n4693) );
  AOI22_X1 U5186 ( .A1(n4687), .A2(keyinput23), .B1(n4686), .B2(keyinput11), 
        .ZN(n4685) );
  OAI221_X1 U5187 ( .B1(n4687), .B2(keyinput23), .C1(n4686), .C2(keyinput11), 
        .A(n4685), .ZN(n4692) );
  INV_X1 U5188 ( .A(DATAI_3_), .ZN(n4690) );
  AOI22_X1 U5189 ( .A1(n4690), .A2(keyinput63), .B1(n4689), .B2(keyinput39), 
        .ZN(n4688) );
  OAI221_X1 U5190 ( .B1(n4690), .B2(keyinput63), .C1(n4689), .C2(keyinput39), 
        .A(n4688), .ZN(n4691) );
  NOR4_X1 U5191 ( .A1(n4694), .A2(n4693), .A3(n4692), .A4(n4691), .ZN(n4735)
         );
  AOI22_X1 U5192 ( .A1(n4613), .A2(keyinput35), .B1(keyinput47), .B2(n4696), 
        .ZN(n4695) );
  OAI221_X1 U5193 ( .B1(n4613), .B2(keyinput35), .C1(n4696), .C2(keyinput47), 
        .A(n4695), .ZN(n4706) );
  INV_X1 U5194 ( .A(DATAI_28_), .ZN(n4699) );
  INV_X1 U5195 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5196 ( .A1(n4699), .A2(keyinput59), .B1(keyinput51), .B2(n4698), 
        .ZN(n4697) );
  OAI221_X1 U5197 ( .B1(n4699), .B2(keyinput59), .C1(n4698), .C2(keyinput51), 
        .A(n4697), .ZN(n4705) );
  XNOR2_X1 U5198 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput55), .ZN(n4703) );
  XNOR2_X1 U5199 ( .A(IR_REG_24__SCAN_IN), .B(keyinput43), .ZN(n4702) );
  XNOR2_X1 U5200 ( .A(REG1_REG_25__SCAN_IN), .B(keyinput19), .ZN(n4701) );
  XNOR2_X1 U5201 ( .A(IR_REG_15__SCAN_IN), .B(keyinput27), .ZN(n4700) );
  NAND4_X1 U5202 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(n4704)
         );
  NOR3_X1 U5203 ( .A1(n4706), .A2(n4705), .A3(n4704), .ZN(n4734) );
  AOI22_X1 U5204 ( .A1(n4708), .A2(keyinput16), .B1(keyinput17), .B2(n2539), 
        .ZN(n4707) );
  OAI221_X1 U5205 ( .B1(n4708), .B2(keyinput16), .C1(n2539), .C2(keyinput17), 
        .A(n4707), .ZN(n4718) );
  AOI22_X1 U5206 ( .A1(n4711), .A2(keyinput21), .B1(keyinput18), .B2(n4710), 
        .ZN(n4709) );
  OAI221_X1 U5207 ( .B1(n4711), .B2(keyinput21), .C1(n4710), .C2(keyinput18), 
        .A(n4709), .ZN(n4717) );
  XNOR2_X1 U5208 ( .A(IR_REG_1__SCAN_IN), .B(keyinput14), .ZN(n4715) );
  XNOR2_X1 U5209 ( .A(IR_REG_20__SCAN_IN), .B(keyinput12), .ZN(n4714) );
  XNOR2_X1 U5210 ( .A(D_REG_0__SCAN_IN), .B(keyinput13), .ZN(n4713) );
  XNOR2_X1 U5211 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput10), .ZN(n4712) );
  NAND4_X1 U5212 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4716)
         );
  NOR3_X1 U5213 ( .A1(n4718), .A2(n4717), .A3(n4716), .ZN(n4733) );
  AOI22_X1 U5214 ( .A1(n4721), .A2(keyinput5), .B1(n4720), .B2(keyinput2), 
        .ZN(n4719) );
  OAI221_X1 U5215 ( .B1(n4721), .B2(keyinput5), .C1(n4720), .C2(keyinput2), 
        .A(n4719), .ZN(n4731) );
  XNOR2_X1 U5216 ( .A(keyinput1), .B(n4722), .ZN(n4730) );
  XNOR2_X1 U5217 ( .A(keyinput9), .B(n4723), .ZN(n4729) );
  XNOR2_X1 U5218 ( .A(REG3_REG_11__SCAN_IN), .B(keyinput8), .ZN(n4727) );
  XNOR2_X1 U5219 ( .A(IR_REG_26__SCAN_IN), .B(keyinput0), .ZN(n4726) );
  XNOR2_X1 U5220 ( .A(IR_REG_30__SCAN_IN), .B(keyinput4), .ZN(n4725) );
  XNOR2_X1 U5221 ( .A(keyinput6), .B(D_REG_6__SCAN_IN), .ZN(n4724) );
  NAND4_X1 U5222 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4728)
         );
  NOR4_X1 U5223 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4732)
         );
  NAND4_X1 U5224 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n4736)
         );
  AOI211_X1 U5225 ( .C1(n4739), .C2(n4738), .A(n4737), .B(n4736), .ZN(n4740)
         );
  XNOR2_X1 U5226 ( .A(n4741), .B(n4740), .ZN(U3294) );
  CLKBUF_X1 U2324 ( .A(n2437), .Z(n2440) );
  CLKBUF_X1 U2474 ( .A(n3584), .Z(n3811) );
endmodule

