

module b22_C_AntiSAT_k_256_4 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631;

  INV_X4 U7386 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7387 ( .A1(n12107), .A2(n12106), .ZN(n12634) );
  INV_X2 U7389 ( .A(n6646), .ZN(n11698) );
  INV_X1 U7390 ( .A(n12236), .ZN(n12069) );
  INV_X2 U7391 ( .A(n10521), .ZN(n6646) );
  NAND2_X1 U7392 ( .A1(n9379), .A2(n9378), .ZN(n11094) );
  INV_X2 U7393 ( .A(n12397), .ZN(n12409) );
  AND3_X1 U7394 ( .A1(n7949), .A2(n7948), .A3(n7944), .ZN(n8214) );
  CLKBUF_X2 U7395 ( .A(n8514), .Z(n12024) );
  CLKBUF_X2 U7396 ( .A(n10884), .Z(n6639) );
  NAND4_X1 U7397 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(n13156)
         );
  CLKBUF_X2 U7398 ( .A(n8723), .Z(n11169) );
  INV_X2 U7399 ( .A(n11363), .ZN(n11358) );
  INV_X1 U7400 ( .A(n11612), .ZN(n11897) );
  CLKBUF_X2 U7401 ( .A(n11333), .Z(n11318) );
  AND3_X1 U7402 ( .A1(n8958), .A2(n8957), .A3(n8956), .ZN(n15137) );
  CLKBUF_X2 U7403 ( .A(n9114), .Z(n6640) );
  AND4_X1 U7404 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .ZN(n11728)
         );
  INV_X1 U7405 ( .A(n11578), .ZN(n11528) );
  XNOR2_X1 U7406 ( .A(n7131), .B(n8105), .ZN(n8106) );
  INV_X2 U7407 ( .A(n6642), .ZN(n6644) );
  XNOR2_X1 U7408 ( .A(n8171), .B(n14357), .ZN(n8173) );
  NAND2_X1 U7409 ( .A1(n7766), .A2(n7705), .ZN(n7809) );
  INV_X1 U7410 ( .A(n11737), .ZN(n11898) );
  INV_X1 U7411 ( .A(n14719), .ZN(n7433) );
  AND2_X1 U7412 ( .A1(n8129), .A2(n12992), .ZN(n12223) );
  NAND2_X1 U7413 ( .A1(n11980), .A2(n12370), .ZN(n12755) );
  NAND2_X1 U7414 ( .A1(n12271), .A2(n12283), .ZN(n15126) );
  NAND2_X1 U7415 ( .A1(n13670), .A2(n8333), .ZN(n8729) );
  INV_X1 U7417 ( .A(n11680), .ZN(n11696) );
  INV_X1 U7418 ( .A(n11878), .ZN(n6642) );
  INV_X1 U7419 ( .A(n10977), .ZN(n12222) );
  XNOR2_X1 U7420 ( .A(n10073), .B(n10089), .ZN(n14983) );
  AND2_X1 U7421 ( .A1(n12406), .A2(n12640), .ZN(n12651) );
  AND2_X1 U7422 ( .A1(n7824), .A2(n7825), .ZN(n8475) );
  NAND2_X1 U7424 ( .A1(n13666), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8329) );
  INV_X1 U7425 ( .A(n11881), .ZN(n11885) );
  INV_X1 U7426 ( .A(n11787), .ZN(n14582) );
  NAND2_X1 U7427 ( .A1(n10296), .A2(n10295), .ZN(n12076) );
  NAND2_X1 U7428 ( .A1(n12992), .A2(n12990), .ZN(n10977) );
  AND4_X1 U7429 ( .A1(n9607), .A2(n9606), .A3(n9605), .A4(n9604), .ZN(n9849)
         );
  NAND2_X1 U7430 ( .A1(n12306), .A2(n12307), .ZN(n12310) );
  NAND2_X1 U7431 ( .A1(n7696), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U7432 ( .A1(n8903), .A2(n8902), .ZN(n11068) );
  NAND2_X1 U7433 ( .A1(n8894), .A2(n8893), .ZN(n14926) );
  NAND2_X2 U7434 ( .A1(n11273), .A2(n11272), .ZN(n13547) );
  OAI21_X1 U7435 ( .B1(n13374), .B2(n13435), .A(n13373), .ZN(n13551) );
  INV_X1 U7436 ( .A(n14694), .ZN(n14200) );
  AOI21_X1 U7437 ( .B1(n12425), .B2(n12424), .A(n6867), .ZN(n12433) );
  XNOR2_X1 U7438 ( .A(n7697), .B(n7690), .ZN(n10474) );
  XNOR2_X1 U7439 ( .A(n8489), .B(n8488), .ZN(n12601) );
  INV_X4 U7440 ( .A(n11898), .ZN(n6808) );
  XNOR2_X1 U7441 ( .A(n8240), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9114) );
  AND2_X1 U7442 ( .A1(n8129), .A2(n8128), .ZN(n8514) );
  INV_X2 U7443 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8341) );
  NOR2_X4 U7444 ( .A1(n7104), .A2(n8234), .ZN(n7674) );
  NAND2_X2 U7445 ( .A1(n8028), .A2(n8027), .ZN(n8032) );
  NAND2_X2 U7446 ( .A1(n8009), .A2(n8008), .ZN(n8028) );
  NAND2_X4 U7447 ( .A1(n11637), .A2(n11636), .ZN(n14030) );
  NAND2_X2 U7448 ( .A1(n14545), .A2(n10691), .ZN(n10952) );
  NAND2_X2 U7449 ( .A1(n8168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7975) );
  OAI21_X2 U7450 ( .B1(n11895), .B2(n11894), .A(n7312), .ZN(n7311) );
  NAND4_X2 U7451 ( .A1(n7658), .A2(n15477), .A3(n7657), .A4(n8803), .ZN(n8234)
         );
  OR2_X4 U7452 ( .A1(n7790), .A2(n7183), .ZN(n8744) );
  AOI22_X2 U7453 ( .A1(n13859), .A2(n13860), .B1(n13870), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n8046) );
  INV_X2 U7454 ( .A(n12634), .ZN(n12641) );
  INV_X2 U7455 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15496) );
  AND2_X2 U7456 ( .A1(n7684), .A2(n7805), .ZN(n7505) );
  OAI21_X2 U7457 ( .B1(n9632), .B2(n9631), .A(n9634), .ZN(n9825) );
  AND2_X2 U7458 ( .A1(n13308), .A2(n13309), .ZN(n13367) );
  NAND2_X2 U7459 ( .A1(n15036), .A2(n10078), .ZN(n10079) );
  XNOR2_X2 U7460 ( .A(n14712), .B(n13829), .ZN(n11922) );
  XNOR2_X2 U7461 ( .A(n12476), .B(n12484), .ZN(n12456) );
  NAND2_X1 U7462 ( .A1(n8275), .A2(n11908), .ZN(n14676) );
  NOR2_X2 U7463 ( .A1(n10436), .A2(n10437), .ZN(n10441) );
  NOR2_X2 U7464 ( .A1(n10174), .A2(n10175), .ZN(n10436) );
  NAND2_X1 U7465 ( .A1(n10477), .A2(n12313), .ZN(n10531) );
  XNOR2_X2 U7466 ( .A(n11094), .B(n11096), .ZN(n11409) );
  NOR2_X2 U7467 ( .A1(n15629), .A2(n14429), .ZN(n14433) );
  NAND3_X2 U7468 ( .A1(n7069), .A2(n7067), .A3(n7065), .ZN(n14653) );
  OAI21_X2 U7469 ( .B1(n13090), .B2(n13005), .A(n13088), .ZN(n13094) );
  NOR2_X2 U7470 ( .A1(n10955), .A2(n10956), .ZN(n13090) );
  AND2_X2 U7471 ( .A1(n13024), .A2(n6756), .ZN(n7352) );
  AOI211_X1 U7472 ( .C1(n11107), .C2(n13128), .A(n9901), .B(n9900), .ZN(n9902)
         );
  NOR3_X2 U7473 ( .A1(n12464), .A2(n12463), .A3(n12462), .ZN(n12482) );
  INV_X2 U7474 ( .A(n8335), .ZN(n13670) );
  XNOR2_X2 U7475 ( .A(n8329), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8335) );
  AOI21_X2 U7476 ( .B1(n7265), .B2(n7269), .A(n7263), .ZN(n7262) );
  NOR2_X2 U7477 ( .A1(n10503), .A2(n7266), .ZN(n7265) );
  INV_X4 U7478 ( .A(n10289), .ZN(n12117) );
  INV_X4 U7479 ( .A(n8753), .ZN(n10289) );
  NOR2_X2 U7480 ( .A1(n14487), .A2(n14486), .ZN(n14485) );
  NAND2_X2 U7481 ( .A1(n9085), .A2(n9084), .ZN(n9153) );
  NAND4_X2 U7482 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7454) );
  OAI21_X2 U7483 ( .B1(n10771), .B2(n10770), .A(n10772), .ZN(n11963) );
  NAND2_X2 U7484 ( .A1(n10584), .A2(n10583), .ZN(n10771) );
  AOI211_X2 U7485 ( .C1(n14938), .C2(n13553), .A(n13552), .B(n13551), .ZN(
        n13634) );
  AND2_X1 U7486 ( .A1(n8172), .A2(n8173), .ZN(n11878) );
  NOR2_X2 U7487 ( .A1(n15062), .A2(n15061), .ZN(n15060) );
  NOR2_X2 U7488 ( .A1(n15043), .A2(n10143), .ZN(n15062) );
  INV_X1 U7489 ( .A(n7737), .ZN(n11345) );
  OAI222_X1 U7490 ( .A1(n12985), .A2(n13000), .B1(P3_U3151), .B2(n12998), .C1(
        n12997), .C2(n12996), .ZN(P3_U3267) );
  NAND2_X2 U7491 ( .A1(n6802), .A2(n6800), .ZN(n12998) );
  XNOR2_X2 U7492 ( .A(n8239), .B(n8238), .ZN(n11315) );
  OAI21_X2 U7493 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10073) );
  BUF_X8 U7494 ( .A(n12223), .Z(n6638) );
  NAND2_X2 U7495 ( .A1(n14988), .A2(n10136), .ZN(n7182) );
  AOI21_X2 U7496 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14436), .A(n15625), .ZN(
        n15618) );
  OR2_X1 U7497 ( .A1(n9695), .A2(n11409), .ZN(n10234) );
  NAND4_X2 U7498 ( .A1(n8791), .A2(n8790), .A3(n8789), .A4(n8788), .ZN(n13154)
         );
  AOI21_X2 U7499 ( .B1(n6906), .B2(n7346), .A(n7345), .ZN(n14381) );
  XNOR2_X2 U7500 ( .A(n10434), .B(n10435), .ZN(n10174) );
  AND2_X2 U7501 ( .A1(n7165), .A2(n7166), .ZN(n10434) );
  OR2_X2 U7502 ( .A1(n15079), .A2(n6778), .ZN(n7166) );
  OAI22_X4 U7503 ( .A1(n13112), .A2(n13110), .B1(n13023), .B2(n13022), .ZN(
        n13024) );
  XNOR2_X2 U7504 ( .A(n13020), .B(n13021), .ZN(n13112) );
  NAND4_X2 U7505 ( .A1(n8857), .A2(n8856), .A3(n8855), .A4(n8854), .ZN(n13831)
         );
  OAI21_X2 U7506 ( .B1(n12460), .B2(n10445), .A(n12455), .ZN(n12476) );
  AOI22_X2 U7507 ( .A1(n11865), .A2(n11864), .B1(n11863), .B2(n11862), .ZN(
        n11868) );
  NOR2_X2 U7508 ( .A1(n15147), .A2(n8700), .ZN(n15144) );
  OAI21_X2 U7509 ( .B1(n10662), .B2(n6744), .A(n7440), .ZN(n13770) );
  OAI22_X2 U7510 ( .A1(n10661), .A2(n10660), .B1(n10659), .B2(n7418), .ZN(
        n10662) );
  OAI21_X2 U7511 ( .B1(n9960), .B2(n9959), .A(n9961), .ZN(n10466) );
  XNOR2_X2 U7512 ( .A(n7903), .B(P2_IR_REG_2__SCAN_IN), .ZN(n14760) );
  BUF_X8 U7513 ( .A(n11345), .Z(n6641) );
  XNOR2_X1 U7514 ( .A(n11107), .B(n13001), .ZN(n9922) );
  INV_X1 U7515 ( .A(n6642), .ZN(n6643) );
  INV_X2 U7516 ( .A(n6642), .ZN(n6645) );
  INV_X2 U7517 ( .A(n11984), .ZN(n12235) );
  XOR2_X2 U7518 ( .A(n12577), .B(n12575), .Z(n12578) );
  XNOR2_X2 U7519 ( .A(n6828), .B(n12527), .ZN(n12500) );
  NAND2_X2 U7520 ( .A1(n7180), .A2(n7179), .ZN(n6828) );
  INV_X8 U7521 ( .A(n12426), .ZN(n6648) );
  NOR2_X2 U7522 ( .A1(n14485), .A2(n14434), .ZN(n15627) );
  XNOR2_X2 U7523 ( .A(n7176), .B(n15051), .ZN(n15044) );
  NAND2_X2 U7524 ( .A1(n7178), .A2(n7177), .ZN(n7176) );
  XNOR2_X1 U7525 ( .A(n14443), .B(n14793), .ZN(n14490) );
  NAND2_X2 U7526 ( .A1(n15619), .A2(n14442), .ZN(n14443) );
  NOR3_X2 U7527 ( .A1(n10455), .A2(n10454), .A3(n10453), .ZN(n12464) );
  NOR2_X2 U7528 ( .A1(n10186), .A2(n10185), .ZN(n10455) );
  OAI21_X1 U7529 ( .B1(n14649), .B2(n14648), .A(n7294), .ZN(n7293) );
  OAI21_X1 U7530 ( .B1(n13281), .B2(n13282), .A(n13284), .ZN(n13497) );
  OAI21_X1 U7531 ( .B1(n10901), .B2(n10900), .A(n10903), .ZN(n13281) );
  NAND2_X1 U7532 ( .A1(n14638), .A2(n14640), .ZN(n14645) );
  OR2_X1 U7533 ( .A1(n10441), .A2(n10440), .ZN(n12452) );
  NOR2_X1 U7534 ( .A1(n10084), .A2(n10085), .ZN(n10176) );
  AOI21_X1 U7535 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15068), .A(n15060), .ZN(
        n10146) );
  NAND2_X1 U7536 ( .A1(n15105), .A2(n10209), .ZN(n12307) );
  INV_X2 U7537 ( .A(n11730), .ZN(n11727) );
  NAND2_X1 U7538 ( .A1(n12292), .A2(n12296), .ZN(n12246) );
  INV_X1 U7539 ( .A(n13155), .ZN(n9283) );
  INV_X1 U7540 ( .A(n13154), .ZN(n9296) );
  INV_X1 U7541 ( .A(n15131), .ZN(n12448) );
  INV_X1 U7542 ( .A(n9359), .ZN(n15150) );
  INV_X1 U7543 ( .A(n15129), .ZN(n12447) );
  XNOR2_X2 U7544 ( .A(n13067), .B(n6820), .ZN(n8735) );
  INV_X4 U7545 ( .A(n11053), .ZN(n11338) );
  INV_X2 U7546 ( .A(n11067), .ZN(n11053) );
  AND2_X1 U7548 ( .A1(n11315), .A2(n11429), .ZN(n14958) );
  INV_X2 U7549 ( .A(n13227), .ZN(n11168) );
  NAND2_X2 U7550 ( .A1(n11008), .A2(n14653), .ZN(n11578) );
  AND2_X2 U7551 ( .A1(n9095), .A2(n7649), .ZN(n7974) );
  INV_X2 U7552 ( .A(n7737), .ZN(n8346) );
  AND4_X2 U7553 ( .A1(n7715), .A2(n7713), .A3(n7714), .A4(n7511), .ZN(n9095)
         );
  INV_X1 U7554 ( .A(n7809), .ZN(n7715) );
  INV_X2 U7555 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7132) );
  NOR2_X4 U7556 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7766) );
  CLKBUF_X2 U7557 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14654) );
  AND2_X1 U7558 ( .A1(n14232), .A2(n14231), .ZN(n14324) );
  OR2_X1 U7559 ( .A1(n11448), .A2(n7479), .ZN(n7478) );
  AND2_X1 U7560 ( .A1(n7213), .A2(n12239), .ZN(n12418) );
  NOR2_X1 U7561 ( .A1(n13987), .A2(n13986), .ZN(n14232) );
  OR2_X1 U7562 ( .A1(n12240), .A2(n12619), .ZN(n7213) );
  NAND2_X1 U7563 ( .A1(n12652), .A2(n12651), .ZN(n12650) );
  NAND2_X1 U7564 ( .A1(n12052), .A2(n12403), .ZN(n12652) );
  XNOR2_X1 U7565 ( .A(n13233), .B(n13239), .ZN(n11438) );
  AND2_X1 U7566 ( .A1(n11855), .A2(n11854), .ZN(n11859) );
  NAND2_X1 U7567 ( .A1(n12071), .A2(n12070), .ZN(n12161) );
  AND2_X1 U7568 ( .A1(n7060), .A2(n6786), .ZN(n14314) );
  AND2_X1 U7569 ( .A1(n11877), .A2(n11876), .ZN(n14318) );
  NAND2_X1 U7570 ( .A1(n11311), .A2(n11310), .ZN(n13246) );
  OAI21_X1 U7571 ( .B1(n12068), .B2(n11967), .A(n11968), .ZN(n12218) );
  NAND2_X1 U7572 ( .A1(n7056), .A2(n7055), .ZN(n13539) );
  OAI211_X1 U7573 ( .C1(n11357), .C2(n11356), .A(n11355), .B(n11354), .ZN(
        n13665) );
  NAND2_X1 U7574 ( .A1(n12055), .A2(n12054), .ZN(n12657) );
  INV_X1 U7575 ( .A(n7527), .ZN(n7526) );
  NAND2_X1 U7576 ( .A1(n11329), .A2(n11328), .ZN(n13534) );
  XNOR2_X1 U7577 ( .A(n11309), .B(n11308), .ZN(n13669) );
  OR2_X1 U7578 ( .A1(n12683), .A2(n12684), .ZN(n12681) );
  NAND2_X1 U7579 ( .A1(n11871), .A2(n11870), .ZN(n13961) );
  NAND2_X1 U7580 ( .A1(n11965), .A2(n11964), .ZN(n12068) );
  NAND2_X1 U7581 ( .A1(n12044), .A2(n12043), .ZN(n12861) );
  AND2_X2 U7582 ( .A1(n11686), .A2(n11685), .ZN(n14323) );
  AND2_X1 U7583 ( .A1(n13354), .A2(n6705), .ZN(n7055) );
  NOR2_X1 U7584 ( .A1(n13404), .A2(n7395), .ZN(n6920) );
  NAND2_X2 U7585 ( .A1(n11365), .A2(n11364), .ZN(n13336) );
  BUF_X1 U7586 ( .A(n13404), .Z(n6836) );
  NAND2_X1 U7587 ( .A1(n13406), .A2(n13405), .ZN(n13404) );
  NAND2_X1 U7588 ( .A1(n7113), .A2(n7112), .ZN(n13377) );
  XNOR2_X1 U7589 ( .A(n11327), .B(n11326), .ZN(n13672) );
  NAND2_X1 U7590 ( .A1(n11668), .A2(n11667), .ZN(n13991) );
  NAND2_X1 U7591 ( .A1(n6972), .A2(n14070), .ZN(n14069) );
  OAI21_X1 U7592 ( .B1(n11007), .B2(n11006), .A(n11304), .ZN(n11684) );
  INV_X1 U7593 ( .A(n13393), .ZN(n7113) );
  INV_X1 U7594 ( .A(n14018), .ZN(n6647) );
  NAND2_X1 U7595 ( .A1(n11007), .A2(n11006), .ZN(n11304) );
  NAND2_X1 U7596 ( .A1(n12021), .A2(n12020), .ZN(n12700) );
  AND2_X1 U7597 ( .A1(n11652), .A2(n11651), .ZN(n14007) );
  NAND2_X1 U7598 ( .A1(n7115), .A2(n7114), .ZN(n13393) );
  NAND2_X1 U7599 ( .A1(n14089), .A2(n14066), .ZN(n6972) );
  NAND2_X1 U7600 ( .A1(n7417), .A2(n13299), .ZN(n13416) );
  AOI21_X1 U7601 ( .B1(n12708), .B2(n12099), .A(n6695), .ZN(n12692) );
  NAND2_X1 U7602 ( .A1(n11251), .A2(n11250), .ZN(n13379) );
  NAND2_X1 U7603 ( .A1(n14110), .A2(n13921), .ZN(n14089) );
  OAI21_X1 U7604 ( .B1(n14517), .B2(n14516), .A(n6909), .ZN(n6819) );
  NAND2_X1 U7605 ( .A1(n7032), .A2(n7031), .ZN(n7246) );
  AND2_X1 U7606 ( .A1(n7331), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U7607 ( .A1(n7211), .A2(n10471), .ZN(n10561) );
  NAND2_X1 U7608 ( .A1(n7293), .A2(n14647), .ZN(n14517) );
  CLKBUF_X1 U7609 ( .A(n13497), .Z(n6916) );
  NAND2_X1 U7610 ( .A1(n7064), .A2(n10749), .ZN(n10934) );
  OAI21_X1 U7611 ( .B1(n14645), .B2(n14644), .A(n15524), .ZN(n6864) );
  AND2_X1 U7612 ( .A1(n10933), .A2(n7467), .ZN(n7064) );
  OAI21_X1 U7613 ( .B1(n14169), .B2(n7545), .A(n7543), .ZN(n14150) );
  OR2_X1 U7614 ( .A1(n10748), .A2(SI_24_), .ZN(n10749) );
  NAND2_X1 U7615 ( .A1(n10748), .A2(SI_24_), .ZN(n10933) );
  NAND2_X1 U7616 ( .A1(n7210), .A2(n7209), .ZN(n9647) );
  AND2_X1 U7617 ( .A1(n14375), .A2(n11578), .ZN(n14263) );
  AND2_X1 U7618 ( .A1(n14147), .A2(n14160), .ZN(n11913) );
  NAND2_X1 U7619 ( .A1(n11531), .A2(n11530), .ZN(n14133) );
  INV_X1 U7620 ( .A(n14284), .ZN(n14147) );
  AND2_X1 U7621 ( .A1(n14284), .A2(n13915), .ZN(n11814) );
  AND2_X1 U7622 ( .A1(n10545), .A2(n7046), .ZN(n6873) );
  AOI21_X1 U7623 ( .B1(n12818), .B2(n12085), .A(n12084), .ZN(n12805) );
  OAI21_X1 U7624 ( .B1(n10711), .B2(n10642), .A(n10643), .ZN(n10830) );
  NAND2_X1 U7625 ( .A1(n11516), .A2(n11515), .ZN(n14284) );
  NAND2_X1 U7626 ( .A1(n9924), .A2(n9905), .ZN(n9908) );
  OAI21_X1 U7627 ( .B1(n14604), .B2(n11915), .A(n10825), .ZN(n13909) );
  OR2_X1 U7628 ( .A1(n10315), .A2(SI_22_), .ZN(n10316) );
  NAND2_X1 U7629 ( .A1(n10315), .A2(SI_22_), .ZN(n10545) );
  XNOR2_X1 U7630 ( .A(n9405), .B(n9593), .ZN(n9404) );
  OR2_X1 U7631 ( .A1(n11514), .A2(n11612), .ZN(n11516) );
  NAND2_X1 U7632 ( .A1(n9776), .A2(n9440), .ZN(n11514) );
  NAND2_X1 U7633 ( .A1(n10925), .A2(n12335), .ZN(n11973) );
  NOR2_X2 U7634 ( .A1(n10713), .A2(n13618), .ZN(n10712) );
  NAND2_X1 U7635 ( .A1(n10236), .A2(n10235), .ZN(n10355) );
  XNOR2_X1 U7636 ( .A(n6907), .B(n14464), .ZN(n14633) );
  NAND2_X1 U7637 ( .A1(n6915), .A2(n9577), .ZN(n9776) );
  NAND2_X1 U7638 ( .A1(n10234), .A2(n10233), .ZN(n10236) );
  NAND2_X1 U7639 ( .A1(n7304), .A2(n7305), .ZN(n6907) );
  AND2_X1 U7640 ( .A1(n13936), .A2(n11809), .ZN(n13934) );
  NAND2_X1 U7641 ( .A1(n9586), .A2(SI_20_), .ZN(n9935) );
  OR2_X1 U7642 ( .A1(n10518), .A2(n6753), .ZN(n7420) );
  OR2_X1 U7643 ( .A1(n9583), .A2(n9578), .ZN(n9775) );
  NAND2_X1 U7644 ( .A1(n7108), .A2(n7107), .ZN(n10360) );
  OAI21_X1 U7645 ( .B1(n9673), .B2(n9672), .A(n9674), .ZN(n9694) );
  AND2_X1 U7646 ( .A1(n11490), .A2(n11489), .ZN(n14181) );
  NAND2_X1 U7647 ( .A1(n10248), .A2(n10247), .ZN(n11787) );
  AND2_X1 U7648 ( .A1(n7167), .A2(n6779), .ZN(n7165) );
  NAND3_X1 U7649 ( .A1(n9132), .A2(n6928), .A3(n7382), .ZN(n9266) );
  OAI211_X1 U7650 ( .C1(n7075), .C2(n9315), .A(n7074), .B(n9314), .ZN(n9320)
         );
  NAND2_X1 U7651 ( .A1(n14491), .A2(n14456), .ZN(n14458) );
  NAND2_X1 U7652 ( .A1(n15071), .A2(n10081), .ZN(n10082) );
  NAND2_X1 U7653 ( .A1(n9518), .A2(n9517), .ZN(n14715) );
  NAND2_X2 U7654 ( .A1(n9011), .A2(n9010), .ZN(n11075) );
  OR2_X2 U7655 ( .A1(n9310), .A2(n11236), .ZN(n9011) );
  INV_X1 U7656 ( .A(n9627), .ZN(n7606) );
  NAND2_X1 U7657 ( .A1(n9278), .A2(n9277), .ZN(n9557) );
  NAND2_X1 U7658 ( .A1(n7954), .A2(n7925), .ZN(n9310) );
  INV_X2 U7659 ( .A(n15162), .ZN(n12846) );
  NAND2_X2 U7660 ( .A1(n13954), .A2(n14683), .ZN(n14686) );
  XNOR2_X1 U7661 ( .A(n7182), .B(n15016), .ZN(n15008) );
  CLKBUF_X1 U7662 ( .A(n13159), .Z(n6917) );
  NAND2_X1 U7663 ( .A1(n8732), .A2(n6876), .ZN(n13155) );
  BUF_X1 U7664 ( .A(n11037), .Z(n11034) );
  OR2_X1 U7665 ( .A1(n14991), .A2(n14990), .ZN(n14988) );
  NAND2_X2 U7666 ( .A1(n8758), .A2(n15149), .ZN(n12202) );
  INV_X1 U7667 ( .A(n9849), .ZN(n15105) );
  INV_X1 U7668 ( .A(n11728), .ZN(n14196) );
  NAND4_X1 U7669 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n13832)
         );
  AND2_X1 U7670 ( .A1(n7471), .A2(n7053), .ZN(n7052) );
  AND4_X1 U7671 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(n9506)
         );
  OR2_X2 U7672 ( .A1(n6658), .A2(n8349), .ZN(n8350) );
  INV_X1 U7673 ( .A(n8729), .ZN(n9136) );
  AND4_X2 U7674 ( .A1(n8762), .A2(n8761), .A3(n8759), .A4(n8760), .ZN(n9359)
         );
  AND4_X1 U7675 ( .A1(n8967), .A2(n8966), .A3(n8965), .A4(n8964), .ZN(n15129)
         );
  INV_X1 U7676 ( .A(n11318), .ZN(n11372) );
  AND2_X2 U7677 ( .A1(n11901), .A2(n8208), .ZN(n10521) );
  OR2_X2 U7678 ( .A1(n14676), .A2(n11907), .ZN(n14719) );
  CLKBUF_X3 U7679 ( .A(n8729), .Z(n6658) );
  NAND2_X1 U7680 ( .A1(n7832), .A2(n7831), .ZN(n9708) );
  NAND2_X2 U7681 ( .A1(n10270), .A2(n6641), .ZN(n12236) );
  NAND2_X1 U7682 ( .A1(n8344), .A2(n13227), .ZN(n14949) );
  CLKBUF_X3 U7683 ( .A(n8852), .Z(n11656) );
  XNOR2_X1 U7684 ( .A(n14386), .B(n15435), .ZN(n14439) );
  AND2_X1 U7685 ( .A1(n11168), .A2(n11427), .ZN(n11429) );
  INV_X1 U7686 ( .A(n6899), .ZN(n14386) );
  NAND2_X2 U7687 ( .A1(n8175), .A2(n8176), .ZN(n11704) );
  NAND2_X2 U7688 ( .A1(n8172), .A2(n8175), .ZN(n11881) );
  NAND2_X1 U7689 ( .A1(n7476), .A2(n8410), .ZN(n7475) );
  AND2_X1 U7690 ( .A1(n7971), .A2(n7970), .ZN(n8279) );
  NAND2_X1 U7691 ( .A1(n6792), .A2(n7741), .ZN(n7749) );
  XNOR2_X1 U7692 ( .A(n7723), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7949) );
  INV_X1 U7693 ( .A(n8333), .ZN(n13674) );
  OR2_X1 U7694 ( .A1(n8103), .A2(n8104), .ZN(n6802) );
  XNOR2_X1 U7695 ( .A(n8185), .B(n8184), .ZN(n13891) );
  NAND2_X1 U7696 ( .A1(n8324), .A2(n8323), .ZN(n13227) );
  NAND2_X1 U7697 ( .A1(n7730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7723) );
  XNOR2_X1 U7698 ( .A(n8331), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8333) );
  OAI21_X1 U7699 ( .B1(n8102), .B2(n7508), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8103) );
  XNOR2_X1 U7700 ( .A(n8126), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U7701 ( .A1(n7000), .A2(n6999), .ZN(n12992) );
  NAND2_X1 U7702 ( .A1(n6843), .A2(n6713), .ZN(n11000) );
  NOR2_X1 U7703 ( .A1(n14382), .A2(n14383), .ZN(n14385) );
  NAND2_X1 U7704 ( .A1(n12982), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8126) );
  OR2_X1 U7705 ( .A1(n7728), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n7730) );
  OR2_X1 U7706 ( .A1(n8182), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n7970) );
  OR2_X1 U7707 ( .A1(n8330), .A2(n8652), .ZN(n8331) );
  NAND2_X1 U7708 ( .A1(n7974), .A2(n7629), .ZN(n14360) );
  OAI21_X1 U7709 ( .B1(n7694), .B2(n6738), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7131) );
  OAI21_X1 U7710 ( .B1(n8319), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8239) );
  OR3_X1 U7711 ( .A1(n7974), .A2(n7976), .A3(n7917), .ZN(n7069) );
  NAND2_X2 U7712 ( .A1(n6641), .A2(P2_U3088), .ZN(n13675) );
  NAND2_X2 U7713 ( .A1(n6641), .A2(P1_U3086), .ZN(n14370) );
  NAND2_X1 U7714 ( .A1(n7505), .A2(n7502), .ZN(n7694) );
  AND2_X1 U7716 ( .A1(n9095), .A2(n7716), .ZN(n9171) );
  AND4_X1 U7717 ( .A1(n9071), .A2(n8236), .A3(n8235), .A4(n15363), .ZN(n7648)
         );
  INV_X1 U7718 ( .A(n6829), .ZN(n7790) );
  NAND2_X1 U7719 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n14426), .ZN(n14425) );
  AND4_X1 U7720 ( .A1(n7708), .A2(n9162), .A3(n7707), .A4(n7706), .ZN(n7714)
         );
  AND4_X1 U7721 ( .A1(n7712), .A2(n7711), .A3(n7710), .A4(n7709), .ZN(n7713)
         );
  AND2_X1 U7722 ( .A1(n6955), .A2(n6957), .ZN(n6954) );
  XNOR2_X1 U7723 ( .A(n6861), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n14424) );
  NAND2_X1 U7724 ( .A1(n7133), .A2(n7132), .ZN(n6829) );
  AND3_X1 U7725 ( .A1(n7491), .A2(n7006), .A3(n7133), .ZN(n7805) );
  AND2_X1 U7726 ( .A1(n7659), .A2(n7676), .ZN(n7660) );
  INV_X1 U7727 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n7676) );
  NOR2_X1 U7728 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6955) );
  NOR2_X1 U7729 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7680) );
  INV_X4 U7730 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7731 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7732 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6861) );
  INV_X1 U7733 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n15362) );
  INV_X1 U7734 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15447) );
  INV_X1 U7735 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7734) );
  INV_X1 U7736 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7733) );
  INV_X1 U7737 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9162) );
  INV_X1 U7738 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7511) );
  NOR2_X1 U7739 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7709) );
  NOR2_X1 U7740 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n7710) );
  NOR2_X1 U7741 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7711) );
  OR2_X1 U7742 ( .A1(n13334), .A2(n13312), .ZN(n7042) );
  XNOR2_X1 U7743 ( .A(n12127), .B(n6771), .ZN(n12138) );
  NAND2_X1 U7744 ( .A1(n8475), .A2(n7835), .ZN(n7832) );
  XNOR2_X1 U7745 ( .A(n12117), .B(n15137), .ZN(n9038) );
  CLKBUF_X1 U7746 ( .A(n14447), .Z(n6649) );
  CLKBUF_X1 U7747 ( .A(n14488), .Z(n6650) );
  OR2_X2 U7748 ( .A1(n10375), .A2(n11116), .ZN(n10713) );
  INV_X1 U7749 ( .A(n10072), .ZN(n6651) );
  XNOR2_X1 U7750 ( .A(n7792), .B(n7791), .ZN(n10129) );
  NAND2_X1 U7751 ( .A1(n14492), .A2(n14808), .ZN(n14491) );
  XNOR2_X1 U7752 ( .A(n9055), .B(n9054), .ZN(n9056) );
  NAND2_X1 U7753 ( .A1(n6805), .A2(n12271), .ZN(n15114) );
  NAND2_X1 U7754 ( .A1(n10197), .A2(n12300), .ZN(n10213) );
  AOI21_X2 U7755 ( .B1(n12650), .B2(n12408), .A(n12407), .ZN(n12229) );
  NAND2_X1 U7756 ( .A1(n7386), .A2(n6652), .ZN(n13327) );
  AND2_X1 U7757 ( .A1(n7387), .A2(n6653), .ZN(n6652) );
  INV_X1 U7758 ( .A(n13332), .ZN(n6653) );
  NAND2_X1 U7759 ( .A1(n6793), .A2(n6657), .ZN(n6654) );
  AND2_X1 U7760 ( .A1(n6654), .A2(n6655), .ZN(n10836) );
  OR2_X1 U7761 ( .A1(n6656), .A2(n10628), .ZN(n6655) );
  INV_X1 U7762 ( .A(n10833), .ZN(n6656) );
  AND2_X1 U7763 ( .A1(n11412), .A2(n10833), .ZN(n6657) );
  NAND2_X1 U7764 ( .A1(n9136), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8364) );
  OAI21_X2 U7765 ( .B1(n11271), .B2(n10996), .A(n10997), .ZN(n11002) );
  NAND2_X2 U7766 ( .A1(n7468), .A2(n10991), .ZN(n11271) );
  NOR2_X2 U7767 ( .A1(n12473), .A2(n12474), .ZN(n12475) );
  NOR2_X2 U7768 ( .A1(n12453), .A2(n15443), .ZN(n12473) );
  OAI22_X2 U7769 ( .A1(n12420), .A2(n12419), .B1(n12418), .B2(n12417), .ZN(
        n12421) );
  OAI211_X2 U7770 ( .C1(n12236), .C2(n7455), .A(n8748), .B(n8747), .ZN(n15156)
         );
  OR2_X1 U7771 ( .A1(n11984), .A2(n8746), .ZN(n8747) );
  NOR2_X2 U7772 ( .A1(n13439), .A2(n13423), .ZN(n7117) );
  NAND2_X2 U7773 ( .A1(n13460), .A2(n13648), .ZN(n13439) );
  AOI21_X2 U7774 ( .B1(n12587), .B2(n12586), .A(n12585), .ZN(n12596) );
  NOR2_X2 U7775 ( .A1(n15622), .A2(n14451), .ZN(n14454) );
  NAND2_X1 U7776 ( .A1(n11578), .A2(n6641), .ZN(n6659) );
  NAND2_X1 U7777 ( .A1(n11578), .A2(n6641), .ZN(n6660) );
  NAND2_X1 U7778 ( .A1(n11578), .A2(n6641), .ZN(n8839) );
  OAI21_X2 U7779 ( .B1(n13416), .B2(n13420), .A(n13301), .ZN(n13406) );
  NOR2_X2 U7780 ( .A1(n10426), .A2(n11792), .ZN(n14505) );
  NOR2_X2 U7781 ( .A1(n14601), .A2(n14602), .ZN(n6806) );
  NOR2_X2 U7782 ( .A1(n10046), .A2(n11765), .ZN(n10045) );
  XNOR2_X1 U7783 ( .A(n14533), .B(n12155), .ZN(n10290) );
  OR2_X1 U7784 ( .A1(n11972), .A2(n12636), .ZN(n12413) );
  INV_X1 U7785 ( .A(n13272), .ZN(n7241) );
  AND2_X1 U7786 ( .A1(n8279), .A2(n11902), .ZN(n11901) );
  NAND2_X1 U7787 ( .A1(n11868), .A2(n11867), .ZN(n6880) );
  NAND2_X1 U7788 ( .A1(n11873), .A2(n11874), .ZN(n7312) );
  NAND2_X1 U7789 ( .A1(n8176), .A2(n8173), .ZN(n8852) );
  NAND2_X1 U7790 ( .A1(n11071), .A2(n6710), .ZN(n6962) );
  NOR2_X1 U7791 ( .A1(n11071), .A2(n6710), .ZN(n6961) );
  OAI21_X1 U7792 ( .B1(n11064), .B2(n11063), .A(n11062), .ZN(n11072) );
  NAND2_X1 U7793 ( .A1(n6693), .A2(n6946), .ZN(n6944) );
  OR2_X1 U7794 ( .A1(n11101), .A2(n11104), .ZN(n11112) );
  AND2_X1 U7795 ( .A1(n11829), .A2(n11828), .ZN(n6914) );
  NOR2_X1 U7796 ( .A1(n11143), .A2(n11145), .ZN(n7583) );
  AND2_X1 U7797 ( .A1(n11194), .A2(n11195), .ZN(n7593) );
  OR2_X1 U7798 ( .A1(n11184), .A2(n11183), .ZN(n11196) );
  NAND2_X1 U7799 ( .A1(n7567), .A2(n11265), .ZN(n7566) );
  NAND2_X1 U7800 ( .A1(n7571), .A2(n7568), .ZN(n7567) );
  NOR2_X1 U7801 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7491) );
  INV_X1 U7802 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7133) );
  INV_X1 U7803 ( .A(n11633), .ZN(n7089) );
  NAND2_X1 U7804 ( .A1(n8029), .A2(SI_9_), .ZN(n8410) );
  NAND2_X1 U7805 ( .A1(n7290), .A2(n7291), .ZN(n7288) );
  NAND2_X1 U7806 ( .A1(n12104), .A2(n6688), .ZN(n7021) );
  INV_X1 U7807 ( .A(n12651), .ZN(n12104) );
  NAND2_X1 U7808 ( .A1(n12102), .A2(n7023), .ZN(n7022) );
  OR2_X1 U7809 ( .A1(n12657), .A2(n12667), .ZN(n12406) );
  OR2_X1 U7810 ( .A1(n12977), .A2(n11974), .ZN(n12344) );
  NAND2_X1 U7811 ( .A1(n15127), .A2(n15126), .ZN(n9361) );
  AOI21_X1 U7812 ( .B1(n7143), .B2(n12260), .A(n6736), .ZN(n7141) );
  INV_X1 U7813 ( .A(n7143), .ZN(n7142) );
  INV_X1 U7814 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15486) );
  NAND2_X1 U7815 ( .A1(n7966), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U7816 ( .A1(n8724), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7773) );
  INV_X1 U7817 ( .A(n13249), .ZN(n7239) );
  NAND2_X1 U7818 ( .A1(n13311), .A2(n11394), .ZN(n13332) );
  OR2_X1 U7819 ( .A1(n13588), .A2(n13457), .ZN(n7109) );
  AND3_X1 U7820 ( .A1(n8011), .A2(n7674), .A3(n7103), .ZN(n8241) );
  AND2_X1 U7821 ( .A1(n7660), .A2(n7663), .ZN(n7103) );
  INV_X1 U7822 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6956) );
  OR2_X1 U7823 ( .A1(n13730), .A2(n7424), .ZN(n7423) );
  XNOR2_X1 U7824 ( .A(n14314), .B(n11882), .ZN(n11943) );
  AND2_X1 U7825 ( .A1(n13923), .A2(n13922), .ZN(n7636) );
  INV_X1 U7826 ( .A(n8173), .ZN(n8175) );
  AOI21_X1 U7827 ( .B1(n6981), .B2(n6979), .A(n6729), .ZN(n6978) );
  INV_X1 U7828 ( .A(n13911), .ZN(n6979) );
  NOR2_X1 U7829 ( .A1(n9971), .A2(n7523), .ZN(n7522) );
  INV_X1 U7830 ( .A(n9970), .ZN(n7523) );
  NAND2_X1 U7831 ( .A1(n7323), .A2(n7320), .ZN(n11736) );
  NAND2_X1 U7832 ( .A1(n11327), .A2(n11326), .ZN(n11353) );
  INV_X1 U7833 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7736) );
  NAND2_X1 U7834 ( .A1(n7483), .A2(n7482), .ZN(n9588) );
  AOI21_X1 U7835 ( .B1(n7484), .B2(n7487), .A(n6777), .ZN(n7482) );
  AOI21_X1 U7836 ( .B1(n7052), .B2(n7474), .A(n6731), .ZN(n7051) );
  XNOR2_X1 U7837 ( .A(n8801), .B(SI_12_), .ZN(n8798) );
  NAND2_X1 U7838 ( .A1(n8006), .A2(SI_8_), .ZN(n8027) );
  OAI22_X1 U7839 ( .A1(n12206), .A2(n7287), .B1(n7288), .B2(n7285), .ZN(n7284)
         );
  INV_X1 U7840 ( .A(n7290), .ZN(n7287) );
  INV_X1 U7841 ( .A(n12176), .ZN(n7285) );
  INV_X1 U7842 ( .A(n7288), .ZN(n7286) );
  INV_X1 U7843 ( .A(n7265), .ZN(n7264) );
  OR2_X1 U7844 ( .A1(n12126), .A2(n12125), .ZN(n6813) );
  OR2_X1 U7845 ( .A1(n9723), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9832) );
  INV_X1 U7846 ( .A(n10268), .ZN(n7270) );
  INV_X1 U7847 ( .A(n10971), .ZN(n7247) );
  AND2_X1 U7848 ( .A1(n12990), .A2(n8128), .ZN(n10884) );
  INV_X1 U7849 ( .A(n12601), .ZN(n12614) );
  NAND2_X1 U7850 ( .A1(n12635), .A2(n12634), .ZN(n12633) );
  NAND2_X1 U7851 ( .A1(n12809), .A2(n12355), .ZN(n12799) );
  NAND2_X1 U7852 ( .A1(n12088), .A2(n12087), .ZN(n12795) );
  NAND2_X1 U7853 ( .A1(n9504), .A2(n7004), .ZN(n10200) );
  NOR2_X1 U7854 ( .A1(n12297), .A2(n7005), .ZN(n7004) );
  INV_X1 U7855 ( .A(n9503), .ZN(n7005) );
  AND2_X1 U7856 ( .A1(n9700), .A2(n12245), .ZN(n15154) );
  NAND2_X1 U7857 ( .A1(n11970), .A2(n11969), .ZN(n11972) );
  NOR2_X1 U7858 ( .A1(n7508), .A2(n7507), .ZN(n7506) );
  NAND2_X1 U7859 ( .A1(n8104), .A2(n7691), .ZN(n7507) );
  INV_X1 U7860 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8161) );
  AND2_X1 U7861 ( .A1(n8026), .A2(n8025), .ZN(n12484) );
  INV_X1 U7862 ( .A(n7189), .ZN(n7188) );
  OAI21_X1 U7863 ( .B1(n7883), .B2(n7190), .A(n7914), .ZN(n7189) );
  NAND2_X1 U7864 ( .A1(n13025), .A2(n7367), .ZN(n7366) );
  INV_X1 U7865 ( .A(n13026), .ZN(n7367) );
  INV_X1 U7866 ( .A(n9015), .ZN(n6837) );
  NOR2_X1 U7867 ( .A1(n13277), .A2(n7058), .ZN(n7057) );
  INV_X1 U7868 ( .A(n13275), .ZN(n7058) );
  INV_X1 U7869 ( .A(n13484), .ZN(n6903) );
  OR2_X1 U7870 ( .A1(n11116), .A2(n10369), .ZN(n10717) );
  NAND2_X1 U7871 ( .A1(n9669), .A2(n9668), .ZN(n9670) );
  NAND2_X1 U7872 ( .A1(n9281), .A2(n9280), .ZN(n10062) );
  INV_X2 U7873 ( .A(n11236), .ZN(n11362) );
  NAND2_X1 U7874 ( .A1(n7660), .A2(n8242), .ZN(n7554) );
  XNOR2_X1 U7875 ( .A(n8621), .B(n9054), .ZN(n8625) );
  NAND2_X1 U7876 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  OR2_X1 U7877 ( .A1(n7432), .A2(n14694), .ZN(n8619) );
  OAI21_X1 U7878 ( .B1(n6669), .B2(n7442), .A(n11471), .ZN(n7441) );
  INV_X1 U7879 ( .A(n7310), .ZN(n7309) );
  OAI21_X1 U7880 ( .B1(n7311), .B2(n6733), .A(n11896), .ZN(n7310) );
  INV_X1 U7881 ( .A(n13947), .ZN(n14034) );
  NAND2_X1 U7882 ( .A1(n14069), .A2(n7636), .ZN(n14061) );
  INV_X1 U7883 ( .A(n7617), .ZN(n7616) );
  AOI21_X1 U7884 ( .B1(n7617), .B2(n7615), .A(n6726), .ZN(n7614) );
  INV_X1 U7885 ( .A(n10502), .ZN(n7263) );
  NAND2_X1 U7886 ( .A1(n7411), .A2(n7409), .ZN(n13532) );
  AOI21_X1 U7887 ( .B1(n13142), .B2(n13120), .A(n7410), .ZN(n7409) );
  NOR2_X1 U7888 ( .A1(n13313), .A2(n13314), .ZN(n7410) );
  AND4_X1 U7889 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n14219) );
  NAND2_X1 U7890 ( .A1(n6795), .A2(n11753), .ZN(n6794) );
  INV_X1 U7891 ( .A(n11752), .ZN(n6795) );
  OR2_X1 U7892 ( .A1(n11777), .A2(n7344), .ZN(n7342) );
  NAND2_X1 U7893 ( .A1(n11086), .A2(n6763), .ZN(n7577) );
  AND2_X1 U7894 ( .A1(n6700), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U7895 ( .A1(n6700), .A2(n6941), .ZN(n6940) );
  NOR2_X1 U7896 ( .A1(n6693), .A2(n6946), .ZN(n6945) );
  NOR2_X1 U7897 ( .A1(n11913), .A2(n6826), .ZN(n11820) );
  OR2_X1 U7898 ( .A1(n11814), .A2(n6827), .ZN(n6826) );
  AND2_X1 U7899 ( .A1(n13914), .A2(n13913), .ZN(n6827) );
  INV_X1 U7900 ( .A(n6939), .ZN(n7555) );
  OAI21_X1 U7901 ( .B1(n11112), .B2(n11113), .A(n6676), .ZN(n6939) );
  INV_X1 U7902 ( .A(n11120), .ZN(n6950) );
  NAND2_X1 U7903 ( .A1(n6948), .A2(n6947), .ZN(n11136) );
  AOI21_X1 U7904 ( .B1(n6670), .B2(n6952), .A(n6752), .ZN(n6947) );
  AND2_X1 U7905 ( .A1(n11120), .A2(n11121), .ZN(n6952) );
  OAI21_X1 U7906 ( .B1(n11834), .B2(n11833), .A(n11832), .ZN(n11835) );
  NAND2_X1 U7907 ( .A1(n7579), .A2(n6721), .ZN(n6960) );
  INV_X1 U7908 ( .A(n11143), .ZN(n7582) );
  AOI21_X1 U7909 ( .B1(n11213), .B2(n7590), .A(n11211), .ZN(n7589) );
  INV_X1 U7910 ( .A(n7594), .ZN(n7590) );
  OAI21_X1 U7911 ( .B1(n7591), .B2(n6720), .A(n7589), .ZN(n7585) );
  NAND2_X1 U7912 ( .A1(n11213), .A2(n7592), .ZN(n7591) );
  INV_X1 U7913 ( .A(n7595), .ZN(n7592) );
  NAND2_X1 U7914 ( .A1(n7589), .A2(n7587), .ZN(n7586) );
  INV_X1 U7915 ( .A(n7593), .ZN(n7587) );
  NOR2_X1 U7916 ( .A1(n7595), .A2(n6720), .ZN(n7584) );
  NAND2_X1 U7917 ( .A1(n11198), .A2(n6712), .ZN(n7594) );
  INV_X1 U7918 ( .A(n11213), .ZN(n6965) );
  NAND2_X1 U7919 ( .A1(n7570), .A2(n7569), .ZN(n7568) );
  INV_X1 U7920 ( .A(n11247), .ZN(n7569) );
  INV_X1 U7921 ( .A(n11248), .ZN(n7570) );
  OAI21_X1 U7922 ( .B1(n12396), .B2(n12395), .A(n12684), .ZN(n12401) );
  NAND2_X1 U7923 ( .A1(n6926), .A2(n14678), .ZN(n11717) );
  INV_X1 U7924 ( .A(n14195), .ZN(n6926) );
  INV_X1 U7925 ( .A(n9433), .ZN(n7486) );
  NOR2_X1 U7926 ( .A1(n9582), .A2(n7489), .ZN(n7488) );
  INV_X1 U7927 ( .A(n9437), .ZN(n7489) );
  NAND2_X1 U7928 ( .A1(n9273), .A2(n12275), .ZN(n6849) );
  AOI21_X1 U7929 ( .B1(n7562), .B2(n7566), .A(n6730), .ZN(n7560) );
  NOR2_X1 U7930 ( .A1(n7562), .A2(n7564), .ZN(n7561) );
  AOI21_X1 U7931 ( .B1(n7401), .B2(n6673), .A(n7399), .ZN(n7398) );
  NOR2_X1 U7932 ( .A1(n13472), .A2(n13292), .ZN(n7399) );
  NOR2_X1 U7933 ( .A1(n13354), .A2(n7390), .ZN(n7389) );
  NOR2_X1 U7934 ( .A1(n13308), .A2(n7391), .ZN(n7390) );
  INV_X1 U7935 ( .A(n13309), .ZN(n7391) );
  NAND2_X1 U7936 ( .A1(n11858), .A2(n6825), .ZN(n11860) );
  MUX2_X1 U7937 ( .A(n14676), .B(n11713), .S(n13891), .Z(n11883) );
  OR2_X1 U7938 ( .A1(n8275), .A2(n8279), .ZN(n11713) );
  NOR2_X1 U7939 ( .A1(n6647), .A2(n7530), .ZN(n7529) );
  INV_X1 U7940 ( .A(n7534), .ZN(n7530) );
  NAND2_X1 U7941 ( .A1(n10747), .A2(n10746), .ZN(n10748) );
  NAND2_X1 U7942 ( .A1(n7473), .A2(n7054), .ZN(n7053) );
  INV_X1 U7943 ( .A(n8027), .ZN(n7054) );
  INV_X1 U7944 ( .A(n8410), .ZN(n6971) );
  NOR2_X1 U7945 ( .A1(n8036), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U7946 ( .A1(n6798), .A2(n12641), .ZN(n6797) );
  NAND2_X1 U7947 ( .A1(n12412), .A2(n12406), .ZN(n6798) );
  AOI21_X1 U7948 ( .B1(n12408), .B2(n12409), .A(n12407), .ZN(n6799) );
  INV_X1 U7949 ( .A(n12992), .ZN(n8128) );
  NAND2_X1 U7950 ( .A1(n15000), .A2(n10075), .ZN(n10076) );
  NAND2_X1 U7951 ( .A1(n10177), .A2(n6913), .ZN(n10446) );
  OR2_X1 U7952 ( .A1(n10178), .A2(n15451), .ZN(n6913) );
  OR2_X1 U7953 ( .A1(n12861), .A2(n12680), .ZN(n12402) );
  OR2_X1 U7954 ( .A1(n12945), .A2(n12730), .ZN(n12392) );
  OR2_X1 U7955 ( .A1(n12011), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n12022) );
  INV_X1 U7956 ( .A(n12380), .ZN(n7139) );
  INV_X1 U7957 ( .A(n12379), .ZN(n7135) );
  INV_X1 U7958 ( .A(n12375), .ZN(n7136) );
  OR2_X1 U7959 ( .A1(n12733), .A2(n12742), .ZN(n12382) );
  AOI21_X1 U7960 ( .B1(n9719), .B2(n12235), .A(n6803), .ZN(n10215) );
  NAND2_X1 U7961 ( .A1(n9721), .A2(n9720), .ZN(n6803) );
  AND2_X1 U7962 ( .A1(n12300), .A2(n12302), .ZN(n15101) );
  AND3_X1 U7963 ( .A1(n9233), .A2(n9232), .A3(n9231), .ZN(n9502) );
  INV_X1 U7964 ( .A(n12777), .ZN(n12785) );
  NAND2_X1 U7965 ( .A1(n12799), .A2(n12798), .ZN(n7145) );
  NAND2_X1 U7966 ( .A1(n9272), .A2(n9271), .ZN(n9405) );
  AND2_X1 U7967 ( .A1(n7039), .A2(n7038), .ZN(n7037) );
  INV_X1 U7968 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7038) );
  INV_X1 U7969 ( .A(n7195), .ZN(n7194) );
  OAI21_X1 U7970 ( .B1(n8450), .B2(n7196), .A(n8872), .ZN(n7195) );
  INV_X1 U7971 ( .A(n8821), .ZN(n7196) );
  AND2_X1 U7972 ( .A1(n8453), .A2(n7040), .ZN(n7039) );
  INV_X1 U7973 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U7974 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  AND2_X1 U7975 ( .A1(n7491), .A2(n7790), .ZN(n7802) );
  NOR2_X1 U7976 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7006) );
  OR2_X1 U7977 ( .A1(n13051), .A2(n13010), .ZN(n7380) );
  OR2_X1 U7978 ( .A1(n13547), .A2(n11395), .ZN(n13308) );
  AND2_X1 U7979 ( .A1(n13398), .A2(n13303), .ZN(n7396) );
  INV_X1 U7980 ( .A(n13438), .ZN(n7230) );
  NAND2_X1 U7981 ( .A1(n13656), .A2(n7111), .ZN(n7110) );
  OAI21_X1 U7982 ( .B1(n6666), .B2(n7239), .A(n13251), .ZN(n7238) );
  INV_X1 U7983 ( .A(n9286), .ZN(n7226) );
  AND2_X1 U7984 ( .A1(n9288), .A2(n11402), .ZN(n7225) );
  NAND2_X1 U7985 ( .A1(n9283), .A2(n11056), .ZN(n9295) );
  NOR2_X1 U7986 ( .A1(n13793), .A2(n7101), .ZN(n7100) );
  INV_X1 U7987 ( .A(n13746), .ZN(n7101) );
  NAND2_X1 U7988 ( .A1(n8277), .A2(n8276), .ZN(n9054) );
  INV_X1 U7989 ( .A(n8172), .ZN(n8176) );
  NOR2_X1 U7990 ( .A1(n13961), .A2(n13974), .ZN(n7128) );
  NAND2_X1 U7991 ( .A1(n13974), .A2(n13948), .ZN(n7647) );
  AND2_X1 U7992 ( .A1(n14066), .A2(n11911), .ZN(n14090) );
  NAND2_X1 U7993 ( .A1(n14184), .A2(n13938), .ZN(n7547) );
  INV_X1 U7994 ( .A(n13938), .ZN(n7544) );
  INV_X1 U7995 ( .A(n11814), .ZN(n11914) );
  INV_X1 U7996 ( .A(n11913), .ZN(n13940) );
  OR2_X1 U7997 ( .A1(n13909), .A2(n6980), .ZN(n6976) );
  INV_X1 U7998 ( .A(n6981), .ZN(n6980) );
  INV_X1 U7999 ( .A(n11807), .ZN(n13936) );
  AND2_X1 U8000 ( .A1(n11804), .A2(n11801), .ZN(n11915) );
  AOI21_X1 U8001 ( .B1(n10243), .B2(n6663), .A(n7552), .ZN(n7550) );
  NOR2_X1 U8002 ( .A1(n14582), .A2(n13825), .ZN(n7552) );
  NAND2_X1 U8003 ( .A1(n6908), .A2(n9988), .ZN(n10016) );
  AOI21_X1 U8004 ( .B1(n6662), .B2(n7612), .A(n7608), .ZN(n7607) );
  NAND2_X1 U8005 ( .A1(n6896), .A2(n6895), .ZN(n10020) );
  INV_X1 U8006 ( .A(n11927), .ZN(n6895) );
  INV_X1 U8007 ( .A(n9976), .ZN(n6896) );
  NAND3_X1 U8008 ( .A1(n7603), .A2(n7602), .A3(n9628), .ZN(n9983) );
  NAND2_X1 U8009 ( .A1(n8671), .A2(n11725), .ZN(n11916) );
  NAND2_X1 U8010 ( .A1(n11304), .A2(n11303), .ZN(n11327) );
  AND3_X1 U8011 ( .A1(n7722), .A2(n7721), .A3(n7720), .ZN(n7725) );
  INV_X1 U8012 ( .A(n7465), .ZN(n7469) );
  NAND2_X1 U8013 ( .A1(n9589), .A2(n7063), .ZN(n7062) );
  XNOR2_X1 U8014 ( .A(n9176), .B(SI_16_), .ZN(n9173) );
  AND2_X1 U8015 ( .A1(n8031), .A2(n8645), .ZN(n6967) );
  NOR2_X1 U8016 ( .A1(n6971), .A2(n8645), .ZN(n6970) );
  NAND2_X1 U8017 ( .A1(n8346), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6838) );
  XNOR2_X1 U8018 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15496), .ZN(n14430) );
  OAI21_X1 U8019 ( .B1(n14424), .B2(n14425), .A(n6739), .ZN(n7346) );
  OAI21_X1 U8020 ( .B1(n14423), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6728), .ZN(
        n6899) );
  INV_X1 U8021 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15435) );
  OAI22_X1 U8022 ( .A1(n14444), .A2(n14389), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n15486), .ZN(n14390) );
  AOI21_X1 U8023 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14401), .A(n14400), .ZN(
        n14416) );
  NOR2_X1 U8024 ( .A1(n14461), .A2(n14462), .ZN(n14400) );
  NAND2_X1 U8025 ( .A1(n8141), .A2(n10307), .ZN(n10299) );
  OR2_X1 U8026 ( .A1(n7284), .A2(n12153), .ZN(n7283) );
  INV_X1 U8027 ( .A(n12183), .ZN(n7277) );
  OR2_X1 U8028 ( .A1(n7283), .A2(n7292), .ZN(n7274) );
  INV_X1 U8029 ( .A(n7281), .ZN(n7280) );
  OAI21_X1 U8030 ( .B1(n7284), .B2(n7282), .A(n7289), .ZN(n7281) );
  OR2_X1 U8031 ( .A1(n12153), .A2(n7286), .ZN(n7282) );
  AND2_X1 U8032 ( .A1(n8959), .A2(n8750), .ZN(n7244) );
  NAND2_X1 U8033 ( .A1(n12182), .A2(n12183), .ZN(n7273) );
  AND2_X1 U8034 ( .A1(n7254), .A2(n9228), .ZN(n7253) );
  INV_X1 U8035 ( .A(n9235), .ZN(n7254) );
  INV_X1 U8036 ( .A(n12145), .ZN(n7031) );
  AND2_X1 U8037 ( .A1(n10292), .A2(n10619), .ZN(n7271) );
  NAND2_X1 U8038 ( .A1(n7257), .A2(n12752), .ZN(n7256) );
  INV_X1 U8039 ( .A(n12123), .ZN(n7257) );
  OR2_X1 U8040 ( .A1(n9861), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10273) );
  OR2_X1 U8041 ( .A1(n10299), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8226) );
  AND4_X1 U8042 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n10479)
         );
  AND4_X1 U8043 ( .A1(n9244), .A2(n9243), .A3(n9242), .A4(n9241), .ZN(n10198)
         );
  OAI21_X1 U8044 ( .B1(n8744), .B2(n8293), .A(n8540), .ZN(n8294) );
  AND2_X1 U8045 ( .A1(n10133), .A2(n14979), .ZN(n10134) );
  OR2_X1 U8046 ( .A1(n15027), .A2(n15026), .ZN(n7178) );
  NAND2_X1 U8047 ( .A1(n15033), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7177) );
  OR2_X1 U8048 ( .A1(n7168), .A2(n10148), .ZN(n7167) );
  OR2_X1 U8049 ( .A1(n15079), .A2(n10486), .ZN(n7169) );
  XNOR2_X1 U8050 ( .A(n10446), .B(n10435), .ZN(n10179) );
  NAND2_X1 U8051 ( .A1(n12452), .A2(n12451), .ZN(n7181) );
  OR2_X1 U8052 ( .A1(n12475), .A2(n12485), .ZN(n7180) );
  NAND2_X1 U8053 ( .A1(n12507), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7179) );
  OAI21_X1 U8054 ( .B1(n12525), .B2(n7174), .A(n7173), .ZN(n12583) );
  NAND2_X1 U8055 ( .A1(n12542), .A2(n12571), .ZN(n7173) );
  NAND2_X1 U8056 ( .A1(n7171), .A2(n12571), .ZN(n7174) );
  NAND2_X1 U8057 ( .A1(n12102), .A2(n12105), .ZN(n7019) );
  NAND2_X1 U8058 ( .A1(n7021), .A2(n12105), .ZN(n7018) );
  NAND2_X1 U8059 ( .A1(n9766), .A2(n9765), .ZN(n12045) );
  INV_X1 U8060 ( .A(n7016), .ZN(n7015) );
  OAI21_X1 U8061 ( .B1(n6692), .B2(n7017), .A(n12754), .ZN(n7016) );
  INV_X1 U8062 ( .A(n12093), .ZN(n7017) );
  AND2_X1 U8063 ( .A1(n6687), .A2(n12726), .ZN(n12743) );
  NAND2_X1 U8064 ( .A1(n7140), .A2(n12373), .ZN(n12757) );
  INV_X1 U8065 ( .A(n12755), .ZN(n7140) );
  NAND2_X1 U8066 ( .A1(n12774), .A2(n6692), .ZN(n12763) );
  OR2_X1 U8067 ( .A1(n12791), .A2(n12091), .ZN(n12767) );
  NAND2_X1 U8068 ( .A1(n12090), .A2(n7500), .ZN(n12774) );
  NOR2_X1 U8069 ( .A1(n12777), .A2(n7501), .ZN(n7500) );
  INV_X1 U8070 ( .A(n12089), .ZN(n7501) );
  AND2_X1 U8071 ( .A1(n12767), .A2(n12364), .ZN(n12777) );
  AND4_X1 U8072 ( .A1(n8231), .A2(n8230), .A3(n8229), .A4(n8228), .ZN(n12836)
         );
  INV_X1 U8073 ( .A(n11973), .ZN(n7153) );
  AOI21_X1 U8074 ( .B1(n7157), .B2(n12321), .A(n7155), .ZN(n7154) );
  INV_X1 U8075 ( .A(n7157), .ZN(n7156) );
  INV_X1 U8076 ( .A(n12328), .ZN(n7155) );
  AND2_X1 U8077 ( .A1(n10759), .A2(n10758), .ZN(n10760) );
  NOR2_X1 U8078 ( .A1(n10730), .A2(n7158), .ZN(n7157) );
  INV_X1 U8079 ( .A(n10735), .ZN(n7158) );
  NAND2_X1 U8080 ( .A1(n10537), .A2(n12321), .ZN(n10729) );
  OR2_X1 U8081 ( .A1(n9424), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9602) );
  INV_X1 U8082 ( .A(n10200), .ZN(n7497) );
  INV_X1 U8083 ( .A(n10199), .ZN(n7496) );
  NAND2_X1 U8084 ( .A1(n10200), .A2(n7498), .ZN(n15103) );
  AND2_X1 U8085 ( .A1(n10201), .A2(n10199), .ZN(n7498) );
  INV_X1 U8086 ( .A(n15101), .ZN(n10201) );
  OAI21_X1 U8087 ( .B1(n9361), .B2(n7494), .A(n7002), .ZN(n9504) );
  INV_X1 U8088 ( .A(n9363), .ZN(n7494) );
  NOR2_X1 U8089 ( .A1(n6691), .A2(n7003), .ZN(n7002) );
  NAND2_X1 U8090 ( .A1(n6780), .A2(n9362), .ZN(n15116) );
  AND3_X1 U8091 ( .A1(n9043), .A2(n9042), .A3(n9041), .ZN(n15120) );
  INV_X1 U8092 ( .A(n12697), .ZN(n15146) );
  NAND2_X1 U8093 ( .A1(n10877), .A2(n10876), .ZN(n12902) );
  NAND2_X1 U8094 ( .A1(n10669), .A2(n10668), .ZN(n12906) );
  OR2_X1 U8095 ( .A1(n10667), .A2(n11984), .ZN(n10669) );
  AND2_X1 U8096 ( .A1(n8506), .A2(n8498), .ZN(n8713) );
  AND2_X1 U8097 ( .A1(n8520), .A2(n12409), .ZN(n15149) );
  OAI21_X1 U8098 ( .B1(n12218), .B2(n12217), .A(n12219), .ZN(n12232) );
  NAND2_X1 U8099 ( .A1(n8124), .A2(n12981), .ZN(n7001) );
  INV_X1 U8100 ( .A(n8106), .ZN(n12426) );
  NOR2_X1 U8101 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7685) );
  AND2_X1 U8102 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  NOR2_X1 U8103 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7688) );
  NOR2_X1 U8104 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7687) );
  NAND2_X1 U8105 ( .A1(n9647), .A2(n9646), .ZN(n9960) );
  OR2_X1 U8106 ( .A1(n8493), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8107) );
  AND2_X1 U8107 ( .A1(n7037), .A2(n7036), .ZN(n7035) );
  INV_X1 U8108 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U8109 ( .A1(n8448), .A2(n8447), .ZN(n8451) );
  NAND2_X1 U8110 ( .A1(n8451), .A2(n8450), .ZN(n8822) );
  INV_X1 U8111 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U8112 ( .A1(n8454), .A2(n7039), .ZN(n8824) );
  NAND2_X1 U8113 ( .A1(n8020), .A2(n10779), .ZN(n7201) );
  AND2_X1 U8114 ( .A1(n7943), .A2(n8023), .ZN(n12460) );
  AND2_X1 U8115 ( .A1(n7932), .A2(n7913), .ZN(n7914) );
  INV_X1 U8116 ( .A(n7911), .ZN(n7190) );
  OR2_X1 U8117 ( .A1(n7851), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7908) );
  AND2_X1 U8118 ( .A1(n7911), .A2(n7882), .ZN(n7883) );
  NAND2_X1 U8119 ( .A1(n7881), .A2(n7880), .ZN(n7884) );
  NAND2_X1 U8120 ( .A1(n7884), .A2(n7883), .ZN(n7912) );
  NAND2_X1 U8121 ( .A1(n7848), .A2(n7847), .ZN(n7881) );
  NAND2_X1 U8122 ( .A1(n7926), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U8123 ( .A1(n7869), .A2(n7841), .ZN(n7890) );
  AND2_X1 U8124 ( .A1(n7843), .A2(n7842), .ZN(n7889) );
  AND2_X1 U8125 ( .A1(n7208), .A2(n7889), .ZN(n7207) );
  NAND2_X1 U8126 ( .A1(n7866), .A2(n7841), .ZN(n7208) );
  OR2_X1 U8127 ( .A1(n7867), .A2(n7866), .ZN(n7869) );
  NAND2_X1 U8128 ( .A1(n7781), .A2(n7780), .ZN(n7837) );
  NAND2_X1 U8129 ( .A1(n6829), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7792) );
  AND2_X1 U8130 ( .A1(n7773), .A2(n7772), .ZN(n7788) );
  AND2_X1 U8131 ( .A1(n9130), .A2(n8923), .ZN(n6929) );
  INV_X1 U8132 ( .A(n7380), .ZN(n6937) );
  NAND2_X1 U8133 ( .A1(n8979), .A2(n8900), .ZN(n6930) );
  NAND2_X1 U8134 ( .A1(n9266), .A2(n9265), .ZN(n9376) );
  NAND2_X1 U8135 ( .A1(n11013), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n11187) );
  INV_X1 U8136 ( .A(n11173), .ZN(n11013) );
  OR2_X1 U8137 ( .A1(n11187), .A2(n13105), .ZN(n11189) );
  NAND2_X1 U8138 ( .A1(n13012), .A2(n13011), .ZN(n7378) );
  NAND2_X1 U8139 ( .A1(n9020), .A2(n9130), .ZN(n9021) );
  NOR2_X1 U8140 ( .A1(n7352), .A2(n7353), .ZN(n13132) );
  OAI21_X1 U8141 ( .B1(n13024), .B2(n7355), .A(n6737), .ZN(n7353) );
  NOR2_X1 U8142 ( .A1(n11452), .A2(n11449), .ZN(n7479) );
  INV_X1 U8143 ( .A(n7481), .ZN(n7480) );
  NOR2_X1 U8144 ( .A1(n11386), .A2(n11385), .ZN(n11447) );
  CLKBUF_X1 U8145 ( .A(n11016), .Z(n11371) );
  CLKBUF_X1 U8146 ( .A(n11337), .Z(n6847) );
  NAND2_X1 U8147 ( .A1(n8335), .A2(n13674), .ZN(n8786) );
  NAND2_X1 U8148 ( .A1(n8335), .A2(n8333), .ZN(n11337) );
  NOR2_X1 U8149 ( .A1(n8435), .A2(n8434), .ZN(n8433) );
  OR2_X1 U8150 ( .A1(n8433), .A2(n6989), .ZN(n6988) );
  AND2_X1 U8151 ( .A1(n8901), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6989) );
  AND2_X1 U8152 ( .A1(n6988), .A2(n6987), .ZN(n14782) );
  INV_X1 U8153 ( .A(n14783), .ZN(n6987) );
  NOR2_X1 U8154 ( .A1(n8879), .A2(n6997), .ZN(n14797) );
  AND2_X1 U8155 ( .A1(n9121), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6997) );
  NOR2_X1 U8156 ( .A1(n14797), .A2(n14796), .ZN(n14795) );
  OR2_X1 U8157 ( .A1(n13206), .A2(n6994), .ZN(n6993) );
  AND2_X1 U8158 ( .A1(n13207), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8159 ( .A1(n6993), .A2(n6992), .ZN(n6991) );
  INV_X1 U8160 ( .A(n14849), .ZN(n6992) );
  NAND2_X1 U8161 ( .A1(n13273), .A2(n7241), .ZN(n7049) );
  NAND2_X1 U8162 ( .A1(n7242), .A2(n13273), .ZN(n7048) );
  NOR2_X1 U8163 ( .A1(n13398), .A2(n7243), .ZN(n7242) );
  INV_X1 U8164 ( .A(n13269), .ZN(n7243) );
  NAND2_X1 U8165 ( .A1(n7117), .A2(n7116), .ZN(n13409) );
  NAND2_X1 U8166 ( .A1(n6836), .A2(n7396), .ZN(n13389) );
  AOI21_X1 U8167 ( .B1(n13257), .B2(n7234), .A(n7233), .ZN(n7232) );
  NOR2_X1 U8168 ( .A1(n13652), .A2(n13259), .ZN(n7233) );
  NOR2_X1 U8169 ( .A1(n13256), .A2(n13260), .ZN(n7234) );
  NAND2_X1 U8170 ( .A1(n13257), .A2(n7236), .ZN(n7235) );
  INV_X1 U8171 ( .A(n13260), .ZN(n7236) );
  AND2_X1 U8172 ( .A1(n13293), .A2(n13432), .ZN(n13452) );
  NAND2_X1 U8173 ( .A1(n7406), .A2(n6690), .ZN(n7405) );
  INV_X1 U8174 ( .A(n6916), .ZN(n7406) );
  NAND2_X1 U8175 ( .A1(n10695), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11159) );
  INV_X1 U8176 ( .A(n10696), .ZN(n10695) );
  NAND2_X1 U8177 ( .A1(n10895), .A2(n6666), .ZN(n13250) );
  NAND2_X1 U8178 ( .A1(n9909), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10633) );
  NOR2_X1 U8179 ( .A1(n11411), .A2(n7415), .ZN(n7414) );
  INV_X1 U8180 ( .A(n10367), .ZN(n7415) );
  NAND2_X1 U8181 ( .A1(n7106), .A2(n7105), .ZN(n10375) );
  INV_X1 U8182 ( .A(n10360), .ZN(n7106) );
  AOI21_X1 U8183 ( .B1(n11409), .B2(n7217), .A(n6722), .ZN(n7216) );
  INV_X1 U8184 ( .A(n9686), .ZN(n7217) );
  INV_X1 U8185 ( .A(n11409), .ZN(n7218) );
  OR2_X1 U8186 ( .A1(n9139), .A2(n9138), .ZN(n9384) );
  NAND2_X1 U8187 ( .A1(n9540), .A2(n9539), .ZN(n9542) );
  OR2_X1 U8188 ( .A1(n11363), .A2(n8724), .ZN(n8725) );
  NAND2_X1 U8189 ( .A1(n13334), .A2(n6689), .ZN(n13538) );
  AND2_X1 U8190 ( .A1(n13329), .A2(n13328), .ZN(n13537) );
  NAND2_X1 U8191 ( .A1(n11171), .A2(n11170), .ZN(n13588) );
  NAND3_X1 U8192 ( .A1(n7648), .A2(n7385), .A3(n8317), .ZN(n8323) );
  OR2_X1 U8193 ( .A1(n8233), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9070) );
  NOR2_X1 U8194 ( .A1(n9070), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U8195 ( .A1(n6953), .A2(n6955), .ZN(n7416) );
  AOI21_X1 U8196 ( .B1(n6671), .B2(n7424), .A(n6742), .ZN(n7421) );
  NOR2_X1 U8197 ( .A1(n7437), .A2(n7099), .ZN(n7096) );
  INV_X1 U8198 ( .A(n7438), .ZN(n7437) );
  INV_X1 U8199 ( .A(n11543), .ZN(n7436) );
  NAND2_X1 U8200 ( .A1(n7096), .A2(n7094), .ZN(n7093) );
  INV_X1 U8201 ( .A(n7100), .ZN(n7094) );
  NAND2_X1 U8202 ( .A1(n14561), .A2(n6887), .ZN(n11485) );
  OR2_X1 U8203 ( .A1(n11479), .A2(n11478), .ZN(n6887) );
  AND2_X1 U8204 ( .A1(n13695), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U8205 ( .A1(n7429), .A2(n11594), .ZN(n7428) );
  INV_X1 U8206 ( .A(n13784), .ZN(n7429) );
  INV_X1 U8207 ( .A(n11594), .ZN(n7430) );
  AOI21_X1 U8208 ( .B1(n11680), .B2(n14195), .A(n8213), .ZN(n8217) );
  NAND2_X1 U8209 ( .A1(n8212), .A2(n8211), .ZN(n8213) );
  NAND2_X1 U8210 ( .A1(n10521), .A2(n14678), .ZN(n8212) );
  AOI21_X1 U8211 ( .B1(n13712), .B2(n11543), .A(n7439), .ZN(n7438) );
  INV_X1 U8212 ( .A(n13763), .ZN(n7439) );
  INV_X1 U8213 ( .A(n10866), .ZN(n7445) );
  NAND2_X1 U8214 ( .A1(n8611), .A2(n7431), .ZN(n9057) );
  NAND2_X1 U8215 ( .A1(n11680), .A2(n14196), .ZN(n7431) );
  XNOR2_X1 U8216 ( .A(n7091), .B(n9054), .ZN(n9059) );
  AOI22_X1 U8217 ( .A1(n14196), .A2(n10521), .B1(n11699), .B2(n11730), .ZN(
        n7091) );
  NAND2_X1 U8218 ( .A1(n13705), .A2(n7083), .ZN(n7073) );
  NAND2_X1 U8219 ( .A1(n7079), .A2(n7081), .ZN(n7077) );
  INV_X1 U8220 ( .A(n7078), .ZN(n7071) );
  AND3_X1 U8221 ( .A1(n11943), .A2(n13965), .A3(n7059), .ZN(n11939) );
  OAI211_X1 U8222 ( .C1(n13901), .C2(n13900), .A(n11900), .B(n6807), .ZN(
        n11944) );
  NAND2_X1 U8223 ( .A1(n13901), .A2(n6808), .ZN(n6807) );
  AOI21_X1 U8224 ( .B1(n7309), .B2(n7311), .A(n6743), .ZN(n7308) );
  AND4_X1 U8225 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n13912) );
  OR2_X1 U8226 ( .A1(n11704), .A2(n13833), .ZN(n8177) );
  INV_X1 U8227 ( .A(n6644), .ZN(n11888) );
  NOR2_X1 U8228 ( .A1(n13965), .A2(n7646), .ZN(n7645) );
  INV_X1 U8229 ( .A(n13931), .ZN(n7646) );
  INV_X1 U8230 ( .A(n7633), .ZN(n7632) );
  AOI21_X1 U8231 ( .B1(n14034), .B2(n13925), .A(n13926), .ZN(n7633) );
  AND2_X1 U8232 ( .A1(n7537), .A2(n14058), .ZN(n7534) );
  OR2_X1 U8233 ( .A1(n7535), .A2(n7532), .ZN(n7531) );
  INV_X1 U8234 ( .A(n7537), .ZN(n7532) );
  AND2_X1 U8235 ( .A1(n13947), .A2(n6706), .ZN(n7535) );
  NAND2_X1 U8236 ( .A1(n14123), .A2(n7541), .ZN(n14108) );
  AOI21_X1 U8237 ( .B1(n7623), .B2(n7621), .A(n6672), .ZN(n7620) );
  INV_X1 U8238 ( .A(n13913), .ZN(n7621) );
  NAND2_X1 U8239 ( .A1(n6976), .A2(n6974), .ZN(n7622) );
  NOR2_X1 U8240 ( .A1(n7624), .A2(n6975), .ZN(n6974) );
  INV_X1 U8241 ( .A(n6978), .ZN(n6975) );
  NAND2_X1 U8242 ( .A1(n6976), .A2(n6978), .ZN(n14155) );
  OR2_X1 U8243 ( .A1(n14169), .A2(n14184), .ZN(n14167) );
  NAND2_X1 U8244 ( .A1(n10783), .A2(n10782), .ZN(n11798) );
  AND2_X1 U8245 ( .A1(n7618), .A2(n14502), .ZN(n7617) );
  NAND2_X1 U8246 ( .A1(n11928), .A2(n10824), .ZN(n7618) );
  AND4_X1 U8247 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n13773) );
  OR2_X1 U8248 ( .A1(n11904), .A2(n8636), .ZN(n14141) );
  AOI21_X1 U8249 ( .B1(n10243), .B2(n7599), .A(n6725), .ZN(n7598) );
  INV_X1 U8250 ( .A(n10017), .ZN(n7599) );
  NAND2_X1 U8251 ( .A1(n7551), .A2(n7600), .ZN(n10258) );
  INV_X1 U8252 ( .A(n10021), .ZN(n7551) );
  INV_X1 U8253 ( .A(n7522), .ZN(n7521) );
  NAND2_X1 U8254 ( .A1(n8861), .A2(n9053), .ZN(n8936) );
  OR2_X1 U8255 ( .A1(n14193), .A2(n8670), .ZN(n14202) );
  INV_X1 U8256 ( .A(n13891), .ZN(n14677) );
  OR2_X1 U8257 ( .A1(n14195), .A2(n14678), .ZN(n8281) );
  OR2_X1 U8258 ( .A1(n9515), .A2(n11612), .ZN(n9518) );
  OR2_X1 U8259 ( .A1(n11612), .A2(n8614), .ZN(n8617) );
  AND2_X1 U8260 ( .A1(n7973), .A2(n7976), .ZN(n7630) );
  AND2_X1 U8261 ( .A1(n7973), .A2(n7976), .ZN(n7068) );
  INV_X1 U8262 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7976) );
  OAI21_X1 U8263 ( .B1(n7976), .B2(n7973), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7066) );
  NAND2_X1 U8264 ( .A1(n9096), .A2(n6723), .ZN(n8182) );
  INV_X1 U8265 ( .A(n7062), .ZN(n7061) );
  AND2_X1 U8266 ( .A1(n7716), .A2(n7717), .ZN(n7447) );
  INV_X1 U8267 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7717) );
  INV_X1 U8268 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8184) );
  OAI21_X1 U8269 ( .B1(n8032), .B2(n7475), .A(n7473), .ZN(n8799) );
  INV_X1 U8270 ( .A(n7462), .ZN(n7461) );
  OAI21_X1 U8271 ( .B1(n7923), .B2(n7463), .A(n7957), .ZN(n7462) );
  INV_X1 U8272 ( .A(n7953), .ZN(n7463) );
  NAND2_X1 U8273 ( .A1(n7924), .A2(n7923), .ZN(n7954) );
  NAND2_X1 U8274 ( .A1(n7448), .A2(SI_1_), .ZN(n7748) );
  OAI21_X1 U8275 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14396), .A(n14395), .ZN(
        n14418) );
  OAI21_X1 U8276 ( .B1(n14635), .B2(n14636), .A(n6898), .ZN(n6897) );
  INV_X1 U8277 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6898) );
  OR2_X1 U8278 ( .A1(n10269), .A2(n7264), .ZN(n7259) );
  AND2_X1 U8279 ( .A1(n7260), .A2(n10505), .ZN(n6848) );
  NAND2_X1 U8280 ( .A1(n7262), .A2(n7264), .ZN(n7260) );
  AND3_X1 U8281 ( .A1(n8818), .A2(n8817), .A3(n8816), .ZN(n12741) );
  NOR2_X1 U8282 ( .A1(n12193), .A2(n12194), .ZN(n12192) );
  NAND2_X1 U8283 ( .A1(n11983), .A2(n11982), .ZN(n12753) );
  AND4_X1 U8284 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10922) );
  AND4_X1 U8285 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n12779) );
  INV_X1 U8286 ( .A(n12418), .ZN(n12267) );
  AND3_X1 U8287 ( .A1(n6869), .A2(n7212), .A3(n12418), .ZN(n12268) );
  INV_X1 U8288 ( .A(n12741), .ZN(n12764) );
  XNOR2_X1 U8289 ( .A(n7181), .B(n12477), .ZN(n12453) );
  NAND2_X1 U8290 ( .A1(n12480), .A2(n12486), .ZN(n12502) );
  NOR2_X1 U8291 ( .A1(n12583), .A2(n7175), .ZN(n12566) );
  AND2_X1 U8292 ( .A1(n12565), .A2(n7170), .ZN(n7175) );
  NOR2_X1 U8293 ( .A1(n12571), .A2(n12542), .ZN(n7170) );
  NAND2_X1 U8294 ( .A1(n12566), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12587) );
  XNOR2_X1 U8295 ( .A(n6789), .B(n12606), .ZN(n12581) );
  NAND2_X1 U8296 ( .A1(n12655), .A2(n6835), .ZN(n12857) );
  OR2_X1 U8297 ( .A1(n12656), .A2(n15154), .ZN(n6835) );
  NAND2_X1 U8298 ( .A1(n12625), .A2(n14537), .ZN(n7026) );
  OAI21_X1 U8299 ( .B1(n12114), .B2(n15154), .A(n12113), .ZN(n12626) );
  NOR2_X1 U8300 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  OAI21_X1 U8301 ( .B1(n12626), .B2(n7160), .A(n7163), .ZN(n6885) );
  OR2_X1 U8302 ( .A1(n15217), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7163) );
  OR2_X1 U8303 ( .A1(n14537), .A2(n15215), .ZN(n7160) );
  INV_X1 U8304 ( .A(n12626), .ZN(n7162) );
  XNOR2_X1 U8305 ( .A(n12229), .B(n7164), .ZN(n12625) );
  INV_X1 U8306 ( .A(n12266), .ZN(n7164) );
  INV_X1 U8307 ( .A(n11972), .ZN(n12627) );
  NOR2_X1 U8308 ( .A1(n12857), .A2(n6834), .ZN(n12930) );
  AND2_X1 U8309 ( .A1(n12858), .A2(n15206), .ZN(n6834) );
  NAND2_X1 U8310 ( .A1(n11979), .A2(n11978), .ZN(n12963) );
  NAND2_X1 U8311 ( .A1(n10501), .A2(n10500), .ZN(n12977) );
  NAND2_X1 U8312 ( .A1(n8125), .A2(n8124), .ZN(n12982) );
  NOR2_X1 U8313 ( .A1(n8125), .A2(n6801), .ZN(n6800) );
  NOR2_X1 U8314 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6801) );
  XNOR2_X1 U8315 ( .A(n8108), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12429) );
  NAND2_X1 U8316 ( .A1(n8107), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8108) );
  INV_X1 U8317 ( .A(n7376), .ZN(n7370) );
  INV_X1 U8318 ( .A(n7372), .ZN(n7371) );
  OAI21_X1 U8319 ( .B1(n7376), .B2(n7374), .A(n7373), .ZN(n7372) );
  AOI21_X1 U8320 ( .B1(n13070), .B2(n7375), .A(n14552), .ZN(n7373) );
  OR2_X1 U8321 ( .A1(n13070), .A2(n7375), .ZN(n7374) );
  NAND2_X1 U8322 ( .A1(n13132), .A2(n13131), .ZN(n13130) );
  NAND2_X1 U8323 ( .A1(n11011), .A2(n11010), .ZN(n13442) );
  NAND2_X1 U8324 ( .A1(n6932), .A2(n7366), .ZN(n6931) );
  NAND2_X1 U8325 ( .A1(n7362), .A2(n7361), .ZN(n6932) );
  NAND2_X1 U8326 ( .A1(n6930), .A2(n8923), .ZN(n9016) );
  OR2_X1 U8327 ( .A1(n11613), .A2(n11236), .ZN(n11239) );
  NAND2_X1 U8328 ( .A1(n11186), .A2(n11185), .ZN(n13457) );
  NAND2_X1 U8329 ( .A1(n11153), .A2(n11152), .ZN(n13289) );
  NAND2_X1 U8330 ( .A1(n10693), .A2(n10692), .ZN(n11133) );
  NOR2_X1 U8331 ( .A1(n14810), .A2(n6996), .ZN(n9653) );
  AND2_X1 U8332 ( .A1(n14815), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6996) );
  NOR2_X1 U8333 ( .A1(n13183), .A2(n13182), .ZN(n13206) );
  NAND2_X1 U8334 ( .A1(n11456), .A2(n8369), .ZN(n13515) );
  NAND2_X1 U8335 ( .A1(n11360), .A2(n11359), .ZN(n13233) );
  INV_X1 U8336 ( .A(n13533), .ZN(n7119) );
  AND2_X1 U8337 ( .A1(n7045), .A2(n6764), .ZN(n7118) );
  NAND2_X1 U8338 ( .A1(n14560), .A2(n6812), .ZN(n14561) );
  AND2_X1 U8339 ( .A1(n14562), .A2(n14559), .ZN(n6812) );
  INV_X1 U8340 ( .A(n14337), .ZN(n13700) );
  INV_X1 U8341 ( .A(n14342), .ZN(n14100) );
  NAND2_X1 U8342 ( .A1(n7446), .A2(n7444), .ZN(n11472) );
  INV_X1 U8343 ( .A(n14181), .ZN(n14300) );
  INV_X1 U8344 ( .A(n10659), .ZN(n7419) );
  NAND2_X1 U8345 ( .A1(n14236), .A2(n13798), .ZN(n6810) );
  INV_X1 U8346 ( .A(n14574), .ZN(n14567) );
  INV_X1 U8347 ( .A(n13773), .ZN(n14578) );
  AND2_X1 U8348 ( .A1(n14061), .A2(n13925), .ZN(n14033) );
  AND2_X1 U8349 ( .A1(n7516), .A2(n7514), .ZN(n14319) );
  AND2_X1 U8350 ( .A1(n11917), .A2(n11901), .ZN(n11723) );
  MUX2_X1 U8351 ( .A(n11719), .B(n11718), .S(n11737), .Z(n11724) );
  NAND2_X1 U8352 ( .A1(n11752), .A2(n7325), .ZN(n7326) );
  OAI21_X1 U8353 ( .B1(n11050), .B2(n11049), .A(n11048), .ZN(n11059) );
  NAND2_X1 U8354 ( .A1(n11762), .A2(n11764), .ZN(n7315) );
  NAND2_X1 U8355 ( .A1(n12279), .A2(n12397), .ZN(n6892) );
  NAND2_X1 U8356 ( .A1(n12278), .A2(n12409), .ZN(n6893) );
  INV_X1 U8357 ( .A(n6763), .ZN(n7576) );
  AOI21_X1 U8358 ( .B1(n11079), .B2(n11078), .A(n11076), .ZN(n11077) );
  NAND2_X1 U8359 ( .A1(n7301), .A2(n7299), .ZN(n7298) );
  NAND2_X1 U8360 ( .A1(n11799), .A2(n7303), .ZN(n7301) );
  NAND2_X1 U8361 ( .A1(n11793), .A2(n11794), .ZN(n7299) );
  NAND2_X1 U8362 ( .A1(n7340), .A2(n7341), .ZN(n11796) );
  NAND2_X1 U8363 ( .A1(n11788), .A2(n11790), .ZN(n7341) );
  INV_X1 U8364 ( .A(n6891), .ZN(n6890) );
  OAI21_X1 U8365 ( .B1(n12409), .B2(n12291), .A(n12289), .ZN(n6891) );
  NAND2_X1 U8366 ( .A1(n11091), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U8367 ( .A1(n11097), .A2(n6678), .ZN(n7572) );
  NAND2_X1 U8368 ( .A1(n11800), .A2(n7302), .ZN(n7300) );
  NAND2_X1 U8369 ( .A1(n12298), .A2(n6889), .ZN(n12294) );
  AND2_X1 U8370 ( .A1(n12297), .A2(n12292), .ZN(n6889) );
  AOI21_X1 U8371 ( .B1(n7654), .B2(n6674), .A(n6741), .ZN(n7319) );
  NAND2_X1 U8372 ( .A1(n7556), .A2(n7558), .ZN(n11122) );
  NAND2_X1 U8373 ( .A1(n6694), .A2(n7559), .ZN(n7558) );
  NAND2_X1 U8374 ( .A1(n11111), .A2(n11110), .ZN(n7557) );
  NAND2_X1 U8375 ( .A1(n6951), .A2(n6950), .ZN(n6949) );
  INV_X1 U8376 ( .A(n11121), .ZN(n6951) );
  INV_X1 U8377 ( .A(n11128), .ZN(n7578) );
  INV_X1 U8378 ( .A(n11836), .ZN(n7339) );
  AOI21_X1 U8379 ( .B1(n6823), .B2(n12255), .A(n6821), .ZN(n12330) );
  NAND2_X1 U8380 ( .A1(n12254), .A2(n6822), .ZN(n6821) );
  NAND2_X1 U8381 ( .A1(n12323), .A2(n12322), .ZN(n6823) );
  INV_X1 U8382 ( .A(n12327), .ZN(n6822) );
  INV_X1 U8383 ( .A(n11840), .ZN(n7334) );
  INV_X1 U8384 ( .A(n11841), .ZN(n7338) );
  NAND2_X1 U8385 ( .A1(n7339), .A2(n11839), .ZN(n7336) );
  INV_X1 U8386 ( .A(n7335), .ZN(n7333) );
  OR2_X1 U8387 ( .A1(n7335), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U8388 ( .A1(n7337), .A2(n7336), .ZN(n7332) );
  NOR2_X1 U8389 ( .A1(n7339), .A2(n11839), .ZN(n7337) );
  OAI22_X1 U8390 ( .A1(n6959), .A2(n6958), .B1(n11165), .B2(n6686), .ZN(n11182) );
  NOR2_X1 U8391 ( .A1(n11198), .A2(n6712), .ZN(n7595) );
  NAND2_X1 U8392 ( .A1(n6883), .A2(n6882), .ZN(n11848) );
  INV_X1 U8393 ( .A(n11848), .ZN(n11853) );
  NAND2_X1 U8394 ( .A1(n6964), .A2(n11214), .ZN(n11230) );
  OAI21_X1 U8395 ( .B1(n11196), .B2(n7586), .A(n7585), .ZN(n11212) );
  AND2_X1 U8396 ( .A1(n11247), .A2(n11248), .ZN(n7571) );
  NOR2_X1 U8397 ( .A1(n7565), .A2(n11265), .ZN(n7564) );
  INV_X1 U8398 ( .A(n7568), .ZN(n7565) );
  OAI21_X1 U8399 ( .B1(n7566), .B2(n7568), .A(n11268), .ZN(n7563) );
  AND2_X1 U8400 ( .A1(n11315), .A2(n6640), .ZN(n6963) );
  INV_X1 U8401 ( .A(n8798), .ZN(n7472) );
  INV_X1 U8402 ( .A(n12101), .ZN(n7023) );
  NOR2_X1 U8403 ( .A1(n7360), .A2(n13095), .ZN(n7359) );
  INV_X1 U8404 ( .A(n13080), .ZN(n7360) );
  INV_X1 U8405 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7657) );
  AND2_X1 U8406 ( .A1(n14355), .A2(n14590), .ZN(n11807) );
  INV_X1 U8407 ( .A(n7601), .ZN(n7604) );
  NAND2_X1 U8408 ( .A1(n7465), .A2(n10991), .ZN(n7464) );
  NAND2_X1 U8409 ( .A1(n10991), .A2(n7467), .ZN(n7466) );
  NAND2_X1 U8410 ( .A1(n10933), .A2(n7470), .ZN(n7465) );
  INV_X1 U8411 ( .A(n10992), .ZN(n7470) );
  AND2_X1 U8412 ( .A1(n7485), .A2(n9581), .ZN(n7484) );
  NAND2_X1 U8413 ( .A1(n7488), .A2(n7486), .ZN(n7485) );
  INV_X1 U8414 ( .A(n7488), .ZN(n7487) );
  NAND2_X1 U8415 ( .A1(n9086), .A2(SI_15_), .ZN(n9089) );
  INV_X1 U8416 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14384) );
  NAND2_X1 U8417 ( .A1(n12132), .A2(n12680), .ZN(n7290) );
  AND2_X1 U8418 ( .A1(n9854), .A2(n7030), .ZN(n7029) );
  INV_X1 U8419 ( .A(n9857), .ZN(n7030) );
  INV_X1 U8420 ( .A(n8743), .ZN(n7033) );
  OAI21_X1 U8421 ( .B1(n9708), .B2(n6850), .A(n6849), .ZN(n8743) );
  NAND2_X1 U8422 ( .A1(n9413), .A2(n9364), .ZN(n6850) );
  NAND2_X1 U8423 ( .A1(n12552), .A2(n12553), .ZN(n12575) );
  NAND2_X1 U8424 ( .A1(n8140), .A2(n8139), .ZN(n10297) );
  INV_X1 U8425 ( .A(n10273), .ZN(n8140) );
  NAND2_X1 U8426 ( .A1(n9363), .A2(n7493), .ZN(n7492) );
  INV_X1 U8427 ( .A(n9360), .ZN(n7493) );
  AND2_X1 U8428 ( .A1(n12284), .A2(n12291), .ZN(n15113) );
  NOR2_X1 U8429 ( .A1(n12785), .A2(n7144), .ZN(n7143) );
  INV_X1 U8430 ( .A(n12360), .ZN(n7144) );
  INV_X1 U8431 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n15334) );
  INV_X1 U8432 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n15477) );
  NAND2_X1 U8433 ( .A1(n8105), .A2(n7509), .ZN(n7508) );
  AND2_X1 U8434 ( .A1(n6709), .A2(n7503), .ZN(n7502) );
  AND2_X1 U8435 ( .A1(n7689), .A2(n7690), .ZN(n7503) );
  INV_X1 U8436 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7941) );
  INV_X1 U8437 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7785) );
  INV_X1 U8438 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7679) );
  INV_X1 U8439 ( .A(n7841), .ZN(n7205) );
  NAND2_X1 U8440 ( .A1(n7907), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U8441 ( .A1(n6677), .A2(n6772), .ZN(n7356) );
  INV_X1 U8442 ( .A(n13040), .ZN(n7365) );
  NAND2_X1 U8443 ( .A1(n13080), .A2(n7358), .ZN(n7357) );
  INV_X1 U8444 ( .A(n7366), .ZN(n7358) );
  NAND2_X1 U8445 ( .A1(n7359), .A2(n7364), .ZN(n7355) );
  NAND2_X1 U8446 ( .A1(n11291), .A2(n11290), .ZN(n11384) );
  OR2_X1 U8447 ( .A1(n11289), .A2(n11288), .ZN(n11290) );
  NAND2_X1 U8448 ( .A1(n11287), .A2(n11286), .ZN(n11291) );
  OR2_X1 U8449 ( .A1(n13336), .A2(n13315), .ZN(n13311) );
  INV_X1 U8450 ( .A(n13305), .ZN(n7395) );
  INV_X1 U8451 ( .A(n7402), .ZN(n7401) );
  OAI21_X1 U8452 ( .B1(n7403), .B2(n6690), .A(n13290), .ZN(n7402) );
  AOI21_X1 U8453 ( .B1(n7389), .B2(n7391), .A(n6715), .ZN(n7387) );
  INV_X1 U8454 ( .A(n7117), .ZN(n13421) );
  AND2_X1 U8455 ( .A1(n9114), .A2(n11427), .ZN(n11024) );
  INV_X1 U8456 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6855) );
  INV_X1 U8457 ( .A(n11650), .ZN(n7424) );
  OR2_X1 U8458 ( .A1(n13755), .A2(n7089), .ZN(n7088) );
  NAND2_X1 U8459 ( .A1(n6702), .A2(n7089), .ZN(n7086) );
  NAND2_X1 U8460 ( .A1(n9056), .A2(n7084), .ZN(n7083) );
  INV_X1 U8461 ( .A(n9060), .ZN(n7084) );
  NOR2_X1 U8462 ( .A1(n13983), .A2(n11937), .ZN(n7059) );
  NOR2_X1 U8463 ( .A1(n7635), .A2(n13926), .ZN(n7634) );
  INV_X1 U8464 ( .A(n7636), .ZN(n7635) );
  NOR2_X1 U8465 ( .A1(n14170), .A2(n7122), .ZN(n14097) );
  NAND2_X1 U8466 ( .A1(n14347), .A2(n7123), .ZN(n7122) );
  NOR2_X1 U8467 ( .A1(n7124), .A2(n11912), .ZN(n7123) );
  OR2_X1 U8468 ( .A1(n14133), .A2(n13823), .ZN(n13917) );
  INV_X1 U8469 ( .A(n13914), .ZN(n7625) );
  NAND2_X1 U8470 ( .A1(n14147), .A2(n14292), .ZN(n7124) );
  NOR2_X1 U8471 ( .A1(n11503), .A2(n11502), .ZN(n11517) );
  OR2_X1 U8472 ( .A1(n10808), .A2(n10807), .ZN(n11503) );
  INV_X1 U8473 ( .A(n10824), .ZN(n7615) );
  NOR2_X1 U8474 ( .A1(n8940), .A2(n8939), .ZN(n9199) );
  NAND2_X1 U8475 ( .A1(n11728), .A2(n11727), .ZN(n11725) );
  NAND2_X1 U8476 ( .A1(n14049), .A2(n7529), .ZN(n7528) );
  OAI21_X1 U8477 ( .B1(n6647), .B2(n7531), .A(n6704), .ZN(n7527) );
  INV_X1 U8478 ( .A(n10750), .ZN(n7467) );
  INV_X1 U8479 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U8480 ( .A1(n9178), .A2(n9177), .ZN(n9434) );
  INV_X1 U8481 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7707) );
  INV_X1 U8482 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7706) );
  INV_X1 U8483 ( .A(n8532), .ZN(n7476) );
  NAND2_X1 U8484 ( .A1(n8411), .A2(n8410), .ZN(n8646) );
  OR2_X1 U8485 ( .A1(n8015), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U8486 ( .A1(n6986), .A2(SI_3_), .ZN(n7814) );
  NAND2_X1 U8487 ( .A1(n7737), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7452) );
  AND2_X1 U8488 ( .A1(n14380), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7345) );
  INV_X1 U8489 ( .A(n14430), .ZN(n6906) );
  XNOR2_X1 U8490 ( .A(n14385), .B(n14384), .ZN(n14423) );
  NOR2_X1 U8491 ( .A1(n14392), .A2(n14391), .ZN(n14452) );
  NOR2_X1 U8492 ( .A1(n14450), .A2(n14449), .ZN(n14391) );
  AOI21_X1 U8493 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14394), .A(n14393), .ZN(
        n14421) );
  NOR2_X1 U8494 ( .A1(n14452), .A2(n14453), .ZN(n14393) );
  OAI22_X1 U8495 ( .A1(n14406), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n14414), 
        .B2(n14405), .ZN(n14468) );
  XNOR2_X1 U8496 ( .A(n12117), .B(n15120), .ZN(n9227) );
  NOR2_X1 U8497 ( .A1(n12192), .A2(n7258), .ZN(n12167) );
  AND2_X1 U8498 ( .A1(n12122), .A2(n12764), .ZN(n7258) );
  INV_X1 U8499 ( .A(n11988), .ZN(n9762) );
  INV_X1 U8500 ( .A(n9832), .ZN(n8138) );
  NAND2_X1 U8501 ( .A1(n10269), .A2(n10268), .ZN(n10617) );
  OR2_X1 U8502 ( .A1(n9859), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U8503 ( .A1(n7244), .A2(n8752), .ZN(n8960) );
  OR2_X1 U8504 ( .A1(n12130), .A2(n12437), .ZN(n7291) );
  NOR2_X1 U8505 ( .A1(n12266), .A2(n12265), .ZN(n7212) );
  AND2_X1 U8506 ( .A1(n6799), .A2(n6797), .ZN(n12415) );
  NAND2_X1 U8507 ( .A1(n12421), .A2(n9701), .ZN(n6824) );
  AND2_X1 U8508 ( .A1(n12228), .A2(n12227), .ZN(n12619) );
  OR2_X1 U8509 ( .A1(n8289), .A2(n15218), .ZN(n8545) );
  INV_X1 U8510 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U8511 ( .A1(n15002), .A2(n15001), .ZN(n15000) );
  INV_X1 U8512 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9423) );
  XNOR2_X1 U8513 ( .A(n10079), .B(n10141), .ZN(n15055) );
  AND2_X1 U8514 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  NOR2_X1 U8515 ( .A1(n10449), .A2(n10450), .ZN(n12454) );
  NAND2_X1 U8516 ( .A1(n12531), .A2(n12530), .ZN(n12552) );
  NAND2_X1 U8517 ( .A1(n8454), .A2(n7037), .ZN(n8869) );
  NAND2_X1 U8518 ( .A1(n7495), .A2(n12103), .ZN(n12649) );
  NAND2_X1 U8519 ( .A1(n12666), .A2(n12102), .ZN(n7495) );
  OAI21_X1 U8520 ( .B1(n12681), .B2(n7024), .A(n7020), .ZN(n12647) );
  INV_X1 U8521 ( .A(n7021), .ZN(n7020) );
  NAND2_X1 U8522 ( .A1(n12681), .A2(n12101), .ZN(n12666) );
  AND2_X1 U8523 ( .A1(n12065), .A2(n12064), .ZN(n12667) );
  INV_X1 U8524 ( .A(n12665), .ZN(n12663) );
  NAND2_X1 U8525 ( .A1(n9764), .A2(n9763), .ZN(n12034) );
  AND2_X1 U8526 ( .A1(n12398), .A2(n12399), .ZN(n12684) );
  INV_X1 U8527 ( .A(n12097), .ZN(n12710) );
  AOI21_X1 U8528 ( .B1(n7015), .B2(n7017), .A(n6751), .ZN(n7014) );
  INV_X1 U8529 ( .A(n7138), .ZN(n7137) );
  AOI21_X1 U8530 ( .B1(n7138), .B2(n7136), .A(n7135), .ZN(n7134) );
  AOI21_X1 U8531 ( .B1(n12754), .B2(n12375), .A(n7139), .ZN(n7138) );
  AND2_X1 U8532 ( .A1(n12382), .A2(n12383), .ZN(n12732) );
  NAND2_X1 U8533 ( .A1(n8814), .A2(n8813), .ZN(n10974) );
  OR2_X1 U8534 ( .A1(n10974), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n11988) );
  NAND2_X1 U8535 ( .A1(n10675), .A2(n8812), .ZN(n10882) );
  NAND2_X1 U8536 ( .A1(n8225), .A2(n8224), .ZN(n10572) );
  INV_X1 U8537 ( .A(n8226), .ZN(n8225) );
  INV_X1 U8538 ( .A(n12086), .ZN(n12811) );
  AOI21_X1 U8539 ( .B1(n7149), .B2(n12339), .A(n7148), .ZN(n7147) );
  INV_X1 U8540 ( .A(n12344), .ZN(n7148) );
  OR2_X1 U8541 ( .A1(n7150), .A2(n12339), .ZN(n12342) );
  OAI21_X1 U8542 ( .B1(n10204), .B2(n7011), .A(n7007), .ZN(n7012) );
  AOI21_X1 U8543 ( .B1(n12249), .B2(n7010), .A(n6732), .ZN(n7007) );
  NAND2_X1 U8544 ( .A1(n10217), .A2(n7010), .ZN(n10480) );
  NOR2_X1 U8545 ( .A1(n7009), .A2(n7008), .ZN(n10218) );
  INV_X1 U8546 ( .A(n10216), .ZN(n7008) );
  INV_X1 U8547 ( .A(n10217), .ZN(n7009) );
  NAND2_X1 U8548 ( .A1(n10204), .A2(n12310), .ZN(n10217) );
  NAND2_X1 U8549 ( .A1(n8137), .A2(n9722), .ZN(n9723) );
  INV_X1 U8550 ( .A(n9602), .ZN(n8137) );
  INV_X1 U8551 ( .A(n10215), .ZN(n10209) );
  NAND2_X1 U8552 ( .A1(n8136), .A2(n9423), .ZN(n9424) );
  INV_X1 U8553 ( .A(n9238), .ZN(n8136) );
  OR2_X1 U8554 ( .A1(n11984), .A2(n9596), .ZN(n9597) );
  AND2_X1 U8555 ( .A1(n12299), .A2(n12293), .ZN(n12297) );
  AND4_X1 U8556 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n10195)
         );
  NAND2_X1 U8557 ( .A1(n15121), .A2(n9237), .ZN(n9238) );
  INV_X1 U8558 ( .A(n15113), .ZN(n9362) );
  NAND2_X1 U8559 ( .A1(n12272), .A2(n12282), .ZN(n15145) );
  NAND2_X1 U8560 ( .A1(n12633), .A2(n6699), .ZN(n12108) );
  NAND2_X1 U8561 ( .A1(n12238), .A2(n12237), .ZN(n12240) );
  NAND2_X1 U8562 ( .A1(n12413), .A2(n12410), .ZN(n12266) );
  NAND2_X1 U8563 ( .A1(n11987), .A2(n11986), .ZN(n12164) );
  OR2_X1 U8564 ( .A1(n11985), .A2(n11984), .ZN(n11987) );
  NAND2_X1 U8565 ( .A1(n7145), .A2(n7143), .ZN(n12898) );
  NAND2_X1 U8566 ( .A1(n7145), .A2(n12360), .ZN(n12786) );
  OR2_X1 U8567 ( .A1(n10565), .A2(n11984), .ZN(n10567) );
  OR2_X1 U8568 ( .A1(n12697), .A2(n15206), .ZN(n14537) );
  INV_X1 U8569 ( .A(n9409), .ZN(n7209) );
  INV_X1 U8570 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7701) );
  AOI21_X1 U8571 ( .B1(n7194), .B2(n7196), .A(n7192), .ZN(n7191) );
  INV_X1 U8572 ( .A(n8874), .ZN(n7192) );
  NAND2_X1 U8573 ( .A1(n8382), .A2(n8381), .ZN(n8385) );
  NAND2_X1 U8574 ( .A1(n8385), .A2(n8384), .ZN(n8448) );
  NAND2_X1 U8575 ( .A1(n7198), .A2(n7201), .ZN(n8166) );
  AND2_X1 U8576 ( .A1(n8381), .A2(n8164), .ZN(n8165) );
  NAND2_X1 U8577 ( .A1(n8166), .A2(n8165), .ZN(n8382) );
  AOI21_X1 U8578 ( .B1(n7188), .B2(n7190), .A(n7186), .ZN(n7185) );
  INV_X1 U8579 ( .A(n7932), .ZN(n7186) );
  AND2_X1 U8580 ( .A1(n8018), .A2(n7934), .ZN(n7935) );
  NAND2_X1 U8581 ( .A1(n7878), .A2(n7845), .ZN(n7848) );
  OAI21_X1 U8582 ( .B1(n7867), .B2(n7206), .A(n7203), .ZN(n7876) );
  AOI21_X1 U8583 ( .B1(n7207), .B2(n7205), .A(n7204), .ZN(n7203) );
  INV_X1 U8584 ( .A(n7207), .ZN(n7206) );
  INV_X1 U8585 ( .A(n7843), .ZN(n7204) );
  AND2_X1 U8586 ( .A1(n7845), .A2(n7844), .ZN(n7875) );
  NAND2_X1 U8587 ( .A1(n7876), .A2(n7875), .ZN(n7878) );
  OR2_X1 U8588 ( .A1(n7939), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7886) );
  AND2_X1 U8589 ( .A1(n7780), .A2(n7779), .ZN(n7800) );
  NAND2_X1 U8590 ( .A1(n7807), .A2(n7806), .ZN(n14997) );
  OR3_X1 U8591 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U8592 ( .A1(n7774), .A2(n7773), .ZN(n7795) );
  NAND2_X1 U8593 ( .A1(n6661), .A2(n6935), .ZN(n6934) );
  AOI22_X1 U8594 ( .A1(n11358), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n11169), 
        .B2(n8773), .ZN(n8775) );
  NOR2_X1 U8595 ( .A1(n13064), .A2(n13033), .ZN(n7376) );
  XNOR2_X1 U8596 ( .A(n8719), .B(n8735), .ZN(n8354) );
  INV_X1 U8597 ( .A(n8780), .ZN(n7350) );
  OR2_X1 U8598 ( .A1(n13123), .A2(n7380), .ZN(n7379) );
  INV_X1 U8599 ( .A(n11189), .ZN(n11014) );
  NOR2_X1 U8600 ( .A1(n9384), .A2(n9382), .ZN(n9747) );
  INV_X1 U8601 ( .A(n6847), .ZN(n11370) );
  CLKBUF_X1 U8602 ( .A(n9136), .Z(n11277) );
  OR2_X1 U8603 ( .A1(n11337), .A2(n8332), .ZN(n8339) );
  OR2_X1 U8604 ( .A1(n11333), .A2(n8334), .ZN(n8338) );
  XNOR2_X1 U8605 ( .A(n14760), .B(n8389), .ZN(n14755) );
  AND2_X1 U8606 ( .A1(n14756), .A2(n14755), .ZN(n14758) );
  NOR2_X1 U8607 ( .A1(n14758), .A2(n6998), .ZN(n8424) );
  AND2_X1 U8608 ( .A1(n14760), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U8609 ( .A1(n14768), .A2(n6717), .ZN(n8435) );
  NOR2_X1 U8610 ( .A1(n9651), .A2(n6776), .ZN(n14812) );
  NOR2_X1 U8611 ( .A1(n14812), .A2(n14811), .ZN(n14810) );
  XNOR2_X1 U8612 ( .A(n13179), .B(n13178), .ZN(n13172) );
  NOR2_X1 U8613 ( .A1(n14835), .A2(n6995), .ZN(n13179) );
  AND2_X1 U8614 ( .A1(n13171), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6995) );
  NOR2_X1 U8615 ( .A1(n13172), .A2(n13614), .ZN(n13180) );
  NAND2_X1 U8616 ( .A1(n14853), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8617 ( .A1(n11274), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U8618 ( .A1(n7388), .A2(n13309), .ZN(n13343) );
  NAND2_X1 U8619 ( .A1(n13358), .A2(n13308), .ZN(n7388) );
  INV_X1 U8620 ( .A(n13558), .ZN(n7114) );
  INV_X1 U8621 ( .A(n13409), .ZN(n7115) );
  NAND2_X1 U8622 ( .A1(n6836), .A2(n13303), .ZN(n13387) );
  OR2_X1 U8623 ( .A1(n11202), .A2(n13115), .ZN(n11217) );
  AOI21_X1 U8624 ( .B1(n7232), .B2(n7235), .A(n7230), .ZN(n7229) );
  NAND2_X1 U8625 ( .A1(n7397), .A2(n7401), .ZN(n13475) );
  NAND2_X1 U8626 ( .A1(n6916), .A2(n7404), .ZN(n7397) );
  OR2_X1 U8627 ( .A1(n11159), .A2(n11012), .ZN(n11173) );
  INV_X1 U8628 ( .A(n7238), .ZN(n7237) );
  OR2_X1 U8629 ( .A1(n10633), .A2(n10632), .ZN(n10696) );
  NAND2_X1 U8630 ( .A1(n10630), .A2(n10629), .ZN(n11125) );
  AND2_X1 U8631 ( .A1(n9747), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9892) );
  NAND2_X1 U8632 ( .A1(n7216), .A2(n7218), .ZN(n7214) );
  INV_X1 U8633 ( .A(n10231), .ZN(n7108) );
  OR2_X1 U8634 ( .A1(n9024), .A2(n9146), .ZN(n9139) );
  NAND2_X1 U8635 ( .A1(n7223), .A2(n7224), .ZN(n9289) );
  NAND2_X1 U8636 ( .A1(n6746), .A2(n9288), .ZN(n7223) );
  NAND2_X1 U8637 ( .A1(n9462), .A2(n7225), .ZN(n7224) );
  NOR2_X2 U8638 ( .A1(n9484), .A2(n11075), .ZN(n9543) );
  INV_X1 U8639 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8904) );
  OR2_X1 U8640 ( .A1(n11449), .A2(n8374), .ZN(n8594) );
  INV_X1 U8641 ( .A(n9275), .ZN(n11399) );
  OAI211_X1 U8642 ( .C1(n11236), .C2(n8614), .A(n7393), .B(n7392), .ZN(n11040)
         );
  NAND2_X1 U8643 ( .A1(n8723), .A2(n14748), .ZN(n7392) );
  OR2_X1 U8644 ( .A1(n11363), .A2(n8347), .ZN(n7393) );
  NAND2_X1 U8645 ( .A1(n11201), .A2(n11200), .ZN(n13423) );
  NOR2_X1 U8646 ( .A1(n13501), .A2(n13599), .ZN(n13489) );
  NAND2_X1 U8647 ( .A1(n10325), .A2(n10324), .ZN(n13618) );
  NAND2_X1 U8648 ( .A1(n9687), .A2(n9686), .ZN(n10230) );
  INV_X1 U8649 ( .A(n14953), .ZN(n14927) );
  OR2_X1 U8650 ( .A1(n8374), .A2(n11455), .ZN(n14953) );
  OR2_X1 U8651 ( .A1(n7671), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n7668) );
  INV_X1 U8652 ( .A(n10318), .ZN(n7046) );
  NAND3_X1 U8653 ( .A1(n7648), .A2(n7385), .A3(n8237), .ZN(n8319) );
  OR2_X1 U8654 ( .A1(n7905), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7897) );
  AND2_X1 U8655 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n11687), .ZN(n11688) );
  NAND2_X1 U8656 ( .A1(n7097), .A2(n7098), .ZN(n13713) );
  NAND2_X1 U8657 ( .A1(n6866), .A2(n7100), .ZN(n7097) );
  INV_X1 U8658 ( .A(n11580), .ZN(n11581) );
  NAND2_X1 U8659 ( .A1(n13783), .A2(n13784), .ZN(n13782) );
  NOR2_X1 U8660 ( .A1(n8625), .A2(n8624), .ZN(n8627) );
  CLKBUF_X1 U8661 ( .A(n13747), .Z(n6866) );
  AND4_X1 U8662 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n13924) );
  AND2_X1 U8663 ( .A1(n11556), .A2(n11555), .ZN(n13920) );
  AND4_X1 U8664 ( .A1(n10805), .A2(n10804), .A3(n10803), .A4(n10802), .ZN(
        n10806) );
  AND4_X1 U8665 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(n11775)
         );
  OR2_X1 U8666 ( .A1(n11656), .A2(n15504), .ZN(n8633) );
  INV_X1 U8667 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14379) );
  OR2_X1 U8668 ( .A1(n8643), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9165) );
  NOR2_X1 U8669 ( .A1(n7129), .A2(n7127), .ZN(n7126) );
  INV_X1 U8670 ( .A(n7128), .ZN(n7127) );
  NAND2_X1 U8671 ( .A1(n7637), .A2(n7643), .ZN(n7642) );
  NOR2_X2 U8672 ( .A1(n13991), .A2(n14004), .ZN(n13978) );
  AND4_X1 U8673 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n14021) );
  NOR2_X1 U8674 ( .A1(n6685), .A2(n14030), .ZN(n14027) );
  AND2_X1 U8675 ( .A1(n7536), .A2(n6706), .ZN(n14035) );
  NAND2_X1 U8676 ( .A1(n14049), .A2(n14058), .ZN(n7536) );
  OR2_X1 U8677 ( .A1(n14100), .A2(n14261), .ZN(n14066) );
  NOR2_X1 U8678 ( .A1(n14098), .A2(n14263), .ZN(n14065) );
  INV_X1 U8679 ( .A(n13943), .ZN(n7540) );
  AND2_X1 U8680 ( .A1(n14085), .A2(n7539), .ZN(n7538) );
  NAND2_X1 U8681 ( .A1(n7542), .A2(n13943), .ZN(n7539) );
  NAND2_X1 U8682 ( .A1(n14108), .A2(n13943), .ZN(n14086) );
  NOR3_X1 U8683 ( .A1(n14170), .A2(n14133), .A3(n7124), .ZN(n14129) );
  OR2_X1 U8684 ( .A1(n11532), .A2(n13716), .ZN(n11548) );
  NOR2_X1 U8685 ( .A1(n14170), .A2(n7124), .ZN(n14138) );
  NOR2_X1 U8686 ( .A1(n14170), .A2(n14158), .ZN(n14157) );
  INV_X1 U8687 ( .A(n7546), .ZN(n7545) );
  AOI21_X1 U8688 ( .B1(n7546), .B2(n7544), .A(n6711), .ZN(n7543) );
  AND2_X1 U8689 ( .A1(n7547), .A2(n13939), .ZN(n7546) );
  OR2_X1 U8690 ( .A1(n14172), .A2(n14300), .ZN(n14170) );
  NAND2_X1 U8691 ( .A1(n6806), .A2(n14355), .ZN(n14172) );
  INV_X1 U8692 ( .A(n11915), .ZN(n14603) );
  NAND2_X1 U8693 ( .A1(n10788), .A2(n10787), .ZN(n14602) );
  NAND2_X1 U8694 ( .A1(n14505), .A2(n14619), .ZN(n14601) );
  NOR2_X1 U8695 ( .A1(n10414), .A2(n15476), .ZN(n10789) );
  OR2_X1 U8696 ( .A1(n10251), .A2(n10250), .ZN(n10414) );
  AND4_X1 U8697 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n13772) );
  AND2_X1 U8698 ( .A1(n7550), .A2(n11928), .ZN(n7548) );
  NAND2_X1 U8699 ( .A1(n7125), .A2(n14582), .ZN(n10426) );
  NAND2_X1 U8700 ( .A1(n10018), .A2(n10017), .ZN(n10244) );
  INV_X1 U8701 ( .A(n7125), .ZN(n10261) );
  NOR2_X1 U8702 ( .A1(n9802), .A2(n10523), .ZN(n10007) );
  OR2_X1 U8703 ( .A1(n9528), .A2(n9527), .ZN(n9802) );
  INV_X1 U8704 ( .A(n9984), .ZN(n7611) );
  INV_X1 U8705 ( .A(n11924), .ZN(n7612) );
  OR2_X1 U8706 ( .A1(n9324), .A2(n9323), .ZN(n9528) );
  NAND2_X1 U8707 ( .A1(n9985), .A2(n9984), .ZN(n10034) );
  NAND2_X1 U8708 ( .A1(n7524), .A2(n9970), .ZN(n10033) );
  NAND2_X1 U8709 ( .A1(n9968), .A2(n11922), .ZN(n7524) );
  NAND2_X1 U8710 ( .A1(n7121), .A2(n7525), .ZN(n10046) );
  INV_X1 U8711 ( .A(n10031), .ZN(n7121) );
  NOR2_X1 U8712 ( .A1(n9818), .A2(n11751), .ZN(n9624) );
  NAND2_X1 U8713 ( .A1(n9624), .A2(n9623), .ZN(n10031) );
  OR2_X1 U8714 ( .A1(n8936), .A2(n11743), .ZN(n9818) );
  NAND2_X1 U8715 ( .A1(n8935), .A2(n11736), .ZN(n9632) );
  AND2_X1 U8716 ( .A1(n14694), .A2(n14189), .ZN(n14191) );
  AND2_X1 U8717 ( .A1(n14191), .A2(n11727), .ZN(n8861) );
  INV_X1 U8718 ( .A(n14719), .ZN(n14504) );
  NAND2_X1 U8719 ( .A1(n11678), .A2(n8278), .ZN(n14289) );
  NAND2_X1 U8720 ( .A1(n11353), .A2(n11343), .ZN(n11309) );
  XNOR2_X1 U8721 ( .A(n11002), .B(n10999), .ZN(n11666) );
  AND2_X1 U8722 ( .A1(n7731), .A2(n7730), .ZN(n7944) );
  NAND2_X1 U8723 ( .A1(n10933), .A2(n10749), .ZN(n10751) );
  NAND2_X1 U8724 ( .A1(n10545), .A2(n10316), .ZN(n11576) );
  NAND2_X1 U8725 ( .A1(n7970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7968) );
  AOI21_X1 U8726 ( .B1(n8030), .B2(n6970), .A(n6748), .ZN(n6968) );
  INV_X1 U8727 ( .A(n6970), .ZN(n6969) );
  AND2_X1 U8728 ( .A1(n8039), .A2(n8419), .ZN(n9965) );
  NAND2_X1 U8729 ( .A1(n8032), .A2(n8031), .ZN(n8411) );
  AOI21_X1 U8730 ( .B1(n7461), .B2(n7463), .A(n7460), .ZN(n7459) );
  INV_X1 U8731 ( .A(n8004), .ZN(n7460) );
  AND2_X1 U8732 ( .A1(n7856), .A2(n7855), .ZN(n7964) );
  OR2_X1 U8733 ( .A1(n7809), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n7811) );
  NOR2_X1 U8734 ( .A1(n7811), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7856) );
  OAI21_X1 U8735 ( .B1(SI_3_), .B2(n6986), .A(n7814), .ZN(n7754) );
  OAI21_X1 U8736 ( .B1(n8346), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6872), .ZN(
        n7740) );
  OR2_X1 U8737 ( .A1(n7737), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6872) );
  INV_X1 U8738 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14426) );
  XNOR2_X1 U8739 ( .A(n14424), .B(n6910), .ZN(n14427) );
  INV_X1 U8740 ( .A(n14425), .ZN(n6910) );
  INV_X1 U8741 ( .A(n7346), .ZN(n14431) );
  XNOR2_X1 U8742 ( .A(n14381), .B(n15343), .ZN(n14435) );
  XNOR2_X1 U8743 ( .A(n14423), .B(n6862), .ZN(n14437) );
  INV_X1 U8744 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6862) );
  XNOR2_X1 U8745 ( .A(n14439), .B(n7314), .ZN(n14441) );
  INV_X1 U8746 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7314) );
  NOR2_X1 U8747 ( .A1(n14388), .A2(n14387), .ZN(n14444) );
  NOR2_X1 U8748 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14439), .ZN(n14387) );
  AOI21_X1 U8749 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(n14461) );
  INV_X1 U8750 ( .A(n7284), .ZN(n7278) );
  NAND2_X1 U8751 ( .A1(n7273), .A2(n7272), .ZN(n7279) );
  AND2_X1 U8752 ( .A1(n7286), .A2(n7292), .ZN(n7272) );
  NAND2_X1 U8753 ( .A1(n9046), .A2(n9045), .ZN(n9229) );
  INV_X1 U8754 ( .A(n7032), .ZN(n12146) );
  INV_X1 U8755 ( .A(n7246), .ZN(n12144) );
  NAND2_X1 U8756 ( .A1(n7275), .A2(n6724), .ZN(n12157) );
  NOR2_X1 U8757 ( .A1(n7283), .A2(n7277), .ZN(n7276) );
  AND4_X1 U8758 ( .A1(n8265), .A2(n8264), .A3(n8263), .A4(n8262), .ZN(n10757)
         );
  INV_X1 U8759 ( .A(n12436), .ZN(n12680) );
  AND2_X1 U8760 ( .A1(n7273), .A2(n7292), .ZN(n12175) );
  NAND2_X1 U8761 ( .A1(n12033), .A2(n12032), .ZN(n12866) );
  NAND2_X1 U8762 ( .A1(n10674), .A2(n10673), .ZN(n10879) );
  INV_X1 U8763 ( .A(n7253), .ZN(n7252) );
  INV_X1 U8764 ( .A(n9419), .ZN(n7251) );
  NAND2_X1 U8765 ( .A1(n9420), .A2(n9421), .ZN(n9846) );
  AND4_X1 U8766 ( .A1(n10888), .A2(n10887), .A3(n10886), .A4(n10885), .ZN(
        n12091) );
  NAND2_X1 U8767 ( .A1(n10879), .A2(n6814), .ZN(n10881) );
  NAND2_X1 U8768 ( .A1(n10878), .A2(n6815), .ZN(n6814) );
  NAND2_X1 U8769 ( .A1(n10881), .A2(n10880), .ZN(n10967) );
  NAND2_X1 U8770 ( .A1(n9229), .A2(n9228), .ZN(n9236) );
  NAND2_X1 U8771 ( .A1(n9854), .A2(n9855), .ZN(n9856) );
  AND2_X1 U8772 ( .A1(n7246), .A2(n7245), .ZN(n12193) );
  NAND2_X1 U8773 ( .A1(n12121), .A2(n12440), .ZN(n7245) );
  NAND2_X1 U8774 ( .A1(n7267), .A2(n7271), .ZN(n10504) );
  NAND2_X1 U8775 ( .A1(n10269), .A2(n7268), .ZN(n7267) );
  INV_X1 U8776 ( .A(n12125), .ZN(n7255) );
  NAND2_X1 U8777 ( .A1(n11998), .A2(n11997), .ZN(n12733) );
  XNOR2_X1 U8778 ( .A(n9038), .B(n9359), .ZN(n8962) );
  OR2_X1 U8779 ( .A1(n12236), .A2(SI_2_), .ZN(n8958) );
  OR2_X1 U8780 ( .A1(n11984), .A2(n8955), .ZN(n8957) );
  AND2_X1 U8781 ( .A1(n12041), .A2(n12040), .ZN(n12695) );
  AND2_X1 U8782 ( .A1(n8522), .A2(n8521), .ZN(n12212) );
  OAI21_X1 U8783 ( .B1(n12175), .B2(n12176), .A(n7291), .ZN(n6919) );
  INV_X1 U8784 ( .A(n12206), .ZN(n6918) );
  AND2_X1 U8785 ( .A1(n12228), .A2(n9789), .ZN(n12636) );
  INV_X1 U8786 ( .A(n12667), .ZN(n12435) );
  INV_X1 U8787 ( .A(n12695), .ZN(n12437) );
  INV_X1 U8788 ( .A(n12091), .ZN(n12796) );
  INV_X1 U8789 ( .A(n10757), .ZN(n10761) );
  INV_X1 U8790 ( .A(n10195), .ZN(n12446) );
  INV_X1 U8791 ( .A(n7178), .ZN(n15025) );
  INV_X1 U8792 ( .A(n7176), .ZN(n10142) );
  AND2_X1 U8793 ( .A1(n7169), .A2(n7168), .ZN(n10149) );
  NAND2_X1 U8794 ( .A1(n7167), .A2(n7166), .ZN(n10172) );
  AND2_X1 U8795 ( .A1(n15093), .A2(n10083), .ZN(n10084) );
  NAND2_X1 U8796 ( .A1(n12478), .A2(n12479), .ZN(n12480) );
  INV_X1 U8797 ( .A(n7181), .ZN(n12472) );
  INV_X1 U8798 ( .A(n7180), .ZN(n12499) );
  INV_X1 U8799 ( .A(n6828), .ZN(n12519) );
  NAND2_X1 U8800 ( .A1(n7499), .A2(n12094), .ZN(n12739) );
  OAI21_X1 U8801 ( .B1(n12774), .B2(n7017), .A(n7015), .ZN(n7499) );
  NAND2_X1 U8802 ( .A1(n12757), .A2(n12375), .ZN(n12744) );
  NAND2_X1 U8803 ( .A1(n12763), .A2(n12093), .ZN(n12750) );
  NAND2_X1 U8804 ( .A1(n12090), .A2(n12089), .ZN(n12776) );
  NAND2_X1 U8805 ( .A1(n10965), .A2(n10964), .ZN(n12791) );
  OR2_X1 U8806 ( .A1(n10963), .A2(n11984), .ZN(n10965) );
  NAND2_X1 U8807 ( .A1(n7151), .A2(n7149), .ZN(n12838) );
  NAND2_X1 U8808 ( .A1(n7153), .A2(n7152), .ZN(n7151) );
  OR2_X1 U8809 ( .A1(n10286), .A2(n11984), .ZN(n10288) );
  INV_X1 U8810 ( .A(n12787), .ZN(n12844) );
  NAND2_X1 U8811 ( .A1(n10729), .A2(n10728), .ZN(n10732) );
  NAND2_X1 U8812 ( .A1(n7159), .A2(n7157), .ZN(n10755) );
  NAND2_X1 U8813 ( .A1(n10734), .A2(n12255), .ZN(n7159) );
  NOR2_X1 U8814 ( .A1(n7497), .A2(n7496), .ZN(n10202) );
  AND3_X1 U8815 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(n9512) );
  OR2_X1 U8816 ( .A1(n11984), .A2(n9415), .ZN(n9417) );
  NAND2_X1 U8817 ( .A1(n15116), .A2(n9363), .ZN(n9365) );
  INV_X1 U8818 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15121) );
  INV_X1 U8819 ( .A(n12782), .ZN(n15157) );
  INV_X1 U8820 ( .A(n12240), .ZN(n12921) );
  NAND2_X1 U8821 ( .A1(n12221), .A2(n12220), .ZN(n12922) );
  INV_X1 U8822 ( .A(n12161), .ZN(n12929) );
  NAND2_X1 U8823 ( .A1(n12010), .A2(n12009), .ZN(n12945) );
  AND2_X1 U8824 ( .A1(n8112), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8506) );
  NAND2_X1 U8825 ( .A1(n8127), .A2(n6727), .ZN(n6999) );
  AND2_X1 U8826 ( .A1(n12982), .A2(n7001), .ZN(n7000) );
  AND2_X1 U8827 ( .A1(n6709), .A2(n7689), .ZN(n7504) );
  INV_X1 U8828 ( .A(n9404), .ZN(n9403) );
  NAND2_X1 U8829 ( .A1(n7034), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U8830 ( .A1(n8822), .A2(n8821), .ZN(n8873) );
  NAND2_X1 U8831 ( .A1(n8454), .A2(n8453), .ZN(n8456) );
  NAND2_X1 U8832 ( .A1(n8025), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U8833 ( .A1(n7197), .A2(n7201), .ZN(n8163) );
  NAND2_X1 U8834 ( .A1(n7199), .A2(n7201), .ZN(n8021) );
  OAI21_X1 U8835 ( .B1(n7884), .B2(n7190), .A(n7188), .ZN(n7933) );
  NAND2_X1 U8836 ( .A1(n7912), .A2(n7911), .ZN(n7915) );
  NAND2_X1 U8837 ( .A1(n7202), .A2(n7207), .ZN(n7892) );
  NAND2_X1 U8838 ( .A1(n7867), .A2(n7841), .ZN(n7202) );
  INV_X1 U8839 ( .A(n10105), .ZN(n15033) );
  OAI21_X1 U8840 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        n7184), .ZN(n7183) );
  INV_X1 U8841 ( .A(n7384), .ZN(n7383) );
  NAND2_X1 U8842 ( .A1(n10687), .A2(n10686), .ZN(n14547) );
  NAND2_X1 U8843 ( .A1(n8772), .A2(n8771), .ZN(n8781) );
  INV_X1 U8844 ( .A(n7379), .ZN(n13057) );
  OAI22_X1 U8845 ( .A1(n13123), .A2(n6936), .B1(n6675), .B2(n13102), .ZN(
        n13075) );
  NAND2_X1 U8846 ( .A1(n6937), .A2(n6938), .ZN(n6936) );
  NAND2_X1 U8847 ( .A1(n9908), .A2(n9921), .ZN(n10330) );
  NAND2_X1 U8848 ( .A1(n10330), .A2(n6661), .ZN(n10687) );
  AND2_X1 U8849 ( .A1(n10330), .A2(n10329), .ZN(n10337) );
  XNOR2_X1 U8850 ( .A(n8768), .B(n8769), .ZN(n8736) );
  NAND2_X1 U8851 ( .A1(n9016), .A2(n9015), .ZN(n9022) );
  XNOR2_X1 U8852 ( .A(n10952), .B(n10950), .ZN(n10694) );
  NAND2_X1 U8853 ( .A1(n10694), .A2(n6863), .ZN(n10954) );
  AND2_X1 U8854 ( .A1(n13143), .A2(n13030), .ZN(n6863) );
  NAND2_X1 U8855 ( .A1(n6698), .A2(n6851), .ZN(n7477) );
  NAND2_X1 U8856 ( .A1(n11447), .A2(n11393), .ZN(n6851) );
  NAND2_X1 U8857 ( .A1(n11445), .A2(n7652), .ZN(n11446) );
  NAND2_X1 U8858 ( .A1(n11448), .A2(n11450), .ZN(n11445) );
  NAND4_X1 U8859 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n13149)
         );
  NOR2_X1 U8860 ( .A1(n11317), .A2(n10065), .ZN(n6878) );
  OR2_X1 U8861 ( .A1(n11337), .A2(n9570), .ZN(n8363) );
  INV_X1 U8862 ( .A(n6988), .ZN(n14784) );
  NOR2_X1 U8863 ( .A1(n14795), .A2(n6770), .ZN(n8882) );
  NAND2_X1 U8864 ( .A1(n8882), .A2(n8881), .ZN(n9215) );
  NAND2_X1 U8865 ( .A1(n9653), .A2(n9654), .ZN(n13168) );
  INV_X1 U8866 ( .A(n6993), .ZN(n14850) );
  INV_X1 U8867 ( .A(n6991), .ZN(n14848) );
  NOR2_X1 U8868 ( .A1(n7222), .A2(n6667), .ZN(n7044) );
  NAND2_X1 U8869 ( .A1(n7222), .A2(n6667), .ZN(n7043) );
  AND2_X1 U8870 ( .A1(n7056), .A2(n6705), .ZN(n13355) );
  NAND2_X1 U8871 ( .A1(n13276), .A2(n13275), .ZN(n13366) );
  NAND2_X1 U8872 ( .A1(n13389), .A2(n13305), .ZN(n13372) );
  NAND2_X1 U8873 ( .A1(n13557), .A2(n13272), .ZN(n13376) );
  NAND2_X1 U8874 ( .A1(n13270), .A2(n7242), .ZN(n13557) );
  NAND2_X1 U8875 ( .A1(n13270), .A2(n13269), .ZN(n13399) );
  OAI21_X1 U8876 ( .B1(n13468), .B2(n7235), .A(n7232), .ZN(n13437) );
  NAND2_X1 U8877 ( .A1(n7231), .A2(n13257), .ZN(n13450) );
  NAND2_X1 U8878 ( .A1(n13468), .A2(n13256), .ZN(n7231) );
  NAND2_X1 U8879 ( .A1(n7405), .A2(n7407), .ZN(n13482) );
  NAND2_X1 U8880 ( .A1(n13250), .A2(n13249), .ZN(n13506) );
  NAND2_X1 U8881 ( .A1(n10895), .A2(n10894), .ZN(n10898) );
  NAND2_X1 U8882 ( .A1(n10897), .A2(n10896), .ZN(n13603) );
  NAND2_X1 U8883 ( .A1(n10368), .A2(n10367), .ZN(n10371) );
  NAND2_X1 U8884 ( .A1(n9907), .A2(n9906), .ZN(n11116) );
  OAI21_X1 U8885 ( .B1(n9687), .B2(n7218), .A(n7216), .ZN(n10350) );
  NAND2_X1 U8886 ( .A1(n7227), .A2(n9286), .ZN(n9476) );
  NAND2_X1 U8887 ( .A1(n11402), .A2(n9462), .ZN(n7227) );
  CLKBUF_X1 U8888 ( .A(n11040), .Z(n6820) );
  INV_X1 U8889 ( .A(n14868), .ZN(n13517) );
  INV_X1 U8890 ( .A(n13507), .ZN(n14872) );
  NAND2_X1 U8891 ( .A1(n14968), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6859) );
  INV_X1 U8892 ( .A(n6922), .ZN(n6921) );
  NAND2_X1 U8893 ( .A1(n13336), .A2(n6902), .ZN(n6901) );
  NAND2_X1 U8894 ( .A1(n8782), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14907) );
  NAND2_X1 U8895 ( .A1(n8244), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8896 ( .A1(n7648), .A2(n7385), .ZN(n8321) );
  INV_X1 U8897 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9443) );
  INV_X1 U8898 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9181) );
  INV_X1 U8899 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9093) );
  INV_X1 U8900 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9160) );
  INV_X1 U8901 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8535) );
  NOR2_X1 U8902 ( .A1(n8656), .A2(n8655), .ZN(n14815) );
  INV_X1 U8903 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8418) );
  INV_X1 U8904 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8035) );
  INV_X1 U8905 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8014) );
  INV_X1 U8906 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7962) );
  INV_X1 U8907 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7931) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n15518) );
  INV_X1 U8909 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7901) );
  INV_X1 U8910 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7907) );
  INV_X1 U8911 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8724) );
  INV_X1 U8912 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U8913 ( .A1(n9519), .A2(n6816), .ZN(n9525) );
  NAND2_X1 U8914 ( .A1(n6818), .A2(n6817), .ZN(n6816) );
  INV_X1 U8915 ( .A(n9521), .ZN(n6817) );
  INV_X1 U8916 ( .A(n9520), .ZN(n6818) );
  NAND2_X1 U8917 ( .A1(n13782), .A2(n11594), .ZN(n13694) );
  AND2_X1 U8918 ( .A1(n13706), .A2(n13703), .ZN(n6865) );
  OR2_X1 U8919 ( .A1(n13713), .A2(n13712), .ZN(n13714) );
  INV_X1 U8920 ( .A(n7096), .ZN(n7095) );
  AOI21_X1 U8921 ( .B1(n7438), .B2(n7436), .A(n6707), .ZN(n7435) );
  AND2_X1 U8922 ( .A1(n7075), .A2(n7082), .ZN(n9316) );
  NAND2_X1 U8923 ( .A1(n7073), .A2(n7081), .ZN(n7082) );
  AOI21_X1 U8924 ( .B1(n7427), .B2(n7430), .A(n6740), .ZN(n7426) );
  OAI211_X1 U8925 ( .C1(n13705), .C2(n7081), .A(n7079), .B(n7076), .ZN(n9185)
         );
  NAND2_X1 U8926 ( .A1(n13705), .A2(n7078), .ZN(n7076) );
  NAND2_X1 U8927 ( .A1(n13714), .A2(n11543), .ZN(n13764) );
  NAND2_X1 U8928 ( .A1(n7434), .A2(n7438), .ZN(n13762) );
  NAND2_X1 U8929 ( .A1(n13713), .A2(n11543), .ZN(n7434) );
  INV_X1 U8930 ( .A(n7441), .ZN(n7440) );
  INV_X1 U8931 ( .A(n10663), .ZN(n7090) );
  INV_X1 U8932 ( .A(n10861), .ZN(n7443) );
  NAND2_X1 U8933 ( .A1(n9065), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14588) );
  AOI21_X1 U8934 ( .B1(n6866), .B2(n13746), .A(n11513), .ZN(n13792) );
  NAND2_X1 U8935 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  NOR2_X1 U8936 ( .A1(n9315), .A2(n9183), .ZN(n7072) );
  AND2_X1 U8937 ( .A1(n9063), .A2(n8187), .ZN(n11957) );
  AND2_X1 U8938 ( .A1(n8637), .A2(n8636), .ZN(n14262) );
  AOI21_X1 U8939 ( .B1(n11949), .B2(n11948), .A(n11947), .ZN(n11950) );
  OAI21_X1 U8940 ( .B1(n11875), .B2(n7311), .A(n7309), .ZN(n11953) );
  OR2_X1 U8941 ( .A1(n11881), .A2(n8174), .ZN(n8178) );
  AND2_X1 U8942 ( .A1(n8207), .A2(n8205), .ZN(n6927) );
  OR2_X1 U8943 ( .A1(n13964), .A2(n6985), .ZN(n14227) );
  AOI21_X1 U8944 ( .B1(n13932), .B2(n13931), .A(n13933), .ZN(n6985) );
  NAND2_X1 U8945 ( .A1(n14019), .A2(n14018), .ZN(n14017) );
  NAND2_X1 U8946 ( .A1(n7533), .A2(n7531), .ZN(n14019) );
  NAND2_X1 U8947 ( .A1(n14049), .A2(n7534), .ZN(n7533) );
  AND2_X1 U8948 ( .A1(n14061), .A2(n14060), .ZN(n14256) );
  NAND2_X1 U8949 ( .A1(n14069), .A2(n13922), .ZN(n14059) );
  AND4_X1 U8950 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n14080) );
  AND2_X1 U8951 ( .A1(n14123), .A2(n13942), .ZN(n14109) );
  NAND2_X1 U8952 ( .A1(n7622), .A2(n7620), .ZN(n14134) );
  NAND2_X1 U8953 ( .A1(n7626), .A2(n13914), .ZN(n14137) );
  NAND2_X1 U8954 ( .A1(n14155), .A2(n13913), .ZN(n7626) );
  NAND2_X1 U8955 ( .A1(n14167), .A2(n13938), .ZN(n14154) );
  NAND2_X1 U8956 ( .A1(n6977), .A2(n6981), .ZN(n14183) );
  NAND2_X1 U8957 ( .A1(n13909), .A2(n13911), .ZN(n6977) );
  INV_X1 U8958 ( .A(n11798), .ZN(n14619) );
  NAND2_X1 U8959 ( .A1(n7613), .A2(n7617), .ZN(n14501) );
  NAND2_X1 U8960 ( .A1(n10823), .A2(n10824), .ZN(n7613) );
  AND2_X1 U8961 ( .A1(n10411), .A2(n10410), .ZN(n11791) );
  NAND2_X1 U8962 ( .A1(n10258), .A2(n10257), .ZN(n10412) );
  NAND2_X1 U8963 ( .A1(n7597), .A2(n7598), .ZN(n10405) );
  OAI21_X1 U8964 ( .B1(n9968), .B2(n7521), .A(n7520), .ZN(n10042) );
  NAND2_X1 U8965 ( .A1(n7605), .A2(n9627), .ZN(n9816) );
  NAND2_X1 U8966 ( .A1(n9626), .A2(n9625), .ZN(n7605) );
  INV_X1 U8967 ( .A(n14130), .ZN(n14606) );
  INV_X1 U8968 ( .A(n14153), .ZN(n14605) );
  OR2_X1 U8969 ( .A1(n9616), .A2(n9615), .ZN(n14683) );
  AND2_X1 U8970 ( .A1(n8610), .A2(n8608), .ZN(n7092) );
  NAND2_X1 U8971 ( .A1(n13665), .A2(n11897), .ZN(n7060) );
  INV_X1 U8972 ( .A(n13991), .ZN(n14327) );
  INV_X1 U8973 ( .A(n14030), .ZN(n14332) );
  OR2_X1 U8974 ( .A1(n14254), .A2(n14253), .ZN(n14333) );
  AND2_X1 U8975 ( .A1(n11598), .A2(n11597), .ZN(n14337) );
  AND2_X1 U8976 ( .A1(n11563), .A2(n11562), .ZN(n14342) );
  INV_X1 U8977 ( .A(n11791), .ZN(n11792) );
  NAND2_X1 U8978 ( .A1(n6984), .A2(n11897), .ZN(n6983) );
  INV_X1 U8979 ( .A(n9999), .ZN(n6984) );
  NAND2_X1 U8980 ( .A1(n11528), .A2(n13853), .ZN(n7321) );
  OR2_X1 U8981 ( .A1(n6660), .A2(n7775), .ZN(n7322) );
  AND2_X1 U8982 ( .A1(n7630), .A2(n8169), .ZN(n7629) );
  OAI21_X1 U8983 ( .B1(n7976), .B2(P1_IR_REG_31__SCAN_IN), .A(n7066), .ZN(
        n7065) );
  NAND2_X1 U8984 ( .A1(n7974), .A2(n7068), .ZN(n7067) );
  XNOR2_X1 U8985 ( .A(n10745), .B(n10743), .ZN(n11595) );
  INV_X1 U8986 ( .A(n8279), .ZN(n11908) );
  NAND2_X1 U8987 ( .A1(n8183), .A2(n8182), .ZN(n11902) );
  NAND2_X1 U8988 ( .A1(n7061), .A2(n9935), .ZN(n9936) );
  NAND2_X1 U8989 ( .A1(n9589), .A2(n9935), .ZN(n9591) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9179) );
  INV_X1 U8991 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9098) );
  INV_X1 U8992 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9168) );
  INV_X1 U8993 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8538) );
  INV_X1 U8994 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n15391) );
  INV_X1 U8995 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8421) );
  INV_X1 U8996 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8040) );
  INV_X1 U8997 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8017) );
  INV_X1 U8998 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7966) );
  OAI21_X1 U8999 ( .B1(n7924), .B2(n7463), .A(n7461), .ZN(n8005) );
  INV_X1 U9000 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7926) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7865) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U9003 ( .A1(n7759), .A2(n7047), .ZN(n7761) );
  INV_X1 U9004 ( .A(n7750), .ZN(n7047) );
  XNOR2_X1 U9005 ( .A(n14427), .B(n14428), .ZN(n15630) );
  XNOR2_X1 U9006 ( .A(n14454), .B(n7327), .ZN(n14492) );
  INV_X1 U9007 ( .A(n14455), .ZN(n7327) );
  NAND2_X1 U9008 ( .A1(n14632), .A2(n14466), .ZN(n14635) );
  INV_X1 U9009 ( .A(n6907), .ZN(n14465) );
  NAND2_X1 U9010 ( .A1(n14635), .A2(n14636), .ZN(n14634) );
  NAND2_X1 U9011 ( .A1(n6864), .A2(n14643), .ZN(n14649) );
  NAND2_X1 U9012 ( .A1(n14649), .A2(n14648), .ZN(n14647) );
  NAND2_X1 U9013 ( .A1(n7259), .A2(n7262), .ZN(n10506) );
  OR2_X1 U9014 ( .A1(n12431), .A2(n12430), .ZN(n6888) );
  AOI21_X1 U9015 ( .B1(n12599), .B2(n12613), .A(n12582), .ZN(n12591) );
  NAND2_X1 U9016 ( .A1(n12617), .A2(n15084), .ZN(n6790) );
  OAI21_X1 U9017 ( .B1(n12626), .B2(n7025), .A(n6683), .ZN(n12115) );
  NAND2_X1 U9018 ( .A1(n7026), .A2(n15227), .ZN(n7025) );
  NAND2_X1 U9019 ( .A1(n6832), .A2(n12878), .ZN(n6830) );
  INV_X1 U9020 ( .A(n6885), .ZN(n6884) );
  NAND2_X1 U9021 ( .A1(n6832), .A2(n12946), .ZN(n6831) );
  NAND2_X1 U9022 ( .A1(n7371), .A2(n7374), .ZN(n7369) );
  XNOR2_X1 U9023 ( .A(n6931), .B(n13080), .ZN(n13084) );
  NAND2_X1 U9024 ( .A1(n13233), .A2(n10558), .ZN(n6886) );
  OR2_X1 U9025 ( .A1(n14970), .A2(n7220), .ZN(n7219) );
  INV_X1 U9026 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U9027 ( .A1(n6860), .A2(n6857), .ZN(P2_U3527) );
  INV_X1 U9028 ( .A(n6858), .ZN(n6857) );
  NAND2_X1 U9029 ( .A1(n13630), .A2(n14970), .ZN(n6860) );
  OAI21_X1 U9030 ( .B1(n13631), .B2(n13616), .A(n6859), .ZN(n6858) );
  OR2_X1 U9031 ( .A1(n14960), .A2(n11334), .ZN(n6874) );
  NAND2_X1 U9032 ( .A1(n6846), .A2(n6844), .ZN(P2_U3495) );
  AND2_X1 U9033 ( .A1(n6901), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U9034 ( .A1(n13630), .A2(n14960), .ZN(n6846) );
  NAND2_X1 U9035 ( .A1(n14959), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6845) );
  AND2_X1 U9036 ( .A1(n13809), .A2(n6810), .ZN(n6809) );
  INV_X1 U9037 ( .A(n6840), .ZN(n6839) );
  OAI22_X1 U9038 ( .A1(n14323), .A2(n14309), .B1(n14741), .B2(n14230), .ZN(
        n6840) );
  OAI21_X1 U9039 ( .B1(n14319), .B2(n14731), .A(n6852), .ZN(P1_U3525) );
  INV_X1 U9040 ( .A(n6853), .ZN(n6852) );
  OAI22_X1 U9041 ( .A1(n14321), .A2(n14354), .B1(n14733), .B2(n14320), .ZN(
        n6853) );
  INV_X1 U9042 ( .A(n6842), .ZN(n6841) );
  OAI22_X1 U9043 ( .A1(n14323), .A2(n14354), .B1(n14733), .B2(n15326), .ZN(
        n6842) );
  XNOR2_X1 U9044 ( .A(n14526), .B(n7348), .ZN(n7347) );
  XNOR2_X1 U9045 ( .A(n6788), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7348) );
  AND2_X1 U9046 ( .A1(n10336), .A2(n10329), .ZN(n6661) );
  AND2_X1 U9047 ( .A1(n7610), .A2(n9987), .ZN(n6662) );
  AND2_X1 U9048 ( .A1(n6697), .A2(n10257), .ZN(n6663) );
  NAND2_X1 U9049 ( .A1(n11429), .A2(n6963), .ZN(n11142) );
  OR2_X2 U9050 ( .A1(n13348), .A2(n13336), .ZN(n6664) );
  AND2_X1 U9051 ( .A1(n12713), .A2(n12392), .ZN(n6665) );
  AND2_X1 U9052 ( .A1(n11416), .A2(n10894), .ZN(n6666) );
  NOR2_X1 U9053 ( .A1(n13631), .A2(n13315), .ZN(n6667) );
  NAND2_X1 U9054 ( .A1(n12127), .A2(n6771), .ZN(n6668) );
  NOR2_X1 U9055 ( .A1(n14572), .A2(n14573), .ZN(n6669) );
  AND2_X1 U9056 ( .A1(n6696), .A2(n6949), .ZN(n6670) );
  NAND2_X1 U9057 ( .A1(n11501), .A2(n11500), .ZN(n14158) );
  AND2_X1 U9058 ( .A1(n13801), .A2(n7423), .ZN(n6671) );
  INV_X1 U9059 ( .A(n13832), .ZN(n7323) );
  AND2_X1 U9060 ( .A1(n7628), .A2(n14160), .ZN(n6672) );
  INV_X1 U9061 ( .A(n7474), .ZN(n7473) );
  AND2_X1 U9062 ( .A1(n6769), .A2(n7403), .ZN(n6673) );
  NAND2_X1 U9063 ( .A1(n11820), .A2(n11813), .ZN(n6674) );
  AND2_X1 U9064 ( .A1(n7378), .A2(n13101), .ZN(n6675) );
  OR2_X1 U9065 ( .A1(n6694), .A2(n7559), .ZN(n6676) );
  INV_X1 U9066 ( .A(n13336), .ZN(n13631) );
  INV_X1 U9067 ( .A(n13233), .ZN(n13625) );
  INV_X1 U9068 ( .A(n11799), .ZN(n7302) );
  NAND2_X1 U9069 ( .A1(n6772), .A2(n13040), .ZN(n6677) );
  AND2_X1 U9070 ( .A1(n11093), .A2(n11092), .ZN(n6678) );
  NAND2_X1 U9071 ( .A1(n7298), .A2(n7300), .ZN(n6679) );
  NAND2_X1 U9072 ( .A1(n12370), .A2(n12371), .ZN(n6680) );
  OR2_X1 U9073 ( .A1(n7370), .A2(n7377), .ZN(n6681) );
  OR2_X1 U9074 ( .A1(n13501), .A2(n7110), .ZN(n6682) );
  INV_X1 U9075 ( .A(n13142), .ZN(n13315) );
  INV_X1 U9076 ( .A(n12933), .ZN(n6832) );
  INV_X1 U9077 ( .A(n9183), .ZN(n7081) );
  INV_X1 U9078 ( .A(n14147), .ZN(n7628) );
  OR2_X1 U9079 ( .A1(n15227), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6683) );
  OR2_X1 U9080 ( .A1(n14741), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6684) );
  OR2_X1 U9081 ( .A1(n14053), .A2(n14045), .ZN(n6685) );
  AND2_X1 U9082 ( .A1(n11167), .A2(n11166), .ZN(n6686) );
  INV_X1 U9083 ( .A(n11925), .ZN(n7608) );
  INV_X1 U9084 ( .A(n13950), .ZN(n7637) );
  INV_X1 U9085 ( .A(n8275), .ZN(n14376) );
  XNOR2_X1 U9086 ( .A(n7968), .B(n7967), .ZN(n8275) );
  BUF_X1 U9087 ( .A(n13067), .Z(n13035) );
  NAND2_X1 U9088 ( .A1(n12164), .A2(n12439), .ZN(n6687) );
  AND2_X1 U9089 ( .A1(n7022), .A2(n12103), .ZN(n6688) );
  OR2_X1 U9090 ( .A1(n13333), .A2(n13332), .ZN(n6689) );
  OR2_X1 U9091 ( .A1(n13599), .A2(n13285), .ZN(n6690) );
  AND2_X1 U9093 ( .A1(n15113), .A2(n9363), .ZN(n6691) );
  AND2_X1 U9094 ( .A1(n6680), .A2(n12092), .ZN(n6692) );
  INV_X1 U9095 ( .A(n12102), .ZN(n7024) );
  AND2_X1 U9096 ( .A1(n11088), .A2(n11087), .ZN(n6693) );
  AND2_X1 U9097 ( .A1(n11115), .A2(n11114), .ZN(n6694) );
  NOR2_X1 U9098 ( .A1(n12098), .A2(n12097), .ZN(n6695) );
  OR2_X1 U9099 ( .A1(n11128), .A2(n11130), .ZN(n6696) );
  OR2_X1 U9100 ( .A1(n11787), .A2(n10859), .ZN(n6697) );
  AND2_X1 U9101 ( .A1(n7478), .A2(n7480), .ZN(n6698) );
  INV_X1 U9102 ( .A(n15156), .ZN(n9355) );
  AND2_X2 U9103 ( .A1(n9701), .A2(n7033), .ZN(n8753) );
  NAND2_X1 U9104 ( .A1(n11147), .A2(n11146), .ZN(n13599) );
  INV_X1 U9105 ( .A(n13599), .ZN(n7111) );
  OR2_X1 U9106 ( .A1(n12929), .A2(n12653), .ZN(n6699) );
  OR2_X1 U9107 ( .A1(n6678), .A2(n11097), .ZN(n6700) );
  AND2_X1 U9108 ( .A1(n7447), .A2(n8184), .ZN(n6701) );
  AND2_X1 U9109 ( .A1(n6671), .A2(n7088), .ZN(n6702) );
  AND2_X1 U9110 ( .A1(n6991), .A2(n6990), .ZN(n6703) );
  NAND2_X1 U9111 ( .A1(n10799), .A2(n10798), .ZN(n13910) );
  INV_X1 U9112 ( .A(n13910), .ZN(n14355) );
  INV_X1 U9113 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14380) );
  OR2_X1 U9114 ( .A1(n14332), .A2(n13999), .ZN(n6704) );
  INV_X1 U9115 ( .A(n12340), .ZN(n7150) );
  INV_X1 U9116 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7917) );
  INV_X1 U9117 ( .A(n9413), .ZN(n12275) );
  XNOR2_X1 U9118 ( .A(n8110), .B(n8109), .ZN(n9413) );
  OR2_X1 U9119 ( .A1(n13547), .A2(n13278), .ZN(n6705) );
  OR2_X1 U9120 ( .A1(n14337), .A2(n14076), .ZN(n6706) );
  INV_X1 U9121 ( .A(n13095), .ZN(n7361) );
  AND3_X1 U9122 ( .A1(n8841), .A2(n7322), .A3(n7321), .ZN(n9053) );
  INV_X1 U9123 ( .A(n9053), .ZN(n7320) );
  INV_X1 U9124 ( .A(n12693), .ZN(n6833) );
  AND2_X1 U9125 ( .A1(n11559), .A2(n11558), .ZN(n6707) );
  OR2_X1 U9126 ( .A1(n8025), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n6708) );
  AND4_X1 U9127 ( .A1(n7686), .A2(n7685), .A3(n8453), .A4(n8161), .ZN(n6709)
         );
  AND2_X1 U9128 ( .A1(n11066), .A2(n11065), .ZN(n6710) );
  AND2_X1 U9129 ( .A1(n14158), .A2(n14140), .ZN(n6711) );
  AND2_X1 U9130 ( .A1(n11023), .A2(n11022), .ZN(n6712) );
  INV_X1 U9131 ( .A(n14318), .ZN(n7129) );
  AND2_X1 U9132 ( .A1(n8327), .A2(n8243), .ZN(n6713) );
  OR2_X1 U9133 ( .A1(n11079), .A2(n11078), .ZN(n6714) );
  AND2_X1 U9134 ( .A1(n11547), .A2(n11546), .ZN(n14272) );
  AND2_X1 U9135 ( .A1(n13541), .A2(n13310), .ZN(n6715) );
  AND2_X1 U9136 ( .A1(n11235), .A2(n11234), .ZN(n6716) );
  AND2_X1 U9137 ( .A1(n14773), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U9138 ( .A1(n13028), .A2(n13029), .ZN(n6718) );
  AND2_X1 U9139 ( .A1(n6940), .A2(n7572), .ZN(n6719) );
  NOR2_X2 U9140 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8237) );
  INV_X1 U9141 ( .A(n7269), .ZN(n7268) );
  OR2_X1 U9142 ( .A1(n10293), .A2(n7270), .ZN(n7269) );
  NOR2_X1 U9143 ( .A1(n11194), .A2(n11195), .ZN(n6720) );
  OR2_X1 U9144 ( .A1(n7582), .A2(n11144), .ZN(n6721) );
  AND2_X1 U9145 ( .A1(n11094), .A2(n13149), .ZN(n6722) );
  AND3_X1 U9146 ( .A1(n7505), .A2(n7506), .A3(n7502), .ZN(n8125) );
  AND2_X1 U9147 ( .A1(n6701), .A2(n7718), .ZN(n6723) );
  AND2_X1 U9148 ( .A1(n7280), .A2(n7274), .ZN(n6724) );
  INV_X1 U9149 ( .A(n7408), .ZN(n7407) );
  NOR2_X1 U9150 ( .A1(n7111), .A2(n13286), .ZN(n7408) );
  INV_X1 U9151 ( .A(n7364), .ZN(n7363) );
  NOR2_X1 U9152 ( .A1(n6772), .A2(n7365), .ZN(n7364) );
  NOR2_X1 U9153 ( .A1(n11778), .A2(n14576), .ZN(n6725) );
  NOR2_X1 U9154 ( .A1(n11798), .A2(n14564), .ZN(n6726) );
  AND2_X1 U9155 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n6727) );
  INV_X1 U9156 ( .A(n7099), .ZN(n7098) );
  OAI21_X1 U9157 ( .B1(n13793), .B2(n7102), .A(n11526), .ZN(n7099) );
  INV_X1 U9158 ( .A(n11416), .ZN(n10904) );
  NAND2_X2 U9159 ( .A1(n11000), .A2(n8249), .ZN(n10321) );
  OR2_X1 U9160 ( .A1(n14385), .A2(n14384), .ZN(n6728) );
  INV_X1 U9161 ( .A(n11753), .ZN(n7325) );
  AND2_X1 U9162 ( .A1(n14181), .A2(n13912), .ZN(n6729) );
  INV_X1 U9163 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8242) );
  AND2_X1 U9164 ( .A1(n7564), .A2(n7571), .ZN(n6730) );
  NAND2_X1 U9165 ( .A1(n8341), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7871) );
  INV_X1 U9166 ( .A(n7624), .ZN(n7623) );
  OR2_X1 U9167 ( .A1(n13916), .A2(n7625), .ZN(n7624) );
  AND2_X1 U9168 ( .A1(n8801), .A2(n8800), .ZN(n6731) );
  AND2_X1 U9169 ( .A1(n10479), .A2(n10478), .ZN(n6732) );
  OR2_X1 U9170 ( .A1(n11873), .A2(n11874), .ZN(n6733) );
  NAND2_X1 U9171 ( .A1(n9096), .A2(n7447), .ZN(n6734) );
  NAND2_X1 U9172 ( .A1(n9096), .A2(n6701), .ZN(n6735) );
  INV_X1 U9173 ( .A(n13070), .ZN(n7377) );
  OAI21_X1 U9174 ( .B1(n7396), .B2(n7395), .A(n13375), .ZN(n7394) );
  NAND2_X1 U9175 ( .A1(n12371), .A2(n12767), .ZN(n6736) );
  AND2_X1 U9176 ( .A1(n7357), .A2(n6718), .ZN(n6737) );
  NAND2_X1 U9177 ( .A1(n7691), .A2(n7509), .ZN(n6738) );
  INV_X1 U9178 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n8606) );
  INV_X1 U9179 ( .A(n7011), .ZN(n7010) );
  NAND2_X1 U9180 ( .A1(n10216), .A2(n10475), .ZN(n7011) );
  NAND2_X1 U9181 ( .A1(n14379), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6739) );
  AND2_X1 U9182 ( .A1(n12328), .A2(n12332), .ZN(n12254) );
  INV_X1 U9183 ( .A(n7444), .ZN(n7442) );
  NOR2_X1 U9184 ( .A1(n10864), .A2(n7445), .ZN(n7444) );
  AND2_X1 U9185 ( .A1(n11611), .A2(n11610), .ZN(n6740) );
  AND2_X1 U9186 ( .A1(n11825), .A2(n13917), .ZN(n6741) );
  AND2_X1 U9187 ( .A1(n11665), .A2(n11664), .ZN(n6742) );
  NAND2_X1 U9188 ( .A1(n11943), .A2(n11946), .ZN(n6743) );
  INV_X1 U9189 ( .A(n11513), .ZN(n7102) );
  NAND2_X1 U9190 ( .A1(n7444), .A2(n7090), .ZN(n6744) );
  AND2_X1 U9191 ( .A1(n8518), .A2(n8515), .ZN(n6745) );
  OR2_X1 U9192 ( .A1(n9287), .A2(n7226), .ZN(n6746) );
  NAND2_X1 U9193 ( .A1(n6686), .A2(n11165), .ZN(n6747) );
  AND2_X1 U9194 ( .A1(n6971), .A2(n8645), .ZN(n6748) );
  OR2_X1 U9195 ( .A1(n12161), .A2(n12653), .ZN(n12107) );
  INV_X1 U9196 ( .A(n14133), .ZN(n14347) );
  AND2_X1 U9197 ( .A1(n7525), .A2(n13828), .ZN(n6749) );
  AND2_X1 U9198 ( .A1(n10688), .A2(n10686), .ZN(n6750) );
  NAND2_X1 U9199 ( .A1(n6687), .A2(n12094), .ZN(n6751) );
  NOR2_X1 U9200 ( .A1(n7578), .A2(n11129), .ZN(n6752) );
  INV_X1 U9201 ( .A(n7542), .ZN(n7541) );
  NAND2_X1 U9202 ( .A1(n14113), .A2(n13942), .ZN(n7542) );
  INV_X1 U9203 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8105) );
  INV_X1 U9204 ( .A(n12419), .ZN(n6869) );
  INV_X1 U9205 ( .A(n13923), .ZN(n14058) );
  INV_X1 U9206 ( .A(n13941), .ZN(n7627) );
  AND2_X1 U9207 ( .A1(n10519), .A2(n10520), .ZN(n6753) );
  AND2_X1 U9208 ( .A1(n12119), .A2(n12796), .ZN(n6754) );
  XNOR2_X1 U9209 ( .A(n13558), .B(n13271), .ZN(n13398) );
  INV_X1 U9210 ( .A(n12339), .ZN(n7152) );
  INV_X1 U9211 ( .A(n13312), .ZN(n7222) );
  XNOR2_X1 U9212 ( .A(n13534), .B(n13141), .ZN(n13312) );
  AND2_X1 U9213 ( .A1(n7379), .A2(n7378), .ZN(n6755) );
  AND2_X1 U9214 ( .A1(n7359), .A2(n7356), .ZN(n6756) );
  AND2_X1 U9215 ( .A1(n10730), .A2(n10728), .ZN(n6757) );
  NOR2_X1 U9216 ( .A1(n12833), .A2(n7150), .ZN(n7149) );
  AND2_X1 U9217 ( .A1(n6911), .A2(n12615), .ZN(n6758) );
  AND2_X1 U9218 ( .A1(n7093), .A2(n7435), .ZN(n6759) );
  AND2_X1 U9219 ( .A1(n7086), .A2(n7421), .ZN(n6760) );
  AND2_X1 U9220 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n6761) );
  OR2_X1 U9221 ( .A1(n11790), .A2(n11788), .ZN(n6762) );
  AND2_X1 U9222 ( .A1(n11082), .A2(n11081), .ZN(n6763) );
  NAND2_X1 U9223 ( .A1(n13534), .A2(n14927), .ZN(n6764) );
  AND2_X1 U9224 ( .A1(n7371), .A2(n6681), .ZN(n6765) );
  INV_X1 U9225 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U9226 ( .A1(n7344), .A2(n11777), .ZN(n6766) );
  NAND2_X1 U9227 ( .A1(n11763), .A2(n7317), .ZN(n6767) );
  AND2_X1 U9228 ( .A1(n6750), .A2(n6934), .ZN(n6768) );
  INV_X1 U9229 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9230 ( .A1(n12129), .A2(n12679), .ZN(n7292) );
  INV_X1 U9231 ( .A(n11413), .ZN(n10379) );
  INV_X1 U9232 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U9233 ( .A1(n7300), .A2(n11793), .ZN(n7297) );
  INV_X1 U9234 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8652) );
  INV_X1 U9235 ( .A(n13379), .ZN(n7112) );
  INV_X1 U9236 ( .A(SI_1_), .ZN(n7455) );
  OR2_X1 U9237 ( .A1(n13588), .A2(n13291), .ZN(n6769) );
  INV_X1 U9238 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7457) );
  AND2_X1 U9239 ( .A1(n14800), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6770) );
  XOR2_X1 U9240 ( .A(n12945), .B(n12117), .Z(n6771) );
  INV_X1 U9241 ( .A(n12439), .ZN(n12752) );
  XOR2_X1 U9242 ( .A(n13568), .B(n13067), .Z(n6772) );
  INV_X1 U9243 ( .A(n15088), .ZN(n10145) );
  NOR2_X1 U9244 ( .A1(n10662), .A2(n10663), .ZN(n10861) );
  OR3_X1 U9245 ( .A1(n13501), .A2(n7110), .A3(n13588), .ZN(n6773) );
  AND4_X1 U9246 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n12825) );
  INV_X1 U9247 ( .A(n12825), .ZN(n6815) );
  INV_X1 U9248 ( .A(n6806), .ZN(n14600) );
  AND2_X1 U9249 ( .A1(n7151), .A2(n12340), .ZN(n6774) );
  INV_X1 U9250 ( .A(n6905), .ZN(n10368) );
  INV_X1 U9251 ( .A(n7404), .ZN(n7403) );
  NOR2_X1 U9252 ( .A1(n13287), .A2(n7408), .ZN(n7404) );
  AND2_X1 U9253 ( .A1(n12774), .A2(n12092), .ZN(n6775) );
  INV_X1 U9254 ( .A(n7446), .ZN(n14571) );
  NAND2_X1 U9255 ( .A1(n7443), .A2(n6669), .ZN(n7446) );
  AND2_X1 U9256 ( .A1(n9733), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6776) );
  INV_X1 U9257 ( .A(n13102), .ZN(n6938) );
  AND2_X1 U9258 ( .A1(n9585), .A2(n11977), .ZN(n6777) );
  OR2_X1 U9259 ( .A1(n10148), .A2(n10486), .ZN(n6778) );
  OR2_X1 U9260 ( .A1(n10178), .A2(n10541), .ZN(n6779) );
  INV_X1 U9261 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7775) );
  XNOR2_X1 U9262 ( .A(n11778), .B(n10654), .ZN(n10243) );
  INV_X1 U9263 ( .A(n10243), .ZN(n7600) );
  INV_X1 U9264 ( .A(n9921), .ZN(n6935) );
  INV_X1 U9265 ( .A(n11107), .ZN(n7105) );
  AND2_X1 U9266 ( .A1(n9361), .A2(n9360), .ZN(n6780) );
  NAND2_X1 U9267 ( .A1(n11216), .A2(n11215), .ZN(n13568) );
  INV_X1 U9268 ( .A(n13568), .ZN(n7116) );
  AND2_X1 U9269 ( .A1(n9504), .A2(n9503), .ZN(n6781) );
  AND2_X1 U9270 ( .A1(n7159), .A2(n10735), .ZN(n6782) );
  AND2_X1 U9271 ( .A1(n7549), .A2(n7550), .ZN(n6783) );
  AND2_X2 U9272 ( .A1(n9305), .A2(n9304), .ZN(n14960) );
  INV_X1 U9273 ( .A(n13662), .ZN(n6902) );
  AND2_X1 U9274 ( .A1(n9210), .A2(n8221), .ZN(n13798) );
  AND2_X2 U9275 ( .A1(n9305), .A2(n8596), .ZN(n14970) );
  INV_X1 U9276 ( .A(n14715), .ZN(n7525) );
  AND2_X2 U9277 ( .A1(n8688), .A2(n8687), .ZN(n14741) );
  INV_X1 U9278 ( .A(n13518), .ZN(n7107) );
  NAND2_X1 U9279 ( .A1(n11429), .A2(n6640), .ZN(n6784) );
  INV_X1 U9280 ( .A(n9701), .ZN(n12422) );
  NAND2_X1 U9281 ( .A1(n12601), .A2(n9273), .ZN(n9701) );
  AND2_X1 U9282 ( .A1(n9229), .A2(n7253), .ZN(n6785) );
  INV_X1 U9283 ( .A(n12524), .ZN(n7171) );
  OR2_X1 U9284 ( .A1(n8839), .A2(n14358), .ZN(n6786) );
  NAND2_X1 U9285 ( .A1(n11962), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6787) );
  AND2_X1 U9286 ( .A1(n8587), .A2(n8586), .ZN(n13435) );
  INV_X1 U9287 ( .A(n13435), .ZN(n13499) );
  XOR2_X1 U9288 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n6788) );
  INV_X1 U9289 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7735) );
  INV_X1 U9290 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6909) );
  INV_X1 U9291 ( .A(n14552), .ZN(n13133) );
  NAND2_X1 U9292 ( .A1(n11745), .A2(n11744), .ZN(n6796) );
  OAI21_X1 U9293 ( .B1(n11724), .B2(n11723), .A(n11722), .ZN(n11732) );
  NAND2_X1 U9294 ( .A1(n14517), .A2(n14516), .ZN(n14515) );
  INV_X1 U9295 ( .A(n12607), .ZN(n6789) );
  NAND3_X1 U9296 ( .A1(n6900), .A2(n6790), .A3(n6758), .ZN(P3_U3201) );
  NAND2_X1 U9297 ( .A1(n12503), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12528) );
  XNOR2_X1 U9298 ( .A(n12526), .B(n12536), .ZN(n12503) );
  NAND2_X1 U9299 ( .A1(n15094), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15093) );
  NAND2_X1 U9300 ( .A1(n15038), .A2(n15037), .ZN(n15036) );
  NAND2_X1 U9301 ( .A1(n15073), .A2(n15072), .ZN(n15071) );
  NAND2_X1 U9302 ( .A1(n12810), .A2(n12811), .ZN(n12809) );
  OAI21_X1 U9303 ( .B1(n12755), .B2(n7137), .A(n7134), .ZN(n12731) );
  NAND2_X1 U9304 ( .A1(n6665), .A2(n6833), .ZN(n12694) );
  OAI22_X1 U9305 ( .A1(n12243), .A2(n12267), .B1(n12921), .B2(n6869), .ZN(
        n12244) );
  NAND2_X1 U9306 ( .A1(n10194), .A2(n12299), .ZN(n15102) );
  NAND2_X1 U9307 ( .A1(n7130), .A2(n12284), .ZN(n9500) );
  NAND2_X1 U9308 ( .A1(n10214), .A2(n12306), .ZN(n10476) );
  NAND2_X1 U9309 ( .A1(n6804), .A2(n12399), .ZN(n12664) );
  NAND2_X2 U9310 ( .A1(n7863), .A2(n7862), .ZN(n7920) );
  XNOR2_X1 U9311 ( .A(n6791), .B(n11168), .ZN(n11426) );
  NAND4_X1 U9312 ( .A1(n11423), .A2(n11424), .A3(n13312), .A4(n11438), .ZN(
        n6791) );
  NOR2_X1 U9313 ( .A1(n7653), .A2(n7477), .ZN(n11461) );
  NAND2_X1 U9314 ( .A1(n7050), .A2(n7051), .ZN(n9081) );
  INV_X1 U9315 ( .A(n7743), .ZN(n6792) );
  NAND2_X1 U9316 ( .A1(n7449), .A2(n6894), .ZN(n7743) );
  OAI21_X2 U9317 ( .B1(n6920), .B2(n7394), .A(n13307), .ZN(n13358) );
  NAND2_X1 U9318 ( .A1(n9561), .A2(n9560), .ZN(n9292) );
  NAND3_X1 U9319 ( .A1(n9560), .A2(n8585), .A3(n8584), .ZN(n9561) );
  NAND2_X1 U9320 ( .A1(n9463), .A2(n9297), .ZN(n9478) );
  NAND2_X1 U9321 ( .A1(n6793), .A2(n11412), .ZN(n10723) );
  NAND2_X1 U9322 ( .A1(n10057), .A2(n9295), .ZN(n9465) );
  OR2_X2 U9323 ( .A1(n13532), .A2(n6925), .ZN(n13629) );
  OAI21_X1 U9324 ( .B1(n13497), .B2(n7400), .A(n7398), .ZN(n13294) );
  NAND2_X1 U9325 ( .A1(n10720), .A2(n10717), .ZN(n6793) );
  XNOR2_X2 U9326 ( .A(n8170), .B(n14356), .ZN(n8172) );
  NAND2_X1 U9327 ( .A1(n9294), .A2(n9293), .ZN(n10057) );
  NAND3_X1 U9328 ( .A1(n6796), .A2(n11750), .A3(n6794), .ZN(n7324) );
  NOR2_X4 U9329 ( .A1(n7416), .A2(n7905), .ZN(n8011) );
  NOR2_X1 U9330 ( .A1(n14523), .A2(n14522), .ZN(n14525) );
  NAND2_X1 U9331 ( .A1(n6819), .A2(n14515), .ZN(n14523) );
  NAND2_X1 U9332 ( .A1(n7118), .A2(n7119), .ZN(n6925) );
  NAND2_X2 U9333 ( .A1(n9285), .A2(n9284), .ZN(n9462) );
  NAND2_X1 U9334 ( .A1(n13334), .A2(n7044), .ZN(n7041) );
  OR2_X2 U9335 ( .A1(n9670), .A2(n11407), .ZN(n9687) );
  NAND2_X1 U9336 ( .A1(n14471), .A2(n14470), .ZN(n14641) );
  NAND2_X1 U9337 ( .A1(n11842), .A2(n11843), .ZN(n11847) );
  NAND2_X1 U9338 ( .A1(n7328), .A2(n7329), .ZN(n11842) );
  NAND2_X1 U9339 ( .A1(n7162), .A2(n15217), .ZN(n7161) );
  NAND2_X1 U9340 ( .A1(n7199), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U9341 ( .A1(n7771), .A2(n7770), .ZN(n7789) );
  NAND2_X1 U9342 ( .A1(n7839), .A2(n7838), .ZN(n7867) );
  NAND2_X1 U9343 ( .A1(n7778), .A2(n7777), .ZN(n7801) );
  OAI21_X1 U9344 ( .B1(n11796), .B2(n7297), .A(n6679), .ZN(n6879) );
  NAND2_X1 U9345 ( .A1(n7200), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7199) );
  OAI21_X1 U9346 ( .B1(n12421), .B2(n12423), .A(n6824), .ZN(n6868) );
  INV_X1 U9347 ( .A(n14441), .ZN(n7313) );
  XNOR2_X1 U9348 ( .A(n12310), .B(n12117), .ZN(n10163) );
  NOR2_X1 U9349 ( .A1(n7248), .A2(n7247), .ZN(n12118) );
  NAND2_X2 U9350 ( .A1(n10270), .A2(n7737), .ZN(n11984) );
  NAND2_X1 U9351 ( .A1(n12678), .A2(n12684), .ZN(n6804) );
  NAND2_X1 U9352 ( .A1(n15125), .A2(n9350), .ZN(n6805) );
  NAND2_X1 U9353 ( .A1(n14065), .A2(n14337), .ZN(n14053) );
  OAI21_X1 U9354 ( .B1(n12799), .B2(n7142), .A(n7141), .ZN(n11980) );
  NAND2_X1 U9355 ( .A1(n14319), .A2(n14741), .ZN(n7513) );
  NAND2_X1 U9356 ( .A1(n7513), .A2(n6684), .ZN(n14223) );
  NAND2_X4 U9357 ( .A1(n7453), .A2(n7454), .ZN(n7737) );
  NAND2_X1 U9358 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  NAND2_X1 U9359 ( .A1(n10745), .A2(n10744), .ZN(n10747) );
  NAND2_X1 U9360 ( .A1(n11349), .A2(n7651), .ZN(n11355) );
  NOR2_X2 U9361 ( .A1(n7740), .A2(n8209), .ZN(n7741) );
  OR2_X1 U9362 ( .A1(n7958), .A2(n7957), .ZN(n7959) );
  NAND2_X2 U9363 ( .A1(n9123), .A2(n9122), .ZN(n11083) );
  NAND2_X1 U9364 ( .A1(n6811), .A2(n6809), .ZN(P1_U3240) );
  NAND2_X1 U9365 ( .A1(n13803), .A2(n14567), .ZN(n6811) );
  INV_X1 U9366 ( .A(n7420), .ZN(n7418) );
  NAND2_X2 U9367 ( .A1(n7425), .A2(n7426), .ZN(n13754) );
  NAND2_X1 U9368 ( .A1(n9525), .A2(n9524), .ZN(n9796) );
  NAND2_X1 U9369 ( .A1(n13811), .A2(n13812), .ZN(n13810) );
  NAND2_X1 U9370 ( .A1(n11571), .A2(n11570), .ZN(n13720) );
  NOR2_X1 U9371 ( .A1(n9799), .A2(n9800), .ZN(n10518) );
  NAND2_X1 U9372 ( .A1(n8660), .A2(n8628), .ZN(n8629) );
  OAI21_X1 U9373 ( .B1(n13747), .B2(n7095), .A(n6759), .ZN(n13722) );
  NAND2_X2 U9374 ( .A1(n13704), .A2(n6865), .ZN(n13705) );
  NAND4_X2 U9375 ( .A1(n15447), .A2(n7736), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U9376 ( .A1(n9380), .A2(n9397), .ZN(n9744) );
  OAI21_X2 U9377 ( .B1(n12198), .B2(n12714), .A(n6813), .ZN(n12127) );
  XNOR2_X2 U9378 ( .A(n12124), .B(n7255), .ZN(n12198) );
  NAND2_X1 U9379 ( .A1(n7279), .A2(n7278), .ZN(n12154) );
  INV_X1 U9380 ( .A(n7198), .ZN(n7197) );
  NAND2_X1 U9381 ( .A1(n7261), .A2(n6848), .ZN(n10568) );
  NAND2_X1 U9382 ( .A1(n8661), .A2(n8662), .ZN(n8660) );
  NAND2_X1 U9383 ( .A1(n7087), .A2(n11633), .ZN(n13731) );
  NAND2_X1 U9384 ( .A1(n11497), .A2(n11496), .ZN(n13747) );
  XNOR2_X1 U9385 ( .A(n14440), .B(n7313), .ZN(n15621) );
  NOR2_X2 U9386 ( .A1(n14497), .A2(n14498), .ZN(n14496) );
  NOR2_X2 U9387 ( .A1(n14493), .A2(n14459), .ZN(n14497) );
  XNOR2_X1 U9388 ( .A(n10146), .B(n10145), .ZN(n15079) );
  NOR2_X2 U9389 ( .A1(n12521), .A2(n12520), .ZN(n12525) );
  NAND2_X4 U9390 ( .A1(n10321), .A2(n7737), .ZN(n11363) );
  NAND3_X2 U9391 ( .A1(n7674), .A2(n8011), .A3(n7553), .ZN(n8327) );
  INV_X1 U9392 ( .A(n7505), .ZN(n8025) );
  AND2_X1 U9393 ( .A1(n7505), .A2(n6709), .ZN(n8490) );
  NAND2_X1 U9394 ( .A1(n12290), .A2(n6890), .ZN(n12298) );
  NAND2_X1 U9395 ( .A1(n6893), .A2(n6892), .ZN(n12280) );
  INV_X1 U9396 ( .A(n11860), .ZN(n11863) );
  NAND2_X1 U9397 ( .A1(n11859), .A2(n11857), .ZN(n6825) );
  INV_X1 U9398 ( .A(n11842), .ZN(n11845) );
  NAND2_X1 U9399 ( .A1(n6761), .A2(n7737), .ZN(n7451) );
  NAND2_X1 U9400 ( .A1(n11834), .A2(n11833), .ZN(n6881) );
  NAND3_X1 U9401 ( .A1(n7456), .A2(n7455), .A3(n7452), .ZN(n6894) );
  NOR2_X1 U9402 ( .A1(n12596), .A2(n12595), .ZN(n12597) );
  NAND2_X1 U9403 ( .A1(n12860), .A2(n6830), .ZN(P3_U3486) );
  NAND2_X1 U9404 ( .A1(n12932), .A2(n6831), .ZN(P3_U3454) );
  NOR2_X2 U9405 ( .A1(n15044), .A2(n10207), .ZN(n15043) );
  NAND2_X1 U9406 ( .A1(n10132), .A2(n6923), .ZN(n14972) );
  NAND2_X1 U9407 ( .A1(n9465), .A2(n9464), .ZN(n9463) );
  NAND2_X1 U9408 ( .A1(n6856), .A2(n11027), .ZN(n9108) );
  NOR2_X2 U9409 ( .A1(n9021), .A2(n6837), .ZN(n7384) );
  NAND2_X1 U9410 ( .A1(n6871), .A2(n6661), .ZN(n6933) );
  OAI21_X2 U9411 ( .B1(n8346), .B2(n8606), .A(n6838), .ZN(n7747) );
  XNOR2_X1 U9412 ( .A(n14715), .B(n9986), .ZN(n11924) );
  OAI21_X1 U9413 ( .B1(n14322), .B2(n14739), .A(n6839), .ZN(P1_U3556) );
  OAI21_X1 U9414 ( .B1(n14322), .B2(n14731), .A(n6841), .ZN(P1_U3524) );
  INV_X1 U9415 ( .A(n13159), .ZN(n6856) );
  XNOR2_X1 U9416 ( .A(n9296), .B(n14926), .ZN(n11402) );
  NAND2_X1 U9417 ( .A1(n7505), .A2(n7504), .ZN(n7696) );
  INV_X1 U9418 ( .A(n7271), .ZN(n7266) );
  XNOR2_X1 U9419 ( .A(n6919), .B(n6918), .ZN(n12215) );
  NAND2_X1 U9420 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  OAI21_X1 U9421 ( .B1(n7652), .B2(n11454), .A(n11453), .ZN(n7481) );
  AOI21_X1 U9422 ( .B1(n7473), .B2(n7475), .A(n7472), .ZN(n7471) );
  NAND2_X1 U9423 ( .A1(n9940), .A2(n9939), .ZN(n10314) );
  NAND3_X1 U9424 ( .A1(n7640), .A2(n7639), .A3(n7638), .ZN(n14216) );
  OAI211_X1 U9425 ( .C1(n10751), .C2(n7466), .A(n10996), .B(n7464), .ZN(n10995) );
  NOR2_X1 U9426 ( .A1(n14221), .A2(n14220), .ZN(n7516) );
  NOR2_X4 U9427 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7902) );
  AND3_X2 U9428 ( .A1(n7894), .A2(n6855), .A3(n6854), .ZN(n6953) );
  INV_X1 U9429 ( .A(n9108), .ZN(n8585) );
  OAI21_X2 U9430 ( .B1(n10895), .B2(n7239), .A(n7237), .ZN(n13253) );
  NAND2_X1 U9431 ( .A1(n6904), .A2(n6903), .ZN(n13487) );
  NAND2_X1 U9432 ( .A1(n10382), .A2(n10381), .ZN(n10641) );
  NOR2_X1 U9433 ( .A1(n15624), .A2(n15623), .ZN(n15622) );
  AOI21_X2 U9434 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n14460), .A(n14496), .ZN(
        n14630) );
  NOR2_X2 U9435 ( .A1(n14490), .A2(n14489), .ZN(n14488) );
  NAND2_X1 U9436 ( .A1(n15621), .A2(n15620), .ZN(n15619) );
  NAND2_X1 U9437 ( .A1(n6897), .A2(n14634), .ZN(n14467) );
  NOR2_X1 U9438 ( .A1(n15630), .A2(n15631), .ZN(n15629) );
  INV_X1 U9439 ( .A(n9908), .ZN(n6871) );
  OAI22_X2 U9440 ( .A1(n13075), .A2(n13074), .B1(n13019), .B2(n13018), .ZN(
        n13020) );
  NAND2_X1 U9441 ( .A1(n8736), .A2(n7351), .ZN(n8772) );
  NAND3_X1 U9442 ( .A1(n7079), .A2(n7071), .A3(n13705), .ZN(n7070) );
  XNOR2_X1 U9443 ( .A(n11485), .B(n11483), .ZN(n13811) );
  NAND2_X1 U9444 ( .A1(n13731), .A2(n13730), .ZN(n7422) );
  NOR2_X1 U9445 ( .A1(n8627), .A2(n8626), .ZN(n8662) );
  NAND2_X1 U9446 ( .A1(n8989), .A2(n8988), .ZN(n9272) );
  OAI21_X1 U9447 ( .B1(n12270), .B2(n12269), .A(n6868), .ZN(n6867) );
  INV_X1 U9448 ( .A(n11963), .ZN(n6870) );
  NAND2_X1 U9449 ( .A1(n6870), .A2(n6787), .ZN(n11965) );
  NAND2_X1 U9450 ( .A1(n8986), .A2(n8985), .ZN(n8989) );
  XNOR2_X2 U9451 ( .A(n8651), .B(n8650), .ZN(n10245) );
  INV_X1 U9452 ( .A(n13722), .ZN(n11571) );
  NAND2_X1 U9453 ( .A1(n8629), .A2(n8630), .ZN(n13704) );
  NAND2_X1 U9454 ( .A1(n7422), .A2(n11650), .ZN(n13802) );
  NAND4_X2 U9455 ( .A1(n8177), .A2(n8178), .A3(n8179), .A4(n8180), .ZN(n14192)
         );
  NAND2_X1 U9456 ( .A1(n13770), .A2(n13771), .ZN(n14560) );
  OR2_X1 U9457 ( .A1(n11333), .A2(n8348), .ZN(n8351) );
  NAND2_X1 U9458 ( .A1(n13629), .A2(n14960), .ZN(n6875) );
  NAND2_X1 U9459 ( .A1(n8731), .A2(n8730), .ZN(n6877) );
  INV_X1 U9460 ( .A(n13485), .ZN(n6904) );
  NAND3_X1 U9461 ( .A1(n7215), .A2(n7214), .A3(n11410), .ZN(n10352) );
  OAI21_X2 U9462 ( .B1(n13270), .B2(n7241), .A(n7240), .ZN(n13276) );
  NOR2_X1 U9463 ( .A1(n15008), .A2(n15009), .ZN(n15007) );
  NAND2_X1 U9464 ( .A1(n10316), .A2(n6873), .ZN(n10546) );
  NOR2_X1 U9465 ( .A1(n10146), .A2(n10145), .ZN(n10147) );
  NOR2_X2 U9466 ( .A1(n12500), .A2(n12501), .ZN(n12520) );
  NAND2_X1 U9467 ( .A1(n12694), .A2(n12390), .ZN(n12678) );
  NAND2_X1 U9468 ( .A1(n7146), .A2(n7147), .ZN(n12827) );
  OAI21_X2 U9469 ( .B1(n10531), .B2(n12318), .A(n12320), .ZN(n10734) );
  NAND2_X1 U9470 ( .A1(n6875), .A2(n6874), .ZN(P2_U3496) );
  OAI22_X1 U9471 ( .A1(n9694), .A2(n9693), .B1(n14945), .B2(n13150), .ZN(n9695) );
  NOR2_X1 U9472 ( .A1(n6878), .A2(n6877), .ZN(n6876) );
  NAND4_X1 U9473 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n13159)
         );
  INV_X1 U9474 ( .A(n6879), .ZN(n7295) );
  AOI21_X1 U9475 ( .B1(n11831), .B2(n11830), .A(n6914), .ZN(n11834) );
  NAND2_X1 U9476 ( .A1(n11835), .A2(n6881), .ZN(n11837) );
  NAND2_X1 U9477 ( .A1(n11845), .A2(n11844), .ZN(n6882) );
  NAND2_X1 U9478 ( .A1(n11847), .A2(n11846), .ZN(n6883) );
  OAI21_X1 U9479 ( .B1(n11859), .B2(n11857), .A(n11856), .ZN(n11858) );
  NAND2_X1 U9480 ( .A1(n11875), .A2(n7309), .ZN(n7307) );
  NAND2_X1 U9481 ( .A1(n11869), .A2(n6880), .ZN(n11875) );
  INV_X1 U9482 ( .A(n8020), .ZN(n7200) );
  NAND2_X1 U9483 ( .A1(n8877), .A2(n8876), .ZN(n8986) );
  NAND2_X1 U9484 ( .A1(n7936), .A2(n7935), .ZN(n8019) );
  OAI21_X1 U9485 ( .B1(n7161), .B2(n12625), .A(n6884), .ZN(n12116) );
  NAND3_X1 U9486 ( .A1(n11773), .A2(n11772), .A3(n6766), .ZN(n7343) );
  OR2_X2 U9487 ( .A1(n10470), .A2(n11237), .ZN(n7211) );
  NAND2_X1 U9488 ( .A1(n13527), .A2(n6886), .ZN(P2_U3530) );
  INV_X2 U9489 ( .A(n11056), .ZN(n14921) );
  OR2_X4 U9490 ( .A1(n10913), .A2(n13603), .ZN(n13501) );
  NOR2_X2 U9491 ( .A1(n6664), .A2(n13534), .ZN(n13317) );
  OR2_X1 U9492 ( .A1(n9482), .A2(n11068), .ZN(n9484) );
  NOR2_X2 U9493 ( .A1(n13377), .A2(n13547), .ZN(n13361) );
  NAND2_X1 U9494 ( .A1(n14645), .A2(n14644), .ZN(n14643) );
  NAND2_X2 U9495 ( .A1(n13720), .A2(n11575), .ZN(n13783) );
  NAND3_X1 U9496 ( .A1(n12347), .A2(n12346), .A3(n12826), .ZN(n12353) );
  NOR2_X1 U9497 ( .A1(n7938), .A2(n7683), .ZN(n7684) );
  OAI21_X1 U9498 ( .B1(n12433), .B2(n12432), .A(n6888), .ZN(P3_U3296) );
  INV_X1 U9499 ( .A(n7694), .ZN(n7692) );
  NAND2_X1 U9500 ( .A1(n7520), .A2(n7521), .ZN(n7518) );
  OR2_X1 U9501 ( .A1(n9310), .A2(n11612), .ZN(n9313) );
  INV_X1 U9502 ( .A(n11922), .ZN(n7517) );
  OAI22_X2 U9503 ( .A1(n13980), .A2(n13983), .B1(n14327), .B2(n14000), .ZN(
        n13966) );
  NAND2_X1 U9504 ( .A1(n14641), .A2(n14642), .ZN(n14638) );
  NAND2_X1 U9505 ( .A1(n6924), .A2(n12588), .ZN(n6900) );
  NAND2_X2 U9506 ( .A1(n13487), .A2(n13255), .ZN(n13468) );
  NAND2_X1 U9507 ( .A1(n13537), .A2(n6921), .ZN(n13630) );
  OAI21_X1 U9508 ( .B1(n13538), .B2(n14931), .A(n13536), .ZN(n6922) );
  NAND2_X1 U9509 ( .A1(n7193), .A2(n7191), .ZN(n8877) );
  NAND2_X1 U9510 ( .A1(n7187), .A2(n7185), .ZN(n7936) );
  INV_X1 U9511 ( .A(n9410), .ZN(n7210) );
  NAND2_X1 U9512 ( .A1(n10368), .A2(n7414), .ZN(n10720) );
  NAND2_X1 U9513 ( .A1(n13629), .A2(n14970), .ZN(n7221) );
  NAND2_X1 U9514 ( .A1(n7412), .A2(n13499), .ZN(n7411) );
  NAND2_X1 U9515 ( .A1(n10723), .A2(n10628), .ZN(n10834) );
  OR2_X1 U9516 ( .A1(n13156), .A2(n14916), .ZN(n10054) );
  NAND2_X1 U9517 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NAND2_X1 U9518 ( .A1(n13327), .A2(n13311), .ZN(n7413) );
  XNOR2_X1 U9519 ( .A(n7413), .B(n7222), .ZN(n7412) );
  NOR2_X1 U9520 ( .A1(n10356), .A2(n10379), .ZN(n6905) );
  NAND2_X1 U9521 ( .A1(n10054), .A2(n9279), .ZN(n9559) );
  NAND2_X1 U9522 ( .A1(n7548), .A2(n7549), .ZN(n10777) );
  AOI22_X2 U9523 ( .A1(n13997), .A2(n13996), .B1(n14021), .B2(n14236), .ZN(
        n13980) );
  NAND2_X1 U9524 ( .A1(n7221), .A2(n7219), .ZN(P2_U3528) );
  XNOR2_X1 U9525 ( .A(n7515), .B(n7637), .ZN(n14222) );
  OAI21_X1 U9526 ( .B1(n14525), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n14524), .ZN(
        n7349) );
  NAND2_X1 U9527 ( .A1(n7596), .A2(n10243), .ZN(n7597) );
  NAND2_X1 U9528 ( .A1(n7607), .A2(n7609), .ZN(n6908) );
  NAND2_X1 U9529 ( .A1(n13929), .A2(n13928), .ZN(n13981) );
  OAI21_X2 U9530 ( .B1(n10823), .B2(n7616), .A(n7614), .ZN(n14604) );
  NAND2_X1 U9531 ( .A1(n7622), .A2(n7619), .ZN(n13918) );
  NAND2_X1 U9532 ( .A1(n7954), .A2(n7953), .ZN(n7958) );
  INV_X1 U9533 ( .A(n14112), .ZN(n6973) );
  NAND2_X1 U9534 ( .A1(n11924), .A2(n7611), .ZN(n7610) );
  NOR2_X1 U9535 ( .A1(n14435), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n14382) );
  XNOR2_X1 U9536 ( .A(n14447), .B(n14448), .ZN(n15624) );
  NOR2_X2 U9537 ( .A1(n14488), .A2(n14446), .ZN(n14447) );
  NAND2_X1 U9538 ( .A1(n14463), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7304) );
  NOR2_X1 U9539 ( .A1(n14495), .A2(n14494), .ZN(n14493) );
  NAND2_X1 U9540 ( .A1(n9092), .A2(n9091), .ZN(n9174) );
  INV_X1 U9541 ( .A(n9439), .ZN(n6915) );
  NAND2_X1 U9542 ( .A1(n7343), .A2(n7342), .ZN(n11781) );
  NAND2_X1 U9543 ( .A1(n7316), .A2(n7315), .ZN(n11768) );
  NAND2_X1 U9544 ( .A1(n6912), .A2(n15095), .ZN(n6911) );
  XNOR2_X1 U9545 ( .A(n12609), .B(n12608), .ZN(n6912) );
  OAI21_X1 U9546 ( .B1(n7456), .B2(n7455), .A(n7451), .ZN(n7450) );
  NAND3_X1 U9547 ( .A1(n9153), .A2(n9089), .A3(n9087), .ZN(n9092) );
  NAND2_X1 U9548 ( .A1(n9081), .A2(n9080), .ZN(n9085) );
  NAND2_X1 U9549 ( .A1(n12165), .A2(n7256), .ZN(n12124) );
  INV_X1 U9550 ( .A(n10970), .ZN(n7248) );
  OAI21_X1 U9551 ( .B1(n7252), .B2(n9045), .A(n7250), .ZN(n9420) );
  NAND2_X1 U9552 ( .A1(n7172), .A2(n7171), .ZN(n12565) );
  NOR2_X1 U9553 ( .A1(n14972), .A2(n10088), .ZN(n14971) );
  OR2_X1 U9554 ( .A1(n10133), .A2(n14979), .ZN(n6923) );
  XNOR2_X1 U9555 ( .A(n12597), .B(n12602), .ZN(n6924) );
  NOR2_X1 U9556 ( .A1(n15007), .A2(n10139), .ZN(n15027) );
  NAND2_X1 U9557 ( .A1(n10836), .A2(n10835), .ZN(n10901) );
  NAND2_X1 U9558 ( .A1(n13297), .A2(n13296), .ZN(n7417) );
  NAND2_X1 U9559 ( .A1(n7510), .A2(n11804), .ZN(n13935) );
  NAND2_X1 U9560 ( .A1(n14506), .A2(n10784), .ZN(n14589) );
  NAND2_X1 U9561 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  NAND2_X2 U9562 ( .A1(n14073), .A2(n13946), .ZN(n14049) );
  OAI21_X2 U9563 ( .B1(n9825), .B2(n9635), .A(n9637), .ZN(n9968) );
  OAI22_X1 U9564 ( .A1(n13966), .A2(n13949), .B1(n14219), .B2(n13974), .ZN(
        n7515) );
  NAND3_X2 U9565 ( .A1(n6927), .A2(n8204), .A3(n8206), .ZN(n14195) );
  NAND2_X1 U9566 ( .A1(n7490), .A2(n9437), .ZN(n9583) );
  OAI21_X1 U9567 ( .B1(n7475), .B2(n8031), .A(n8531), .ZN(n7474) );
  NAND2_X1 U9568 ( .A1(n12167), .A2(n12166), .ZN(n12165) );
  NAND2_X1 U9569 ( .A1(n7028), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U9570 ( .A1(n14633), .A2(n15507), .ZN(n14632) );
  INV_X1 U9571 ( .A(n14628), .ZN(n7305) );
  XNOR2_X1 U9572 ( .A(n7349), .B(n7347), .ZN(SUB_1596_U4) );
  NAND2_X4 U9573 ( .A1(n14949), .A2(n11390), .ZN(n13067) );
  NAND2_X1 U9574 ( .A1(n8319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U9575 ( .A1(n6930), .A2(n6929), .ZN(n6928) );
  NAND2_X1 U9576 ( .A1(n6933), .A2(n6768), .ZN(n14545) );
  NAND2_X1 U9577 ( .A1(n6942), .A2(n6719), .ZN(n11103) );
  AND2_X1 U9578 ( .A1(n6945), .A2(n6944), .ZN(n6941) );
  INV_X1 U9579 ( .A(n11090), .ZN(n6946) );
  NAND2_X1 U9580 ( .A1(n11122), .A2(n6670), .ZN(n6948) );
  NAND2_X2 U9581 ( .A1(n7902), .A2(n6957), .ZN(n7905) );
  NAND4_X1 U9582 ( .A1(n6954), .A2(n6956), .A3(n6953), .A4(n7902), .ZN(n8233)
         );
  INV_X1 U9583 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6957) );
  AOI21_X1 U9584 ( .B1(n6960), .B2(n11151), .A(n11150), .ZN(n6958) );
  OAI21_X1 U9585 ( .B1(n6960), .B2(n11151), .A(n6747), .ZN(n6959) );
  OAI21_X1 U9586 ( .B1(n11072), .B2(n6961), .A(n6962), .ZN(n11079) );
  NAND2_X1 U9587 ( .A1(n8323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8318) );
  NAND3_X1 U9588 ( .A1(n7588), .A2(n7594), .A3(n6965), .ZN(n6964) );
  NAND2_X1 U9589 ( .A1(n8032), .A2(n6967), .ZN(n6966) );
  OAI211_X1 U9590 ( .C1(n8032), .C2(n6969), .A(n6968), .B(n6966), .ZN(n8413)
         );
  INV_X1 U9591 ( .A(n8413), .ZN(n8412) );
  NAND2_X2 U9592 ( .A1(n6973), .A2(n13919), .ZN(n14110) );
  OAI21_X1 U9593 ( .B1(n13909), .B2(n13934), .A(n13911), .ZN(n14185) );
  AOI21_X1 U9594 ( .B1(n13934), .B2(n13911), .A(n6982), .ZN(n6981) );
  INV_X1 U9595 ( .A(n14184), .ZN(n6982) );
  NAND2_X2 U9596 ( .A1(n6983), .A2(n10001), .ZN(n11778) );
  OR2_X2 U9597 ( .A1(n13930), .A2(n13981), .ZN(n13932) );
  MUX2_X1 U9598 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7737), .Z(n6986) );
  NAND2_X1 U9599 ( .A1(n15156), .A2(n15131), .ZN(n12282) );
  AND3_X2 U9600 ( .A1(n6745), .A2(n8517), .A3(n8516), .ZN(n15131) );
  NAND2_X1 U9601 ( .A1(n7492), .A2(n12246), .ZN(n7003) );
  INV_X1 U9602 ( .A(n7012), .ZN(n10481) );
  NAND2_X1 U9603 ( .A1(n12774), .A2(n7015), .ZN(n7013) );
  NAND2_X1 U9604 ( .A1(n7013), .A2(n7014), .ZN(n12727) );
  OAI21_X1 U9605 ( .B1(n12681), .B2(n7019), .A(n7018), .ZN(n12635) );
  NAND2_X1 U9606 ( .A1(n7027), .A2(n9951), .ZN(n7028) );
  NAND2_X1 U9607 ( .A1(n9855), .A2(n7029), .ZN(n7027) );
  NAND2_X1 U9608 ( .A1(n9952), .A2(n9951), .ZN(n10269) );
  NAND2_X1 U9609 ( .A1(n7029), .A2(n9855), .ZN(n9952) );
  OAI21_X2 U9610 ( .B1(n12138), .B2(n12438), .A(n6668), .ZN(n12182) );
  OR2_X2 U9611 ( .A1(n12118), .A2(n6754), .ZN(n7032) );
  XNOR2_X1 U9612 ( .A(n8753), .B(n9355), .ZN(n8749) );
  NAND2_X1 U9613 ( .A1(n8454), .A2(n7035), .ZN(n7034) );
  NAND3_X1 U9614 ( .A1(n7042), .A2(n7041), .A3(n7043), .ZN(n13535) );
  NAND4_X1 U9615 ( .A1(n7042), .A2(n7041), .A3(n7043), .A4(n14938), .ZN(n7045)
         );
  NAND2_X1 U9616 ( .A1(n10546), .A2(n10545), .ZN(n10745) );
  NAND2_X1 U9617 ( .A1(n7048), .A2(n7049), .ZN(n7240) );
  NAND2_X1 U9618 ( .A1(n8028), .A2(n7052), .ZN(n7050) );
  NAND2_X1 U9619 ( .A1(n13276), .A2(n7057), .ZN(n7056) );
  NAND2_X1 U9620 ( .A1(n7062), .A2(n9935), .ZN(n9940) );
  INV_X1 U9621 ( .A(n9590), .ZN(n7063) );
  OAI21_X2 U9622 ( .B1(n11002), .B2(n11001), .A(n11005), .ZN(n11007) );
  NAND2_X1 U9623 ( .A1(n10752), .A2(n10934), .ZN(n11613) );
  OAI211_X1 U9624 ( .C1(n13705), .C2(n7077), .A(n7070), .B(n9184), .ZN(n7075)
         );
  AND2_X1 U9625 ( .A1(n7081), .A2(n7083), .ZN(n7078) );
  NAND2_X1 U9626 ( .A1(n7080), .A2(n9183), .ZN(n7079) );
  INV_X1 U9627 ( .A(n7083), .ZN(n7080) );
  NAND2_X1 U9628 ( .A1(n13754), .A2(n6702), .ZN(n7085) );
  NAND2_X1 U9629 ( .A1(n7085), .A2(n6760), .ZN(n13687) );
  NAND2_X1 U9630 ( .A1(n13754), .A2(n13755), .ZN(n7087) );
  NAND2_X2 U9631 ( .A1(n7092), .A2(n8609), .ZN(n11730) );
  NAND4_X1 U9632 ( .A1(n8237), .A2(n7656), .A3(n8235), .A4(n8236), .ZN(n7104)
         );
  NOR3_X4 U9633 ( .A1(n13501), .A2(n7109), .A3(n7110), .ZN(n13460) );
  AND2_X2 U9634 ( .A1(n8617), .A2(n7120), .ZN(n14694) );
  AND2_X1 U9635 ( .A1(n8618), .A2(n8616), .ZN(n7120) );
  NOR2_X2 U9636 ( .A1(n10002), .A2(n11778), .ZN(n7125) );
  NAND2_X1 U9637 ( .A1(n13978), .A2(n7128), .ZN(n13957) );
  NAND2_X1 U9638 ( .A1(n13978), .A2(n7126), .ZN(n13904) );
  NAND2_X1 U9639 ( .A1(n13978), .A2(n14323), .ZN(n13971) );
  INV_X1 U9640 ( .A(n13957), .ZN(n13905) );
  NAND2_X1 U9641 ( .A1(n15114), .A2(n15113), .ZN(n7130) );
  NAND2_X1 U9642 ( .A1(n11973), .A2(n7149), .ZN(n7146) );
  OAI21_X2 U9643 ( .B1(n10734), .B2(n7156), .A(n7154), .ZN(n10924) );
  INV_X1 U9644 ( .A(n7169), .ZN(n15078) );
  INV_X1 U9645 ( .A(n10147), .ZN(n7168) );
  INV_X1 U9646 ( .A(n12525), .ZN(n7172) );
  INV_X1 U9647 ( .A(n7182), .ZN(n10138) );
  NOR2_X1 U9648 ( .A1(n14971), .A2(n10134), .ZN(n14991) );
  NAND3_X1 U9649 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n7184) );
  NAND2_X1 U9650 ( .A1(n7884), .A2(n7188), .ZN(n7187) );
  NAND2_X1 U9651 ( .A1(n8451), .A2(n7194), .ZN(n7193) );
  OAI21_X2 U9652 ( .B1(n10561), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7211), .ZN(
        n10582) );
  OAI22_X2 U9653 ( .A1(n10641), .A2(n10640), .B1(n11116), .B2(n13146), .ZN(
        n10711) );
  NAND2_X1 U9654 ( .A1(n9687), .A2(n7216), .ZN(n7215) );
  NAND2_X1 U9655 ( .A1(n13468), .A2(n7232), .ZN(n7228) );
  NAND2_X1 U9656 ( .A1(n7228), .A2(n7229), .ZN(n13263) );
  OAI211_X1 U9657 ( .C1(n7244), .C2(n15142), .A(n8960), .B(n8755), .ZN(n8756)
         );
  NAND2_X1 U9658 ( .A1(n7692), .A2(n7691), .ZN(n8102) );
  INV_X1 U9659 ( .A(n9046), .ZN(n7249) );
  AOI21_X1 U9660 ( .B1(n7249), .B2(n7253), .A(n7251), .ZN(n7250) );
  NAND2_X1 U9661 ( .A1(n12182), .A2(n7276), .ZN(n7275) );
  OR2_X1 U9662 ( .A1(n12152), .A2(n12435), .ZN(n7289) );
  NAND2_X1 U9663 ( .A1(n8961), .A2(n8962), .ZN(n9046) );
  OAI21_X1 U9664 ( .B1(n12836), .B2(n10672), .A(n10671), .ZN(n10674) );
  NAND2_X1 U9665 ( .A1(n9358), .A2(n15150), .ZN(n12283) );
  NAND2_X1 U9666 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  NAND2_X1 U9667 ( .A1(n10582), .A2(n10581), .ZN(n10584) );
  NAND2_X1 U9668 ( .A1(n10466), .A2(n10465), .ZN(n10469) );
  NAND2_X1 U9669 ( .A1(n7801), .A2(n7800), .ZN(n7781) );
  OAI22_X1 U9670 ( .A1(n12232), .A2(n12231), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14364), .ZN(n12234) );
  NAND2_X1 U9671 ( .A1(n9501), .A2(n12292), .ZN(n10193) );
  NAND2_X1 U9672 ( .A1(n12711), .A2(n12710), .ZN(n12713) );
  XNOR2_X1 U9673 ( .A(n11075), .B(n13152), .ZN(n11404) );
  NAND2_X1 U9674 ( .A1(n13266), .A2(n13265), .ZN(n13403) );
  NOR2_X1 U9675 ( .A1(n9567), .A2(n11034), .ZN(n10064) );
  NOR2_X2 U9676 ( .A1(n9680), .A2(n11089), .ZN(n9688) );
  NAND2_X1 U9677 ( .A1(n9295), .A2(n9282), .ZN(n11400) );
  OAI21_X1 U9678 ( .B1(n12779), .B2(n10968), .A(n10967), .ZN(n10970) );
  OR2_X2 U9679 ( .A1(n10893), .A2(n11418), .ZN(n10895) );
  OR2_X2 U9680 ( .A1(n13403), .A2(n13267), .ZN(n13270) );
  NAND2_X1 U9681 ( .A1(n9289), .A2(n9301), .ZN(n9540) );
  NAND2_X1 U9682 ( .A1(n10469), .A2(n10468), .ZN(n10470) );
  NAND2_X1 U9683 ( .A1(n9407), .A2(n9406), .ZN(n9410) );
  OR2_X1 U9684 ( .A1(n11337), .A2(n9928), .ZN(n8353) );
  NOR3_X2 U9685 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n7663) );
  INV_X1 U9686 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U9687 ( .A1(n7296), .A2(n7295), .ZN(n11803) );
  NAND2_X1 U9688 ( .A1(n11797), .A2(n7300), .ZN(n7296) );
  INV_X1 U9689 ( .A(n11800), .ZN(n7303) );
  INV_X1 U9690 ( .A(n14467), .ZN(n14471) );
  INV_X1 U9691 ( .A(n14640), .ZN(n14639) );
  NAND2_X1 U9692 ( .A1(n14467), .A2(n7306), .ZN(n14640) );
  INV_X1 U9693 ( .A(n14470), .ZN(n7306) );
  NAND2_X1 U9694 ( .A1(n7307), .A2(n7308), .ZN(n11951) );
  NOR2_X2 U9695 ( .A1(n15616), .A2(n14438), .ZN(n14440) );
  NAND3_X1 U9696 ( .A1(n11761), .A2(n11760), .A3(n6767), .ZN(n7316) );
  INV_X1 U9697 ( .A(n11762), .ZN(n7317) );
  NAND2_X1 U9698 ( .A1(n7318), .A2(n7319), .ZN(n11831) );
  NAND3_X1 U9699 ( .A1(n11810), .A2(n7655), .A3(n7654), .ZN(n7318) );
  INV_X2 U9700 ( .A(n8839), .ZN(n11529) );
  NAND2_X1 U9701 ( .A1(n7324), .A2(n7326), .ZN(n11756) );
  NAND3_X1 U9702 ( .A1(n11837), .A2(n7333), .A3(n7336), .ZN(n7328) );
  OR2_X1 U9703 ( .A1(n7334), .A2(n7338), .ZN(n7330) );
  NOR2_X2 U9704 ( .A1(n11841), .A2(n11840), .ZN(n7335) );
  NAND3_X1 U9705 ( .A1(n11786), .A2(n6762), .A3(n11785), .ZN(n7340) );
  INV_X1 U9706 ( .A(n11776), .ZN(n7344) );
  NAND3_X1 U9707 ( .A1(n8772), .A2(n8771), .A3(n7350), .ZN(n8897) );
  NAND2_X1 U9708 ( .A1(n8722), .A2(n8721), .ZN(n7351) );
  OAI21_X1 U9709 ( .B1(n13024), .B2(n7363), .A(n7354), .ZN(n7362) );
  NAND2_X1 U9710 ( .A1(n13024), .A2(n7356), .ZN(n7354) );
  INV_X1 U9711 ( .A(n7362), .ZN(n13096) );
  XNOR2_X1 U9712 ( .A(n13024), .B(n6772), .ZN(n13041) );
  NAND2_X1 U9713 ( .A1(n13130), .A2(n6765), .ZN(n7368) );
  OAI211_X1 U9714 ( .C1(n13130), .C2(n7369), .A(n7368), .B(n13073), .ZN(
        P2_U3192) );
  NAND2_X1 U9715 ( .A1(n13130), .A2(n13034), .ZN(n13065) );
  NOR2_X1 U9716 ( .A1(n13063), .A2(n13062), .ZN(n7375) );
  NOR2_X2 U9717 ( .A1(n13125), .A2(n13124), .ZN(n13123) );
  OR2_X2 U9718 ( .A1(n9885), .A2(n7381), .ZN(n9924) );
  OR2_X1 U9719 ( .A1(n9889), .A2(n9884), .ZN(n7381) );
  AND2_X2 U9720 ( .A1(n9745), .A2(n9746), .ZN(n9885) );
  AND2_X1 U9721 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  NAND2_X1 U9722 ( .A1(n9016), .A2(n7384), .ZN(n9131) );
  NAND2_X1 U9723 ( .A1(n7383), .A2(n9130), .ZN(n7382) );
  INV_X1 U9724 ( .A(n8233), .ZN(n7385) );
  INV_X1 U9725 ( .A(n13035), .ZN(n13001) );
  NAND2_X1 U9726 ( .A1(n13358), .A2(n7389), .ZN(n7386) );
  NAND2_X1 U9727 ( .A1(n7386), .A2(n7387), .ZN(n13325) );
  INV_X2 U9728 ( .A(n11040), .ZN(n8590) );
  NAND2_X2 U9729 ( .A1(n10321), .A2(n6641), .ZN(n11236) );
  NAND2_X1 U9730 ( .A1(n7401), .A2(n6769), .ZN(n7400) );
  INV_X1 U9731 ( .A(n7663), .ZN(n7664) );
  NAND2_X2 U9732 ( .A1(n9560), .A2(n8584), .ZN(n9275) );
  XNOR2_X2 U9733 ( .A(n7420), .B(n7419), .ZN(n10661) );
  NAND2_X1 U9734 ( .A1(n13783), .A2(n7427), .ZN(n7425) );
  NOR2_X4 U9735 ( .A1(n7433), .A2(n7432), .ZN(n11680) );
  INV_X2 U9736 ( .A(n8605), .ZN(n7432) );
  NOR2_X1 U9737 ( .A1(n14571), .A2(n10864), .ZN(n10867) );
  NAND2_X1 U9738 ( .A1(n7452), .A2(n7456), .ZN(n7448) );
  INV_X1 U9739 ( .A(n7450), .ZN(n7449) );
  NAND3_X1 U9740 ( .A1(n7453), .A2(n7454), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n7456) );
  NAND2_X1 U9741 ( .A1(n7924), .A2(n7461), .ZN(n7458) );
  NAND2_X1 U9742 ( .A1(n7458), .A2(n7459), .ZN(n8009) );
  NAND2_X1 U9743 ( .A1(n10934), .A2(n7469), .ZN(n7468) );
  NAND2_X1 U9744 ( .A1(n10934), .A2(n10933), .ZN(n10993) );
  NAND2_X1 U9745 ( .A1(n9434), .A2(n7484), .ZN(n7483) );
  NAND2_X1 U9746 ( .A1(n9434), .A2(n9433), .ZN(n7490) );
  NAND2_X1 U9747 ( .A1(n12448), .A2(n9355), .ZN(n12272) );
  NAND2_X1 U9748 ( .A1(n15103), .A2(n10203), .ZN(n10204) );
  NAND2_X1 U9749 ( .A1(n10729), .A2(n6757), .ZN(n10759) );
  NAND2_X1 U9750 ( .A1(n13935), .A2(n13934), .ZN(n13937) );
  NAND2_X1 U9751 ( .A1(n14589), .A2(n11801), .ZN(n7510) );
  NAND3_X1 U9752 ( .A1(n7715), .A2(n7714), .A3(n7713), .ZN(n7512) );
  NAND2_X1 U9753 ( .A1(n7512), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U9754 ( .A1(n14222), .A2(n14592), .ZN(n7514) );
  NAND2_X1 U9755 ( .A1(n9968), .A2(n7520), .ZN(n7519) );
  AOI21_X2 U9756 ( .B1(n7522), .B2(n7517), .A(n6749), .ZN(n7520) );
  NAND3_X1 U9757 ( .A1(n7519), .A2(n7608), .A3(n7518), .ZN(n9974) );
  NAND2_X2 U9758 ( .A1(n7528), .A2(n7526), .ZN(n13997) );
  NAND2_X1 U9759 ( .A1(n14252), .A2(n14020), .ZN(n7537) );
  OAI21_X2 U9760 ( .B1(n14123), .B2(n7540), .A(n7538), .ZN(n14084) );
  NAND2_X1 U9761 ( .A1(n10021), .A2(n6663), .ZN(n7549) );
  NAND3_X1 U9762 ( .A1(n7674), .A2(n8011), .A3(n7660), .ZN(n7665) );
  NOR2_X2 U9763 ( .A1(n7554), .A2(n7664), .ZN(n7553) );
  NOR2_X2 U9764 ( .A1(n8327), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U9765 ( .A1(n7557), .A2(n7555), .ZN(n7556) );
  INV_X1 U9766 ( .A(n11117), .ZN(n7559) );
  AOI21_X1 U9767 ( .B1(n11182), .B2(n11181), .A(n11180), .ZN(n11184) );
  OAI21_X1 U9768 ( .B1(n6716), .B2(n7561), .A(n7560), .ZN(n11289) );
  INV_X1 U9769 ( .A(n7563), .ZN(n7562) );
  NAND2_X1 U9770 ( .A1(n7573), .A2(n7577), .ZN(n11091) );
  NAND3_X1 U9771 ( .A1(n7574), .A2(n6714), .A3(n11080), .ZN(n7573) );
  NAND2_X1 U9772 ( .A1(n7576), .A2(n7575), .ZN(n7574) );
  INV_X1 U9773 ( .A(n11086), .ZN(n7575) );
  NAND2_X1 U9774 ( .A1(n7581), .A2(n7580), .ZN(n7579) );
  NOR2_X1 U9775 ( .A1(n11137), .A2(n7583), .ZN(n7580) );
  INV_X1 U9776 ( .A(n11138), .ZN(n7581) );
  OAI21_X1 U9777 ( .B1(n11196), .B2(n7593), .A(n7584), .ZN(n7588) );
  INV_X1 U9778 ( .A(n10018), .ZN(n7596) );
  NAND3_X1 U9779 ( .A1(n7597), .A2(n7598), .A3(n10404), .ZN(n10407) );
  OAI21_X1 U9780 ( .B1(n7606), .B2(n9625), .A(n9815), .ZN(n7601) );
  NAND2_X1 U9781 ( .A1(n7604), .A2(n7606), .ZN(n7602) );
  NAND2_X1 U9782 ( .A1(n9626), .A2(n7604), .ZN(n7603) );
  OAI21_X1 U9783 ( .B1(n9985), .B2(n7612), .A(n6662), .ZN(n10051) );
  NAND2_X1 U9784 ( .A1(n9985), .A2(n6662), .ZN(n7609) );
  OAI21_X1 U9785 ( .B1(n10823), .B2(n11928), .A(n10824), .ZN(n14503) );
  AND2_X1 U9786 ( .A1(n7627), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U9787 ( .A1(n7974), .A2(n7630), .ZN(n8168) );
  NAND2_X1 U9788 ( .A1(n14069), .A2(n7634), .ZN(n7631) );
  NAND2_X1 U9789 ( .A1(n7632), .A2(n7631), .ZN(n14014) );
  AND2_X1 U9790 ( .A1(n13932), .A2(n7645), .ZN(n13964) );
  NAND3_X1 U9791 ( .A1(n13932), .A2(n7637), .A3(n7645), .ZN(n7638) );
  OR2_X2 U9792 ( .A1(n13932), .A2(n7644), .ZN(n7639) );
  INV_X1 U9793 ( .A(n7641), .ZN(n7640) );
  OAI21_X1 U9794 ( .B1(n7645), .B2(n7644), .A(n7642), .ZN(n7641) );
  INV_X1 U9795 ( .A(n7647), .ZN(n7643) );
  NAND2_X1 U9796 ( .A1(n13950), .A2(n7647), .ZN(n7644) );
  INV_X1 U9797 ( .A(n6640), .ZN(n11425) );
  NAND2_X2 U9798 ( .A1(n14958), .A2(n6640), .ZN(n11067) );
  INV_X1 U9799 ( .A(n8129), .ZN(n12990) );
  INV_X1 U9800 ( .A(n11230), .ZN(n11233) );
  OR2_X2 U9801 ( .A1(n13157), .A2(n8590), .ZN(n9560) );
  NAND4_X4 U9802 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n13157)
         );
  OR2_X1 U9803 ( .A1(n11560), .A2(n11236), .ZN(n11011) );
  OR2_X1 U9804 ( .A1(n11199), .A2(n11236), .ZN(n11201) );
  OR2_X1 U9805 ( .A1(n11544), .A2(n11236), .ZN(n11186) );
  OR2_X1 U9806 ( .A1(n11514), .A2(n11236), .ZN(n11153) );
  NAND2_X1 U9807 ( .A1(n11289), .A2(n11288), .ZN(n11287) );
  OR2_X1 U9808 ( .A1(n14192), .A2(n14200), .ZN(n8674) );
  OR2_X1 U9809 ( .A1(n11613), .A2(n11612), .ZN(n11616) );
  NAND4_X2 U9810 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n8507), .ZN(n15147)
         );
  INV_X1 U9811 ( .A(n15227), .ZN(n15231) );
  AND2_X1 U9812 ( .A1(n7725), .A2(n7724), .ZN(n7649) );
  INV_X1 U9813 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7690) );
  OR2_X1 U9814 ( .A1(n12733), .A2(n12714), .ZN(n7650) );
  AND2_X1 U9815 ( .A1(n11350), .A2(n11348), .ZN(n7651) );
  AND2_X1 U9816 ( .A1(n11444), .A2(n11443), .ZN(n7652) );
  NOR2_X1 U9817 ( .A1(n11447), .A2(n11446), .ZN(n7653) );
  AND3_X1 U9818 ( .A1(n11823), .A2(n11822), .A3(n13941), .ZN(n7654) );
  INV_X1 U9819 ( .A(n12254), .ZN(n10730) );
  OR2_X1 U9820 ( .A1(n11809), .A2(n11898), .ZN(n7655) );
  NAND2_X1 U9821 ( .A1(n12083), .A2(n12082), .ZN(n12084) );
  INV_X1 U9822 ( .A(n11144), .ZN(n11145) );
  INV_X1 U9823 ( .A(n11819), .ZN(n11811) );
  INV_X1 U9824 ( .A(n11231), .ZN(n11232) );
  INV_X1 U9825 ( .A(n11285), .ZN(n11286) );
  INV_X1 U9826 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7682) );
  NOR2_X1 U9827 ( .A1(n9577), .A2(SI_18_), .ZN(n9582) );
  INV_X1 U9828 ( .A(n12034), .ZN(n9766) );
  INV_X1 U9829 ( .A(n10572), .ZN(n8811) );
  INV_X1 U9830 ( .A(n12022), .ZN(n9764) );
  INV_X1 U9831 ( .A(n10297), .ZN(n8141) );
  INV_X1 U9832 ( .A(n12056), .ZN(n9768) );
  INV_X1 U9833 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7691) );
  INV_X1 U9834 ( .A(n14548), .ZN(n10688) );
  NAND2_X1 U9835 ( .A1(n9292), .A2(n11397), .ZN(n10055) );
  NAND2_X1 U9836 ( .A1(n8214), .A2(n14654), .ZN(n8211) );
  AND2_X1 U9837 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n11581), .ZN(n11599) );
  AND2_X1 U9838 ( .A1(n11599), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11618) );
  INV_X1 U9839 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9527) );
  INV_X1 U9840 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7973) );
  INV_X1 U9841 ( .A(n8649), .ZN(n8529) );
  INV_X1 U9842 ( .A(n10972), .ZN(n8814) );
  AND2_X1 U9843 ( .A1(n8811), .A2(n8810), .ZN(n10675) );
  OR2_X1 U9844 ( .A1(n12045), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n12056) );
  OR2_X1 U9845 ( .A1(n11999), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U9846 ( .A1(n9768), .A2(n9767), .ZN(n12058) );
  OR2_X1 U9847 ( .A1(n8486), .A2(n8485), .ZN(n8708) );
  OR2_X1 U9848 ( .A1(n9405), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9406) );
  AND2_X1 U9849 ( .A1(n7880), .A2(n7846), .ZN(n7847) );
  NAND2_X1 U9850 ( .A1(n7901), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7780) );
  INV_X1 U9851 ( .A(n11275), .ZN(n11274) );
  OR2_X1 U9852 ( .A1(n11255), .A2(n11252), .ZN(n11275) );
  NAND2_X1 U9853 ( .A1(n11014), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11202) );
  AND2_X1 U9854 ( .A1(n11618), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11638) );
  INV_X1 U9855 ( .A(n11670), .ZN(n11687) );
  NOR2_X1 U9856 ( .A1(n13765), .A2(n11548), .ZN(n11564) );
  NAND2_X1 U9857 ( .A1(n10791), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U9858 ( .A1(n9174), .A2(n9173), .ZN(n9178) );
  OR2_X1 U9859 ( .A1(n14469), .A2(n14468), .ZN(n14407) );
  NAND2_X1 U9860 ( .A1(n9762), .A2(n9761), .ZN(n11999) );
  NAND2_X1 U9861 ( .A1(n8138), .A2(n9858), .ZN(n9859) );
  OR2_X1 U9862 ( .A1(n10882), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n10972) );
  INV_X1 U9863 ( .A(n6638), .ZN(n12062) );
  INV_X1 U9864 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9722) );
  INV_X1 U9865 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9858) );
  OR2_X1 U9866 ( .A1(n12058), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12620) );
  INV_X1 U9867 ( .A(n12715), .ZN(n12679) );
  INV_X1 U9868 ( .A(n12260), .ZN(n12798) );
  INV_X1 U9869 ( .A(n12821), .ZN(n12826) );
  AND2_X1 U9870 ( .A1(n8708), .A2(n8713), .ZN(n8709) );
  INV_X1 U9871 ( .A(n15149), .ZN(n15128) );
  AND2_X1 U9872 ( .A1(n12614), .A2(n9273), .ZN(n12423) );
  AND2_X1 U9873 ( .A1(n7777), .A2(n7776), .ZN(n7794) );
  AND2_X1 U9874 ( .A1(n9892), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9909) );
  AND2_X1 U9875 ( .A1(n11458), .A2(n6640), .ZN(n8366) );
  OR2_X1 U9876 ( .A1(n11217), .A2(n13044), .ZN(n11255) );
  OAI211_X1 U9877 ( .C1(n11236), .C2(n8727), .A(n8726), .B(n8725), .ZN(n11037)
         );
  OR2_X1 U9878 ( .A1(n13512), .A2(n9470), .ZN(n14868) );
  OR2_X1 U9879 ( .A1(n8802), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U9880 ( .A1(n8613), .A2(n8217), .ZN(n8612) );
  AND2_X1 U9881 ( .A1(n8202), .A2(n8267), .ZN(n9612) );
  INV_X1 U9882 ( .A(n11656), .ZN(n11884) );
  INV_X1 U9883 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8939) );
  INV_X1 U9884 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10523) );
  INV_X1 U9885 ( .A(n13933), .ZN(n13965) );
  INV_X1 U9886 ( .A(n11902), .ZN(n11907) );
  INV_X1 U9887 ( .A(n14564), .ZN(n14610) );
  INV_X1 U9888 ( .A(n14201), .ZN(n14180) );
  INV_X1 U9889 ( .A(n14262), .ZN(n14609) );
  INV_X1 U9890 ( .A(n8214), .ZN(n8208) );
  XNOR2_X1 U9891 ( .A(n9436), .B(SI_17_), .ZN(n9433) );
  XNOR2_X1 U9892 ( .A(n9083), .B(SI_13_), .ZN(n9080) );
  INV_X1 U9893 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7705) );
  OAI21_X1 U9894 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14408), .A(n14407), .ZN(
        n14413) );
  INV_X1 U9895 ( .A(n12714), .ZN(n12742) );
  INV_X1 U9896 ( .A(n12209), .ZN(n12199) );
  NAND2_X1 U9897 ( .A1(n9037), .A2(n12432), .ZN(n12207) );
  AND2_X1 U9898 ( .A1(n12017), .A2(n12016), .ZN(n12730) );
  INV_X1 U9899 ( .A(n12616), .ZN(n15095) );
  OAI21_X1 U9900 ( .B1(n12652), .B2(n12651), .A(n12650), .ZN(n12858) );
  INV_X1 U9901 ( .A(n15130), .ZN(n15148) );
  INV_X1 U9902 ( .A(n15154), .ZN(n15133) );
  INV_X1 U9903 ( .A(n12321), .ZN(n12255) );
  INV_X1 U9904 ( .A(n12842), .ZN(n12792) );
  INV_X1 U9905 ( .A(n15209), .ZN(n15155) );
  AND2_X1 U9906 ( .A1(n12423), .A2(n11971), .ZN(n15206) );
  NAND2_X1 U9907 ( .A1(n10954), .A2(n10953), .ZN(n10955) );
  INV_X1 U9908 ( .A(n14558), .ZN(n13121) );
  OR2_X1 U9909 ( .A1(n11368), .A2(n11330), .ZN(n13318) );
  INV_X1 U9910 ( .A(n8399), .ZN(n14773) );
  OR2_X1 U9911 ( .A1(n8248), .A2(n8247), .ZN(n8258) );
  INV_X1 U9912 ( .A(n13225), .ZN(n14847) );
  INV_X1 U9913 ( .A(n14846), .ZN(n14854) );
  AND2_X1 U9914 ( .A1(n11369), .A2(n13318), .ZN(n13331) );
  INV_X1 U9915 ( .A(n13431), .ZN(n13474) );
  INV_X1 U9916 ( .A(n13411), .ZN(n14862) );
  AND2_X1 U9917 ( .A1(n14949), .A2(n8582), .ZN(n14931) );
  INV_X1 U9918 ( .A(n14931), .ZN(n14938) );
  AND2_X1 U9919 ( .A1(n8302), .A2(n8301), .ZN(n14875) );
  AND2_X1 U9920 ( .A1(n8304), .A2(n8303), .ZN(n8592) );
  AND2_X1 U9921 ( .A1(n8326), .A2(n10548), .ZN(n8782) );
  AND2_X1 U9922 ( .A1(n10789), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10791) );
  INV_X1 U9923 ( .A(n14141), .ZN(n14591) );
  AND2_X1 U9924 ( .A1(n14675), .A2(n8218), .ZN(n14717) );
  AND2_X1 U9925 ( .A1(n8688), .A2(n9612), .ZN(n13818) );
  OR2_X1 U9926 ( .A1(n11671), .A2(n14040), .ZN(n11624) );
  OR2_X1 U9927 ( .A1(n14658), .A2(n11956), .ZN(n13886) );
  INV_X1 U9928 ( .A(n13867), .ZN(n14669) );
  INV_X1 U9929 ( .A(n13996), .ZN(n13994) );
  INV_X1 U9930 ( .A(n13919), .ZN(n14113) );
  NAND2_X1 U9931 ( .A1(n14504), .A2(n14677), .ZN(n9616) );
  NAND2_X1 U9932 ( .A1(n8280), .A2(n11714), .ZN(n14592) );
  AND2_X1 U9933 ( .A1(n11957), .A2(n8274), .ZN(n8688) );
  INV_X1 U9934 ( .A(n14592), .ZN(n14704) );
  INV_X1 U9935 ( .A(n14717), .ZN(n14729) );
  INV_X1 U9936 ( .A(n14289), .ZN(n14725) );
  INV_X1 U9937 ( .A(n8274), .ZN(n9613) );
  AND2_X1 U9938 ( .A1(n9103), .A2(n8808), .ZN(n10781) );
  AND2_X1 U9939 ( .A1(n8118), .A2(n8117), .ZN(n15092) );
  NAND2_X1 U9940 ( .A1(n8513), .A2(n8713), .ZN(n12214) );
  AND2_X1 U9941 ( .A1(n12228), .A2(n9784), .ZN(n12241) );
  INV_X1 U9942 ( .A(n12730), .ZN(n12438) );
  INV_X1 U9943 ( .A(n10479), .ZN(n12445) );
  AND2_X1 U9944 ( .A1(n12639), .A2(n12638), .ZN(n12854) );
  NAND2_X1 U9945 ( .A1(n15227), .A2(n15155), .ZN(n12918) );
  AND2_X2 U9946 ( .A1(n8698), .A2(n8713), .ZN(n15217) );
  INV_X1 U9947 ( .A(n15217), .ZN(n15215) );
  INV_X1 U9948 ( .A(SI_10_), .ZN(n9945) );
  INV_X1 U9949 ( .A(n10114), .ZN(n15068) );
  INV_X1 U9950 ( .A(n12979), .ZN(n12997) );
  NAND2_X1 U9951 ( .A1(n8375), .A2(n14953), .ZN(n14552) );
  OR2_X1 U9952 ( .A1(n13512), .A2(n11168), .ZN(n13411) );
  OR2_X1 U9953 ( .A1(n13512), .A2(n9461), .ZN(n13507) );
  INV_X1 U9954 ( .A(n13246), .ZN(n13628) );
  INV_X1 U9955 ( .A(n13289), .ZN(n13656) );
  INV_X1 U9956 ( .A(n14960), .ZN(n14959) );
  NOR2_X1 U9957 ( .A1(n14875), .A2(n14907), .ZN(n14887) );
  CLKBUF_X1 U9958 ( .A(n14887), .Z(n14904) );
  INV_X1 U9959 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10322) );
  INV_X1 U9960 ( .A(n14263), .ZN(n13791) );
  INV_X1 U9961 ( .A(n14080), .ZN(n14261) );
  INV_X1 U9962 ( .A(n10806), .ZN(n14590) );
  OR2_X1 U9963 ( .A1(n14658), .A2(n8636), .ZN(n13885) );
  OR2_X1 U9964 ( .A1(n14658), .A2(n8047), .ZN(n13867) );
  OR3_X1 U9965 ( .A1(n13978), .A2(n13977), .A3(n14719), .ZN(n14231) );
  INV_X1 U9966 ( .A(n14686), .ZN(n14177) );
  NAND2_X1 U9967 ( .A1(n14686), .A2(n13891), .ZN(n14130) );
  INV_X1 U9968 ( .A(n14686), .ZN(n14689) );
  INV_X1 U9969 ( .A(n14741), .ZN(n14739) );
  INV_X1 U9970 ( .A(n13961), .ZN(n14321) );
  INV_X1 U9971 ( .A(n14733), .ZN(n14731) );
  AND3_X2 U9972 ( .A1(n8687), .A2(n11957), .A3(n9613), .ZN(n14733) );
  AND2_X1 U9973 ( .A1(n9062), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8187) );
  INV_X1 U9974 ( .A(n7944), .ZN(n10754) );
  INV_X1 U9975 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9446) );
  INV_X1 U9976 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10779) );
  NOR2_X2 U9977 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8236) );
  NOR2_X2 U9978 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8235) );
  NOR2_X1 U9979 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7656) );
  NOR2_X2 U9980 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7658) );
  INV_X2 U9981 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8803) );
  NOR2_X1 U9982 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7659) );
  OR2_X1 U9983 ( .A1(n7665), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9984 ( .A1(n7668), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7661) );
  MUX2_X1 U9985 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7661), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n7662) );
  INV_X1 U9986 ( .A(n7662), .ZN(n7666) );
  NOR2_X1 U9987 ( .A1(n7666), .A2(n8241), .ZN(n8302) );
  NAND2_X1 U9988 ( .A1(n7671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7667) );
  MUX2_X1 U9989 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7667), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n7669) );
  NAND2_X1 U9990 ( .A1(n7669), .A2(n7668), .ZN(n10935) );
  NAND2_X1 U9991 ( .A1(n7665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7670) );
  MUX2_X1 U9992 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7670), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n7672) );
  NAND2_X1 U9993 ( .A1(n7672), .A2(n7671), .ZN(n10753) );
  NOR2_X1 U9994 ( .A1(n10935), .A2(n10753), .ZN(n7673) );
  NAND2_X1 U9995 ( .A1(n8302), .A2(n7673), .ZN(n8326) );
  INV_X1 U9996 ( .A(n7674), .ZN(n7675) );
  OAI21_X1 U9997 ( .B1(n9070), .B2(n7675), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7677) );
  XNOR2_X1 U9998 ( .A(n7677), .B(n7676), .ZN(n10548) );
  INV_X1 U9999 ( .A(n10548), .ZN(n7678) );
  NOR2_X1 U10000 ( .A1(n8326), .A2(n7678), .ZN(n8247) );
  AND2_X1 U10001 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8247), .ZN(P2_U3947) );
  NOR2_X1 U10002 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7681) );
  NAND4_X1 U10003 ( .A1(n7681), .A2(n7680), .A3(n7679), .A4(n15362), .ZN(n7938) );
  NAND3_X1 U10004 ( .A1(n7785), .A2(n7941), .A3(n7682), .ZN(n7683) );
  NOR2_X1 U10005 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n7686) );
  NAND2_X1 U10006 ( .A1(n8102), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7693) );
  XNOR2_X1 U10007 ( .A(n7693), .B(P3_IR_REG_26__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10008 ( .A1(n7694), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7695) );
  XNOR2_X1 U10009 ( .A(n7695), .B(n7691), .ZN(n10564) );
  INV_X1 U10010 ( .A(n10564), .ZN(n7699) );
  INV_X1 U10011 ( .A(n10474), .ZN(n7698) );
  AND2_X1 U10012 ( .A1(n7699), .A2(n7698), .ZN(n7700) );
  NAND2_X1 U10013 ( .A1(n7825), .A2(n7700), .ZN(n8498) );
  INV_X1 U10014 ( .A(n8498), .ZN(n7704) );
  NAND2_X1 U10015 ( .A1(n8490), .A2(n7701), .ZN(n8493) );
  OAI21_X1 U10016 ( .B1(n8107), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7703) );
  INV_X1 U10017 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U10018 ( .A(n7703), .B(n7702), .ZN(n8112) );
  AND2_X2 U10019 ( .A1(n7704), .A2(n8506), .ZN(P3_U3897) );
  NOR2_X1 U10020 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7708) );
  NOR2_X1 U10021 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7712) );
  INV_X1 U10022 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7718) );
  OAI21_X1 U10023 ( .B1(n7970), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7719) );
  XNOR2_X1 U10024 ( .A(n7719), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7972) );
  INV_X1 U10025 ( .A(n7972), .ZN(n9062) );
  NOR2_X1 U10026 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n7722) );
  NOR2_X1 U10027 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n7721) );
  NOR2_X1 U10028 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n7720) );
  NAND2_X1 U10029 ( .A1(n9171), .A2(n7725), .ZN(n7728) );
  NOR3_X1 U10030 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(P1_IR_REG_24__SCAN_IN), .ZN(n7724) );
  INV_X1 U10031 ( .A(n7974), .ZN(n7726) );
  NAND2_X1 U10032 ( .A1(n7726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7727) );
  XNOR2_X1 U10033 ( .A(n7727), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10034 ( .A1(n7728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7729) );
  MUX2_X1 U10035 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7729), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n7731) );
  AND2_X2 U10036 ( .A1(n8187), .A2(n8214), .ZN(P1_U4016) );
  OAI21_X1 U10037 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(n8341), .A(n7871), .ZN(
        n7738) );
  MUX2_X1 U10038 ( .A(n7738), .B(SI_0_), .S(n6641), .Z(n8511) );
  NAND2_X1 U10039 ( .A1(n8511), .A2(P3_U3151), .ZN(n7739) );
  OAI21_X1 U10040 ( .B1(n7132), .B2(P3_U3151), .A(n7739), .ZN(P3_U3295) );
  NAND2_X1 U10041 ( .A1(n7737), .A2(P2_U3088), .ZN(n13681) );
  INV_X1 U10042 ( .A(SI_0_), .ZN(n8209) );
  INV_X1 U10043 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U10044 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  NAND2_X1 U10045 ( .A1(n7749), .A2(n7744), .ZN(n8614) );
  INV_X1 U10046 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U10047 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7745) );
  XNOR2_X1 U10048 ( .A(n7746), .B(n7745), .ZN(n8395) );
  OAI222_X1 U10049 ( .A1(n13681), .A2(n8347), .B1(n13675), .B2(n8614), .C1(
        n8395), .C2(P2_U3088), .ZN(P2_U3326) );
  AND2_X1 U10050 ( .A1(n7737), .A2(P1_U3086), .ZN(n10551) );
  INV_X2 U10051 ( .A(n10551), .ZN(n14373) );
  NAND2_X1 U10052 ( .A1(n7747), .A2(SI_2_), .ZN(n7752) );
  OAI21_X1 U10053 ( .B1(n7747), .B2(SI_2_), .A(n7752), .ZN(n7759) );
  INV_X1 U10054 ( .A(n7759), .ZN(n7751) );
  NAND2_X1 U10055 ( .A1(n7751), .A2(n7750), .ZN(n7760) );
  NAND2_X1 U10056 ( .A1(n7760), .A2(n7752), .ZN(n7756) );
  INV_X1 U10057 ( .A(n7756), .ZN(n7753) );
  NAND2_X1 U10058 ( .A1(n7753), .A2(n7754), .ZN(n7757) );
  INV_X1 U10059 ( .A(n7754), .ZN(n7755) );
  NAND2_X1 U10060 ( .A1(n7756), .A2(n7755), .ZN(n7815) );
  NAND2_X1 U10061 ( .A1(n7757), .A2(n7815), .ZN(n8840) );
  NAND2_X1 U10062 ( .A1(n7809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7758) );
  XNOR2_X1 U10063 ( .A(n7758), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13853) );
  INV_X1 U10064 ( .A(n13853), .ZN(n8049) );
  OAI222_X1 U10065 ( .A1(n14370), .A2(n7775), .B1(n14373), .B2(n8840), .C1(
        P1_U3086), .C2(n8049), .ZN(P1_U3352) );
  NAND2_X1 U10066 ( .A1(n7761), .A2(n7760), .ZN(n8727) );
  NOR2_X1 U10067 ( .A1(n7766), .A2(n7917), .ZN(n7762) );
  MUX2_X1 U10068 ( .A(n7917), .B(n7762), .S(P1_IR_REG_2__SCAN_IN), .Z(n7763)
         );
  INV_X1 U10069 ( .A(n7763), .ZN(n7764) );
  NAND2_X1 U10070 ( .A1(n7764), .A2(n7809), .ZN(n8607) );
  OAI222_X1 U10071 ( .A1(n14370), .A2(n8606), .B1(n14373), .B2(n8727), .C1(
        P1_U3086), .C2(n8607), .ZN(P1_U3353) );
  NAND2_X1 U10072 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14654), .ZN(n7765) );
  MUX2_X1 U10073 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7765), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7768) );
  INV_X1 U10074 ( .A(n7766), .ZN(n7767) );
  NAND2_X1 U10075 ( .A1(n7768), .A2(n7767), .ZN(n8615) );
  OAI222_X1 U10076 ( .A1(n14370), .A2(n7457), .B1(n14373), .B2(n8614), .C1(
        P1_U3086), .C2(n8615), .ZN(P1_U3354) );
  INV_X1 U10077 ( .A(n7871), .ZN(n7769) );
  XNOR2_X1 U10078 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7872) );
  NAND2_X1 U10079 ( .A1(n7769), .A2(n7872), .ZN(n7771) );
  NAND2_X1 U10080 ( .A1(n8347), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U10081 ( .A1(n8606), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10082 ( .A1(n7789), .A2(n7788), .ZN(n7774) );
  NAND2_X1 U10083 ( .A1(n7775), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10084 ( .A1(n7795), .A2(n7794), .ZN(n7778) );
  NAND2_X1 U10085 ( .A1(n7821), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7779) );
  XNOR2_X1 U10086 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7782) );
  XNOR2_X1 U10087 ( .A(n7837), .B(n7782), .ZN(n9415) );
  NOR2_X1 U10088 ( .A1(n6641), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12979) );
  INV_X1 U10089 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12981) );
  NOR2_X1 U10090 ( .A1(n7805), .A2(n12981), .ZN(n7783) );
  MUX2_X1 U10091 ( .A(n12981), .B(n7783), .S(P3_IR_REG_5__SCAN_IN), .Z(n7784)
         );
  INV_X1 U10092 ( .A(n7784), .ZN(n7786) );
  NAND2_X1 U10093 ( .A1(n7805), .A2(n7785), .ZN(n7939) );
  NAND2_X1 U10094 ( .A1(n7786), .A2(n7939), .ZN(n15016) );
  INV_X1 U10095 ( .A(n15016), .ZN(n10137) );
  AND2_X1 U10096 ( .A1(n6641), .A2(P3_U3151), .ZN(n8458) );
  AOI222_X1 U10097 ( .A1(n9415), .A2(n12979), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10137), .C1(SI_5_), .C2(n8458), .ZN(n7787) );
  INV_X1 U10098 ( .A(n7787), .ZN(P3_U3290) );
  XNOR2_X1 U10099 ( .A(n7789), .B(n7788), .ZN(n8955) );
  INV_X1 U10100 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7791) );
  INV_X1 U10101 ( .A(n10129), .ZN(n10072) );
  AOI222_X1 U10102 ( .A1(n8955), .A2(n12979), .B1(n10072), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n8458), .C2(SI_2_), .ZN(n7793) );
  INV_X1 U10103 ( .A(n7793), .ZN(P3_U3293) );
  XNOR2_X1 U10104 ( .A(n7795), .B(n7794), .ZN(n9040) );
  INV_X1 U10105 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10106 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7796), .ZN(n7797) );
  XNOR2_X1 U10107 ( .A(n7798), .B(n7797), .ZN(n14979) );
  INV_X1 U10108 ( .A(n14979), .ZN(n10089) );
  AOI222_X1 U10109 ( .A1(n9040), .A2(n12979), .B1(n8458), .B2(SI_3_), .C1(
        n10089), .C2(P3_STATE_REG_SCAN_IN), .ZN(n7799) );
  INV_X1 U10110 ( .A(n7799), .ZN(P3_U3292) );
  XNOR2_X1 U10111 ( .A(n7801), .B(n7800), .ZN(n9230) );
  NOR2_X1 U10112 ( .A1(n7802), .A2(n12981), .ZN(n7803) );
  MUX2_X1 U10113 ( .A(n12981), .B(n7803), .S(P3_IR_REG_4__SCAN_IN), .Z(n7804)
         );
  INV_X1 U10114 ( .A(n7804), .ZN(n7807) );
  INV_X1 U10115 ( .A(n7805), .ZN(n7806) );
  INV_X1 U10116 ( .A(n14997), .ZN(n10095) );
  AOI222_X1 U10117 ( .A1(n9230), .A2(n12979), .B1(n10095), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n8458), .ZN(n7808) );
  INV_X1 U10118 ( .A(n7808), .ZN(P3_U3291) );
  NAND2_X1 U10119 ( .A1(n7811), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7810) );
  MUX2_X1 U10120 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7810), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7813) );
  INV_X1 U10121 ( .A(n7856), .ZN(n7812) );
  AND2_X1 U10122 ( .A1(n7813), .A2(n7812), .ZN(n13870) );
  INV_X1 U10123 ( .A(n13870), .ZN(n7822) );
  NAND2_X1 U10124 ( .A1(n7815), .A2(n7814), .ZN(n7819) );
  MUX2_X1 U10125 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6641), .Z(n7816) );
  NAND2_X1 U10126 ( .A1(n7816), .A2(SI_4_), .ZN(n7858) );
  OAI21_X1 U10127 ( .B1(n7816), .B2(SI_4_), .A(n7858), .ZN(n7817) );
  INV_X1 U10128 ( .A(n7817), .ZN(n7818) );
  OR2_X1 U10129 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  NAND2_X1 U10130 ( .A1(n7819), .A2(n7818), .ZN(n7859) );
  AND2_X1 U10131 ( .A1(n7859), .A2(n7820), .ZN(n8931) );
  INV_X1 U10132 ( .A(n8931), .ZN(n7900) );
  OAI222_X1 U10133 ( .A1(P1_U3086), .A2(n7822), .B1(n14373), .B2(n7900), .C1(
        n7821), .C2(n14370), .ZN(P1_U3351) );
  INV_X1 U10134 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n7830) );
  XNOR2_X1 U10135 ( .A(n10474), .B(P3_B_REG_SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10136 ( .A1(n7823), .A2(n10564), .ZN(n7824) );
  NAND2_X1 U10137 ( .A1(n8475), .A2(n7830), .ZN(n7827) );
  INV_X1 U10138 ( .A(n7825), .ZN(n10586) );
  NAND2_X1 U10139 ( .A1(n10586), .A2(n10564), .ZN(n7826) );
  NAND2_X1 U10140 ( .A1(n7827), .A2(n7826), .ZN(n9704) );
  INV_X1 U10141 ( .A(n9704), .ZN(n7828) );
  NAND2_X1 U10142 ( .A1(n7828), .A2(n8506), .ZN(n7829) );
  OAI21_X1 U10143 ( .B1(n8506), .B2(n7830), .A(n7829), .ZN(P3_U3377) );
  INV_X1 U10144 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10145 ( .A1(n10586), .A2(n10474), .ZN(n7831) );
  INV_X1 U10146 ( .A(n9708), .ZN(n7833) );
  NAND2_X1 U10147 ( .A1(n7833), .A2(n8506), .ZN(n7834) );
  OAI21_X1 U10148 ( .B1(n8506), .B2(n7835), .A(n7834), .ZN(P3_U3376) );
  NAND2_X1 U10149 ( .A1(n7865), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10150 ( .A1(n15518), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10151 ( .A1(n7931), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10152 ( .A1(n7841), .A2(n7840), .ZN(n7866) );
  NAND2_X1 U10153 ( .A1(n7962), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U10154 ( .A1(n8017), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10155 ( .A1(n8014), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10156 ( .A1(n8040), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U10157 ( .A1(n8035), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7846) );
  OR2_X1 U10158 ( .A1(n7848), .A2(n7847), .ZN(n7849) );
  AND2_X1 U10159 ( .A1(n7881), .A2(n7849), .ZN(n9829) );
  NOR2_X1 U10160 ( .A1(n7886), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U10161 ( .A1(n7873), .A2(n15362), .ZN(n7851) );
  NAND2_X1 U10162 ( .A1(n7851), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7850) );
  MUX2_X1 U10163 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7850), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7852) );
  NAND2_X1 U10164 ( .A1(n7852), .A2(n7908), .ZN(n15088) );
  AOI222_X1 U10165 ( .A1(n9829), .A2(n12979), .B1(SI_9_), .B2(n8458), .C1(
        n10145), .C2(P3_STATE_REG_SCAN_IN), .ZN(n7853) );
  INV_X1 U10166 ( .A(n7853), .ZN(P3_U3286) );
  NOR2_X1 U10167 ( .A1(n7856), .A2(n7917), .ZN(n7854) );
  MUX2_X1 U10168 ( .A(n7917), .B(n7854), .S(P1_IR_REG_5__SCAN_IN), .Z(n7857)
         );
  INV_X1 U10169 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7855) );
  OR2_X1 U10170 ( .A1(n7857), .A2(n7964), .ZN(n8062) );
  NAND2_X1 U10171 ( .A1(n7859), .A2(n7858), .ZN(n7863) );
  MUX2_X1 U10172 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6641), .Z(n7860) );
  NAND2_X1 U10173 ( .A1(n7860), .A2(SI_5_), .ZN(n7919) );
  OAI21_X1 U10174 ( .B1(n7860), .B2(SI_5_), .A(n7919), .ZN(n7861) );
  INV_X1 U10175 ( .A(n7861), .ZN(n7862) );
  OR2_X1 U10176 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  NAND2_X1 U10177 ( .A1(n7920), .A2(n7864), .ZN(n9186) );
  OAI222_X1 U10178 ( .A1(P1_U3086), .A2(n8062), .B1(n14373), .B2(n9186), .C1(
        n7865), .C2(n14370), .ZN(P1_U3350) );
  NAND2_X1 U10179 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  NAND2_X1 U10180 ( .A1(n7869), .A2(n7868), .ZN(n9596) );
  INV_X1 U10181 ( .A(n8458), .ZN(n12985) );
  INV_X1 U10182 ( .A(SI_6_), .ZN(n9599) );
  NAND2_X1 U10183 ( .A1(n7939), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7870) );
  XNOR2_X1 U10184 ( .A(n7870), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10105) );
  OAI222_X1 U10185 ( .A1(n12997), .A2(n9596), .B1(n12985), .B2(n9599), .C1(
        P3_U3151), .C2(n15033), .ZN(P3_U3289) );
  XNOR2_X1 U10186 ( .A(n7871), .B(n7872), .ZN(n8746) );
  OAI222_X1 U10187 ( .A1(n12997), .A2(n8746), .B1(n12985), .B2(n7455), .C1(
        P3_U3151), .C2(n8744), .ZN(P3_U3294) );
  OR2_X1 U10188 ( .A1(n7873), .A2(n12981), .ZN(n7874) );
  XNOR2_X1 U10189 ( .A(n7874), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10114) );
  INV_X1 U10190 ( .A(SI_8_), .ZN(n9841) );
  OR2_X1 U10191 ( .A1(n7876), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U10192 ( .A1(n7878), .A2(n7877), .ZN(n9838) );
  OAI222_X1 U10193 ( .A1(P3_U3151), .A2(n15068), .B1(n12985), .B2(n9841), .C1(
        n12997), .C2(n9838), .ZN(P3_U3287) );
  NAND2_X1 U10194 ( .A1(n7908), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7879) );
  XNOR2_X1 U10195 ( .A(n7879), .B(P3_IR_REG_10__SCAN_IN), .ZN(n10178) );
  INV_X1 U10196 ( .A(n10178), .ZN(n10173) );
  NAND2_X1 U10197 ( .A1(n8421), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10198 ( .A1(n8418), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7882) );
  OR2_X1 U10199 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X1 U10200 ( .A1(n7912), .A2(n7885), .ZN(n9944) );
  OAI222_X1 U10201 ( .A1(P3_U3151), .A2(n10173), .B1(n12985), .B2(n9945), .C1(
        n12997), .C2(n9944), .ZN(P3_U3285) );
  NAND2_X1 U10202 ( .A1(n7886), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7888) );
  INV_X1 U10203 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U10204 ( .A(n7888), .B(n7887), .ZN(n15051) );
  INV_X1 U10205 ( .A(SI_7_), .ZN(n7893) );
  OR2_X1 U10206 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  NAND2_X1 U10207 ( .A1(n7892), .A2(n7891), .ZN(n9719) );
  OAI222_X1 U10208 ( .A1(P3_U3151), .A2(n15051), .B1(n12985), .B2(n7893), .C1(
        n12997), .C2(n9719), .ZN(P3_U3288) );
  INV_X1 U10209 ( .A(n13681), .ZN(n13677) );
  INV_X1 U10210 ( .A(n13677), .ZN(n11464) );
  INV_X1 U10211 ( .A(n7897), .ZN(n7895) );
  INV_X1 U10212 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10213 ( .A1(n7895), .A2(n7894), .ZN(n7927) );
  NAND2_X1 U10214 ( .A1(n7927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7896) );
  XNOR2_X1 U10215 ( .A(n7896), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8901) );
  INV_X1 U10216 ( .A(n8901), .ZN(n8446) );
  OAI222_X1 U10217 ( .A1(n11464), .A2(n15518), .B1(n13675), .B2(n9186), .C1(
        n8446), .C2(P2_U3088), .ZN(P2_U3322) );
  NAND2_X1 U10218 ( .A1(n7897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7898) );
  MUX2_X1 U10219 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7898), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7899) );
  NAND2_X1 U10220 ( .A1(n7899), .A2(n7927), .ZN(n8399) );
  OAI222_X1 U10221 ( .A1(n13681), .A2(n7901), .B1(n13675), .B2(n7900), .C1(
        n8399), .C2(P2_U3088), .ZN(P2_U3323) );
  OR2_X1 U10222 ( .A1(n7902), .A2(n8652), .ZN(n7903) );
  INV_X1 U10223 ( .A(n14760), .ZN(n7904) );
  OAI222_X1 U10224 ( .A1(n13681), .A2(n8724), .B1(n13675), .B2(n8727), .C1(
        n7904), .C2(P2_U3088), .ZN(P2_U3325) );
  NAND2_X1 U10225 ( .A1(n7905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7906) );
  XNOR2_X1 U10226 ( .A(n7906), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8773) );
  INV_X1 U10227 ( .A(n8773), .ZN(n8432) );
  OAI222_X1 U10228 ( .A1(n13681), .A2(n7907), .B1(n13675), .B2(n8840), .C1(
        n8432), .C2(P2_U3088), .ZN(P2_U3324) );
  OAI21_X1 U10229 ( .B1(n7908), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7910) );
  INV_X1 U10230 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7909) );
  XNOR2_X1 U10231 ( .A(n7910), .B(n7909), .ZN(n10451) );
  INV_X1 U10232 ( .A(SI_11_), .ZN(n8526) );
  NAND2_X1 U10233 ( .A1(n15391), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7932) );
  INV_X1 U10234 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U10235 ( .A1(n8659), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7913) );
  OR2_X1 U10236 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  NAND2_X1 U10237 ( .A1(n7933), .A2(n7916), .ZN(n10272) );
  OAI222_X1 U10238 ( .A1(P3_U3151), .A2(n10451), .B1(n12985), .B2(n8526), .C1(
        n12997), .C2(n10272), .ZN(P3_U3284) );
  OR2_X1 U10239 ( .A1(n7964), .A2(n7917), .ZN(n7918) );
  XNOR2_X1 U10240 ( .A(n7918), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9311) );
  INV_X1 U10241 ( .A(n9311), .ZN(n8101) );
  NAND2_X2 U10242 ( .A1(n7920), .A2(n7919), .ZN(n7924) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6641), .Z(n7921) );
  NAND2_X1 U10244 ( .A1(n7921), .A2(SI_6_), .ZN(n7953) );
  OAI21_X1 U10245 ( .B1(n7921), .B2(SI_6_), .A(n7953), .ZN(n7922) );
  INV_X1 U10246 ( .A(n7922), .ZN(n7923) );
  OR2_X1 U10247 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  OAI222_X1 U10248 ( .A1(P1_U3086), .A2(n8101), .B1(n14373), .B2(n9310), .C1(
        n7926), .C2(n14370), .ZN(P1_U3349) );
  INV_X1 U10249 ( .A(n7927), .ZN(n7928) );
  NAND2_X1 U10250 ( .A1(n7928), .A2(n6854), .ZN(n7960) );
  NAND2_X1 U10251 ( .A1(n7960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7929) );
  XNOR2_X1 U10252 ( .A(n7929), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14787) );
  INV_X1 U10253 ( .A(n14787), .ZN(n7930) );
  OAI222_X1 U10254 ( .A1(n13681), .A2(n7931), .B1(n13675), .B2(n9310), .C1(
        n7930), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U10255 ( .A(SI_12_), .ZN(n8800) );
  NAND2_X1 U10256 ( .A1(n8538), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10257 ( .A1(n8535), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7934) );
  OR2_X1 U10258 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  NAND2_X1 U10259 ( .A1(n8019), .A2(n7937), .ZN(n10286) );
  NOR2_X1 U10260 ( .A1(n7939), .A2(n7938), .ZN(n7942) );
  OR2_X1 U10261 ( .A1(n7942), .A2(n12981), .ZN(n7940) );
  MUX2_X1 U10262 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7940), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7943) );
  NAND2_X1 U10263 ( .A1(n7942), .A2(n7941), .ZN(n8023) );
  INV_X1 U10264 ( .A(n12460), .ZN(n12450) );
  OAI222_X1 U10265 ( .A1(n12985), .A2(n8800), .B1(n12997), .B2(n10286), .C1(
        n12450), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U10266 ( .A1(n8187), .A2(n8208), .ZN(n9615) );
  INV_X1 U10267 ( .A(n7949), .ZN(n10937) );
  NAND3_X1 U10268 ( .A1(n10937), .A2(P1_B_REG_SCAN_IN), .A3(n10754), .ZN(n7946) );
  INV_X1 U10269 ( .A(P1_B_REG_SCAN_IN), .ZN(n13898) );
  INV_X1 U10270 ( .A(n7948), .ZN(n14374) );
  AOI21_X1 U10271 ( .B1(n7944), .B2(n13898), .A(n14374), .ZN(n7945) );
  NAND2_X1 U10272 ( .A1(n7946), .A2(n7945), .ZN(n8270) );
  INV_X1 U10273 ( .A(n8270), .ZN(n7947) );
  OR2_X1 U10274 ( .A1(n9615), .A2(n7947), .ZN(n14691) );
  INV_X1 U10275 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8200) );
  OR2_X1 U10276 ( .A1(n7949), .A2(n7948), .ZN(n8267) );
  INV_X1 U10277 ( .A(n8267), .ZN(n7950) );
  AOI22_X1 U10278 ( .A1(n14691), .A2(n8200), .B1(n8187), .B2(n7950), .ZN(
        P1_U3446) );
  INV_X1 U10279 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10280 ( .A1(n10754), .A2(n14374), .ZN(n8188) );
  INV_X1 U10281 ( .A(n8188), .ZN(n7951) );
  AOI22_X1 U10282 ( .A1(n14691), .A2(n7952), .B1(n8187), .B2(n7951), .ZN(
        P1_U3445) );
  MUX2_X1 U10283 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6641), .Z(n7955) );
  NAND2_X1 U10284 ( .A1(n7955), .A2(SI_7_), .ZN(n8004) );
  OAI21_X1 U10285 ( .B1(n7955), .B2(SI_7_), .A(n8004), .ZN(n7956) );
  INV_X1 U10286 ( .A(n7956), .ZN(n7957) );
  NAND2_X1 U10287 ( .A1(n8005), .A2(n7959), .ZN(n9515) );
  OAI21_X1 U10288 ( .B1(n7960), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U10289 ( .A(n7961), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9121) );
  INV_X1 U10290 ( .A(n9121), .ZN(n8406) );
  OAI222_X1 U10291 ( .A1(n11464), .A2(n7962), .B1(n13675), .B2(n9515), .C1(
        n8406), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U10292 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10293 ( .A1(n7964), .A2(n7963), .ZN(n8015) );
  NAND2_X1 U10294 ( .A1(n8015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7965) );
  XNOR2_X1 U10295 ( .A(n7965), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9516) );
  INV_X1 U10296 ( .A(n9516), .ZN(n8074) );
  OAI222_X1 U10297 ( .A1(P1_U3086), .A2(n8074), .B1(n14373), .B2(n9515), .C1(
        n7966), .C2(n14370), .ZN(P1_U3348) );
  AND2_X1 U10298 ( .A1(n7972), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11954) );
  INV_X1 U10299 ( .A(n11954), .ZN(n11959) );
  NAND2_X1 U10300 ( .A1(n9615), .A2(n11959), .ZN(n8043) );
  INV_X1 U10301 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10302 ( .A1(n8182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7969) );
  MUX2_X1 U10303 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7969), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n7971) );
  NAND2_X1 U10304 ( .A1(n14376), .A2(n8279), .ZN(n11904) );
  OR2_X1 U10305 ( .A1(n11904), .A2(n7972), .ZN(n7977) );
  XNOR2_X2 U10306 ( .A(n7975), .B(n8169), .ZN(n11008) );
  NAND2_X1 U10307 ( .A1(n7977), .A2(n11578), .ZN(n8041) );
  AND2_X1 U10308 ( .A1(n8043), .A2(n8041), .ZN(n14656) );
  NOR2_X1 U10309 ( .A1(n14656), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U10310 ( .A(n8506), .ZN(n7978) );
  OR2_X1 U10311 ( .A1(n7978), .A2(n8475), .ZN(n15233) );
  INV_X2 U10312 ( .A(n15233), .ZN(n8003) );
  INV_X1 U10313 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n7979) );
  NOR2_X1 U10314 ( .A1(n8003), .A2(n7979), .ZN(P3_U3253) );
  INV_X1 U10315 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n7980) );
  NOR2_X1 U10316 ( .A1(n8003), .A2(n7980), .ZN(P3_U3255) );
  INV_X1 U10317 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n7981) );
  NOR2_X1 U10318 ( .A1(n8003), .A2(n7981), .ZN(P3_U3252) );
  INV_X1 U10319 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n7982) );
  NOR2_X1 U10320 ( .A1(n8003), .A2(n7982), .ZN(P3_U3256) );
  INV_X1 U10321 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n7983) );
  NOR2_X1 U10322 ( .A1(n8003), .A2(n7983), .ZN(P3_U3257) );
  INV_X1 U10323 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U10324 ( .A1(n8003), .A2(n15333), .ZN(P3_U3254) );
  INV_X1 U10325 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n7984) );
  NOR2_X1 U10326 ( .A1(n8003), .A2(n7984), .ZN(P3_U3243) );
  INV_X1 U10327 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n7985) );
  NOR2_X1 U10328 ( .A1(n8003), .A2(n7985), .ZN(P3_U3242) );
  INV_X1 U10329 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n7986) );
  NOR2_X1 U10330 ( .A1(n8003), .A2(n7986), .ZN(P3_U3241) );
  INV_X1 U10331 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n7987) );
  NOR2_X1 U10332 ( .A1(n8003), .A2(n7987), .ZN(P3_U3258) );
  INV_X1 U10333 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n7988) );
  NOR2_X1 U10334 ( .A1(n8003), .A2(n7988), .ZN(P3_U3239) );
  INV_X1 U10335 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U10336 ( .A1(n8003), .A2(n15349), .ZN(P3_U3238) );
  INV_X1 U10337 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n7989) );
  NOR2_X1 U10338 ( .A1(n8003), .A2(n7989), .ZN(P3_U3237) );
  INV_X1 U10339 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n7990) );
  NOR2_X1 U10340 ( .A1(n8003), .A2(n7990), .ZN(P3_U3236) );
  INV_X1 U10341 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n7991) );
  NOR2_X1 U10342 ( .A1(n8003), .A2(n7991), .ZN(P3_U3235) );
  INV_X1 U10343 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n7992) );
  NOR2_X1 U10344 ( .A1(n8003), .A2(n7992), .ZN(P3_U3234) );
  INV_X1 U10345 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n7993) );
  NOR2_X1 U10346 ( .A1(n8003), .A2(n7993), .ZN(P3_U3259) );
  INV_X1 U10347 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15406) );
  NOR2_X1 U10348 ( .A1(n8003), .A2(n15406), .ZN(P3_U3260) );
  INV_X1 U10349 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n7994) );
  NOR2_X1 U10350 ( .A1(n8003), .A2(n7994), .ZN(P3_U3261) );
  INV_X1 U10351 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U10352 ( .A1(n8003), .A2(n15377), .ZN(P3_U3263) );
  INV_X1 U10353 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n7995) );
  NOR2_X1 U10354 ( .A1(n8003), .A2(n7995), .ZN(P3_U3251) );
  INV_X1 U10355 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n7996) );
  NOR2_X1 U10356 ( .A1(n8003), .A2(n7996), .ZN(P3_U3250) );
  INV_X1 U10357 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n7997) );
  NOR2_X1 U10358 ( .A1(n8003), .A2(n7997), .ZN(P3_U3249) );
  INV_X1 U10359 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n15321) );
  NOR2_X1 U10360 ( .A1(n8003), .A2(n15321), .ZN(P3_U3248) );
  INV_X1 U10361 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n7998) );
  NOR2_X1 U10362 ( .A1(n8003), .A2(n7998), .ZN(P3_U3247) );
  INV_X1 U10363 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n7999) );
  NOR2_X1 U10364 ( .A1(n8003), .A2(n7999), .ZN(P3_U3246) );
  INV_X1 U10365 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n8000) );
  NOR2_X1 U10366 ( .A1(n8003), .A2(n8000), .ZN(P3_U3245) );
  INV_X1 U10367 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n8001) );
  NOR2_X1 U10368 ( .A1(n8003), .A2(n8001), .ZN(P3_U3244) );
  INV_X1 U10369 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n8002) );
  NOR2_X1 U10370 ( .A1(n8003), .A2(n8002), .ZN(P3_U3262) );
  MUX2_X1 U10371 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6641), .Z(n8006) );
  OAI21_X1 U10372 ( .B1(n8006), .B2(SI_8_), .A(n8027), .ZN(n8007) );
  INV_X1 U10373 ( .A(n8007), .ZN(n8008) );
  OR2_X1 U10374 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  NAND2_X1 U10375 ( .A1(n8028), .A2(n8010), .ZN(n9791) );
  OR2_X1 U10376 ( .A1(n8011), .A2(n8652), .ZN(n8012) );
  XNOR2_X1 U10377 ( .A(n8012), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14800) );
  INV_X1 U10378 ( .A(n14800), .ZN(n8013) );
  OAI222_X1 U10379 ( .A1(n13681), .A2(n8014), .B1(n13675), .B2(n9791), .C1(
        n8013), .C2(P2_U3088), .ZN(P2_U3319) );
  NAND2_X1 U10380 ( .A1(n8036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8016) );
  XNOR2_X1 U10381 ( .A(n8016), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9792) );
  INV_X1 U10382 ( .A(n9792), .ZN(n8082) );
  OAI222_X1 U10383 ( .A1(P1_U3086), .A2(n8082), .B1(n14373), .B2(n9791), .C1(
        n8017), .C2(n14370), .ZN(P1_U3347) );
  INV_X1 U10384 ( .A(SI_13_), .ZN(n9082) );
  NAND2_X1 U10385 ( .A1(n8021), .A2(n10322), .ZN(n8022) );
  NAND2_X1 U10386 ( .A1(n8163), .A2(n8022), .ZN(n10294) );
  NAND2_X1 U10387 ( .A1(n8023), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8024) );
  MUX2_X1 U10388 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8024), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8026) );
  INV_X1 U10389 ( .A(n12484), .ZN(n12477) );
  OAI222_X1 U10390 ( .A1(n12985), .A2(n9082), .B1(n12997), .B2(n10294), .C1(
        n12477), .C2(P3_U3151), .ZN(P3_U3282) );
  MUX2_X1 U10391 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8346), .Z(n8029) );
  OAI21_X1 U10392 ( .B1(n8029), .B2(SI_9_), .A(n8410), .ZN(n8030) );
  INV_X1 U10393 ( .A(n8030), .ZN(n8031) );
  OR2_X1 U10394 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U10395 ( .A1(n8411), .A2(n8033), .ZN(n9964) );
  NAND2_X1 U10396 ( .A1(n8233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8034) );
  XNOR2_X1 U10397 ( .A(n8034), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9377) );
  INV_X1 U10398 ( .A(n9377), .ZN(n8889) );
  OAI222_X1 U10399 ( .A1(n13681), .A2(n8035), .B1(n13675), .B2(n9964), .C1(
        n8889), .C2(P2_U3088), .ZN(P2_U3318) );
  OR2_X1 U10400 ( .A1(n8537), .A2(n7917), .ZN(n8038) );
  INV_X1 U10401 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8037) );
  OR2_X1 U10402 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  NAND2_X1 U10403 ( .A1(n8038), .A2(n8037), .ZN(n8419) );
  INV_X1 U10404 ( .A(n9965), .ZN(n8465) );
  OAI222_X1 U10405 ( .A1(P1_U3086), .A2(n8465), .B1(n14373), .B2(n9964), .C1(
        n8040), .C2(n14370), .ZN(P1_U3346) );
  INV_X1 U10406 ( .A(n8041), .ZN(n8042) );
  NAND2_X1 U10407 ( .A1(n8043), .A2(n8042), .ZN(n14658) );
  INV_X1 U10408 ( .A(n11008), .ZN(n8636) );
  INV_X1 U10409 ( .A(n14653), .ZN(n11956) );
  INV_X1 U10410 ( .A(n13886), .ZN(n14668) );
  INV_X1 U10411 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n8631) );
  INV_X1 U10412 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U10413 ( .A(n8600), .B(P1_REG1_REG_2__SCAN_IN), .S(n8607), .Z(n8574)
         );
  XNOR2_X1 U10414 ( .A(n8615), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13838) );
  AND2_X1 U10415 ( .A1(n14654), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n13837) );
  NAND2_X1 U10416 ( .A1(n13838), .A2(n13837), .ZN(n13836) );
  INV_X1 U10417 ( .A(n8615), .ZN(n13835) );
  NAND2_X1 U10418 ( .A1(n13835), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U10419 ( .A1(n13836), .A2(n8044), .ZN(n8573) );
  NAND2_X1 U10420 ( .A1(n8574), .A2(n8573), .ZN(n8572) );
  OAI21_X1 U10421 ( .B1(n8600), .B2(n8607), .A(n8572), .ZN(n13846) );
  XOR2_X1 U10422 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n13853), .Z(n13847) );
  NAND2_X1 U10423 ( .A1(n13846), .A2(n13847), .ZN(n13845) );
  OAI21_X1 U10424 ( .B1(n8049), .B2(n8631), .A(n13845), .ZN(n13859) );
  XOR2_X1 U10425 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n13870), .Z(n13860) );
  INV_X1 U10426 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8938) );
  MUX2_X1 U10427 ( .A(n8938), .B(P1_REG1_REG_5__SCAN_IN), .S(n8062), .Z(n8045)
         );
  NAND2_X1 U10428 ( .A1(n8046), .A2(n8045), .ZN(n8057) );
  OAI21_X1 U10429 ( .B1(n8046), .B2(n8045), .A(n8057), .ZN(n8054) );
  OR2_X1 U10430 ( .A1(n11008), .A2(n14653), .ZN(n8047) );
  INV_X1 U10431 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8599) );
  MUX2_X1 U10432 ( .A(n8599), .B(P1_REG2_REG_2__SCAN_IN), .S(n8607), .Z(n8571)
         );
  INV_X1 U10433 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14198) );
  MUX2_X1 U10434 ( .A(n14198), .B(P1_REG2_REG_1__SCAN_IN), .S(n8615), .Z(
        n13840) );
  AND2_X1 U10435 ( .A1(n14654), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U10436 ( .A1(n13840), .A2(n13841), .ZN(n13839) );
  NAND2_X1 U10437 ( .A1(n13835), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10438 ( .A1(n13839), .A2(n8048), .ZN(n8570) );
  NAND2_X1 U10439 ( .A1(n8571), .A2(n8570), .ZN(n13850) );
  INV_X1 U10440 ( .A(n8607), .ZN(n8575) );
  NAND2_X1 U10441 ( .A1(n8575), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13849) );
  INV_X1 U10442 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n15504) );
  MUX2_X1 U10443 ( .A(n15504), .B(P1_REG2_REG_3__SCAN_IN), .S(n13853), .Z(
        n13848) );
  AOI21_X1 U10444 ( .B1(n13850), .B2(n13849), .A(n13848), .ZN(n13864) );
  NOR2_X1 U10445 ( .A1(n8049), .A2(n15504), .ZN(n13862) );
  INV_X1 U10446 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8853) );
  MUX2_X1 U10447 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n8853), .S(n13870), .Z(
        n13863) );
  OAI21_X1 U10448 ( .B1(n13864), .B2(n13862), .A(n13863), .ZN(n13861) );
  NAND2_X1 U10449 ( .A1(n13870), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8051) );
  INV_X1 U10450 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n15340) );
  MUX2_X1 U10451 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n15340), .S(n8062), .Z(n8050) );
  AOI21_X1 U10452 ( .B1(n13861), .B2(n8051), .A(n8050), .ZN(n8093) );
  AND3_X1 U10453 ( .A1(n13861), .A2(n8051), .A3(n8050), .ZN(n8052) );
  NOR3_X1 U10454 ( .A1(n13867), .A2(n8093), .A3(n8052), .ZN(n8053) );
  AOI21_X1 U10455 ( .B1(n14668), .B2(n8054), .A(n8053), .ZN(n8056) );
  NOR2_X1 U10456 ( .A1(n8939), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9209) );
  AOI21_X1 U10457 ( .B1(n14656), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9209), .ZN(
        n8055) );
  OAI211_X1 U10458 ( .C1(n8062), .C2(n13885), .A(n8056), .B(n8055), .ZN(
        P1_U3248) );
  INV_X1 U10459 ( .A(n8062), .ZN(n9187) );
  OAI21_X1 U10460 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9187), .A(n8057), .ZN(
        n8088) );
  INV_X1 U10461 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n8058) );
  MUX2_X1 U10462 ( .A(n8058), .B(P1_REG1_REG_6__SCAN_IN), .S(n9311), .Z(n8089)
         );
  NOR2_X1 U10463 ( .A1(n8088), .A2(n8089), .ZN(n8087) );
  AOI21_X1 U10464 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9311), .A(n8087), .ZN(
        n8061) );
  INV_X1 U10465 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8059) );
  MUX2_X1 U10466 ( .A(n8059), .B(P1_REG1_REG_7__SCAN_IN), .S(n9516), .Z(n8060)
         );
  NOR2_X1 U10467 ( .A1(n8061), .A2(n8060), .ZN(n8070) );
  AOI211_X1 U10468 ( .C1(n8061), .C2(n8060), .A(n13886), .B(n8070), .ZN(n8069)
         );
  NOR2_X1 U10469 ( .A1(n8062), .A2(n15340), .ZN(n8092) );
  INV_X1 U10470 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9201) );
  MUX2_X1 U10471 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9201), .S(n9311), .Z(n8091)
         );
  OAI21_X1 U10472 ( .B1(n8093), .B2(n8092), .A(n8091), .ZN(n8090) );
  NAND2_X1 U10473 ( .A1(n9311), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8064) );
  INV_X1 U10474 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8073) );
  MUX2_X1 U10475 ( .A(n8073), .B(P1_REG2_REG_7__SCAN_IN), .S(n9516), .Z(n8063)
         );
  AOI21_X1 U10476 ( .B1(n8090), .B2(n8064), .A(n8063), .ZN(n8077) );
  AND3_X1 U10477 ( .A1(n8090), .A2(n8064), .A3(n8063), .ZN(n8065) );
  NOR3_X1 U10478 ( .A1(n13867), .A2(n8077), .A3(n8065), .ZN(n8068) );
  NAND2_X1 U10479 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9534) );
  NAND2_X1 U10480 ( .A1(n14656), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n8066) );
  OAI211_X1 U10481 ( .C1(n13885), .C2(n8074), .A(n9534), .B(n8066), .ZN(n8067)
         );
  OR3_X1 U10482 ( .A1(n8069), .A2(n8068), .A3(n8067), .ZN(P1_U3250) );
  AOI21_X1 U10483 ( .B1(n9516), .B2(P1_REG1_REG_7__SCAN_IN), .A(n8070), .ZN(
        n8072) );
  INV_X1 U10484 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9526) );
  MUX2_X1 U10485 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9526), .S(n9792), .Z(n8071)
         );
  NAND2_X1 U10486 ( .A1(n8072), .A2(n8071), .ZN(n8152) );
  OAI21_X1 U10487 ( .B1(n8072), .B2(n8071), .A(n8152), .ZN(n8085) );
  NOR2_X1 U10488 ( .A1(n8074), .A2(n8073), .ZN(n8076) );
  INV_X1 U10489 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U10490 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10048), .S(n9792), .Z(n8075) );
  OAI21_X1 U10491 ( .B1(n8077), .B2(n8076), .A(n8075), .ZN(n8150) );
  INV_X1 U10492 ( .A(n8150), .ZN(n8079) );
  NOR3_X1 U10493 ( .A1(n8077), .A2(n8076), .A3(n8075), .ZN(n8078) );
  NOR3_X1 U10494 ( .A1(n8079), .A2(n8078), .A3(n13867), .ZN(n8084) );
  NOR2_X1 U10495 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9527), .ZN(n8080) );
  AOI21_X1 U10496 ( .B1(n14656), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n8080), .ZN(
        n8081) );
  OAI21_X1 U10497 ( .B1(n13885), .B2(n8082), .A(n8081), .ZN(n8083) );
  AOI211_X1 U10498 ( .C1(n8085), .C2(n14668), .A(n8084), .B(n8083), .ZN(n8086)
         );
  INV_X1 U10499 ( .A(n8086), .ZN(P1_U3251) );
  AOI211_X1 U10500 ( .C1(n8089), .C2(n8088), .A(n8087), .B(n13886), .ZN(n8097)
         );
  INV_X1 U10501 ( .A(n8090), .ZN(n8095) );
  NOR3_X1 U10502 ( .A1(n8093), .A2(n8092), .A3(n8091), .ZN(n8094) );
  NOR3_X1 U10503 ( .A1(n13867), .A2(n8095), .A3(n8094), .ZN(n8096) );
  NOR2_X1 U10504 ( .A1(n8097), .A2(n8096), .ZN(n8100) );
  INV_X1 U10505 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9332) );
  NOR2_X1 U10506 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9332), .ZN(n8098) );
  AOI21_X1 U10507 ( .B1(n14656), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n8098), .ZN(
        n8099) );
  OAI211_X1 U10508 ( .C1(n8101), .C2(n13885), .A(n8100), .B(n8099), .ZN(
        P1_U3249) );
  INV_X1 U10509 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8104) );
  INV_X1 U10510 ( .A(n8125), .ZN(n8127) );
  NAND2_X4 U10511 ( .A1(n12998), .A2(n8106), .ZN(n10270) );
  NAND2_X1 U10512 ( .A1(n8493), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8110) );
  INV_X1 U10513 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10515 ( .A1(n12409), .A2(n8112), .ZN(n8111) );
  NAND2_X1 U10516 ( .A1(n10270), .A2(n8111), .ZN(n8117) );
  OR2_X1 U10517 ( .A1(n8112), .A2(P3_U3151), .ZN(n12432) );
  INV_X1 U10518 ( .A(n12432), .ZN(n8113) );
  NOR2_X1 U10519 ( .A1(n8713), .A2(n8113), .ZN(n8116) );
  NOR2_X1 U10520 ( .A1(n8117), .A2(n8116), .ZN(n8119) );
  INV_X1 U10521 ( .A(n12998), .ZN(n12109) );
  NAND2_X1 U10522 ( .A1(n12109), .A2(n12426), .ZN(n8757) );
  INV_X1 U10523 ( .A(n8757), .ZN(n8114) );
  NAND2_X1 U10524 ( .A1(n8119), .A2(n8114), .ZN(n15099) );
  INV_X1 U10525 ( .A(n15099), .ZN(n12588) );
  NAND2_X1 U10526 ( .A1(n8119), .A2(n6648), .ZN(n12616) );
  AND2_X1 U10527 ( .A1(P3_U3897), .A2(n12998), .ZN(n15084) );
  NOR3_X1 U10528 ( .A1(n12588), .A2(n15095), .A3(n15084), .ZN(n8123) );
  MUX2_X1 U10529 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n6648), .Z(n8115) );
  NOR2_X1 U10530 ( .A1(n8115), .A2(n7132), .ZN(n8286) );
  AOI21_X1 U10531 ( .B1(n7132), .B2(n8115), .A(n8286), .ZN(n8122) );
  INV_X1 U10532 ( .A(n8116), .ZN(n8118) );
  AOI22_X1 U10533 ( .A1(n15092), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n8121) );
  MUX2_X1 U10534 ( .A(P3_U3897), .B(n8119), .S(n12998), .Z(n12613) );
  NAND2_X1 U10535 ( .A1(n12613), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8120) );
  OAI211_X1 U10536 ( .C1(n8123), .C2(n8122), .A(n8121), .B(n8120), .ZN(
        P3_U3182) );
  INV_X1 U10537 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n15402) );
  INV_X1 U10538 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10539 ( .A1(n6638), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10540 ( .A1(n10884), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10541 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8130) );
  NAND2_X1 U10542 ( .A1(n9238), .A2(n8130), .ZN(n9370) );
  NAND2_X1 U10543 ( .A1(n8514), .A2(n9370), .ZN(n8132) );
  INV_X1 U10544 ( .A(n10977), .ZN(n9240) );
  NAND2_X1 U10545 ( .A1(n9240), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8131) );
  INV_X1 U10546 ( .A(n9506), .ZN(n15115) );
  NAND2_X1 U10547 ( .A1(n15115), .A2(P3_U3897), .ZN(n8135) );
  OAI21_X1 U10548 ( .B1(P3_U3897), .B2(n15402), .A(n8135), .ZN(P3_U3495) );
  INV_X1 U10549 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15309) );
  NAND2_X1 U10550 ( .A1(n6639), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8146) );
  INV_X1 U10551 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8139) );
  INV_X1 U10552 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U10553 ( .A1(n10299), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10554 ( .A1(n8226), .A2(n8142), .ZN(n12840) );
  NAND2_X1 U10555 ( .A1(n12024), .A2(n12840), .ZN(n8145) );
  NAND2_X1 U10556 ( .A1(n6638), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U10557 ( .A1(n12222), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8143) );
  NAND4_X1 U10558 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n11974) );
  NAND2_X1 U10559 ( .A1(n11974), .A2(P3_U3897), .ZN(n8147) );
  OAI21_X1 U10560 ( .B1(P3_U3897), .B2(n15309), .A(n8147), .ZN(P3_U3505) );
  NAND2_X1 U10561 ( .A1(n9792), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8149) );
  INV_X1 U10562 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8464) );
  MUX2_X1 U10563 ( .A(n8464), .B(P1_REG2_REG_9__SCAN_IN), .S(n9965), .Z(n8148)
         );
  AOI21_X1 U10564 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8468) );
  NAND3_X1 U10565 ( .A1(n8150), .A2(n8149), .A3(n8148), .ZN(n8151) );
  NAND2_X1 U10566 ( .A1(n8151), .A2(n14669), .ZN(n8160) );
  INV_X1 U10567 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9801) );
  MUX2_X1 U10568 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9801), .S(n9965), .Z(n8154)
         );
  OAI21_X1 U10569 ( .B1(n9792), .B2(P1_REG1_REG_8__SCAN_IN), .A(n8152), .ZN(
        n8153) );
  NAND2_X1 U10570 ( .A1(n8153), .A2(n8154), .ZN(n8461) );
  OAI21_X1 U10571 ( .B1(n8154), .B2(n8153), .A(n8461), .ZN(n8155) );
  NAND2_X1 U10572 ( .A1(n8155), .A2(n14668), .ZN(n8159) );
  NOR2_X1 U10573 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10523), .ZN(n8157) );
  NOR2_X1 U10574 ( .A1(n13885), .A2(n8465), .ZN(n8156) );
  AOI211_X1 U10575 ( .C1(n14656), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n8157), .B(
        n8156), .ZN(n8158) );
  OAI211_X1 U10576 ( .C1(n8468), .C2(n8160), .A(n8159), .B(n8158), .ZN(
        P1_U3252) );
  XNOR2_X1 U10577 ( .A(n8162), .B(n8161), .ZN(n12507) );
  INV_X1 U10578 ( .A(SI_14_), .ZN(n10499) );
  INV_X1 U10579 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U10580 ( .A1(n9105), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8381) );
  INV_X1 U10581 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U10582 ( .A1(n9102), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8164) );
  OR2_X1 U10583 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  NAND2_X1 U10584 ( .A1(n8382), .A2(n8167), .ZN(n10498) );
  OAI222_X1 U10585 ( .A1(P3_U3151), .A2(n12507), .B1(n12985), .B2(n10499), 
        .C1(n12997), .C2(n10498), .ZN(P3_U3281) );
  OAI21_X2 U10586 ( .B1(n14360), .B2(P1_IR_REG_29__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8170) );
  INV_X1 U10587 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U10588 ( .A1(n14360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8171) );
  INV_X1 U10589 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U10590 ( .A1(n6643), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8180) );
  OR2_X1 U10591 ( .A1(n8852), .A2(n14198), .ZN(n8179) );
  INV_X1 U10592 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8174) );
  INV_X1 U10593 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13833) );
  NAND2_X1 U10594 ( .A1(n14192), .A2(n14591), .ZN(n14681) );
  INV_X1 U10595 ( .A(n11904), .ZN(n8637) );
  NAND2_X1 U10596 ( .A1(n6735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8181) );
  MUX2_X1 U10597 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8181), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8183) );
  NAND2_X1 U10598 ( .A1(n6734), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U10599 ( .A1(n11902), .A2(n13891), .ZN(n8186) );
  AOI21_X1 U10600 ( .B1(n8637), .B2(n8186), .A(n8214), .ZN(n9063) );
  OR2_X1 U10601 ( .A1(n8270), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8189) );
  AND2_X1 U10602 ( .A1(n8189), .A2(n8188), .ZN(n8274) );
  NOR2_X1 U10603 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .ZN(
        n8193) );
  NOR4_X1 U10604 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n8192) );
  NOR4_X1 U10605 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8191) );
  NOR4_X1 U10606 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n8190) );
  AND4_X1 U10607 ( .A1(n8193), .A2(n8192), .A3(n8191), .A4(n8190), .ZN(n8199)
         );
  NOR4_X1 U10608 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8197) );
  NOR4_X1 U10609 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8196) );
  NOR4_X1 U10610 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n8195) );
  NOR4_X1 U10611 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8194) );
  AND4_X1 U10612 ( .A1(n8197), .A2(n8196), .A3(n8195), .A4(n8194), .ZN(n8198)
         );
  NAND2_X1 U10613 ( .A1(n8199), .A2(n8198), .ZN(n8268) );
  NOR2_X1 U10614 ( .A1(n8268), .A2(n8200), .ZN(n8201) );
  OR2_X1 U10615 ( .A1(n8270), .A2(n8201), .ZN(n8202) );
  INV_X1 U10616 ( .A(n13818), .ZN(n13776) );
  NOR2_X1 U10617 ( .A1(n11901), .A2(n8214), .ZN(n8605) );
  NAND2_X1 U10618 ( .A1(n6644), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8207) );
  INV_X1 U10619 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14682) );
  OR2_X1 U10620 ( .A1(n11704), .A2(n14682), .ZN(n8206) );
  INV_X1 U10621 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8203) );
  OR2_X1 U10622 ( .A1(n8852), .A2(n8203), .ZN(n8205) );
  INV_X1 U10623 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14652) );
  OR2_X1 U10624 ( .A1(n11881), .A2(n14652), .ZN(n8204) );
  INV_X1 U10625 ( .A(n14654), .ZN(n8567) );
  NOR2_X1 U10626 ( .A1(n6641), .A2(n8209), .ZN(n8210) );
  XNOR2_X1 U10627 ( .A(n8210), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14377) );
  MUX2_X1 U10628 ( .A(n8567), .B(n14377), .S(n11578), .Z(n14189) );
  INV_X1 U10629 ( .A(n14189), .ZN(n14678) );
  NAND2_X1 U10630 ( .A1(n14195), .A2(n10521), .ZN(n8216) );
  NAND2_X1 U10631 ( .A1(n8214), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8215) );
  OAI211_X1 U10632 ( .C1(n7432), .C2(n14189), .A(n8216), .B(n8215), .ZN(n8613)
         );
  OAI21_X1 U10633 ( .B1(n8217), .B2(n8613), .A(n8612), .ZN(n8565) );
  INV_X1 U10634 ( .A(n9615), .ZN(n9211) );
  AND3_X1 U10635 ( .A1(n9612), .A2(n8274), .A3(n11904), .ZN(n8219) );
  OR2_X1 U10636 ( .A1(n14676), .A2(n11902), .ZN(n14675) );
  OR2_X1 U10637 ( .A1(n14676), .A2(n13891), .ZN(n8218) );
  NAND3_X1 U10638 ( .A1(n9211), .A2(n8219), .A3(n14717), .ZN(n14574) );
  NAND2_X1 U10639 ( .A1(n8565), .A2(n14567), .ZN(n8223) );
  NAND2_X1 U10640 ( .A1(n9612), .A2(n8274), .ZN(n8220) );
  NAND2_X1 U10641 ( .A1(n9616), .A2(n8220), .ZN(n9210) );
  NOR2_X1 U10642 ( .A1(n14717), .A2(n9615), .ZN(n8221) );
  NAND2_X1 U10643 ( .A1(n9210), .A2(n11957), .ZN(n8663) );
  AOI22_X1 U10644 ( .A1(n13798), .A2(n14678), .B1(n8663), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n8222) );
  OAI211_X1 U10645 ( .C1(n14681), .C2(n13776), .A(n8223), .B(n8222), .ZN(
        P1_U3232) );
  INV_X1 U10646 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15341) );
  NAND2_X1 U10647 ( .A1(n6638), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U10648 ( .A1(n6639), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8230) );
  INV_X1 U10649 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10650 ( .A1(n8226), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10651 ( .A1(n10572), .A2(n8227), .ZN(n12828) );
  NAND2_X1 U10652 ( .A1(n12024), .A2(n12828), .ZN(n8229) );
  NAND2_X1 U10653 ( .A1(n12222), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8228) );
  INV_X1 U10654 ( .A(n12836), .ZN(n12806) );
  NAND2_X1 U10655 ( .A1(n12806), .A2(P3_U3897), .ZN(n8232) );
  OAI21_X1 U10656 ( .B1(P3_U3897), .B2(n15341), .A(n8232), .ZN(P3_U3506) );
  INV_X1 U10657 ( .A(n8234), .ZN(n9071) );
  INV_X1 U10658 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n15363) );
  INV_X1 U10659 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8238) );
  INV_X1 U10660 ( .A(n11315), .ZN(n11458) );
  NOR2_X1 U10661 ( .A1(n8241), .A2(n8652), .ZN(n8244) );
  NAND2_X1 U10662 ( .A1(n8652), .A2(n8242), .ZN(n8243) );
  NAND2_X1 U10663 ( .A1(n8327), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8246) );
  INV_X1 U10664 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8245) );
  XNOR2_X2 U10665 ( .A(n8246), .B(n8245), .ZN(n8249) );
  INV_X1 U10666 ( .A(n10321), .ZN(n8723) );
  AOI21_X1 U10667 ( .B1(n8366), .B2(n10548), .A(n11169), .ZN(n8248) );
  INV_X1 U10668 ( .A(n8249), .ZN(n8360) );
  NOR2_X1 U10669 ( .A1(n8249), .A2(P2_U3088), .ZN(n13676) );
  AND2_X1 U10670 ( .A1(n8258), .A2(n13676), .ZN(n8251) );
  INV_X1 U10671 ( .A(n11000), .ZN(n13235) );
  NAND2_X1 U10672 ( .A1(n8251), .A2(n13235), .ZN(n14802) );
  AND2_X1 U10673 ( .A1(n8251), .A2(n11000), .ZN(n13225) );
  INV_X1 U10674 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U10675 ( .A1(n13225), .A2(n8252), .ZN(n8254) );
  AND2_X1 U10676 ( .A1(n8249), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8253) );
  NAND2_X1 U10677 ( .A1(n8258), .A2(n8253), .ZN(n14846) );
  OAI211_X1 U10678 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14802), .A(n8254), .B(
        n14846), .ZN(n8255) );
  INV_X1 U10679 ( .A(n8255), .ZN(n8257) );
  INV_X1 U10680 ( .A(n14802), .ZN(n14856) );
  AOI22_X1 U10681 ( .A1(n14856), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n13225), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n8256) );
  INV_X1 U10682 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8343) );
  MUX2_X1 U10683 ( .A(n8257), .B(n8256), .S(n8343), .Z(n8260) );
  NOR2_X2 U10684 ( .A1(n8258), .A2(P2_U3088), .ZN(n14840) );
  AOI22_X1 U10685 ( .A1(n14840), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n8259) );
  NAND2_X1 U10686 ( .A1(n8260), .A2(n8259), .ZN(P2_U3214) );
  INV_X1 U10687 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15491) );
  NAND2_X1 U10688 ( .A1(n6638), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10689 ( .A1(n6639), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U10690 ( .A1(n9861), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10691 ( .A1(n10273), .A2(n8261), .ZN(n10737) );
  NAND2_X1 U10692 ( .A1(n12024), .A2(n10737), .ZN(n8263) );
  NAND2_X1 U10693 ( .A1(n12222), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10694 ( .A1(n10761), .A2(P3_U3897), .ZN(n8266) );
  OAI21_X1 U10695 ( .B1(P3_U3897), .B2(n15491), .A(n8266), .ZN(P3_U3502) );
  OAI21_X1 U10696 ( .B1(n8270), .B2(P1_D_REG_1__SCAN_IN), .A(n8267), .ZN(n8272) );
  INV_X1 U10697 ( .A(n8268), .ZN(n8269) );
  OR2_X1 U10698 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  AND2_X1 U10699 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  AND2_X1 U10700 ( .A1(n9616), .A2(n8273), .ZN(n8687) );
  INV_X1 U10701 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15449) );
  INV_X1 U10702 ( .A(n11901), .ZN(n8277) );
  OR2_X1 U10703 ( .A1(n8275), .A2(n14677), .ZN(n8276) );
  NAND2_X1 U10704 ( .A1(n11901), .A2(n14376), .ZN(n8278) );
  OR2_X1 U10705 ( .A1(n8275), .A2(n13891), .ZN(n8280) );
  NAND2_X1 U10706 ( .A1(n8279), .A2(n11907), .ZN(n11714) );
  NAND2_X1 U10707 ( .A1(n14195), .A2(n14678), .ZN(n14203) );
  NAND2_X1 U10708 ( .A1(n14203), .A2(n8281), .ZN(n11917) );
  INV_X1 U10709 ( .A(n11917), .ZN(n8282) );
  OAI21_X1 U10710 ( .B1(n14725), .B2(n14592), .A(n8282), .ZN(n14685) );
  OAI211_X1 U10711 ( .C1(n14189), .C2(n14676), .A(n14685), .B(n14681), .ZN(
        n14310) );
  NAND2_X1 U10712 ( .A1(n14310), .A2(n14733), .ZN(n8283) );
  OAI21_X1 U10713 ( .B1(n14733), .B2(n15449), .A(n8283), .ZN(P1_U3459) );
  INV_X1 U10714 ( .A(n12613), .ZN(n15089) );
  MUX2_X1 U10715 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6648), .Z(n8284) );
  NOR2_X1 U10716 ( .A1(n8284), .A2(n8744), .ZN(n8555) );
  AOI21_X1 U10717 ( .B1(n8284), .B2(n8744), .A(n8555), .ZN(n8285) );
  NAND2_X1 U10718 ( .A1(n8285), .A2(n8286), .ZN(n8561) );
  OAI21_X1 U10719 ( .B1(n8286), .B2(n8285), .A(n8561), .ZN(n8298) );
  AND2_X1 U10720 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n7132), .ZN(n8288) );
  INV_X1 U10721 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8287) );
  OR3_X1 U10722 ( .A1(n8287), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8544) );
  OAI21_X1 U10723 ( .B1(n8744), .B2(n8288), .A(n8544), .ZN(n8289) );
  INV_X1 U10724 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U10725 ( .A1(n8289), .A2(n15218), .ZN(n8290) );
  AND2_X1 U10726 ( .A1(n8545), .A2(n8290), .ZN(n8292) );
  AOI22_X1 U10727 ( .A1(n15092), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n8291) );
  OAI21_X1 U10728 ( .B1(n8292), .B2(n12616), .A(n8291), .ZN(n8297) );
  AND2_X1 U10729 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n7132), .ZN(n8293) );
  NAND2_X1 U10730 ( .A1(n7790), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8540) );
  INV_X1 U10731 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15164) );
  OR2_X1 U10732 ( .A1(n8294), .A2(n15164), .ZN(n8541) );
  NAND2_X1 U10733 ( .A1(n8294), .A2(n15164), .ZN(n8295) );
  AOI21_X1 U10734 ( .B1(n8541), .B2(n8295), .A(n15099), .ZN(n8296) );
  AOI211_X1 U10735 ( .C1(n15084), .C2(n8298), .A(n8297), .B(n8296), .ZN(n8299)
         );
  OAI21_X1 U10736 ( .B1(n8744), .B2(n15089), .A(n8299), .ZN(P3_U3183) );
  INV_X1 U10737 ( .A(P2_B_REG_SCAN_IN), .ZN(n15460) );
  XOR2_X1 U10738 ( .A(n10753), .B(n15460), .Z(n8300) );
  NAND2_X1 U10739 ( .A1(n10935), .A2(n8300), .ZN(n8301) );
  INV_X1 U10740 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14908) );
  NAND2_X1 U10741 ( .A1(n14875), .A2(n14908), .ZN(n8304) );
  INV_X1 U10742 ( .A(n8302), .ZN(n13683) );
  NAND2_X1 U10743 ( .A1(n13683), .A2(n10935), .ZN(n8303) );
  NOR4_X1 U10744 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8313) );
  INV_X1 U10745 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14894) );
  INV_X1 U10746 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15320) );
  INV_X1 U10747 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15478) );
  INV_X1 U10748 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15483) );
  NAND4_X1 U10749 ( .A1(n14894), .A2(n15320), .A3(n15478), .A4(n15483), .ZN(
        n8310) );
  NOR4_X1 U10750 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8308) );
  NOR4_X1 U10751 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n8307) );
  NOR4_X1 U10752 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8306) );
  NOR4_X1 U10753 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8305) );
  NAND4_X1 U10754 ( .A1(n8308), .A2(n8307), .A3(n8306), .A4(n8305), .ZN(n8309)
         );
  NOR4_X1 U10755 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8310), .A4(n8309), .ZN(n8312) );
  NOR4_X1 U10756 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8311) );
  NAND3_X1 U10757 ( .A1(n8313), .A2(n8312), .A3(n8311), .ZN(n8314) );
  NAND2_X1 U10758 ( .A1(n8314), .A2(n14875), .ZN(n8593) );
  NAND2_X1 U10759 ( .A1(n8592), .A2(n8593), .ZN(n8356) );
  INV_X1 U10760 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10761 ( .A1(n14875), .A2(n8315), .ZN(n8316) );
  NAND2_X1 U10762 ( .A1(n13683), .A2(n10753), .ZN(n14903) );
  NAND2_X1 U10763 ( .A1(n8316), .A2(n14903), .ZN(n9304) );
  INV_X1 U10764 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8317) );
  MUX2_X1 U10765 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8318), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8320) );
  NAND2_X1 U10766 ( .A1(n8320), .A2(n8319), .ZN(n11427) );
  NAND2_X1 U10767 ( .A1(n8321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8322) );
  MUX2_X1 U10768 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8322), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n8324) );
  INV_X1 U10769 ( .A(n11429), .ZN(n11449) );
  NAND2_X1 U10770 ( .A1(n11315), .A2(n11425), .ZN(n8374) );
  OAI21_X1 U10771 ( .B1(n8356), .B2(n9304), .A(n8594), .ZN(n8325) );
  NAND2_X1 U10772 ( .A1(n11427), .A2(n13227), .ZN(n11314) );
  NAND2_X1 U10773 ( .A1(n8366), .A2(n11314), .ZN(n9109) );
  NAND2_X1 U10774 ( .A1(n8325), .A2(n9109), .ZN(n8784) );
  OR2_X1 U10775 ( .A1(n8784), .A2(n14907), .ZN(n8741) );
  INV_X1 U10776 ( .A(n8741), .ZN(n8373) );
  INV_X1 U10777 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9928) );
  INV_X1 U10778 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10779 ( .A1(n8330), .A2(n8328), .ZN(n13666) );
  NAND2_X1 U10780 ( .A1(n9136), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8340) );
  INV_X1 U10781 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8332) );
  NAND2_X2 U10782 ( .A1(n13670), .A2(n13674), .ZN(n11333) );
  INV_X1 U10783 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8334) );
  INV_X1 U10784 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8336) );
  OR2_X1 U10785 ( .A1(n8786), .A2(n8336), .ZN(n8337) );
  NAND2_X1 U10786 ( .A1(n6641), .A2(SI_0_), .ZN(n8342) );
  XNOR2_X1 U10787 ( .A(n8342), .B(n8341), .ZN(n13684) );
  MUX2_X1 U10788 ( .A(n8343), .B(n13684), .S(n10321), .Z(n11028) );
  INV_X1 U10789 ( .A(n11028), .ZN(n11027) );
  AND2_X1 U10790 ( .A1(n6917), .A2(n11027), .ZN(n8583) );
  XNOR2_X1 U10791 ( .A(n11024), .B(n11315), .ZN(n8344) );
  INV_X1 U10792 ( .A(n11024), .ZN(n11390) );
  NOR2_X1 U10793 ( .A1(n13067), .A2(n11027), .ZN(n8345) );
  AOI21_X1 U10794 ( .B1(n8583), .B2(n8374), .A(n8345), .ZN(n8355) );
  INV_X1 U10795 ( .A(n8786), .ZN(n11016) );
  NAND2_X1 U10796 ( .A1(n11016), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8352) );
  INV_X1 U10797 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8348) );
  INV_X1 U10798 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8349) );
  INV_X1 U10799 ( .A(n11427), .ZN(n11396) );
  OR2_X2 U10800 ( .A1(n8374), .A2(n11396), .ZN(n13030) );
  NAND2_X1 U10801 ( .A1(n13157), .A2(n13030), .ZN(n8719) );
  NAND2_X1 U10802 ( .A1(n8354), .A2(n8355), .ZN(n8722) );
  OAI21_X1 U10803 ( .B1(n8355), .B2(n8354), .A(n8722), .ZN(n8359) );
  INV_X1 U10804 ( .A(n8356), .ZN(n9112) );
  NOR2_X1 U10805 ( .A1(n14907), .A2(n9304), .ZN(n8357) );
  AND2_X1 U10806 ( .A1(n9112), .A2(n8357), .ZN(n8368) );
  INV_X1 U10807 ( .A(n8368), .ZN(n8358) );
  NOR2_X1 U10808 ( .A1(n8358), .A2(n8366), .ZN(n8375) );
  INV_X1 U10809 ( .A(n11314), .ZN(n11455) );
  NAND2_X1 U10810 ( .A1(n8359), .A2(n13133), .ZN(n8372) );
  AND2_X2 U10811 ( .A1(n8366), .A2(n8360), .ZN(n13120) );
  INV_X1 U10812 ( .A(n13120), .ZN(n13316) );
  INV_X1 U10813 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8361) );
  OR2_X1 U10814 ( .A1(n11333), .A2(n8361), .ZN(n8365) );
  INV_X1 U10815 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9570) );
  INV_X1 U10816 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9571) );
  OR2_X1 U10817 ( .A1(n8786), .A2(n9571), .ZN(n8362) );
  INV_X1 U10818 ( .A(n13156), .ZN(n8367) );
  AND2_X2 U10819 ( .A1(n8366), .A2(n8249), .ZN(n13237) );
  INV_X1 U10820 ( .A(n13237), .ZN(n13135) );
  OAI22_X1 U10821 ( .A1(n6856), .A2(n13316), .B1(n8367), .B2(n13135), .ZN(
        n8588) );
  NAND2_X1 U10822 ( .A1(n8368), .A2(n11455), .ZN(n14554) );
  INV_X1 U10823 ( .A(n14554), .ZN(n13137) );
  INV_X1 U10824 ( .A(n8374), .ZN(n8377) );
  AND2_X1 U10825 ( .A1(n8377), .A2(n11396), .ZN(n9469) );
  NAND2_X1 U10826 ( .A1(n8368), .A2(n9469), .ZN(n8370) );
  INV_X1 U10827 ( .A(n14907), .ZN(n11456) );
  INV_X1 U10828 ( .A(n8594), .ZN(n8369) );
  NAND2_X1 U10829 ( .A1(n8370), .A2(n13515), .ZN(n13128) );
  AOI22_X1 U10830 ( .A1(n8588), .A2(n13137), .B1(n6820), .B2(n13128), .ZN(
        n8371) );
  OAI211_X1 U10831 ( .C1(n8373), .C2(n9928), .A(n8372), .B(n8371), .ZN(
        P2_U3194) );
  INV_X1 U10832 ( .A(n13128), .ZN(n14550) );
  NAND2_X1 U10833 ( .A1(n8375), .A2(n8374), .ZN(n13048) );
  NAND2_X1 U10834 ( .A1(n6917), .A2(n11028), .ZN(n9107) );
  NAND2_X1 U10835 ( .A1(n13157), .A2(n13237), .ZN(n9115) );
  OAI22_X1 U10836 ( .A1(n13048), .A2(n9107), .B1(n14554), .B2(n9115), .ZN(
        n8376) );
  AOI21_X1 U10837 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n8741), .A(n8376), .ZN(
        n8379) );
  NAND2_X1 U10838 ( .A1(n11027), .A2(n8377), .ZN(n9117) );
  INV_X1 U10839 ( .A(n9117), .ZN(n14910) );
  OAI21_X1 U10840 ( .B1(n8585), .B2(n14910), .A(n13133), .ZN(n8378) );
  OAI211_X1 U10841 ( .C1(n14550), .C2(n11028), .A(n8379), .B(n8378), .ZN(
        P2_U3204) );
  NAND2_X1 U10842 ( .A1(n6708), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8380) );
  XNOR2_X1 U10843 ( .A(n8380), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12536) );
  INV_X1 U10844 ( .A(n12536), .ZN(n12527) );
  INV_X1 U10845 ( .A(SI_15_), .ZN(n9088) );
  NAND2_X1 U10846 ( .A1(n9168), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10847 ( .A1(n9160), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8383) );
  AND2_X1 U10848 ( .A1(n8447), .A2(n8383), .ZN(n8384) );
  OR2_X1 U10849 ( .A1(n8385), .A2(n8384), .ZN(n8386) );
  NAND2_X1 U10850 ( .A1(n8448), .A2(n8386), .ZN(n10565) );
  OAI222_X1 U10851 ( .A1(P3_U3151), .A2(n12527), .B1(n12985), .B2(n9088), .C1(
        n12997), .C2(n10565), .ZN(P3_U3280) );
  XNOR2_X1 U10852 ( .A(n8395), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U10853 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14746) );
  INV_X1 U10854 ( .A(n14746), .ZN(n8387) );
  NAND2_X1 U10855 ( .A1(n14742), .A2(n8387), .ZN(n14743) );
  INV_X1 U10856 ( .A(n8395), .ZN(n14748) );
  NAND2_X1 U10857 ( .A1(n14748), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10858 ( .A1(n14743), .A2(n8388), .ZN(n14756) );
  INV_X1 U10859 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8389) );
  XNOR2_X1 U10860 ( .A(n8773), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n8423) );
  NOR2_X1 U10861 ( .A1(n8424), .A2(n8423), .ZN(n8422) );
  AOI21_X1 U10862 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n8773), .A(n8422), .ZN(
        n14770) );
  XNOR2_X1 U10863 ( .A(n14773), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n14769) );
  NOR2_X1 U10864 ( .A1(n14770), .A2(n14769), .ZN(n14768) );
  XNOR2_X1 U10865 ( .A(n8901), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n8434) );
  INV_X1 U10866 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8390) );
  MUX2_X1 U10867 ( .A(n8390), .B(P2_REG1_REG_6__SCAN_IN), .S(n14787), .Z(
        n14783) );
  AOI21_X1 U10868 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n14787), .A(n14782), .ZN(
        n8393) );
  INV_X1 U10869 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8391) );
  MUX2_X1 U10870 ( .A(n8391), .B(P2_REG1_REG_7__SCAN_IN), .S(n9121), .Z(n8392)
         );
  NOR2_X1 U10871 ( .A1(n8393), .A2(n8392), .ZN(n8879) );
  AOI211_X1 U10872 ( .C1(n8393), .C2(n8392), .A(n14847), .B(n8879), .ZN(n8409)
         );
  INV_X1 U10873 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9481) );
  XOR2_X1 U10874 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n14760), .Z(n14761) );
  INV_X1 U10875 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8394) );
  OR2_X1 U10876 ( .A1(n8395), .A2(n8394), .ZN(n8397) );
  NAND2_X1 U10877 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  AND2_X1 U10878 ( .A1(n8397), .A2(n8396), .ZN(n14751) );
  AND2_X1 U10879 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14750) );
  NAND2_X1 U10880 ( .A1(n14751), .A2(n14750), .ZN(n14749) );
  NAND2_X1 U10881 ( .A1(n14749), .A2(n8397), .ZN(n14762) );
  AOI22_X1 U10882 ( .A1(n14761), .A2(n14762), .B1(n14760), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n8427) );
  INV_X1 U10883 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10065) );
  MUX2_X1 U10884 ( .A(n10065), .B(P2_REG2_REG_3__SCAN_IN), .S(n8773), .Z(n8426) );
  NOR2_X1 U10885 ( .A1(n8427), .A2(n8426), .ZN(n8425) );
  AOI21_X1 U10886 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n8773), .A(n8425), .ZN(
        n14776) );
  INV_X1 U10887 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8398) );
  MUX2_X1 U10888 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n8398), .S(n8399), .Z(n14775) );
  NOR2_X1 U10889 ( .A1(n14776), .A2(n14775), .ZN(n14774) );
  NOR2_X1 U10890 ( .A1(n8399), .A2(n8398), .ZN(n8438) );
  MUX2_X1 U10891 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9481), .S(n8901), .Z(n8437)
         );
  OAI21_X1 U10892 ( .B1(n14774), .B2(n8438), .A(n8437), .ZN(n8436) );
  OAI21_X1 U10893 ( .B1(n9481), .B2(n8446), .A(n8436), .ZN(n14790) );
  INV_X1 U10894 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9492) );
  MUX2_X1 U10895 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9492), .S(n14787), .Z(
        n14789) );
  NAND2_X1 U10896 ( .A1(n14790), .A2(n14789), .ZN(n14788) );
  NAND2_X1 U10897 ( .A1(n14787), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8402) );
  INV_X1 U10898 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8400) );
  MUX2_X1 U10899 ( .A(n8400), .B(P2_REG2_REG_7__SCAN_IN), .S(n9121), .Z(n8401)
         );
  AOI21_X1 U10900 ( .B1(n14788), .B2(n8402), .A(n8401), .ZN(n8883) );
  AND3_X1 U10901 ( .A1(n14788), .A2(n8402), .A3(n8401), .ZN(n8403) );
  NOR3_X1 U10902 ( .A1(n8883), .A2(n8403), .A3(n14802), .ZN(n8408) );
  INV_X1 U10903 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9146) );
  NOR2_X1 U10904 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9146), .ZN(n8404) );
  AOI21_X1 U10905 ( .B1(n14840), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8404), .ZN(
        n8405) );
  OAI21_X1 U10906 ( .B1(n8406), .B2(n14846), .A(n8405), .ZN(n8407) );
  OR3_X1 U10907 ( .A1(n8409), .A2(n8408), .A3(n8407), .ZN(P2_U3221) );
  MUX2_X1 U10908 ( .A(n8421), .B(n8418), .S(n6641), .Z(n8527) );
  NAND2_X1 U10909 ( .A1(n8412), .A2(SI_10_), .ZN(n8648) );
  NAND2_X1 U10910 ( .A1(n8413), .A2(n9945), .ZN(n8414) );
  NAND2_X1 U10911 ( .A1(n8648), .A2(n8414), .ZN(n9999) );
  NAND2_X1 U10912 ( .A1(n9070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8415) );
  MUX2_X1 U10913 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8415), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n8417) );
  INV_X1 U10914 ( .A(n8653), .ZN(n8416) );
  NAND2_X1 U10915 ( .A1(n8417), .A2(n8416), .ZN(n9650) );
  OAI222_X1 U10916 ( .A1(n13681), .A2(n8418), .B1(n13675), .B2(n9999), .C1(
        n9650), .C2(P2_U3088), .ZN(P2_U3317) );
  NAND2_X1 U10917 ( .A1(n8419), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8420) );
  XNOR2_X1 U10918 ( .A(n8420), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10000) );
  INV_X1 U10919 ( .A(n10000), .ZN(n8829) );
  OAI222_X1 U10920 ( .A1(P1_U3086), .A2(n8829), .B1(n14373), .B2(n9999), .C1(
        n8421), .C2(n14370), .ZN(P1_U3345) );
  AOI211_X1 U10921 ( .C1(n8424), .C2(n8423), .A(n8422), .B(n14847), .ZN(n8429)
         );
  AOI211_X1 U10922 ( .C1(n8427), .C2(n8426), .A(n8425), .B(n14802), .ZN(n8428)
         );
  NOR2_X1 U10923 ( .A1(n8429), .A2(n8428), .ZN(n8431) );
  AOI22_X1 U10924 ( .A1(n14840), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3088), .ZN(n8430) );
  OAI211_X1 U10925 ( .C1(n8432), .C2(n14846), .A(n8431), .B(n8430), .ZN(
        P2_U3217) );
  AOI211_X1 U10926 ( .C1(n8435), .C2(n8434), .A(n14847), .B(n8433), .ZN(n8442)
         );
  INV_X1 U10927 ( .A(n8436), .ZN(n8440) );
  NOR3_X1 U10928 ( .A1(n14774), .A2(n8438), .A3(n8437), .ZN(n8439) );
  NOR3_X1 U10929 ( .A1(n8440), .A2(n8439), .A3(n14802), .ZN(n8441) );
  NOR2_X1 U10930 ( .A1(n8442), .A2(n8441), .ZN(n8445) );
  AND2_X1 U10931 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8443) );
  AOI21_X1 U10932 ( .B1(n14840), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8443), .ZN(
        n8444) );
  OAI211_X1 U10933 ( .C1(n8446), .C2(n14846), .A(n8445), .B(n8444), .ZN(
        P2_U3219) );
  NAND2_X1 U10934 ( .A1(n9098), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U10935 ( .A1(n9093), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8449) );
  AND2_X1 U10936 ( .A1(n8821), .A2(n8449), .ZN(n8450) );
  OR2_X1 U10937 ( .A1(n8451), .A2(n8450), .ZN(n8452) );
  NAND2_X1 U10938 ( .A1(n8822), .A2(n8452), .ZN(n10667) );
  INV_X1 U10939 ( .A(n6708), .ZN(n8454) );
  NAND2_X1 U10940 ( .A1(n8456), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8455) );
  MUX2_X1 U10941 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8455), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8457) );
  AND2_X1 U10942 ( .A1(n8457), .A2(n8824), .ZN(n12541) );
  AOI22_X1 U10943 ( .A1(n12541), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_16_), .B2(
        n8458), .ZN(n8459) );
  OAI21_X1 U10944 ( .B1(n10667), .B2(n12997), .A(n8459), .ZN(P3_U3279) );
  INV_X1 U10945 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8460) );
  MUX2_X1 U10946 ( .A(n8460), .B(P1_REG1_REG_10__SCAN_IN), .S(n10000), .Z(
        n8463) );
  OAI21_X1 U10947 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9965), .A(n8461), .ZN(
        n8462) );
  NOR2_X1 U10948 ( .A1(n8462), .A2(n8463), .ZN(n8830) );
  AOI211_X1 U10949 ( .C1(n8463), .C2(n8462), .A(n13886), .B(n8830), .ZN(n8474)
         );
  NOR2_X1 U10950 ( .A1(n8465), .A2(n8464), .ZN(n8467) );
  INV_X1 U10951 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U10952 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9978), .S(n10000), .Z(
        n8466) );
  OAI21_X1 U10953 ( .B1(n8468), .B2(n8467), .A(n8466), .ZN(n8828) );
  OR3_X1 U10954 ( .A1(n8468), .A2(n8467), .A3(n8466), .ZN(n8469) );
  NAND3_X1 U10955 ( .A1(n8828), .A2(n14669), .A3(n8469), .ZN(n8472) );
  NAND2_X1 U10956 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10650)
         );
  INV_X1 U10957 ( .A(n10650), .ZN(n8470) );
  AOI21_X1 U10958 ( .B1(n14656), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n8470), .ZN(
        n8471) );
  OAI211_X1 U10959 ( .C1(n13885), .C2(n8829), .A(n8472), .B(n8471), .ZN(n8473)
         );
  OR2_X1 U10960 ( .A1(n8474), .A2(n8473), .ZN(P1_U3253) );
  OR2_X1 U10961 ( .A1(n9708), .A2(n9704), .ZN(n8710) );
  INV_X1 U10962 ( .A(n8710), .ZN(n8487) );
  INV_X1 U10963 ( .A(n8475), .ZN(n8486) );
  NOR4_X1 U10964 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8484) );
  OR4_X1 U10965 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_3__SCAN_IN), .ZN(n8481) );
  NOR4_X1 U10966 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8479) );
  NOR4_X1 U10967 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8478) );
  NOR4_X1 U10968 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8477) );
  NOR4_X1 U10969 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n8476) );
  NAND4_X1 U10970 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n8480)
         );
  NOR4_X1 U10971 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8481), .A4(n8480), .ZN(n8483) );
  NOR4_X1 U10972 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8482) );
  AND3_X1 U10973 ( .A1(n8484), .A2(n8483), .A3(n8482), .ZN(n8485) );
  NAND2_X1 U10974 ( .A1(n8487), .A2(n8708), .ZN(n8697) );
  INV_X1 U10975 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10976 ( .A1(n12601), .A2(n9413), .ZN(n8497) );
  INV_X1 U10977 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U10978 ( .A1(n8491), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8492) );
  MUX2_X1 U10979 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8492), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8494) );
  NAND2_X1 U10980 ( .A1(n8494), .A2(n8493), .ZN(n9273) );
  AND2_X1 U10981 ( .A1(n9413), .A2(n9273), .ZN(n9702) );
  INV_X1 U10982 ( .A(n9702), .ZN(n8495) );
  XNOR2_X1 U10983 ( .A(n12429), .B(n8495), .ZN(n8496) );
  NAND2_X1 U10984 ( .A1(n8497), .A2(n8496), .ZN(n9352) );
  NAND2_X1 U10985 ( .A1(n8697), .A2(n9352), .ZN(n8502) );
  NAND3_X1 U10986 ( .A1(n9708), .A2(n9704), .A3(n8708), .ZN(n8694) );
  NAND2_X1 U10987 ( .A1(n12614), .A2(n12429), .ZN(n9700) );
  INV_X1 U10988 ( .A(n9273), .ZN(n9364) );
  NAND2_X1 U10989 ( .A1(n9413), .A2(n9364), .ZN(n12269) );
  OR2_X1 U10990 ( .A1(n9700), .A2(n12269), .ZN(n8693) );
  INV_X1 U10991 ( .A(n8693), .ZN(n8500) );
  NAND2_X1 U10992 ( .A1(n9701), .A2(n12409), .ZN(n9707) );
  NAND2_X1 U10993 ( .A1(n9707), .A2(n8498), .ZN(n8499) );
  AOI21_X1 U10994 ( .B1(n8694), .B2(n8500), .A(n8499), .ZN(n8501) );
  NAND2_X1 U10995 ( .A1(n8502), .A2(n8501), .ZN(n8505) );
  INV_X1 U10996 ( .A(n8713), .ZN(n12428) );
  OR2_X1 U10997 ( .A1(n9701), .A2(n12397), .ZN(n12427) );
  NOR2_X1 U10998 ( .A1(n12428), .A2(n12427), .ZN(n8503) );
  AND2_X1 U10999 ( .A1(n8694), .A2(n8503), .ZN(n8504) );
  AOI21_X1 U11000 ( .B1(n8505), .B2(P3_STATE_REG_SCAN_IN), .A(n8504), .ZN(
        n9037) );
  AND2_X1 U11001 ( .A1(n9037), .A2(n8506), .ZN(n8972) );
  INV_X1 U11002 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11003 ( .A1(n10884), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U11004 ( .A1(n8514), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U11005 ( .A1(n9240), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U11006 ( .A1(n6638), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8507) );
  MUX2_X1 U11007 ( .A(P3_IR_REG_0__SCAN_IN), .B(n8511), .S(n10270), .Z(n9714)
         );
  INV_X1 U11008 ( .A(n9714), .ZN(n8700) );
  NAND2_X1 U11009 ( .A1(n15147), .A2(n8700), .ZN(n12274) );
  INV_X1 U11010 ( .A(n12274), .ZN(n12273) );
  NOR2_X1 U11011 ( .A1(n15144), .A2(n12273), .ZN(n12250) );
  INV_X1 U11012 ( .A(n12250), .ZN(n8524) );
  INV_X1 U11013 ( .A(n12429), .ZN(n11971) );
  NAND2_X1 U11014 ( .A1(n11971), .A2(n9413), .ZN(n15209) );
  NAND2_X1 U11015 ( .A1(n9352), .A2(n15209), .ZN(n8512) );
  OAI22_X1 U11016 ( .A1(n8697), .A2(n8512), .B1(n8693), .B2(n8694), .ZN(n8513)
         );
  INV_X1 U11017 ( .A(n12214), .ZN(n12168) );
  NAND2_X1 U11018 ( .A1(n8514), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U11019 ( .A1(n9240), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U11020 ( .A1(n6638), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U11021 ( .A1(n10884), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U11022 ( .A1(n12422), .A2(n8713), .ZN(n8519) );
  NOR2_X1 U11023 ( .A1(n8694), .A2(n8519), .ZN(n8758) );
  NAND2_X1 U11024 ( .A1(n8757), .A2(n10270), .ZN(n8520) );
  INV_X1 U11025 ( .A(n12423), .ZN(n15158) );
  NAND2_X1 U11026 ( .A1(n8697), .A2(n15158), .ZN(n8522) );
  AND2_X1 U11027 ( .A1(n8713), .A2(n15155), .ZN(n8521) );
  INV_X1 U11028 ( .A(n12212), .ZN(n12174) );
  OAI22_X1 U11029 ( .A1(n15131), .A2(n12202), .B1(n8700), .B2(n12174), .ZN(
        n8523) );
  AOI21_X1 U11030 ( .B1(n8524), .B2(n12168), .A(n8523), .ZN(n8525) );
  OAI21_X1 U11031 ( .B1(n8972), .B2(n8715), .A(n8525), .ZN(P3_U3172) );
  MUX2_X1 U11032 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6641), .Z(n8649) );
  OAI22_X1 U11033 ( .A1(n8527), .A2(n9945), .B1(n8529), .B2(n8526), .ZN(n8532)
         );
  INV_X1 U11034 ( .A(n8527), .ZN(n8645) );
  OAI21_X1 U11035 ( .B1(n8645), .B2(SI_10_), .A(SI_11_), .ZN(n8530) );
  NOR2_X1 U11036 ( .A1(SI_11_), .A2(SI_10_), .ZN(n8528) );
  AOI22_X1 U11037 ( .A1(n8530), .A2(n8529), .B1(n8528), .B2(n8527), .ZN(n8531)
         );
  MUX2_X1 U11038 ( .A(n8538), .B(n8535), .S(n6641), .Z(n8801) );
  XNOR2_X1 U11039 ( .A(n8799), .B(n8798), .ZN(n10408) );
  INV_X1 U11040 ( .A(n10408), .ZN(n8539) );
  INV_X1 U11041 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U11042 ( .A1(n8653), .A2(n8533), .ZN(n8802) );
  NAND2_X1 U11043 ( .A1(n8802), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8534) );
  XNOR2_X1 U11044 ( .A(n8534), .B(P2_IR_REG_12__SCAN_IN), .ZN(n13169) );
  INV_X1 U11045 ( .A(n13169), .ZN(n13161) );
  OAI222_X1 U11046 ( .A1(n11464), .A2(n8535), .B1(n13675), .B2(n8539), .C1(
        n13161), .C2(P2_U3088), .ZN(P2_U3315) );
  NOR2_X1 U11047 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8536) );
  NAND2_X1 U11048 ( .A1(n8537), .A2(n8536), .ZN(n8643) );
  NAND2_X1 U11049 ( .A1(n9165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8805) );
  XNOR2_X1 U11050 ( .A(n8805), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10409) );
  INV_X1 U11051 ( .A(n10409), .ZN(n9005) );
  OAI222_X1 U11052 ( .A1(P1_U3086), .A2(n9005), .B1(n14373), .B2(n8539), .C1(
        n8538), .C2(n14370), .ZN(P1_U3343) );
  INV_X1 U11053 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15141) );
  XNOR2_X1 U11054 ( .A(n10129), .B(n15141), .ZN(n8543) );
  NAND2_X1 U11055 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U11056 ( .A1(n8542), .A2(n8543), .ZN(n10131) );
  OAI21_X1 U11057 ( .B1(n8543), .B2(n8542), .A(n10131), .ZN(n8554) );
  INV_X1 U11058 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10071) );
  MUX2_X1 U11059 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10071), .S(n10129), .Z(
        n8547) );
  NAND2_X1 U11060 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  NAND2_X1 U11061 ( .A1(n8547), .A2(n8546), .ZN(n10070) );
  OAI21_X1 U11062 ( .B1(n8547), .B2(n8546), .A(n10070), .ZN(n8548) );
  INV_X1 U11063 ( .A(n8548), .ZN(n8551) );
  INV_X1 U11064 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n8971) );
  NOR2_X1 U11065 ( .A1(n8971), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8549) );
  AOI21_X1 U11066 ( .B1(n15092), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n8549), .ZN(
        n8550) );
  OAI21_X1 U11067 ( .B1(n12616), .B2(n8551), .A(n8550), .ZN(n8553) );
  NOR2_X1 U11068 ( .A1(n15089), .A2(n6651), .ZN(n8552) );
  AOI211_X1 U11069 ( .C1(n12588), .C2(n8554), .A(n8553), .B(n8552), .ZN(n8564)
         );
  INV_X1 U11070 ( .A(n8555), .ZN(n8560) );
  MUX2_X1 U11071 ( .A(n15141), .B(n10071), .S(n6648), .Z(n8556) );
  NAND2_X1 U11072 ( .A1(n8556), .A2(n10072), .ZN(n10086) );
  INV_X1 U11073 ( .A(n8556), .ZN(n8557) );
  NAND2_X1 U11074 ( .A1(n8557), .A2(n6651), .ZN(n8558) );
  NAND2_X1 U11075 ( .A1(n10086), .A2(n8558), .ZN(n8559) );
  AOI21_X1 U11076 ( .B1(n8561), .B2(n8560), .A(n8559), .ZN(n14975) );
  AND3_X1 U11077 ( .A1(n8561), .A2(n8560), .A3(n8559), .ZN(n8562) );
  OAI21_X1 U11078 ( .B1(n14975), .B2(n8562), .A(n15084), .ZN(n8563) );
  NAND2_X1 U11079 ( .A1(n8564), .A2(n8563), .ZN(P3_U3184) );
  INV_X1 U11080 ( .A(n13841), .ZN(n8566) );
  MUX2_X1 U11081 ( .A(n8566), .B(n8565), .S(n14653), .Z(n8569) );
  OAI21_X1 U11082 ( .B1(n14653), .B2(P1_REG2_REG_0__SCAN_IN), .A(n8636), .ZN(
        n14651) );
  NAND2_X1 U11083 ( .A1(n14651), .A2(n8567), .ZN(n8568) );
  OAI211_X1 U11084 ( .C1(n8569), .C2(n11008), .A(P1_U4016), .B(n8568), .ZN(
        n13874) );
  INV_X1 U11085 ( .A(n13874), .ZN(n8581) );
  OAI211_X1 U11086 ( .C1(n8571), .C2(n8570), .A(n14669), .B(n13850), .ZN(n8579) );
  OAI211_X1 U11087 ( .C1(n8574), .C2(n8573), .A(n14668), .B(n8572), .ZN(n8578)
         );
  AOI22_X1 U11088 ( .A1(n14656), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n8577) );
  INV_X1 U11089 ( .A(n13885), .ZN(n14665) );
  NAND2_X1 U11090 ( .A1(n14665), .A2(n8575), .ZN(n8576) );
  NAND4_X1 U11091 ( .A1(n8579), .A2(n8578), .A3(n8577), .A4(n8576), .ZN(n8580)
         );
  OR2_X1 U11092 ( .A1(n8581), .A2(n8580), .ZN(P1_U3245) );
  INV_X1 U11093 ( .A(n14958), .ZN(n8582) );
  INV_X1 U11094 ( .A(n8583), .ZN(n9276) );
  NAND2_X1 U11095 ( .A1(n13157), .A2(n8590), .ZN(n8584) );
  XNOR2_X1 U11096 ( .A(n9275), .B(n9276), .ZN(n9931) );
  OAI21_X1 U11097 ( .B1(n11399), .B2(n8585), .A(n9561), .ZN(n8589) );
  OR2_X1 U11098 ( .A1(n11315), .A2(n13227), .ZN(n8587) );
  NAND2_X1 U11099 ( .A1(n6640), .A2(n11396), .ZN(n8586) );
  AOI21_X1 U11100 ( .B1(n8589), .B2(n13499), .A(n8588), .ZN(n9934) );
  NAND2_X1 U11101 ( .A1(n8590), .A2(n11028), .ZN(n9567) );
  OAI211_X1 U11102 ( .C1(n8590), .C2(n11028), .A(n13488), .B(n9567), .ZN(n9927) );
  OAI211_X1 U11103 ( .C1(n8590), .C2(n14953), .A(n9934), .B(n9927), .ZN(n8591)
         );
  AOI21_X1 U11104 ( .B1(n14938), .B2(n9931), .A(n8591), .ZN(n14912) );
  NOR2_X1 U11105 ( .A1(n8592), .A2(n14907), .ZN(n14906) );
  AND3_X1 U11106 ( .A1(n9109), .A2(n8594), .A3(n8593), .ZN(n8595) );
  AND2_X1 U11107 ( .A1(n14906), .A2(n8595), .ZN(n9305) );
  INV_X1 U11108 ( .A(n9304), .ZN(n8596) );
  INV_X2 U11109 ( .A(n14970), .ZN(n14968) );
  NAND2_X1 U11110 ( .A1(n14968), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8597) );
  OAI21_X1 U11111 ( .B1(n14912), .B2(n14968), .A(n8597), .ZN(P2_U3500) );
  NAND2_X1 U11112 ( .A1(n6645), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8604) );
  INV_X1 U11113 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8598) );
  OR2_X1 U11114 ( .A1(n11704), .A2(n8598), .ZN(n8603) );
  OR2_X1 U11115 ( .A1(n8852), .A2(n8599), .ZN(n8602) );
  OR2_X1 U11116 ( .A1(n11881), .A2(n8600), .ZN(n8601) );
  NAND2_X2 U11117 ( .A1(n11578), .A2(n7737), .ZN(n11612) );
  OR2_X1 U11118 ( .A1(n8727), .A2(n11612), .ZN(n8610) );
  OR2_X1 U11119 ( .A1(n6660), .A2(n8606), .ZN(n8609) );
  OR2_X1 U11120 ( .A1(n11578), .A2(n8607), .ZN(n8608) );
  NAND2_X1 U11121 ( .A1(n11730), .A2(n10521), .ZN(n8611) );
  XNOR2_X1 U11122 ( .A(n9059), .B(n9057), .ZN(n8630) );
  OAI21_X1 U11123 ( .B1(n9192), .B2(n8613), .A(n8612), .ZN(n8661) );
  NAND2_X1 U11124 ( .A1(n14192), .A2(n10521), .ZN(n8620) );
  OR2_X1 U11125 ( .A1(n6659), .A2(n7457), .ZN(n8618) );
  OR2_X1 U11126 ( .A1(n11578), .A2(n8615), .ZN(n8616) );
  NAND2_X1 U11127 ( .A1(n11680), .A2(n14192), .ZN(n8623) );
  NAND2_X1 U11128 ( .A1(n14200), .A2(n10521), .ZN(n8622) );
  NAND2_X1 U11129 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  AND2_X1 U11130 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  INV_X1 U11131 ( .A(n8627), .ZN(n8628) );
  OAI21_X1 U11132 ( .B1(n8630), .B2(n8629), .A(n13704), .ZN(n8641) );
  NAND2_X1 U11133 ( .A1(n6645), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8635) );
  OR2_X1 U11134 ( .A1(n11881), .A2(n8631), .ZN(n8634) );
  OR2_X1 U11135 ( .A1(n11704), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11136 ( .A1(n13818), .A2(n14591), .ZN(n13806) );
  AND2_X1 U11137 ( .A1(n13818), .A2(n14262), .ZN(n14577) );
  NAND2_X1 U11138 ( .A1(n14577), .A2(n14192), .ZN(n8639) );
  AOI22_X1 U11139 ( .A1(n13798), .A2(n11730), .B1(n8663), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8638) );
  OAI211_X1 U11140 ( .C1(n7323), .C2(n13806), .A(n8639), .B(n8638), .ZN(n8640)
         );
  AOI21_X1 U11141 ( .B1(n8641), .B2(n14567), .A(n8640), .ZN(n8642) );
  INV_X1 U11142 ( .A(n8642), .ZN(P1_U3237) );
  NAND2_X1 U11143 ( .A1(n8643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8644) );
  XNOR2_X1 U11144 ( .A(n8644), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10246) );
  INV_X1 U11145 ( .A(n10246), .ZN(n8997) );
  NAND2_X1 U11146 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  NAND2_X1 U11147 ( .A1(n8648), .A2(n8647), .ZN(n8651) );
  XNOR2_X1 U11148 ( .A(n8649), .B(SI_11_), .ZN(n8650) );
  INV_X1 U11149 ( .A(n10245), .ZN(n8658) );
  OAI222_X1 U11150 ( .A1(n8997), .A2(P1_U3086), .B1(n14373), .B2(n8658), .C1(
        n15391), .C2(n14370), .ZN(P1_U3344) );
  NOR2_X1 U11151 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  MUX2_X1 U11152 ( .A(n8652), .B(n8654), .S(P2_IR_REG_11__SCAN_IN), .Z(n8656)
         );
  INV_X1 U11153 ( .A(n8802), .ZN(n8655) );
  INV_X1 U11154 ( .A(n14815), .ZN(n8657) );
  OAI222_X1 U11155 ( .A1(n13681), .A2(n8659), .B1(n13675), .B2(n8658), .C1(
        P2_U3088), .C2(n8657), .ZN(P2_U3316) );
  OAI21_X1 U11156 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8667) );
  NAND2_X1 U11157 ( .A1(n14577), .A2(n14195), .ZN(n8665) );
  AOI22_X1 U11158 ( .A1(n13798), .A2(n14200), .B1(n8663), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8664) );
  OAI211_X1 U11159 ( .C1(n11728), .C2(n13806), .A(n8665), .B(n8664), .ZN(n8666) );
  AOI21_X1 U11160 ( .B1(n8667), .B2(n14567), .A(n8666), .ZN(n8668) );
  INV_X1 U11161 ( .A(n8668), .ZN(P1_U3222) );
  NAND2_X1 U11162 ( .A1(n14192), .A2(n14200), .ZN(n8669) );
  NAND2_X1 U11163 ( .A1(n8674), .A2(n8669), .ZN(n14193) );
  INV_X1 U11164 ( .A(n14203), .ZN(n8670) );
  NAND2_X1 U11165 ( .A1(n14202), .A2(n8674), .ZN(n8673) );
  NAND2_X1 U11166 ( .A1(n14196), .A2(n11730), .ZN(n8671) );
  INV_X1 U11167 ( .A(n11916), .ZN(n8672) );
  NAND2_X1 U11168 ( .A1(n8673), .A2(n8672), .ZN(n8844) );
  NAND3_X1 U11169 ( .A1(n14202), .A2(n8674), .A3(n11916), .ZN(n8675) );
  NAND2_X1 U11170 ( .A1(n8844), .A2(n8675), .ZN(n8676) );
  NAND2_X1 U11171 ( .A1(n8676), .A2(n14725), .ZN(n8681) );
  INV_X1 U11172 ( .A(n11717), .ZN(n8677) );
  NAND2_X1 U11173 ( .A1(n14192), .A2(n14694), .ZN(n11720) );
  NAND2_X1 U11174 ( .A1(n8677), .A2(n11720), .ZN(n11719) );
  OR2_X1 U11175 ( .A1(n14192), .A2(n14694), .ZN(n11721) );
  NAND2_X1 U11176 ( .A1(n11719), .A2(n11721), .ZN(n8847) );
  XNOR2_X1 U11177 ( .A(n8847), .B(n11916), .ZN(n8678) );
  NAND2_X1 U11178 ( .A1(n8678), .A2(n14592), .ZN(n8680) );
  AOI22_X1 U11179 ( .A1(n14262), .A2(n14192), .B1(n13832), .B2(n14591), .ZN(
        n8679) );
  NAND3_X1 U11180 ( .A1(n8681), .A2(n8680), .A3(n8679), .ZN(n10982) );
  OAI21_X1 U11181 ( .B1(n14191), .B2(n11727), .A(n14504), .ZN(n8682) );
  OR2_X1 U11182 ( .A1(n8861), .A2(n8682), .ZN(n10985) );
  INV_X1 U11183 ( .A(n10985), .ZN(n8683) );
  NOR2_X1 U11184 ( .A1(n10982), .A2(n8683), .ZN(n8690) );
  NAND2_X1 U11185 ( .A1(n14733), .A2(n14729), .ZN(n14354) );
  INV_X1 U11186 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8684) );
  OAI22_X1 U11187 ( .A1(n14354), .A2(n11727), .B1(n14733), .B2(n8684), .ZN(
        n8685) );
  INV_X1 U11188 ( .A(n8685), .ZN(n8686) );
  OAI21_X1 U11189 ( .B1(n8690), .B2(n14731), .A(n8686), .ZN(P1_U3465) );
  NAND2_X1 U11190 ( .A1(n14741), .A2(n14729), .ZN(n14309) );
  INV_X1 U11191 ( .A(n14309), .ZN(n10515) );
  AOI22_X1 U11192 ( .A1(n10515), .A2(n11730), .B1(n14739), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n8689) );
  OAI21_X1 U11193 ( .B1(n8690), .B2(n14739), .A(n8689), .ZN(P1_U3530) );
  INV_X1 U11194 ( .A(n12427), .ZN(n8691) );
  NOR3_X1 U11195 ( .A1(n12250), .A2(n15155), .A3(n8691), .ZN(n8692) );
  AOI21_X1 U11196 ( .B1(n15149), .B2(n12448), .A(n8692), .ZN(n9716) );
  AND2_X1 U11197 ( .A1(n12427), .A2(n8693), .ZN(n8696) );
  INV_X1 U11198 ( .A(n9352), .ZN(n8695) );
  OAI22_X1 U11199 ( .A1(n8697), .A2(n8696), .B1(n8695), .B2(n8694), .ZN(n8698)
         );
  NAND2_X1 U11200 ( .A1(n15217), .A2(n15155), .ZN(n12978) );
  INV_X1 U11201 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8699) );
  OAI22_X1 U11202 ( .A1(n12978), .A2(n8700), .B1(n15217), .B2(n8699), .ZN(
        n8701) );
  INV_X1 U11203 ( .A(n8701), .ZN(n8702) );
  OAI21_X1 U11204 ( .B1(n9716), .B2(n15215), .A(n8702), .ZN(P3_U3390) );
  INV_X1 U11205 ( .A(n9707), .ZN(n8704) );
  AND2_X1 U11206 ( .A1(n12429), .A2(n9364), .ZN(n8703) );
  NAND2_X1 U11207 ( .A1(n12601), .A2(n8703), .ZN(n9353) );
  NAND2_X1 U11208 ( .A1(n9353), .A2(n12397), .ZN(n9706) );
  OAI21_X1 U11209 ( .B1(n8704), .B2(n9708), .A(n9706), .ZN(n8707) );
  INV_X1 U11210 ( .A(n9706), .ZN(n8705) );
  NAND2_X1 U11211 ( .A1(n8705), .A2(n9704), .ZN(n8706) );
  AND2_X1 U11212 ( .A1(n8707), .A2(n8706), .ZN(n8712) );
  NAND2_X1 U11213 ( .A1(n8710), .A2(n8709), .ZN(n9713) );
  INV_X1 U11214 ( .A(n9713), .ZN(n8711) );
  NAND2_X1 U11215 ( .A1(n8712), .A2(n8711), .ZN(n8714) );
  NAND3_X1 U11216 ( .A1(n8713), .A2(n15155), .A3(n12423), .ZN(n12782) );
  NAND2_X2 U11217 ( .A1(n8714), .A2(n12782), .ZN(n15162) );
  OR2_X1 U11218 ( .A1(n8714), .A2(n12423), .ZN(n10928) );
  INV_X1 U11219 ( .A(n10928), .ZN(n15122) );
  NAND2_X1 U11220 ( .A1(n15122), .A2(n15155), .ZN(n12842) );
  INV_X1 U11221 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n8716) );
  OAI22_X1 U11222 ( .A1(n15162), .A2(n8716), .B1(n8715), .B2(n12782), .ZN(
        n8717) );
  AOI21_X1 U11223 ( .B1(n12792), .B2(n9714), .A(n8717), .ZN(n8718) );
  OAI21_X1 U11224 ( .B1(n9716), .B2(n12846), .A(n8718), .ZN(P3_U3233) );
  INV_X1 U11225 ( .A(n8735), .ZN(n8720) );
  NAND2_X1 U11226 ( .A1(n8720), .A2(n8719), .ZN(n8721) );
  NAND2_X1 U11227 ( .A1(n8723), .A2(n14760), .ZN(n8726) );
  XNOR2_X1 U11228 ( .A(n13067), .B(n11034), .ZN(n8768) );
  NAND2_X1 U11229 ( .A1(n13156), .A2(n13030), .ZN(n8769) );
  INV_X1 U11230 ( .A(n11037), .ZN(n14916) );
  NAND2_X1 U11231 ( .A1(n13157), .A2(n13120), .ZN(n8734) );
  NAND2_X1 U11232 ( .A1(n11372), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8732) );
  OR2_X1 U11233 ( .A1(n11337), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8731) );
  INV_X1 U11234 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8728) );
  OR2_X1 U11235 ( .A1(n6658), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U11236 ( .A1(n13155), .A2(n13237), .ZN(n8733) );
  AND2_X1 U11237 ( .A1(n8734), .A2(n8733), .ZN(n9564) );
  OAI22_X1 U11238 ( .A1(n14550), .A2(n14916), .B1(n9564), .B2(n14554), .ZN(
        n8740) );
  INV_X1 U11239 ( .A(n13048), .ZN(n13111) );
  AOI22_X1 U11240 ( .A1(n13111), .A2(n13157), .B1(n13133), .B2(n8735), .ZN(
        n8738) );
  INV_X1 U11241 ( .A(n8722), .ZN(n8737) );
  NOR3_X1 U11242 ( .A1(n8738), .A2(n8737), .A3(n8736), .ZN(n8739) );
  AOI211_X1 U11243 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n8741), .A(n8740), .B(
        n8739), .ZN(n8742) );
  OAI21_X1 U11244 ( .B1(n8772), .B2(n14552), .A(n8742), .ZN(P2_U3209) );
  INV_X1 U11245 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n8767) );
  INV_X1 U11246 ( .A(n8744), .ZN(n8745) );
  NAND2_X1 U11247 ( .A1(n10875), .A2(n8745), .ZN(n8748) );
  NAND3_X1 U11248 ( .A1(n12448), .A2(n8753), .A3(n15156), .ZN(n8750) );
  NAND2_X1 U11249 ( .A1(n15131), .A2(n8749), .ZN(n8959) );
  NAND2_X1 U11250 ( .A1(n15147), .A2(n9714), .ZN(n15142) );
  NAND2_X1 U11251 ( .A1(n15144), .A2(n12272), .ZN(n9349) );
  NAND2_X1 U11252 ( .A1(n15142), .A2(n12117), .ZN(n8751) );
  NAND2_X1 U11253 ( .A1(n9349), .A2(n8751), .ZN(n8752) );
  INV_X1 U11254 ( .A(n15144), .ZN(n8754) );
  NAND3_X1 U11255 ( .A1(n8754), .A2(n15145), .A3(n10289), .ZN(n8755) );
  NAND2_X1 U11256 ( .A1(n8756), .A2(n12168), .ZN(n8766) );
  INV_X1 U11257 ( .A(n15147), .ZN(n8763) );
  NAND3_X1 U11258 ( .A1(n8757), .A2(n12409), .A3(n10270), .ZN(n15130) );
  NAND2_X1 U11259 ( .A1(n8758), .A2(n15148), .ZN(n12209) );
  NAND2_X1 U11260 ( .A1(n8514), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11261 ( .A1(n10884), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U11262 ( .A1(n9240), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11263 ( .A1(n6638), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8759) );
  OAI22_X1 U11264 ( .A1(n8763), .A2(n12209), .B1(n9359), .B2(n12202), .ZN(
        n8764) );
  AOI21_X1 U11265 ( .B1(n12212), .B2(n15156), .A(n8764), .ZN(n8765) );
  OAI211_X1 U11266 ( .C1(n8972), .C2(n8767), .A(n8766), .B(n8765), .ZN(
        P3_U3162) );
  INV_X1 U11267 ( .A(n8768), .ZN(n8770) );
  NAND2_X1 U11268 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  OR2_X1 U11269 ( .A1(n8840), .A2(n11236), .ZN(n8774) );
  NAND2_X1 U11270 ( .A1(n8775), .A2(n8774), .ZN(n11056) );
  XNOR2_X1 U11271 ( .A(n13067), .B(n11056), .ZN(n8776) );
  AND2_X1 U11272 ( .A1(n13155), .A2(n13030), .ZN(n8777) );
  NAND2_X1 U11273 ( .A1(n8776), .A2(n8777), .ZN(n8895) );
  INV_X1 U11274 ( .A(n8776), .ZN(n8973) );
  INV_X1 U11275 ( .A(n8777), .ZN(n8778) );
  NAND2_X1 U11276 ( .A1(n8973), .A2(n8778), .ZN(n8779) );
  NAND2_X1 U11277 ( .A1(n8895), .A2(n8779), .ZN(n8780) );
  INV_X1 U11278 ( .A(n8897), .ZN(n8975) );
  AOI211_X1 U11279 ( .C1(n8781), .C2(n8780), .A(n14552), .B(n8975), .ZN(n8797)
         );
  INV_X1 U11280 ( .A(n8782), .ZN(n8783) );
  OR2_X1 U11281 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  NAND2_X1 U11282 ( .A1(n8785), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14558) );
  MUX2_X1 U11283 ( .A(n13121), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n8796) );
  NAND2_X1 U11284 ( .A1(n13156), .A2(n13120), .ZN(n8793) );
  NAND2_X1 U11285 ( .A1(n9136), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8791) );
  OR2_X1 U11286 ( .A1(n11317), .A2(n8398), .ZN(n8790) );
  NAND2_X1 U11287 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8905) );
  OAI21_X1 U11288 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8905), .ZN(n9471) );
  OR2_X1 U11289 ( .A1(n11337), .A2(n9471), .ZN(n8789) );
  INV_X1 U11290 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8787) );
  OR2_X1 U11291 ( .A1(n11318), .A2(n8787), .ZN(n8788) );
  NAND2_X1 U11292 ( .A1(n13154), .A2(n13237), .ZN(n8792) );
  NAND2_X1 U11293 ( .A1(n8793), .A2(n8792), .ZN(n10058) );
  INV_X1 U11294 ( .A(n10058), .ZN(n8794) );
  OAI22_X1 U11295 ( .A1(n14550), .A2(n14921), .B1(n8794), .B2(n14554), .ZN(
        n8795) );
  OR3_X1 U11296 ( .A1(n8797), .A2(n8796), .A3(n8795), .ZN(P2_U3190) );
  MUX2_X1 U11297 ( .A(n10779), .B(n10322), .S(n6641), .Z(n9083) );
  XNOR2_X1 U11298 ( .A(n9081), .B(n9080), .ZN(n10778) );
  INV_X1 U11299 ( .A(n10778), .ZN(n8809) );
  NAND2_X1 U11300 ( .A1(n9100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8804) );
  XNOR2_X1 U11301 ( .A(n8804), .B(n8803), .ZN(n14833) );
  OAI222_X1 U11302 ( .A1(n13681), .A2(n10322), .B1(n13675), .B2(n8809), .C1(
        n14833), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U11303 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11304 ( .A1(n8805), .A2(n9163), .ZN(n8806) );
  NAND2_X1 U11305 ( .A1(n8806), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11306 ( .A1(n8807), .A2(n9162), .ZN(n9103) );
  OR2_X1 U11307 ( .A1(n8807), .A2(n9162), .ZN(n8808) );
  INV_X1 U11308 ( .A(n10781), .ZN(n9451) );
  OAI222_X1 U11309 ( .A1(P1_U3086), .A2(n9451), .B1(n14373), .B2(n8809), .C1(
        n10779), .C2(n14370), .ZN(P1_U3342) );
  INV_X1 U11310 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n8820) );
  INV_X1 U11311 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8810) );
  INV_X1 U11312 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8812) );
  INV_X1 U11313 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11314 ( .A1(n10974), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U11315 ( .A1(n11988), .A2(n8815), .ZN(n12758) );
  NAND2_X1 U11316 ( .A1(n12758), .A2(n12024), .ZN(n8818) );
  AOI22_X1 U11317 ( .A1(n6639), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n12222), 
        .B2(P3_REG0_REG_20__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11318 ( .A1(n6638), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11319 ( .A1(n12764), .A2(P3_U3897), .ZN(n8819) );
  OAI21_X1 U11320 ( .B1(P3_U3897), .B2(n8820), .A(n8819), .ZN(P3_U3511) );
  INV_X1 U11321 ( .A(SI_17_), .ZN(n9435) );
  NAND2_X1 U11322 ( .A1(n9179), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11323 ( .A1(n9181), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U11324 ( .A1(n8874), .A2(n8823), .ZN(n8871) );
  XNOR2_X1 U11325 ( .A(n8873), .B(n8871), .ZN(n10874) );
  INV_X1 U11326 ( .A(n10874), .ZN(n8827) );
  NAND2_X1 U11327 ( .A1(n8824), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8825) );
  MUX2_X1 U11328 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8825), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8826) );
  AND2_X1 U11329 ( .A1(n8826), .A2(n8869), .ZN(n12577) );
  INV_X1 U11330 ( .A(n12577), .ZN(n12571) );
  OAI222_X1 U11331 ( .A1(n12985), .A2(n9435), .B1(n12997), .B2(n8827), .C1(
        P3_U3151), .C2(n12571), .ZN(P3_U3278) );
  INV_X1 U11332 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8996) );
  MUX2_X1 U11333 ( .A(n8996), .B(P1_REG2_REG_11__SCAN_IN), .S(n10246), .Z(
        n8992) );
  OAI21_X1 U11334 ( .B1(n9978), .B2(n8829), .A(n8828), .ZN(n8994) );
  XOR2_X1 U11335 ( .A(n8992), .B(n8994), .Z(n8838) );
  AOI21_X1 U11336 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n10000), .A(n8830), .ZN(
        n8832) );
  INV_X1 U11337 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10009) );
  MUX2_X1 U11338 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10009), .S(n10246), .Z(
        n8831) );
  NAND2_X1 U11339 ( .A1(n8832), .A2(n8831), .ZN(n9001) );
  OAI21_X1 U11340 ( .B1(n8832), .B2(n8831), .A(n9001), .ZN(n8833) );
  NAND2_X1 U11341 ( .A1(n8833), .A2(n14668), .ZN(n8837) );
  NAND2_X1 U11342 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14585)
         );
  INV_X1 U11343 ( .A(n14585), .ZN(n8835) );
  NOR2_X1 U11344 ( .A1(n13885), .A2(n8997), .ZN(n8834) );
  AOI211_X1 U11345 ( .C1(n14656), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8835), .B(
        n8834), .ZN(n8836) );
  OAI211_X1 U11346 ( .C1(n13867), .C2(n8838), .A(n8837), .B(n8836), .ZN(
        P1_U3254) );
  NAND2_X1 U11347 ( .A1(n8844), .A2(n11725), .ZN(n8842) );
  OR2_X1 U11348 ( .A1(n8840), .A2(n11612), .ZN(n8841) );
  NAND2_X1 U11349 ( .A1(n13832), .A2(n9053), .ZN(n11735) );
  NAND2_X1 U11350 ( .A1(n11736), .A2(n11735), .ZN(n8843) );
  NAND2_X1 U11351 ( .A1(n8842), .A2(n8843), .ZN(n8930) );
  INV_X1 U11352 ( .A(n8843), .ZN(n11918) );
  NAND3_X1 U11353 ( .A1(n8844), .A2(n11918), .A3(n11725), .ZN(n8845) );
  NAND2_X1 U11354 ( .A1(n8930), .A2(n8845), .ZN(n8846) );
  NAND2_X1 U11355 ( .A1(n8846), .A2(n14725), .ZN(n8860) );
  NAND2_X1 U11356 ( .A1(n8847), .A2(n11916), .ZN(n8849) );
  NAND2_X1 U11357 ( .A1(n11728), .A2(n11730), .ZN(n8848) );
  NAND2_X1 U11358 ( .A1(n8849), .A2(n8848), .ZN(n8934) );
  XNOR2_X1 U11359 ( .A(n8934), .B(n11918), .ZN(n8850) );
  NAND2_X1 U11360 ( .A1(n8850), .A2(n14592), .ZN(n8859) );
  NAND2_X1 U11361 ( .A1(n6644), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8857) );
  INV_X1 U11362 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8851) );
  OR2_X1 U11363 ( .A1(n11881), .A2(n8851), .ZN(n8856) );
  NAND2_X1 U11364 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8940) );
  OAI21_X1 U11365 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8940), .ZN(n9066) );
  OR2_X1 U11366 ( .A1(n11671), .A2(n9066), .ZN(n8855) );
  OR2_X1 U11367 ( .A1(n11656), .A2(n8853), .ZN(n8854) );
  AOI22_X1 U11368 ( .A1(n14196), .A2(n14262), .B1(n14591), .B2(n13831), .ZN(
        n8858) );
  NAND3_X1 U11369 ( .A1(n8860), .A2(n8859), .A3(n8858), .ZN(n9617) );
  INV_X1 U11370 ( .A(n9617), .ZN(n8862) );
  OAI211_X1 U11371 ( .C1(n8861), .C2(n9053), .A(n14504), .B(n8936), .ZN(n9622)
         );
  NAND2_X1 U11372 ( .A1(n8862), .A2(n9622), .ZN(n8867) );
  INV_X1 U11373 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8863) );
  OAI22_X1 U11374 ( .A1(n14354), .A2(n9053), .B1(n14733), .B2(n8863), .ZN(
        n8864) );
  AOI21_X1 U11375 ( .B1(n8867), .B2(n14733), .A(n8864), .ZN(n8865) );
  INV_X1 U11376 ( .A(n8865), .ZN(P1_U3468) );
  OAI22_X1 U11377 ( .A1(n14309), .A2(n9053), .B1(n14741), .B2(n8631), .ZN(
        n8866) );
  AOI21_X1 U11378 ( .B1(n8867), .B2(n14741), .A(n8866), .ZN(n8868) );
  INV_X1 U11379 ( .A(n8868), .ZN(P1_U3531) );
  NAND2_X1 U11380 ( .A1(n8869), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8870) );
  XNOR2_X1 U11381 ( .A(n8870), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12599) );
  INV_X1 U11382 ( .A(n12599), .ZN(n12605) );
  INV_X1 U11383 ( .A(SI_18_), .ZN(n9578) );
  INV_X1 U11384 ( .A(n8871), .ZN(n8872) );
  NAND2_X1 U11385 ( .A1(n9446), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11386 ( .A1(n9443), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8875) );
  AND2_X1 U11387 ( .A1(n8985), .A2(n8875), .ZN(n8876) );
  OR2_X1 U11388 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  NAND2_X1 U11389 ( .A1(n8986), .A2(n8878), .ZN(n10963) );
  OAI222_X1 U11390 ( .A1(P3_U3151), .A2(n12605), .B1(n12985), .B2(n9578), .C1(
        n12997), .C2(n10963), .ZN(P3_U3277) );
  INV_X1 U11391 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8880) );
  MUX2_X1 U11392 ( .A(n8880), .B(P2_REG1_REG_8__SCAN_IN), .S(n14800), .Z(
        n14796) );
  INV_X1 U11393 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9254) );
  MUX2_X1 U11394 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9254), .S(n9377), .Z(n8881)
         );
  OAI21_X1 U11395 ( .B1(n8882), .B2(n8881), .A(n9215), .ZN(n8891) );
  AOI21_X1 U11396 ( .B1(n9121), .B2(P2_REG2_REG_7__SCAN_IN), .A(n8883), .ZN(
        n14804) );
  MUX2_X1 U11397 ( .A(n9141), .B(P2_REG2_REG_8__SCAN_IN), .S(n14800), .Z(
        n14803) );
  NOR2_X1 U11398 ( .A1(n14804), .A2(n14803), .ZN(n14801) );
  AOI21_X1 U11399 ( .B1(n14800), .B2(P2_REG2_REG_8__SCAN_IN), .A(n14801), .ZN(
        n8885) );
  INV_X1 U11400 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n15485) );
  MUX2_X1 U11401 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n15485), .S(n9377), .Z(n8884) );
  NAND2_X1 U11402 ( .A1(n8885), .A2(n8884), .ZN(n9218) );
  OAI21_X1 U11403 ( .B1(n8885), .B2(n8884), .A(n9218), .ZN(n8886) );
  NAND2_X1 U11404 ( .A1(n8886), .A2(n14856), .ZN(n8888) );
  INV_X1 U11405 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9383) );
  NOR2_X1 U11406 ( .A1(n9383), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9394) );
  AOI21_X1 U11407 ( .B1(n14840), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9394), .ZN(
        n8887) );
  OAI211_X1 U11408 ( .C1(n14846), .C2(n8889), .A(n8888), .B(n8887), .ZN(n8890)
         );
  AOI21_X1 U11409 ( .B1(n8891), .B2(n13225), .A(n8890), .ZN(n8892) );
  INV_X1 U11410 ( .A(n8892), .ZN(P2_U3223) );
  NAND2_X1 U11411 ( .A1(n8931), .A2(n11362), .ZN(n8894) );
  AOI22_X1 U11412 ( .A1(n11358), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11169), 
        .B2(n14773), .ZN(n8893) );
  XNOR2_X1 U11413 ( .A(n14926), .B(n13067), .ZN(n8922) );
  NAND2_X1 U11414 ( .A1(n13154), .A2(n13030), .ZN(n8898) );
  XNOR2_X1 U11415 ( .A(n8922), .B(n8898), .ZN(n8983) );
  AND2_X1 U11416 ( .A1(n8983), .A2(n8895), .ZN(n8896) );
  NAND2_X1 U11417 ( .A1(n8897), .A2(n8896), .ZN(n8979) );
  INV_X1 U11418 ( .A(n8922), .ZN(n8899) );
  NAND2_X1 U11419 ( .A1(n8899), .A2(n8898), .ZN(n8900) );
  OR2_X1 U11420 ( .A1(n9186), .A2(n11236), .ZN(n8903) );
  AOI22_X1 U11421 ( .A1(n11358), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11169), 
        .B2(n8901), .ZN(n8902) );
  XNOR2_X1 U11422 ( .A(n11068), .B(n13067), .ZN(n9012) );
  NAND2_X1 U11423 ( .A1(n9136), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8911) );
  OR2_X1 U11424 ( .A1(n11317), .A2(n9481), .ZN(n8910) );
  AND2_X1 U11425 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  NOR2_X1 U11426 ( .A1(n8905), .A2(n8904), .ZN(n8912) );
  OR2_X1 U11427 ( .A1(n8906), .A2(n8912), .ZN(n9485) );
  OR2_X1 U11428 ( .A1(n6847), .A2(n9485), .ZN(n8909) );
  INV_X1 U11429 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8907) );
  OR2_X1 U11430 ( .A1(n11318), .A2(n8907), .ZN(n8908) );
  NAND4_X1 U11431 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n13153) );
  NAND2_X1 U11432 ( .A1(n13153), .A2(n13030), .ZN(n9013) );
  XNOR2_X1 U11433 ( .A(n9012), .B(n9013), .ZN(n8923) );
  NAND2_X1 U11434 ( .A1(n13154), .A2(n13120), .ZN(n8920) );
  NAND2_X1 U11435 ( .A1(n9136), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8918) );
  OR2_X1 U11436 ( .A1(n11317), .A2(n9492), .ZN(n8917) );
  NAND2_X1 U11437 ( .A1(n8912), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9024) );
  OR2_X1 U11438 ( .A1(n8912), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U11439 ( .A1(n9024), .A2(n8913), .ZN(n9493) );
  OR2_X1 U11440 ( .A1(n6847), .A2(n9493), .ZN(n8916) );
  INV_X1 U11441 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8914) );
  OR2_X1 U11442 ( .A1(n11318), .A2(n8914), .ZN(n8915) );
  NAND4_X1 U11443 ( .A1(n8918), .A2(n8917), .A3(n8916), .A4(n8915), .ZN(n13152) );
  NAND2_X1 U11444 ( .A1(n13152), .A2(n13237), .ZN(n8919) );
  NAND2_X1 U11445 ( .A1(n8920), .A2(n8919), .ZN(n9479) );
  AOI22_X1 U11446 ( .A1(n13137), .A2(n9479), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3088), .ZN(n8921) );
  OAI21_X1 U11447 ( .B1(n9485), .B2(n14558), .A(n8921), .ZN(n8927) );
  INV_X1 U11448 ( .A(n8979), .ZN(n8925) );
  AOI22_X1 U11449 ( .A1(n13111), .A2(n13154), .B1(n13133), .B2(n8922), .ZN(
        n8924) );
  NOR3_X1 U11450 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n8926) );
  AOI211_X1 U11451 ( .C1(n11068), .C2(n13128), .A(n8927), .B(n8926), .ZN(n8928) );
  OAI21_X1 U11452 ( .B1(n9016), .B2(n14552), .A(n8928), .ZN(P2_U3199) );
  NAND2_X1 U11453 ( .A1(n7323), .A2(n9053), .ZN(n8929) );
  NAND2_X1 U11454 ( .A1(n8930), .A2(n8929), .ZN(n9626) );
  NAND2_X1 U11455 ( .A1(n8931), .A2(n11897), .ZN(n8933) );
  AOI22_X1 U11456 ( .A1(n11529), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11528), 
        .B2(n13870), .ZN(n8932) );
  NAND2_X1 U11457 ( .A1(n8933), .A2(n8932), .ZN(n11743) );
  XNOR2_X1 U11458 ( .A(n11743), .B(n13831), .ZN(n11919) );
  XNOR2_X1 U11459 ( .A(n9626), .B(n11919), .ZN(n9880) );
  NAND2_X1 U11460 ( .A1(n8934), .A2(n11918), .ZN(n8935) );
  XNOR2_X1 U11461 ( .A(n9632), .B(n11919), .ZN(n9878) );
  AOI21_X1 U11462 ( .B1(n8936), .B2(n11743), .A(n14719), .ZN(n8937) );
  AND2_X1 U11463 ( .A1(n9818), .A2(n8937), .ZN(n9871) );
  NAND2_X1 U11464 ( .A1(n13832), .A2(n14262), .ZN(n8947) );
  NAND2_X1 U11465 ( .A1(n6644), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8945) );
  OR2_X1 U11466 ( .A1(n11881), .A2(n8938), .ZN(n8944) );
  AND2_X1 U11467 ( .A1(n8940), .A2(n8939), .ZN(n8941) );
  OR2_X1 U11468 ( .A1(n8941), .A2(n9199), .ZN(n9820) );
  OR2_X1 U11469 ( .A1(n11704), .A2(n9820), .ZN(n8943) );
  OR2_X1 U11470 ( .A1(n11656), .A2(n15340), .ZN(n8942) );
  NAND4_X1 U11471 ( .A1(n8945), .A2(n8944), .A3(n8943), .A4(n8942), .ZN(n13830) );
  NAND2_X1 U11472 ( .A1(n13830), .A2(n14591), .ZN(n8946) );
  NAND2_X1 U11473 ( .A1(n8947), .A2(n8946), .ZN(n9870) );
  AOI211_X1 U11474 ( .C1(n9878), .C2(n14592), .A(n9871), .B(n9870), .ZN(n8948)
         );
  OAI21_X1 U11475 ( .B1(n14289), .B2(n9880), .A(n8948), .ZN(n8953) );
  INV_X1 U11476 ( .A(n11743), .ZN(n9633) );
  OAI22_X1 U11477 ( .A1(n14309), .A2(n9633), .B1(n14741), .B2(n8851), .ZN(
        n8949) );
  AOI21_X1 U11478 ( .B1(n8953), .B2(n14741), .A(n8949), .ZN(n8950) );
  INV_X1 U11479 ( .A(n8950), .ZN(P1_U3532) );
  INV_X1 U11480 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8951) );
  OAI22_X1 U11481 ( .A1(n14354), .A2(n9633), .B1(n14733), .B2(n8951), .ZN(
        n8952) );
  AOI21_X1 U11482 ( .B1(n8953), .B2(n14733), .A(n8952), .ZN(n8954) );
  INV_X1 U11483 ( .A(n8954), .ZN(P1_U3471) );
  INV_X2 U11484 ( .A(n10270), .ZN(n10875) );
  NAND2_X1 U11485 ( .A1(n10875), .A2(n6651), .ZN(n8956) );
  NAND2_X1 U11486 ( .A1(n8960), .A2(n8959), .ZN(n8961) );
  OAI21_X1 U11487 ( .B1(n8962), .B2(n8961), .A(n9046), .ZN(n8963) );
  NAND2_X1 U11488 ( .A1(n8963), .A2(n12168), .ZN(n8970) );
  NAND2_X1 U11489 ( .A1(n8514), .A2(n15121), .ZN(n8967) );
  NAND2_X1 U11490 ( .A1(n9240), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11491 ( .A1(n6638), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U11492 ( .A1(n10884), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8964) );
  OAI22_X1 U11493 ( .A1(n15131), .A2(n12209), .B1(n15129), .B2(n12202), .ZN(
        n8968) );
  AOI21_X1 U11494 ( .B1(n15137), .B2(n12212), .A(n8968), .ZN(n8969) );
  OAI211_X1 U11495 ( .C1(n8972), .C2(n8971), .A(n8970), .B(n8969), .ZN(
        P3_U3177) );
  NOR3_X1 U11496 ( .A1(n13048), .A2(n8973), .A3(n9283), .ZN(n8974) );
  AOI21_X1 U11497 ( .B1(n8975), .B2(n13133), .A(n8974), .ZN(n8984) );
  NAND2_X1 U11498 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14767) );
  NAND2_X1 U11499 ( .A1(n13155), .A2(n13120), .ZN(n8977) );
  NAND2_X1 U11500 ( .A1(n13153), .A2(n13237), .ZN(n8976) );
  NAND2_X1 U11501 ( .A1(n8977), .A2(n8976), .ZN(n9466) );
  NAND2_X1 U11502 ( .A1(n13137), .A2(n9466), .ZN(n8978) );
  OAI211_X1 U11503 ( .C1(n14558), .C2(n9471), .A(n14767), .B(n8978), .ZN(n8981) );
  NOR2_X1 U11504 ( .A1(n8979), .A2(n14552), .ZN(n8980) );
  AOI211_X1 U11505 ( .C1(n14926), .C2(n13128), .A(n8981), .B(n8980), .ZN(n8982) );
  OAI21_X1 U11506 ( .B1(n8984), .B2(n8983), .A(n8982), .ZN(P2_U3202) );
  INV_X1 U11507 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9779) );
  NAND2_X1 U11508 ( .A1(n9779), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9271) );
  INV_X1 U11509 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11463) );
  NAND2_X1 U11510 ( .A1(n11463), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8987) );
  AND2_X1 U11511 ( .A1(n9271), .A2(n8987), .ZN(n8988) );
  OR2_X1 U11512 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  NAND2_X1 U11513 ( .A1(n9272), .A2(n8990), .ZN(n11976) );
  INV_X1 U11514 ( .A(SI_19_), .ZN(n11977) );
  OAI222_X1 U11515 ( .A1(n12997), .A2(n11976), .B1(n12985), .B2(n11977), .C1(
        P3_U3151), .C2(n12601), .ZN(P3_U3276) );
  INV_X1 U11516 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8991) );
  AOI22_X1 U11517 ( .A1(n10409), .A2(n8991), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9005), .ZN(n8999) );
  INV_X1 U11518 ( .A(n8992), .ZN(n8993) );
  NAND2_X1 U11519 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  OAI21_X1 U11520 ( .B1(n8997), .B2(n8996), .A(n8995), .ZN(n8998) );
  NOR2_X1 U11521 ( .A1(n8999), .A2(n8998), .ZN(n9344) );
  AOI21_X1 U11522 ( .B1(n8999), .B2(n8998), .A(n9344), .ZN(n9009) );
  INV_X1 U11523 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9000) );
  AOI22_X1 U11524 ( .A1(n10409), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9000), 
        .B2(n9005), .ZN(n9003) );
  OAI21_X1 U11525 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10246), .A(n9001), .ZN(
        n9002) );
  NAND2_X1 U11526 ( .A1(n9003), .A2(n9002), .ZN(n9338) );
  OAI21_X1 U11527 ( .B1(n9003), .B2(n9002), .A(n9338), .ZN(n9007) );
  NAND2_X1 U11528 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10868)
         );
  NAND2_X1 U11529 ( .A1(n14656), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n9004) );
  OAI211_X1 U11530 ( .C1(n13885), .C2(n9005), .A(n10868), .B(n9004), .ZN(n9006) );
  AOI21_X1 U11531 ( .B1(n9007), .B2(n14668), .A(n9006), .ZN(n9008) );
  OAI21_X1 U11532 ( .B1(n9009), .B2(n13867), .A(n9008), .ZN(P1_U3255) );
  AOI22_X1 U11533 ( .A1(n11358), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11169), 
        .B2(n14787), .ZN(n9010) );
  INV_X1 U11534 ( .A(n11075), .ZN(n9494) );
  INV_X1 U11535 ( .A(n9012), .ZN(n9014) );
  NAND2_X1 U11536 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  XNOR2_X1 U11537 ( .A(n11075), .B(n13067), .ZN(n9017) );
  AND2_X1 U11538 ( .A1(n13152), .A2(n13030), .ZN(n9018) );
  NAND2_X1 U11539 ( .A1(n9017), .A2(n9018), .ZN(n9130) );
  INV_X1 U11540 ( .A(n9017), .ZN(n9129) );
  INV_X1 U11541 ( .A(n9018), .ZN(n9019) );
  NAND2_X1 U11542 ( .A1(n9129), .A2(n9019), .ZN(n9020) );
  AOI21_X1 U11543 ( .B1(n9022), .B2(n9021), .A(n14552), .ZN(n9023) );
  NAND2_X1 U11544 ( .A1(n9023), .A2(n9131), .ZN(n9036) );
  INV_X1 U11545 ( .A(n9493), .ZN(n9034) );
  NAND2_X1 U11546 ( .A1(n13153), .A2(n13120), .ZN(n9032) );
  NAND2_X1 U11547 ( .A1(n9136), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9030) );
  OR2_X1 U11548 ( .A1(n11317), .A2(n8400), .ZN(n9029) );
  NAND2_X1 U11549 ( .A1(n9024), .A2(n9146), .ZN(n9025) );
  NAND2_X1 U11550 ( .A1(n9139), .A2(n9025), .ZN(n9135) );
  OR2_X1 U11551 ( .A1(n6847), .A2(n9135), .ZN(n9028) );
  INV_X1 U11552 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9026) );
  OR2_X1 U11553 ( .A1(n11318), .A2(n9026), .ZN(n9027) );
  NAND4_X1 U11554 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n13151) );
  NAND2_X1 U11555 ( .A1(n13151), .A2(n13237), .ZN(n9031) );
  AND2_X1 U11556 ( .A1(n9032), .A2(n9031), .ZN(n9302) );
  NAND2_X1 U11557 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n14781) );
  OAI21_X1 U11558 ( .B1(n9302), .B2(n14554), .A(n14781), .ZN(n9033) );
  AOI21_X1 U11559 ( .B1(n13121), .B2(n9034), .A(n9033), .ZN(n9035) );
  OAI211_X1 U11560 ( .C1(n9494), .C2(n14550), .A(n9036), .B(n9035), .ZN(
        P2_U3211) );
  INV_X1 U11561 ( .A(n12207), .ZN(n9958) );
  INV_X1 U11562 ( .A(n9038), .ZN(n9039) );
  NAND2_X1 U11563 ( .A1(n9359), .A2(n9039), .ZN(n9044) );
  AND2_X1 U11564 ( .A1(n9046), .A2(n9044), .ZN(n9048) );
  OR2_X1 U11565 ( .A1(n12236), .A2(SI_3_), .ZN(n9043) );
  OR2_X1 U11566 ( .A1(n11984), .A2(n9040), .ZN(n9042) );
  NAND2_X1 U11567 ( .A1(n10875), .A2(n14979), .ZN(n9041) );
  XNOR2_X1 U11568 ( .A(n9227), .B(n15129), .ZN(n9047) );
  AND2_X1 U11569 ( .A1(n9047), .A2(n9044), .ZN(n9045) );
  OAI211_X1 U11570 ( .C1(n9048), .C2(n9047), .A(n12168), .B(n9229), .ZN(n9051)
         );
  NOR2_X1 U11571 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15121), .ZN(n14981) );
  INV_X1 U11572 ( .A(n15120), .ZN(n9351) );
  OAI22_X1 U11573 ( .A1(n9506), .A2(n12202), .B1(n12174), .B2(n9351), .ZN(
        n9049) );
  AOI211_X1 U11574 ( .C1(n12199), .C2(n15150), .A(n14981), .B(n9049), .ZN(
        n9050) );
  OAI211_X1 U11575 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n9958), .A(n9051), .B(
        n9050), .ZN(P3_U3158) );
  AOI22_X1 U11576 ( .A1(n11680), .A2(n13832), .B1(n10521), .B2(n7320), .ZN(
        n9060) );
  NAND2_X1 U11577 ( .A1(n13832), .A2(n10521), .ZN(n9052) );
  OAI21_X1 U11578 ( .B1(n9053), .B2(n7432), .A(n9052), .ZN(n9055) );
  INV_X1 U11579 ( .A(n9054), .ZN(n9192) );
  XNOR2_X1 U11580 ( .A(n9056), .B(n9060), .ZN(n13706) );
  INV_X1 U11581 ( .A(n9057), .ZN(n9058) );
  NAND2_X1 U11582 ( .A1(n9059), .A2(n9058), .ZN(n13703) );
  AOI22_X1 U11583 ( .A1(n11680), .A2(n13831), .B1(n11743), .B2(n10521), .ZN(
        n9183) );
  AOI22_X1 U11584 ( .A1(n11743), .A2(n11699), .B1(n13831), .B2(n10521), .ZN(
        n9061) );
  XOR2_X1 U11585 ( .A(n11678), .B(n9061), .Z(n9184) );
  XNOR2_X1 U11586 ( .A(n9185), .B(n9184), .ZN(n9069) );
  AND2_X1 U11587 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13858) );
  AOI21_X1 U11588 ( .B1(n13798), .B2(n11743), .A(n13858), .ZN(n9068) );
  AND2_X1 U11589 ( .A1(n9063), .A2(n9062), .ZN(n9064) );
  NAND2_X1 U11590 ( .A1(n9210), .A2(n9064), .ZN(n9065) );
  INV_X1 U11591 ( .A(n14588), .ZN(n13778) );
  INV_X1 U11592 ( .A(n9066), .ZN(n9872) );
  AOI22_X1 U11593 ( .A1(n13818), .A2(n9870), .B1(n13778), .B2(n9872), .ZN(
        n9067) );
  OAI211_X1 U11594 ( .C1(n9069), .C2(n14574), .A(n9068), .B(n9067), .ZN(
        P1_U3230) );
  INV_X1 U11595 ( .A(n9070), .ZN(n9072) );
  NAND2_X1 U11596 ( .A1(n9072), .A2(n9071), .ZN(n9151) );
  NOR2_X1 U11597 ( .A1(n9151), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9077) );
  INV_X1 U11598 ( .A(n9077), .ZN(n9073) );
  NAND2_X1 U11599 ( .A1(n9073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9074) );
  MUX2_X1 U11600 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9074), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9075) );
  INV_X1 U11601 ( .A(n9075), .ZN(n9079) );
  INV_X1 U11602 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11603 ( .A1(n9077), .A2(n9076), .ZN(n9441) );
  INV_X1 U11604 ( .A(n9441), .ZN(n9078) );
  NOR2_X1 U11605 ( .A1(n9079), .A2(n9078), .ZN(n13207) );
  INV_X1 U11606 ( .A(n13207), .ZN(n13201) );
  NAND2_X1 U11607 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  MUX2_X1 U11608 ( .A(n9168), .B(n9160), .S(n6641), .Z(n9157) );
  INV_X1 U11609 ( .A(n9157), .ZN(n9086) );
  MUX2_X1 U11610 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6641), .Z(n9155) );
  NAND2_X1 U11611 ( .A1(n9155), .A2(SI_14_), .ZN(n9087) );
  NOR2_X1 U11612 ( .A1(n9155), .A2(SI_14_), .ZN(n9090) );
  AOI22_X1 U11613 ( .A1(n9090), .A2(n9089), .B1(n9157), .B2(n9088), .ZN(n9091)
         );
  MUX2_X1 U11614 ( .A(n9098), .B(n9093), .S(n6641), .Z(n9176) );
  XNOR2_X1 U11615 ( .A(n9174), .B(n9173), .ZN(n11487) );
  INV_X1 U11616 ( .A(n11487), .ZN(n9099) );
  OAI222_X1 U11617 ( .A1(P2_U3088), .A2(n13201), .B1(n13675), .B2(n9099), .C1(
        n9093), .C2(n13681), .ZN(P2_U3311) );
  MUX2_X1 U11618 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9094), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9097) );
  INV_X1 U11619 ( .A(n9096), .ZN(n9169) );
  AND2_X1 U11620 ( .A1(n9097), .A2(n9169), .ZN(n11488) );
  INV_X1 U11621 ( .A(n11488), .ZN(n10400) );
  OAI222_X1 U11622 ( .A1(P1_U3086), .A2(n10400), .B1(n14373), .B2(n9099), .C1(
        n9098), .C2(n14370), .ZN(P1_U3339) );
  XNOR2_X1 U11623 ( .A(n9153), .B(n10499), .ZN(n9156) );
  XNOR2_X1 U11624 ( .A(n9156), .B(n9155), .ZN(n10785) );
  INV_X1 U11625 ( .A(n10785), .ZN(n9106) );
  OAI21_X1 U11626 ( .B1(n9100), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9101) );
  XNOR2_X1 U11627 ( .A(n9101), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13171) );
  INV_X1 U11628 ( .A(n13171), .ZN(n14845) );
  OAI222_X1 U11629 ( .A1(n11464), .A2(n9102), .B1(n13675), .B2(n9106), .C1(
        n14845), .C2(P2_U3088), .ZN(P2_U3313) );
  NAND2_X1 U11630 ( .A1(n9103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9104) );
  XNOR2_X1 U11631 ( .A(n9104), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10786) );
  INV_X1 U11632 ( .A(n10786), .ZN(n9457) );
  OAI222_X1 U11633 ( .A1(P1_U3086), .A2(n9457), .B1(n14373), .B2(n9106), .C1(
        n9105), .C2(n14370), .ZN(P1_U3341) );
  NAND2_X1 U11634 ( .A1(n9108), .A2(n9107), .ZN(n14911) );
  INV_X1 U11635 ( .A(n14911), .ZN(n11398) );
  NAND2_X1 U11636 ( .A1(n9304), .A2(n9109), .ZN(n9110) );
  NOR2_X1 U11637 ( .A1(n9110), .A2(n14907), .ZN(n9111) );
  NAND2_X1 U11638 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  AND2_X2 U11639 ( .A1(n9113), .A2(n13515), .ZN(n13512) );
  OR2_X1 U11640 ( .A1(n13512), .A2(n6784), .ZN(n9685) );
  INV_X1 U11641 ( .A(n14949), .ZN(n9558) );
  OAI21_X1 U11642 ( .B1(n9558), .B2(n13499), .A(n14911), .ZN(n9116) );
  NAND2_X1 U11643 ( .A1(n9116), .A2(n9115), .ZN(n14909) );
  NOR2_X1 U11644 ( .A1(n9117), .A2(n11429), .ZN(n9118) );
  OAI21_X1 U11645 ( .B1(n14909), .B2(n9118), .A(n13471), .ZN(n9120) );
  INV_X1 U11646 ( .A(n13515), .ZN(n14864) );
  AOI22_X1 U11647 ( .A1(n13512), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n14864), .ZN(n9119) );
  OAI211_X1 U11648 ( .C1(n11398), .C2(n9685), .A(n9120), .B(n9119), .ZN(
        P2_U3265) );
  OR2_X1 U11649 ( .A1(n9515), .A2(n11236), .ZN(n9123) );
  AOI22_X1 U11650 ( .A1(n11358), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11169), 
        .B2(n9121), .ZN(n9122) );
  INV_X1 U11651 ( .A(n11083), .ZN(n14869) );
  XNOR2_X1 U11652 ( .A(n11083), .B(n13067), .ZN(n9124) );
  AND2_X1 U11653 ( .A1(n13151), .A2(n13030), .ZN(n9125) );
  NAND2_X1 U11654 ( .A1(n9124), .A2(n9125), .ZN(n9264) );
  INV_X1 U11655 ( .A(n9124), .ZN(n9249) );
  INV_X1 U11656 ( .A(n9125), .ZN(n9126) );
  NAND2_X1 U11657 ( .A1(n9249), .A2(n9126), .ZN(n9127) );
  AND2_X1 U11658 ( .A1(n9264), .A2(n9127), .ZN(n9132) );
  INV_X1 U11659 ( .A(n9132), .ZN(n9128) );
  AOI21_X1 U11660 ( .B1(n9131), .B2(n9128), .A(n14552), .ZN(n9134) );
  INV_X1 U11661 ( .A(n13152), .ZN(n9547) );
  NOR3_X1 U11662 ( .A1(n9129), .A2(n9547), .A3(n13048), .ZN(n9133) );
  OAI21_X1 U11663 ( .B1(n9134), .B2(n9133), .A(n9266), .ZN(n9150) );
  INV_X1 U11664 ( .A(n9135), .ZN(n14865) );
  NAND2_X1 U11665 ( .A1(n11277), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9145) );
  INV_X1 U11666 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9137) );
  OR2_X1 U11667 ( .A1(n11318), .A2(n9137), .ZN(n9144) );
  INV_X1 U11668 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11669 ( .A1(n9139), .A2(n9138), .ZN(n9140) );
  NAND2_X1 U11670 ( .A1(n9384), .A2(n9140), .ZN(n9681) );
  OR2_X1 U11671 ( .A1(n6847), .A2(n9681), .ZN(n9143) );
  INV_X1 U11672 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9141) );
  OR2_X1 U11673 ( .A1(n11317), .A2(n9141), .ZN(n9142) );
  NAND4_X1 U11674 ( .A1(n9145), .A2(n9144), .A3(n9143), .A4(n9142), .ZN(n13150) );
  INV_X1 U11675 ( .A(n13150), .ZN(n9692) );
  OAI22_X1 U11676 ( .A1(n9692), .A2(n13135), .B1(n9547), .B2(n13316), .ZN(
        n9550) );
  INV_X1 U11677 ( .A(n9550), .ZN(n9147) );
  OAI22_X1 U11678 ( .A1(n9147), .A2(n14554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9146), .ZN(n9148) );
  AOI21_X1 U11679 ( .B1(n14865), .B2(n13121), .A(n9148), .ZN(n9149) );
  OAI211_X1 U11680 ( .C1(n14869), .C2(n14550), .A(n9150), .B(n9149), .ZN(
        P2_U3185) );
  NAND2_X1 U11681 ( .A1(n9151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9152) );
  XNOR2_X1 U11682 ( .A(n9152), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13185) );
  INV_X1 U11683 ( .A(n13185), .ZN(n13178) );
  INV_X1 U11684 ( .A(n9153), .ZN(n9154) );
  OAI22_X1 U11685 ( .A1(n9156), .A2(n9155), .B1(n9154), .B2(SI_14_), .ZN(n9159) );
  XNOR2_X1 U11686 ( .A(n9157), .B(SI_15_), .ZN(n9158) );
  XNOR2_X1 U11687 ( .A(n9159), .B(n9158), .ZN(n10797) );
  INV_X1 U11688 ( .A(n10797), .ZN(n9167) );
  OAI222_X1 U11689 ( .A1(P2_U3088), .A2(n13178), .B1(n13675), .B2(n9167), .C1(
        n9160), .C2(n11464), .ZN(P2_U3312) );
  INV_X1 U11690 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9161) );
  NAND3_X1 U11691 ( .A1(n9163), .A2(n9162), .A3(n9161), .ZN(n9164) );
  OAI21_X1 U11692 ( .B1(n9165), .B2(n9164), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9166) );
  XNOR2_X1 U11693 ( .A(n9166), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14666) );
  INV_X1 U11694 ( .A(n14666), .ZN(n10394) );
  OAI222_X1 U11695 ( .A1(n14370), .A2(n9168), .B1(n14373), .B2(n9167), .C1(
        P1_U3086), .C2(n10394), .ZN(P1_U3340) );
  NAND2_X1 U11696 ( .A1(n9169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9170) );
  MUX2_X1 U11697 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9170), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9172) );
  INV_X1 U11698 ( .A(n9171), .ZN(n9444) );
  NAND2_X1 U11699 ( .A1(n9172), .A2(n9444), .ZN(n10939) );
  INV_X1 U11700 ( .A(SI_16_), .ZN(n9175) );
  NAND2_X1 U11701 ( .A1(n9176), .A2(n9175), .ZN(n9177) );
  MUX2_X1 U11702 ( .A(n9179), .B(n9181), .S(n6641), .Z(n9436) );
  XNOR2_X1 U11703 ( .A(n9434), .B(n9433), .ZN(n11498) );
  INV_X1 U11704 ( .A(n11498), .ZN(n9182) );
  OAI222_X1 U11705 ( .A1(P1_U3086), .A2(n10939), .B1(n14373), .B2(n9182), .C1(
        n9179), .C2(n14370), .ZN(P1_U3338) );
  NAND2_X1 U11706 ( .A1(n9441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9180) );
  XNOR2_X1 U11707 ( .A(n9180), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14853) );
  INV_X1 U11708 ( .A(n14853), .ZN(n13202) );
  OAI222_X1 U11709 ( .A1(P2_U3088), .A2(n13202), .B1(n13675), .B2(n9182), .C1(
        n9181), .C2(n11464), .ZN(P2_U3310) );
  OR2_X1 U11710 ( .A1(n9186), .A2(n11612), .ZN(n9189) );
  AOI22_X1 U11711 ( .A1(n11529), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11528), 
        .B2(n9187), .ZN(n9188) );
  NAND2_X1 U11712 ( .A1(n9189), .A2(n9188), .ZN(n11751) );
  NAND2_X1 U11713 ( .A1(n11751), .A2(n11699), .ZN(n9191) );
  NAND2_X1 U11714 ( .A1(n13830), .A2(n11698), .ZN(n9190) );
  NAND2_X1 U11715 ( .A1(n9191), .A2(n9190), .ZN(n9193) );
  XNOR2_X1 U11716 ( .A(n9193), .B(n9192), .ZN(n9195) );
  AOI22_X1 U11717 ( .A1(n11751), .A2(n11698), .B1(n11680), .B2(n13830), .ZN(
        n9194) );
  AND2_X1 U11718 ( .A1(n9195), .A2(n9194), .ZN(n9315) );
  INV_X1 U11719 ( .A(n9315), .ZN(n9196) );
  OR2_X1 U11720 ( .A1(n9195), .A2(n9194), .ZN(n9314) );
  NAND2_X1 U11721 ( .A1(n9196), .A2(n9314), .ZN(n9197) );
  XNOR2_X1 U11722 ( .A(n9316), .B(n9197), .ZN(n9214) );
  NAND2_X1 U11723 ( .A1(n13831), .A2(n14262), .ZN(n9207) );
  NAND2_X1 U11724 ( .A1(n11885), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9205) );
  INV_X1 U11725 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9198) );
  OR2_X1 U11726 ( .A1(n11888), .A2(n9198), .ZN(n9204) );
  NAND2_X1 U11727 ( .A1(n9199), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9324) );
  OR2_X1 U11728 ( .A1(n9199), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U11729 ( .A1(n9324), .A2(n9200), .ZN(n9321) );
  OR2_X1 U11730 ( .A1(n11704), .A2(n9321), .ZN(n9203) );
  OR2_X1 U11731 ( .A1(n11656), .A2(n9201), .ZN(n9202) );
  NAND4_X1 U11732 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n13829) );
  NAND2_X1 U11733 ( .A1(n13829), .A2(n14591), .ZN(n9206) );
  NAND2_X1 U11734 ( .A1(n9207), .A2(n9206), .ZN(n14700) );
  NOR2_X1 U11735 ( .A1(n14588), .A2(n9820), .ZN(n9208) );
  AOI211_X1 U11736 ( .C1(n13818), .C2(n14700), .A(n9209), .B(n9208), .ZN(n9213) );
  INV_X1 U11737 ( .A(n11751), .ZN(n9817) );
  NOR2_X1 U11738 ( .A1(n9817), .A2(n14717), .ZN(n14701) );
  NAND3_X1 U11739 ( .A1(n14701), .A2(n9211), .A3(n9210), .ZN(n9212) );
  OAI211_X1 U11740 ( .C1(n9214), .C2(n14574), .A(n9213), .B(n9212), .ZN(
        P1_U3227) );
  INV_X1 U11741 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9381) );
  MUX2_X1 U11742 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9381), .S(n9650), .Z(n9217) );
  OAI21_X1 U11743 ( .B1(n9377), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9215), .ZN(
        n9216) );
  NOR2_X1 U11744 ( .A1(n9216), .A2(n9217), .ZN(n9651) );
  AOI211_X1 U11745 ( .C1(n9217), .C2(n9216), .A(n14847), .B(n9651), .ZN(n9226)
         );
  OAI21_X1 U11746 ( .B1(n9377), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9218), .ZN(
        n9221) );
  INV_X1 U11747 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9219) );
  MUX2_X1 U11748 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n9219), .S(n9650), .Z(n9220) );
  NOR2_X1 U11749 ( .A1(n9221), .A2(n9220), .ZN(n9655) );
  AOI211_X1 U11750 ( .C1(n9221), .C2(n9220), .A(n14802), .B(n9655), .ZN(n9225)
         );
  AND2_X1 U11751 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9222) );
  AOI21_X1 U11752 ( .B1(n14840), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9222), .ZN(
        n9223) );
  OAI21_X1 U11753 ( .B1(n9650), .B2(n14846), .A(n9223), .ZN(n9224) );
  OR3_X1 U11754 ( .A1(n9226), .A2(n9225), .A3(n9224), .ZN(P2_U3224) );
  NAND2_X1 U11755 ( .A1(n12447), .A2(n9227), .ZN(n9228) );
  OR2_X1 U11756 ( .A1(n12236), .A2(SI_4_), .ZN(n9233) );
  OR2_X1 U11757 ( .A1(n11984), .A2(n9230), .ZN(n9232) );
  NAND2_X1 U11758 ( .A1(n10875), .A2(n14997), .ZN(n9231) );
  XNOR2_X1 U11759 ( .A(n9502), .B(n10289), .ZN(n9234) );
  NAND2_X1 U11760 ( .A1(n9506), .A2(n9234), .ZN(n9419) );
  OAI21_X1 U11761 ( .B1(n9506), .B2(n9234), .A(n9419), .ZN(n9235) );
  AOI21_X1 U11762 ( .B1(n9236), .B2(n9235), .A(n6785), .ZN(n9248) );
  NOR2_X1 U11763 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9237), .ZN(n14999) );
  NAND2_X1 U11764 ( .A1(n6639), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U11765 ( .A1(n6638), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11766 ( .A1(n9238), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11767 ( .A1(n9424), .A2(n9239), .ZN(n9414) );
  NAND2_X1 U11768 ( .A1(n12024), .A2(n9414), .ZN(n9242) );
  NAND2_X1 U11769 ( .A1(n12222), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9241) );
  INV_X1 U11770 ( .A(n9502), .ZN(n9369) );
  OAI22_X1 U11771 ( .A1(n10198), .A2(n12202), .B1(n9369), .B2(n12174), .ZN(
        n9245) );
  AOI211_X1 U11772 ( .C1(n12199), .C2(n12447), .A(n14999), .B(n9245), .ZN(
        n9247) );
  NAND2_X1 U11773 ( .A1(n12207), .A2(n9370), .ZN(n9246) );
  OAI211_X1 U11774 ( .C1(n9248), .C2(n12214), .A(n9247), .B(n9246), .ZN(
        P3_U3170) );
  INV_X1 U11775 ( .A(n9266), .ZN(n9251) );
  INV_X1 U11776 ( .A(n13151), .ZN(n11085) );
  NOR3_X1 U11777 ( .A1(n9249), .A2(n11085), .A3(n13048), .ZN(n9250) );
  AOI21_X1 U11778 ( .B1(n9251), .B2(n13133), .A(n9250), .ZN(n9270) );
  OR2_X1 U11779 ( .A1(n9791), .A2(n11236), .ZN(n9253) );
  AOI22_X1 U11780 ( .A1(n11358), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11169), 
        .B2(n14800), .ZN(n9252) );
  NAND2_X2 U11781 ( .A1(n9253), .A2(n9252), .ZN(n11089) );
  XNOR2_X1 U11782 ( .A(n11089), .B(n13067), .ZN(n9396) );
  NAND2_X1 U11783 ( .A1(n13150), .A2(n13066), .ZN(n9373) );
  XNOR2_X1 U11784 ( .A(n9396), .B(n9373), .ZN(n9269) );
  NOR2_X1 U11785 ( .A1(n14558), .A2(n9681), .ZN(n9263) );
  NAND2_X1 U11786 ( .A1(n13151), .A2(n13120), .ZN(n9261) );
  NAND2_X1 U11787 ( .A1(n11371), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9259) );
  OR2_X1 U11788 ( .A1(n6658), .A2(n9254), .ZN(n9258) );
  XNOR2_X1 U11789 ( .A(n9384), .B(n9383), .ZN(n9689) );
  OR2_X1 U11790 ( .A1(n6847), .A2(n9689), .ZN(n9257) );
  INV_X1 U11791 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9255) );
  OR2_X1 U11792 ( .A1(n11318), .A2(n9255), .ZN(n9256) );
  NAND2_X1 U11793 ( .A1(n13149), .A2(n13237), .ZN(n9260) );
  AND2_X1 U11794 ( .A1(n9261), .A2(n9260), .ZN(n9678) );
  NAND2_X1 U11795 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14794) );
  OAI21_X1 U11796 ( .B1(n9678), .B2(n14554), .A(n14794), .ZN(n9262) );
  AOI211_X1 U11797 ( .C1(n11089), .C2(n13128), .A(n9263), .B(n9262), .ZN(n9268) );
  AND2_X1 U11798 ( .A1(n9269), .A2(n9264), .ZN(n9265) );
  INV_X1 U11799 ( .A(n9376), .ZN(n9399) );
  NAND2_X1 U11800 ( .A1(n9399), .A2(n13133), .ZN(n9267) );
  OAI211_X1 U11801 ( .C1(n9270), .C2(n9269), .A(n9268), .B(n9267), .ZN(
        P2_U3193) );
  INV_X1 U11802 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11545) );
  XNOR2_X1 U11803 ( .A(n9403), .B(n11545), .ZN(n11981) );
  INV_X1 U11804 ( .A(n11981), .ZN(n9274) );
  INV_X1 U11805 ( .A(SI_20_), .ZN(n9587) );
  OAI222_X1 U11806 ( .A1(n12997), .A2(n9274), .B1(n12985), .B2(n9587), .C1(
        P3_U3151), .C2(n9273), .ZN(P3_U3275) );
  NAND2_X1 U11807 ( .A1(n9276), .A2(n9275), .ZN(n9278) );
  OR2_X1 U11808 ( .A1(n13157), .A2(n6820), .ZN(n9277) );
  NAND2_X1 U11809 ( .A1(n13156), .A2(n14916), .ZN(n9279) );
  NAND2_X1 U11810 ( .A1(n9557), .A2(n9559), .ZN(n9281) );
  OR2_X1 U11811 ( .A1(n13156), .A2(n11034), .ZN(n9280) );
  NAND2_X1 U11812 ( .A1(n13155), .A2(n14921), .ZN(n9282) );
  NAND2_X1 U11813 ( .A1(n10062), .A2(n11400), .ZN(n9285) );
  NAND2_X1 U11814 ( .A1(n9283), .A2(n14921), .ZN(n9284) );
  OR2_X1 U11815 ( .A1(n14926), .A2(n13154), .ZN(n9286) );
  NOR2_X1 U11816 ( .A1(n11068), .A2(n13153), .ZN(n9287) );
  NAND2_X1 U11817 ( .A1(n11068), .A2(n13153), .ZN(n9288) );
  INV_X1 U11818 ( .A(n11404), .ZN(n9301) );
  OAI21_X1 U11819 ( .B1(n9289), .B2(n9301), .A(n9540), .ZN(n9489) );
  NAND2_X1 U11820 ( .A1(n10064), .A2(n14921), .ZN(n10063) );
  OR2_X1 U11821 ( .A1(n10063), .A2(n14926), .ZN(n9482) );
  NAND2_X1 U11822 ( .A1(n9484), .A2(n11075), .ZN(n9290) );
  NAND2_X1 U11823 ( .A1(n9290), .A2(n13488), .ZN(n9291) );
  NOR2_X1 U11824 ( .A1(n9543), .A2(n9291), .ZN(n9496) );
  INV_X1 U11825 ( .A(n9559), .ZN(n11397) );
  NAND2_X1 U11826 ( .A1(n10055), .A2(n10054), .ZN(n9294) );
  INV_X1 U11827 ( .A(n11400), .ZN(n9293) );
  INV_X1 U11828 ( .A(n11402), .ZN(n9464) );
  NAND2_X1 U11829 ( .A1(n9296), .A2(n14926), .ZN(n9297) );
  INV_X1 U11830 ( .A(n11068), .ZN(n14936) );
  NAND2_X1 U11831 ( .A1(n14936), .A2(n13153), .ZN(n9298) );
  NAND2_X1 U11832 ( .A1(n9478), .A2(n9298), .ZN(n9300) );
  INV_X1 U11833 ( .A(n13153), .ZN(n11070) );
  NAND2_X1 U11834 ( .A1(n11068), .A2(n11070), .ZN(n9299) );
  NAND2_X1 U11835 ( .A1(n9300), .A2(n9299), .ZN(n9546) );
  XNOR2_X1 U11836 ( .A(n9546), .B(n9301), .ZN(n9303) );
  OAI21_X1 U11837 ( .B1(n9303), .B2(n13435), .A(n9302), .ZN(n9490) );
  AOI211_X1 U11838 ( .C1(n14938), .C2(n9489), .A(n9496), .B(n9490), .ZN(n9309)
         );
  NAND2_X1 U11839 ( .A1(n14960), .A2(n14927), .ZN(n13662) );
  NOR2_X1 U11840 ( .A1(n14960), .A2(n8914), .ZN(n9306) );
  AOI21_X1 U11841 ( .B1(n6902), .B2(n11075), .A(n9306), .ZN(n9307) );
  OAI21_X1 U11842 ( .B1(n9309), .B2(n14959), .A(n9307), .ZN(P2_U3448) );
  NAND2_X1 U11843 ( .A1(n14970), .A2(n14927), .ZN(n13616) );
  INV_X1 U11844 ( .A(n13616), .ZN(n10558) );
  AOI22_X1 U11845 ( .A1(n10558), .A2(n11075), .B1(n14968), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n9308) );
  OAI21_X1 U11846 ( .B1(n9309), .B2(n14968), .A(n9308), .ZN(P2_U3505) );
  AOI22_X1 U11847 ( .A1(n11529), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11528), 
        .B2(n9311), .ZN(n9312) );
  NAND2_X1 U11848 ( .A1(n9313), .A2(n9312), .ZN(n14712) );
  INV_X1 U11849 ( .A(n14712), .ZN(n9623) );
  INV_X1 U11850 ( .A(n13798), .ZN(n14581) );
  INV_X1 U11851 ( .A(n13829), .ZN(n9969) );
  NOR2_X1 U11852 ( .A1(n9969), .A2(n11696), .ZN(n9317) );
  AOI21_X1 U11853 ( .B1(n14712), .B2(n11698), .A(n9317), .ZN(n9521) );
  AOI22_X1 U11854 ( .A1(n14712), .A2(n11699), .B1(n11698), .B2(n13829), .ZN(
        n9318) );
  XNOR2_X1 U11855 ( .A(n9318), .B(n11678), .ZN(n9520) );
  XOR2_X1 U11856 ( .A(n9521), .B(n9520), .Z(n9319) );
  NAND2_X1 U11857 ( .A1(n9320), .A2(n9319), .ZN(n9519) );
  OAI211_X1 U11858 ( .C1(n9320), .C2(n9319), .A(n9519), .B(n14567), .ZN(n9335)
         );
  INV_X1 U11859 ( .A(n9321), .ZN(n9643) );
  NAND2_X1 U11860 ( .A1(n13830), .A2(n14262), .ZN(n9331) );
  NAND2_X1 U11861 ( .A1(n11885), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9329) );
  INV_X1 U11862 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9322) );
  OR2_X1 U11863 ( .A1(n11888), .A2(n9322), .ZN(n9328) );
  INV_X1 U11864 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11865 ( .A1(n9324), .A2(n9323), .ZN(n9325) );
  NAND2_X1 U11866 ( .A1(n9528), .A2(n9325), .ZN(n10032) );
  OR2_X1 U11867 ( .A1(n11671), .A2(n10032), .ZN(n9327) );
  OR2_X1 U11868 ( .A1(n11656), .A2(n8073), .ZN(n9326) );
  NAND4_X1 U11869 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n13828) );
  NAND2_X1 U11870 ( .A1(n13828), .A2(n14591), .ZN(n9330) );
  AND2_X1 U11871 ( .A1(n9331), .A2(n9330), .ZN(n9639) );
  OAI22_X1 U11872 ( .A1(n13776), .A2(n9639), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9332), .ZN(n9333) );
  AOI21_X1 U11873 ( .B1(n9643), .B2(n13778), .A(n9333), .ZN(n9334) );
  OAI211_X1 U11874 ( .C1(n9623), .C2(n14581), .A(n9335), .B(n9334), .ZN(
        P1_U3239) );
  INV_X1 U11875 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n15476) );
  NOR2_X1 U11876 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15476), .ZN(n9336) );
  AOI21_X1 U11877 ( .B1(n14656), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9336), .ZN(
        n9337) );
  INV_X1 U11878 ( .A(n9337), .ZN(n9342) );
  OAI21_X1 U11879 ( .B1(n10409), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9338), .ZN(
        n9340) );
  INV_X1 U11880 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10418) );
  MUX2_X1 U11881 ( .A(n10418), .B(P1_REG1_REG_13__SCAN_IN), .S(n10781), .Z(
        n9339) );
  NOR2_X1 U11882 ( .A1(n9340), .A2(n9339), .ZN(n9447) );
  AOI211_X1 U11883 ( .C1(n9340), .C2(n9339), .A(n9447), .B(n13886), .ZN(n9341)
         );
  AOI211_X1 U11884 ( .C1(n14665), .C2(n10781), .A(n9342), .B(n9341), .ZN(n9348) );
  NOR2_X1 U11885 ( .A1(n10409), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9343) );
  NOR2_X1 U11886 ( .A1(n9344), .A2(n9343), .ZN(n9346) );
  INV_X1 U11887 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10417) );
  MUX2_X1 U11888 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n10417), .S(n10781), .Z(
        n9345) );
  NAND2_X1 U11889 ( .A1(n9345), .A2(n9346), .ZN(n9450) );
  OAI211_X1 U11890 ( .C1(n9346), .C2(n9345), .A(n14669), .B(n9450), .ZN(n9347)
         );
  NAND2_X1 U11891 ( .A1(n9348), .A2(n9347), .ZN(P1_U3256) );
  NAND2_X1 U11892 ( .A1(n9349), .A2(n12282), .ZN(n15125) );
  NAND2_X1 U11893 ( .A1(n9359), .A2(n15137), .ZN(n12271) );
  INV_X1 U11894 ( .A(n15137), .ZN(n9358) );
  INV_X1 U11895 ( .A(n15126), .ZN(n9350) );
  NAND2_X1 U11896 ( .A1(n15129), .A2(n15120), .ZN(n12284) );
  NAND2_X1 U11897 ( .A1(n12447), .A2(n9351), .ZN(n12291) );
  NAND2_X1 U11898 ( .A1(n9506), .A2(n9502), .ZN(n12292) );
  NAND2_X1 U11899 ( .A1(n15115), .A2(n9369), .ZN(n12296) );
  XNOR2_X1 U11900 ( .A(n9500), .B(n12246), .ZN(n15179) );
  AND2_X1 U11901 ( .A1(n12423), .A2(n12275), .ZN(n15136) );
  AND2_X1 U11902 ( .A1(n15162), .A2(n15136), .ZN(n12704) );
  INV_X1 U11903 ( .A(n12704), .ZN(n12723) );
  INV_X1 U11904 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10094) );
  NAND3_X1 U11905 ( .A1(n9352), .A2(n12422), .A3(n15209), .ZN(n9354) );
  NAND2_X1 U11906 ( .A1(n9354), .A2(n9353), .ZN(n12697) );
  INV_X1 U11907 ( .A(n10198), .ZN(n15104) );
  AOI22_X1 U11908 ( .A1(n15149), .A2(n15104), .B1(n12447), .B2(n15148), .ZN(
        n9367) );
  NAND2_X1 U11909 ( .A1(n15145), .A2(n15142), .ZN(n9357) );
  NAND2_X1 U11910 ( .A1(n15131), .A2(n9355), .ZN(n9356) );
  NAND2_X1 U11911 ( .A1(n9357), .A2(n9356), .ZN(n15127) );
  NAND2_X1 U11912 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  NAND2_X1 U11913 ( .A1(n12447), .A2(n15120), .ZN(n9363) );
  NAND2_X1 U11914 ( .A1(n12275), .A2(n9364), .ZN(n12245) );
  OAI211_X1 U11915 ( .C1(n9365), .C2(n12246), .A(n9504), .B(n15133), .ZN(n9366) );
  OAI211_X1 U11916 ( .C1(n15179), .C2(n15146), .A(n9367), .B(n9366), .ZN(
        n15180) );
  INV_X1 U11917 ( .A(n15180), .ZN(n9368) );
  MUX2_X1 U11918 ( .A(n10094), .B(n9368), .S(n15162), .Z(n9372) );
  NOR2_X1 U11919 ( .A1(n9369), .A2(n15209), .ZN(n15181) );
  AOI22_X1 U11920 ( .A1(n15181), .A2(n15122), .B1(n15157), .B2(n9370), .ZN(
        n9371) );
  OAI211_X1 U11921 ( .C1(n15179), .C2(n12723), .A(n9372), .B(n9371), .ZN(
        P3_U3229) );
  INV_X1 U11922 ( .A(n9396), .ZN(n9374) );
  NAND2_X1 U11923 ( .A1(n9374), .A2(n9373), .ZN(n9375) );
  NAND2_X1 U11924 ( .A1(n9376), .A2(n9375), .ZN(n9380) );
  OR2_X1 U11925 ( .A1(n9964), .A2(n11236), .ZN(n9379) );
  AOI22_X1 U11926 ( .A1(n11358), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n11169), 
        .B2(n9377), .ZN(n9378) );
  XNOR2_X1 U11927 ( .A(n11094), .B(n13035), .ZN(n9740) );
  NAND2_X1 U11928 ( .A1(n13149), .A2(n13066), .ZN(n9741) );
  XNOR2_X1 U11929 ( .A(n9740), .B(n9741), .ZN(n9397) );
  NAND2_X1 U11930 ( .A1(n13150), .A2(n13120), .ZN(n9393) );
  NAND2_X1 U11931 ( .A1(n11371), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9391) );
  OR2_X1 U11932 ( .A1(n6658), .A2(n9381), .ZN(n9390) );
  NAND2_X1 U11933 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n9382) );
  INV_X1 U11934 ( .A(n9747), .ZN(n9386) );
  INV_X1 U11935 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9756) );
  OAI21_X1 U11936 ( .B1(n9384), .B2(n9383), .A(n9756), .ZN(n9385) );
  NAND2_X1 U11937 ( .A1(n9386), .A2(n9385), .ZN(n13514) );
  OR2_X1 U11938 ( .A1(n6847), .A2(n13514), .ZN(n9389) );
  INV_X1 U11939 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9387) );
  OR2_X1 U11940 ( .A1(n11318), .A2(n9387), .ZN(n9388) );
  NAND4_X1 U11941 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n13148) );
  NAND2_X1 U11942 ( .A1(n13148), .A2(n13237), .ZN(n9392) );
  NAND2_X1 U11943 ( .A1(n9393), .A2(n9392), .ZN(n9696) );
  AOI21_X1 U11944 ( .B1(n13137), .B2(n9696), .A(n9394), .ZN(n9395) );
  OAI21_X1 U11945 ( .B1(n9689), .B2(n14558), .A(n9395), .ZN(n9401) );
  AOI22_X1 U11946 ( .A1(n9396), .A2(n13133), .B1(n13111), .B2(n13150), .ZN(
        n9398) );
  NOR3_X1 U11947 ( .A1(n9399), .A2(n9398), .A3(n9397), .ZN(n9400) );
  AOI211_X1 U11948 ( .C1(n11094), .C2(n13128), .A(n9401), .B(n9400), .ZN(n9402) );
  OAI21_X1 U11949 ( .B1(n9744), .B2(n14552), .A(n9402), .ZN(P2_U3203) );
  INV_X1 U11950 ( .A(SI_21_), .ZN(n9412) );
  NAND2_X1 U11951 ( .A1(n9404), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9407) );
  INV_X1 U11952 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U11953 ( .A1(n11561), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9646) );
  INV_X1 U11954 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U11955 ( .A1(n11009), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9408) );
  NAND2_X1 U11956 ( .A1(n9646), .A2(n9408), .ZN(n9409) );
  NAND2_X1 U11957 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U11958 ( .A1(n9647), .A2(n9411), .ZN(n11985) );
  OAI222_X1 U11959 ( .A1(P3_U3151), .A2(n9413), .B1(n12985), .B2(n9412), .C1(
        n12997), .C2(n11985), .ZN(P3_U3274) );
  INV_X1 U11960 ( .A(n9414), .ZN(n9510) );
  OR2_X1 U11961 ( .A1(n12236), .A2(SI_5_), .ZN(n9418) );
  NAND2_X1 U11962 ( .A1(n10875), .A2(n15016), .ZN(n9416) );
  XNOR2_X1 U11963 ( .A(n12117), .B(n9512), .ZN(n9594) );
  XNOR2_X1 U11964 ( .A(n9594), .B(n10198), .ZN(n9421) );
  OAI21_X1 U11965 ( .B1(n9421), .B2(n9420), .A(n9846), .ZN(n9422) );
  NAND2_X1 U11966 ( .A1(n9422), .A2(n12168), .ZN(n9432) );
  NOR2_X1 U11967 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9423), .ZN(n15018) );
  NAND2_X1 U11968 ( .A1(n6638), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U11969 ( .A1(n6639), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11970 ( .A1(n9424), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11971 ( .A1(n9602), .A2(n9425), .ZN(n15110) );
  NAND2_X1 U11972 ( .A1(n12024), .A2(n15110), .ZN(n9427) );
  NAND2_X1 U11973 ( .A1(n12222), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9426) );
  INV_X1 U11974 ( .A(n9512), .ZN(n15184) );
  OAI22_X1 U11975 ( .A1(n10195), .A2(n12202), .B1(n15184), .B2(n12174), .ZN(
        n9430) );
  AOI211_X1 U11976 ( .C1(n12199), .C2(n15115), .A(n15018), .B(n9430), .ZN(
        n9431) );
  OAI211_X1 U11977 ( .C1(n9510), .C2(n9958), .A(n9432), .B(n9431), .ZN(
        P3_U3167) );
  NAND2_X1 U11978 ( .A1(n9436), .A2(n9435), .ZN(n9437) );
  NAND2_X1 U11979 ( .A1(n9583), .A2(n9578), .ZN(n9438) );
  NAND2_X1 U11980 ( .A1(n9775), .A2(n9438), .ZN(n9439) );
  MUX2_X1 U11981 ( .A(n9446), .B(n9443), .S(n6641), .Z(n9579) );
  NAND2_X1 U11982 ( .A1(n9439), .A2(n9579), .ZN(n9440) );
  OAI21_X1 U11983 ( .B1(n9441), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9442) );
  XNOR2_X1 U11984 ( .A(n9442), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13218) );
  INV_X1 U11985 ( .A(n13218), .ZN(n13213) );
  OAI222_X1 U11986 ( .A1(n11464), .A2(n9443), .B1(n13675), .B2(n11514), .C1(
        n13213), .C2(P2_U3088), .ZN(P2_U3309) );
  NAND2_X1 U11987 ( .A1(n9444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9445) );
  XNOR2_X1 U11988 ( .A(n9445), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13875) );
  INV_X1 U11989 ( .A(n13875), .ZN(n10945) );
  OAI222_X1 U11990 ( .A1(P1_U3086), .A2(n10945), .B1(n14373), .B2(n11514), 
        .C1(n9446), .C2(n14370), .ZN(P1_U3337) );
  INV_X1 U11991 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10792) );
  MUX2_X1 U11992 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10792), .S(n10786), .Z(
        n9449) );
  AOI21_X1 U11993 ( .B1(n10781), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9447), .ZN(
        n9448) );
  NAND2_X1 U11994 ( .A1(n9449), .A2(n9448), .ZN(n10393) );
  OAI21_X1 U11995 ( .B1(n9449), .B2(n9448), .A(n10393), .ZN(n9459) );
  INV_X1 U11996 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14596) );
  MUX2_X1 U11997 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14596), .S(n10786), .Z(
        n9453) );
  OAI21_X1 U11998 ( .B1(n9451), .B2(n10417), .A(n9450), .ZN(n9452) );
  NAND2_X1 U11999 ( .A1(n9453), .A2(n9452), .ZN(n10385) );
  OAI211_X1 U12000 ( .C1(n9453), .C2(n9452), .A(n14669), .B(n10385), .ZN(n9456) );
  NAND2_X1 U12001 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14569)
         );
  INV_X1 U12002 ( .A(n14569), .ZN(n9454) );
  AOI21_X1 U12003 ( .B1(n14656), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9454), .ZN(
        n9455) );
  OAI211_X1 U12004 ( .C1(n13885), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9458)
         );
  AOI21_X1 U12005 ( .B1(n14668), .B2(n9459), .A(n9458), .ZN(n9460) );
  INV_X1 U12006 ( .A(n9460), .ZN(P1_U3257) );
  AND2_X1 U12007 ( .A1(n14949), .A2(n6784), .ZN(n9461) );
  XNOR2_X1 U12008 ( .A(n9464), .B(n9462), .ZN(n14930) );
  OAI21_X1 U12009 ( .B1(n9465), .B2(n9464), .A(n9463), .ZN(n9467) );
  AOI21_X1 U12010 ( .B1(n9467), .B2(n13499), .A(n9466), .ZN(n14928) );
  INV_X2 U12011 ( .A(n13512), .ZN(n13471) );
  MUX2_X1 U12012 ( .A(n8398), .B(n14928), .S(n13471), .Z(n9475) );
  INV_X1 U12013 ( .A(n9482), .ZN(n9468) );
  AOI211_X1 U12014 ( .C1(n14926), .C2(n10063), .A(n13066), .B(n9468), .ZN(
        n14925) );
  INV_X1 U12015 ( .A(n9469), .ZN(n9470) );
  INV_X1 U12016 ( .A(n14926), .ZN(n9472) );
  OAI22_X1 U12017 ( .A1(n14868), .A2(n9472), .B1(n9471), .B2(n13515), .ZN(
        n9473) );
  AOI21_X1 U12018 ( .B1(n14925), .B2(n14862), .A(n9473), .ZN(n9474) );
  OAI211_X1 U12019 ( .C1(n13507), .C2(n14930), .A(n9475), .B(n9474), .ZN(
        P2_U3261) );
  XNOR2_X1 U12020 ( .A(n11068), .B(n11070), .ZN(n11403) );
  INV_X1 U12021 ( .A(n11403), .ZN(n9477) );
  XNOR2_X1 U12022 ( .A(n9476), .B(n9477), .ZN(n14933) );
  XNOR2_X1 U12023 ( .A(n9478), .B(n9477), .ZN(n9480) );
  AOI21_X1 U12024 ( .B1(n9480), .B2(n13499), .A(n9479), .ZN(n14941) );
  MUX2_X1 U12025 ( .A(n9481), .B(n14941), .S(n13471), .Z(n9488) );
  AOI21_X1 U12026 ( .B1(n9482), .B2(n11068), .A(n13066), .ZN(n9483) );
  AND2_X1 U12027 ( .A1(n9484), .A2(n9483), .ZN(n14934) );
  OAI22_X1 U12028 ( .A1(n14868), .A2(n14936), .B1(n13515), .B2(n9485), .ZN(
        n9486) );
  AOI21_X1 U12029 ( .B1(n14934), .B2(n14862), .A(n9486), .ZN(n9487) );
  OAI211_X1 U12030 ( .C1(n13507), .C2(n14933), .A(n9488), .B(n9487), .ZN(
        P2_U3260) );
  INV_X1 U12031 ( .A(n9489), .ZN(n9499) );
  INV_X1 U12032 ( .A(n9490), .ZN(n9491) );
  MUX2_X1 U12033 ( .A(n9492), .B(n9491), .S(n13471), .Z(n9498) );
  OAI22_X1 U12034 ( .A1(n9494), .A2(n14868), .B1(n13515), .B2(n9493), .ZN(
        n9495) );
  AOI21_X1 U12035 ( .B1(n9496), .B2(n14862), .A(n9495), .ZN(n9497) );
  OAI211_X1 U12036 ( .C1(n13507), .C2(n9499), .A(n9498), .B(n9497), .ZN(
        P2_U3259) );
  NAND2_X1 U12037 ( .A1(n10198), .A2(n9512), .ZN(n12299) );
  NAND2_X1 U12038 ( .A1(n15104), .A2(n15184), .ZN(n12293) );
  INV_X1 U12039 ( .A(n12246), .ZN(n12289) );
  NAND2_X1 U12040 ( .A1(n9500), .A2(n12289), .ZN(n9501) );
  XOR2_X1 U12041 ( .A(n10193), .B(n12297), .Z(n15186) );
  NAND2_X1 U12042 ( .A1(n15115), .A2(n9502), .ZN(n9503) );
  INV_X1 U12043 ( .A(n12297), .ZN(n9505) );
  OAI21_X1 U12044 ( .B1(n6781), .B2(n9505), .A(n10200), .ZN(n9508) );
  OAI22_X1 U12045 ( .A1(n10195), .A2(n15128), .B1(n9506), .B2(n15130), .ZN(
        n9507) );
  AOI21_X1 U12046 ( .B1(n9508), .B2(n15133), .A(n9507), .ZN(n9509) );
  OAI21_X1 U12047 ( .B1(n15186), .B2(n15146), .A(n9509), .ZN(n15188) );
  NAND2_X1 U12048 ( .A1(n15188), .A2(n15162), .ZN(n9514) );
  INV_X1 U12049 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15009) );
  OAI22_X1 U12050 ( .A1(n15162), .A2(n15009), .B1(n9510), .B2(n12782), .ZN(
        n9511) );
  AOI21_X1 U12051 ( .B1(n12792), .B2(n9512), .A(n9511), .ZN(n9513) );
  OAI211_X1 U12052 ( .C1(n15186), .C2(n12723), .A(n9514), .B(n9513), .ZN(
        P3_U3228) );
  AOI22_X1 U12053 ( .A1(n11529), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11528), 
        .B2(n9516), .ZN(n9517) );
  INV_X1 U12054 ( .A(n13828), .ZN(n9986) );
  NOR2_X1 U12055 ( .A1(n9986), .A2(n11696), .ZN(n9522) );
  AOI21_X1 U12056 ( .B1(n14715), .B2(n11698), .A(n9522), .ZN(n9798) );
  AOI22_X1 U12057 ( .A1(n14715), .A2(n11699), .B1(n11698), .B2(n13828), .ZN(
        n9523) );
  INV_X2 U12058 ( .A(n9192), .ZN(n11678) );
  XNOR2_X1 U12059 ( .A(n9523), .B(n11678), .ZN(n9797) );
  XOR2_X1 U12060 ( .A(n9798), .B(n9797), .Z(n9524) );
  OAI211_X1 U12061 ( .C1(n9525), .C2(n9524), .A(n9796), .B(n14567), .ZN(n9538)
         );
  INV_X1 U12062 ( .A(n13806), .ZN(n14579) );
  NAND2_X1 U12063 ( .A1(n6644), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9533) );
  OR2_X1 U12064 ( .A1(n11881), .A2(n9526), .ZN(n9532) );
  NAND2_X1 U12065 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  NAND2_X1 U12066 ( .A1(n9802), .A2(n9529), .ZN(n10047) );
  OR2_X1 U12067 ( .A1(n11704), .A2(n10047), .ZN(n9531) );
  OR2_X1 U12068 ( .A1(n11656), .A2(n10048), .ZN(n9530) );
  NAND4_X1 U12069 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n13827) );
  NAND2_X1 U12070 ( .A1(n14577), .A2(n13829), .ZN(n9535) );
  OAI211_X1 U12071 ( .C1(n14588), .C2(n10032), .A(n9535), .B(n9534), .ZN(n9536) );
  AOI21_X1 U12072 ( .B1(n14579), .B2(n13827), .A(n9536), .ZN(n9537) );
  OAI211_X1 U12073 ( .C1(n7525), .C2(n14581), .A(n9538), .B(n9537), .ZN(
        P1_U3213) );
  OR2_X1 U12074 ( .A1(n11075), .A2(n13152), .ZN(n9539) );
  XNOR2_X1 U12075 ( .A(n11083), .B(n13151), .ZN(n11405) );
  INV_X1 U12076 ( .A(n11405), .ZN(n9541) );
  NAND2_X1 U12077 ( .A1(n9542), .A2(n9541), .ZN(n9669) );
  OAI21_X1 U12078 ( .B1(n9542), .B2(n9541), .A(n9669), .ZN(n14871) );
  INV_X1 U12079 ( .A(n9543), .ZN(n9545) );
  NAND2_X1 U12080 ( .A1(n9543), .A2(n14869), .ZN(n9680) );
  INV_X1 U12081 ( .A(n9680), .ZN(n9544) );
  AOI211_X1 U12082 ( .C1(n11083), .C2(n9545), .A(n13066), .B(n9544), .ZN(
        n14863) );
  NAND2_X1 U12083 ( .A1(n9546), .A2(n11404), .ZN(n9549) );
  NAND2_X1 U12084 ( .A1(n11075), .A2(n9547), .ZN(n9548) );
  NAND2_X1 U12085 ( .A1(n9549), .A2(n9548), .ZN(n9673) );
  XNOR2_X1 U12086 ( .A(n9673), .B(n11405), .ZN(n9551) );
  AOI21_X1 U12087 ( .B1(n9551), .B2(n13499), .A(n9550), .ZN(n14874) );
  INV_X1 U12088 ( .A(n14874), .ZN(n9552) );
  AOI211_X1 U12089 ( .C1(n14938), .C2(n14871), .A(n14863), .B(n9552), .ZN(
        n9556) );
  AOI22_X1 U12090 ( .A1(n11083), .A2(n10558), .B1(n14968), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n9553) );
  OAI21_X1 U12091 ( .B1(n9556), .B2(n14968), .A(n9553), .ZN(P2_U3506) );
  OAI22_X1 U12092 ( .A1(n14869), .A2(n13662), .B1(n14960), .B2(n9026), .ZN(
        n9554) );
  INV_X1 U12093 ( .A(n9554), .ZN(n9555) );
  OAI21_X1 U12094 ( .B1(n9556), .B2(n14959), .A(n9555), .ZN(P2_U3451) );
  XNOR2_X1 U12095 ( .A(n9557), .B(n9559), .ZN(n14913) );
  INV_X1 U12096 ( .A(n14913), .ZN(n9576) );
  NAND2_X1 U12097 ( .A1(n14913), .A2(n9558), .ZN(n9566) );
  NAND3_X1 U12098 ( .A1(n9561), .A2(n9560), .A3(n9559), .ZN(n9562) );
  NAND2_X1 U12099 ( .A1(n10055), .A2(n9562), .ZN(n9563) );
  NAND2_X1 U12100 ( .A1(n9563), .A2(n13499), .ZN(n9565) );
  NAND3_X1 U12101 ( .A1(n9566), .A2(n9565), .A3(n9564), .ZN(n14918) );
  NAND2_X1 U12102 ( .A1(n14918), .A2(n13471), .ZN(n9575) );
  NAND2_X1 U12103 ( .A1(n9567), .A2(n11034), .ZN(n9568) );
  NAND2_X1 U12104 ( .A1(n9568), .A2(n13488), .ZN(n9569) );
  OR2_X1 U12105 ( .A1(n10064), .A2(n9569), .ZN(n14914) );
  NOR2_X1 U12106 ( .A1(n13411), .A2(n14914), .ZN(n9573) );
  OAI22_X1 U12107 ( .A1(n13471), .A2(n9571), .B1(n9570), .B2(n13515), .ZN(
        n9572) );
  AOI211_X1 U12108 ( .C1(n13517), .C2(n11034), .A(n9573), .B(n9572), .ZN(n9574) );
  OAI211_X1 U12109 ( .C1(n9576), .C2(n9685), .A(n9575), .B(n9574), .ZN(
        P2_U3263) );
  INV_X1 U12110 ( .A(n9579), .ZN(n9577) );
  MUX2_X1 U12111 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6641), .Z(n9584) );
  XNOR2_X1 U12112 ( .A(n9584), .B(SI_19_), .ZN(n9777) );
  NOR2_X1 U12113 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  NOR2_X1 U12114 ( .A1(n9777), .A2(n9580), .ZN(n9581) );
  INV_X1 U12115 ( .A(n9584), .ZN(n9585) );
  INV_X1 U12116 ( .A(n9588), .ZN(n9586) );
  NAND2_X1 U12117 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  INV_X1 U12118 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9593) );
  MUX2_X1 U12119 ( .A(n11545), .B(n9593), .S(n6641), .Z(n9590) );
  NAND2_X1 U12120 ( .A1(n9591), .A2(n9590), .ZN(n9592) );
  NAND2_X1 U12121 ( .A1(n9936), .A2(n9592), .ZN(n11544) );
  OAI222_X1 U12122 ( .A1(P1_U3086), .A2(n11902), .B1(n14373), .B2(n11544), 
        .C1(n11545), .C2(n14370), .ZN(P1_U3335) );
  OAI222_X1 U12123 ( .A1(n11464), .A2(n9593), .B1(P2_U3088), .B2(n11427), .C1(
        n13675), .C2(n11544), .ZN(P2_U3307) );
  INV_X1 U12124 ( .A(n15110), .ZN(n9611) );
  INV_X1 U12125 ( .A(n9594), .ZN(n9595) );
  NAND2_X1 U12126 ( .A1(n10198), .A2(n9595), .ZN(n9843) );
  AND2_X1 U12127 ( .A1(n9846), .A2(n9843), .ZN(n9601) );
  NAND2_X1 U12128 ( .A1(n10875), .A2(n10105), .ZN(n9598) );
  OAI211_X1 U12129 ( .C1(n12236), .C2(n9599), .A(n9598), .B(n9597), .ZN(n15109) );
  XNOR2_X1 U12130 ( .A(n10289), .B(n15109), .ZN(n9842) );
  XNOR2_X1 U12131 ( .A(n12446), .B(n9842), .ZN(n9600) );
  NAND2_X1 U12132 ( .A1(n9601), .A2(n9600), .ZN(n9718) );
  OAI211_X1 U12133 ( .C1(n9601), .C2(n9600), .A(n9718), .B(n12168), .ZN(n9610)
         );
  AND2_X1 U12134 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U12135 ( .A1(n10884), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U12136 ( .A1(n6638), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U12137 ( .A1(n9602), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U12138 ( .A1(n9723), .A2(n9603), .ZN(n10210) );
  NAND2_X1 U12139 ( .A1(n8514), .A2(n10210), .ZN(n9605) );
  NAND2_X1 U12140 ( .A1(n9240), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9604) );
  INV_X1 U12141 ( .A(n15109), .ZN(n10196) );
  OAI22_X1 U12142 ( .A1(n9849), .A2(n12202), .B1(n10196), .B2(n12174), .ZN(
        n9608) );
  AOI211_X1 U12143 ( .C1(n12199), .C2(n15104), .A(n15035), .B(n9608), .ZN(
        n9609) );
  OAI211_X1 U12144 ( .C1(n9611), .C2(n9958), .A(n9610), .B(n9609), .ZN(
        P3_U3179) );
  AND2_X1 U12145 ( .A1(n9613), .A2(n9612), .ZN(n9614) );
  NAND2_X1 U12146 ( .A1(n11957), .A2(n9614), .ZN(n13954) );
  MUX2_X1 U12147 ( .A(n9617), .B(P1_REG2_REG_3__SCAN_IN), .S(n14689), .Z(n9618) );
  INV_X1 U12148 ( .A(n9618), .ZN(n9621) );
  NOR2_X2 U12149 ( .A1(n14177), .A2(n14675), .ZN(n14201) );
  INV_X1 U12150 ( .A(n14683), .ZN(n14199) );
  INV_X1 U12151 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9619) );
  AOI22_X1 U12152 ( .A1(n14201), .A2(n7320), .B1(n14199), .B2(n9619), .ZN(
        n9620) );
  OAI211_X1 U12153 ( .C1(n14130), .C2(n9622), .A(n9621), .B(n9620), .ZN(
        P1_U3290) );
  OAI211_X1 U12154 ( .C1(n9624), .C2(n9623), .A(n10031), .B(n14504), .ZN(
        n14709) );
  NAND2_X1 U12155 ( .A1(n11743), .A2(n13831), .ZN(n9625) );
  OR2_X1 U12156 ( .A1(n11743), .A2(n13831), .ZN(n9627) );
  XNOR2_X1 U12157 ( .A(n11751), .B(n13830), .ZN(n11920) );
  INV_X1 U12158 ( .A(n11920), .ZN(n9815) );
  INV_X1 U12159 ( .A(n13830), .ZN(n9636) );
  NAND2_X1 U12160 ( .A1(n9817), .A2(n9636), .ZN(n9628) );
  XNOR2_X1 U12161 ( .A(n9983), .B(n7517), .ZN(n9629) );
  NAND2_X1 U12162 ( .A1(n9629), .A2(n14725), .ZN(n9641) );
  INV_X1 U12163 ( .A(n13831), .ZN(n9630) );
  AND2_X1 U12164 ( .A1(n9630), .A2(n11743), .ZN(n9631) );
  NAND2_X1 U12165 ( .A1(n9633), .A2(n13831), .ZN(n9634) );
  NOR2_X1 U12166 ( .A1(n11751), .A2(n9636), .ZN(n9635) );
  NAND2_X1 U12167 ( .A1(n11751), .A2(n9636), .ZN(n9637) );
  XNOR2_X1 U12168 ( .A(n9968), .B(n11922), .ZN(n9638) );
  NAND2_X1 U12169 ( .A1(n9638), .A2(n14592), .ZN(n9640) );
  NAND3_X1 U12170 ( .A1(n9641), .A2(n9640), .A3(n9639), .ZN(n14710) );
  MUX2_X1 U12171 ( .A(n14710), .B(P1_REG2_REG_6__SCAN_IN), .S(n14689), .Z(
        n9642) );
  INV_X1 U12172 ( .A(n9642), .ZN(n9645) );
  AOI22_X1 U12173 ( .A1(n14201), .A2(n14712), .B1(n14199), .B2(n9643), .ZN(
        n9644) );
  OAI211_X1 U12174 ( .C1(n14130), .C2(n14709), .A(n9645), .B(n9644), .ZN(
        P1_U3287) );
  INV_X1 U12175 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10320) );
  XNOR2_X1 U12176 ( .A(n10320), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9959) );
  XNOR2_X1 U12177 ( .A(n9960), .B(n9959), .ZN(n11996) );
  INV_X1 U12178 ( .A(n11996), .ZN(n9649) );
  OAI22_X1 U12179 ( .A1(n12429), .A2(P3_U3151), .B1(SI_22_), .B2(n12985), .ZN(
        n9648) );
  AOI21_X1 U12180 ( .B1(n9649), .B2(n12979), .A(n9648), .ZN(P3_U3273) );
  INV_X1 U12181 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9891) );
  XNOR2_X1 U12182 ( .A(n13169), .B(n9891), .ZN(n9654) );
  INV_X1 U12183 ( .A(n9650), .ZN(n9733) );
  INV_X1 U12184 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9652) );
  MUX2_X1 U12185 ( .A(n9652), .B(P2_REG1_REG_11__SCAN_IN), .S(n14815), .Z(
        n14811) );
  OAI21_X1 U12186 ( .B1(n9654), .B2(n9653), .A(n13168), .ZN(n9666) );
  AOI21_X1 U12187 ( .B1(n9733), .B2(P2_REG2_REG_10__SCAN_IN), .A(n9655), .ZN(
        n14817) );
  INV_X1 U12188 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9656) );
  MUX2_X1 U12189 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9656), .S(n14815), .Z(
        n14818) );
  NAND2_X1 U12190 ( .A1(n14817), .A2(n14818), .ZN(n14816) );
  OR2_X1 U12191 ( .A1(n14815), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9659) );
  INV_X1 U12192 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9657) );
  MUX2_X1 U12193 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n9657), .S(n13169), .Z(
        n9658) );
  INV_X1 U12194 ( .A(n9658), .ZN(n9660) );
  AOI21_X1 U12195 ( .B1(n14816), .B2(n9659), .A(n9660), .ZN(n13160) );
  INV_X1 U12196 ( .A(n13160), .ZN(n9662) );
  NAND3_X1 U12197 ( .A1(n14816), .A2(n9660), .A3(n9659), .ZN(n9661) );
  AOI21_X1 U12198 ( .B1(n9662), .B2(n9661), .A(n14802), .ZN(n9665) );
  NAND2_X1 U12199 ( .A1(n14840), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12200 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9919) );
  OAI211_X1 U12201 ( .C1(n14846), .C2(n13161), .A(n9663), .B(n9919), .ZN(n9664) );
  AOI211_X1 U12202 ( .C1(n9666), .C2(n13225), .A(n9665), .B(n9664), .ZN(n9667)
         );
  INV_X1 U12203 ( .A(n9667), .ZN(P2_U3226) );
  OR2_X1 U12204 ( .A1(n11083), .A2(n13151), .ZN(n9668) );
  XNOR2_X1 U12205 ( .A(n11089), .B(n13150), .ZN(n11407) );
  NAND2_X1 U12206 ( .A1(n9670), .A2(n11407), .ZN(n9671) );
  NAND2_X1 U12207 ( .A1(n9687), .A2(n9671), .ZN(n14942) );
  AND2_X1 U12208 ( .A1(n11083), .A2(n11085), .ZN(n9672) );
  OR2_X1 U12209 ( .A1(n11083), .A2(n11085), .ZN(n9674) );
  INV_X1 U12210 ( .A(n11407), .ZN(n9675) );
  XNOR2_X1 U12211 ( .A(n9694), .B(n9675), .ZN(n9676) );
  NAND2_X1 U12212 ( .A1(n9676), .A2(n13499), .ZN(n9677) );
  OAI211_X1 U12213 ( .C1(n14942), .C2(n14949), .A(n9678), .B(n9677), .ZN(
        n14946) );
  MUX2_X1 U12214 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14946), .S(n13471), .Z(
        n9679) );
  INV_X1 U12215 ( .A(n9679), .ZN(n9684) );
  AOI211_X1 U12216 ( .C1(n11089), .C2(n9680), .A(n13066), .B(n9688), .ZN(
        n14943) );
  INV_X1 U12217 ( .A(n11089), .ZN(n14945) );
  OAI22_X1 U12218 ( .A1(n14945), .A2(n14868), .B1(n9681), .B2(n13515), .ZN(
        n9682) );
  AOI21_X1 U12219 ( .B1(n14943), .B2(n14862), .A(n9682), .ZN(n9683) );
  OAI211_X1 U12220 ( .C1(n14942), .C2(n9685), .A(n9684), .B(n9683), .ZN(
        P2_U3257) );
  INV_X1 U12221 ( .A(n13149), .ZN(n11096) );
  NAND2_X1 U12222 ( .A1(n11089), .A2(n13150), .ZN(n9686) );
  XOR2_X1 U12223 ( .A(n11409), .B(n10230), .Z(n14957) );
  INV_X1 U12224 ( .A(n14957), .ZN(n14950) );
  INV_X1 U12225 ( .A(n11094), .ZN(n14954) );
  NAND2_X1 U12226 ( .A1(n14954), .A2(n9688), .ZN(n10231) );
  OAI211_X1 U12227 ( .C1(n14954), .C2(n9688), .A(n13488), .B(n10231), .ZN(
        n14951) );
  INV_X1 U12228 ( .A(n14951), .ZN(n9691) );
  OAI22_X1 U12229 ( .A1(n14954), .A2(n14868), .B1(n13515), .B2(n9689), .ZN(
        n9690) );
  AOI21_X1 U12230 ( .B1(n9691), .B2(n14862), .A(n9690), .ZN(n9699) );
  NOR2_X1 U12231 ( .A1(n11089), .A2(n9692), .ZN(n9693) );
  AOI21_X1 U12232 ( .B1(n9695), .B2(n11409), .A(n13435), .ZN(n9697) );
  AOI21_X1 U12233 ( .B1(n9697), .B2(n10234), .A(n9696), .ZN(n14952) );
  MUX2_X1 U12234 ( .A(n15485), .B(n14952), .S(n13471), .Z(n9698) );
  OAI211_X1 U12235 ( .C1(n14950), .C2(n13507), .A(n9699), .B(n9698), .ZN(
        P2_U3256) );
  OAI211_X1 U12236 ( .C1(n12429), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9703)
         );
  NAND2_X1 U12237 ( .A1(n9703), .A2(n12397), .ZN(n9705) );
  NAND2_X1 U12238 ( .A1(n9705), .A2(n9704), .ZN(n9711) );
  NAND2_X1 U12239 ( .A1(n9707), .A2(n9706), .ZN(n9709) );
  NAND2_X1 U12240 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  NAND2_X1 U12241 ( .A1(n9711), .A2(n9710), .ZN(n9712) );
  NOR2_X4 U12242 ( .A1(n9713), .A2(n9712), .ZN(n15227) );
  INV_X1 U12243 ( .A(n12918), .ZN(n12878) );
  AOI22_X1 U12244 ( .A1(n12878), .A2(n9714), .B1(n15231), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n9715) );
  OAI21_X1 U12245 ( .B1(n9716), .B2(n15231), .A(n9715), .ZN(P3_U3459) );
  INV_X1 U12246 ( .A(n9842), .ZN(n9717) );
  NAND2_X1 U12247 ( .A1(n12446), .A2(n9717), .ZN(n9847) );
  NAND2_X1 U12248 ( .A1(n9718), .A2(n9847), .ZN(n10164) );
  OR2_X1 U12249 ( .A1(n12236), .A2(SI_7_), .ZN(n9721) );
  NAND2_X1 U12250 ( .A1(n10875), .A2(n15051), .ZN(n9720) );
  NAND2_X1 U12251 ( .A1(n9849), .A2(n10215), .ZN(n12306) );
  XNOR2_X1 U12252 ( .A(n10164), .B(n10163), .ZN(n9732) );
  NOR2_X1 U12253 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9722), .ZN(n15053) );
  NAND2_X1 U12254 ( .A1(n6639), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U12255 ( .A1(n6638), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U12256 ( .A1(n9723), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12257 ( .A1(n9832), .A2(n9724), .ZN(n10224) );
  NAND2_X1 U12258 ( .A1(n12024), .A2(n10224), .ZN(n9726) );
  NAND2_X1 U12259 ( .A1(n12222), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9725) );
  OAI22_X1 U12260 ( .A1(n10479), .A2(n12202), .B1(n12174), .B2(n10209), .ZN(
        n9729) );
  AOI211_X1 U12261 ( .C1(n12199), .C2(n12446), .A(n15053), .B(n9729), .ZN(
        n9731) );
  NAND2_X1 U12262 ( .A1(n12207), .A2(n10210), .ZN(n9730) );
  OAI211_X1 U12263 ( .C1(n9732), .C2(n12214), .A(n9731), .B(n9730), .ZN(
        P3_U3153) );
  OR2_X1 U12264 ( .A1(n9999), .A2(n11236), .ZN(n9735) );
  AOI22_X1 U12265 ( .A1(n11358), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11169), 
        .B2(n9733), .ZN(n9734) );
  NAND2_X2 U12266 ( .A1(n9735), .A2(n9734), .ZN(n13518) );
  XNOR2_X1 U12267 ( .A(n13518), .B(n13035), .ZN(n9886) );
  AND2_X1 U12268 ( .A1(n13148), .A2(n13030), .ZN(n9736) );
  NAND2_X1 U12269 ( .A1(n9886), .A2(n9736), .ZN(n9883) );
  INV_X1 U12270 ( .A(n9886), .ZN(n9738) );
  INV_X1 U12271 ( .A(n9736), .ZN(n9737) );
  NAND2_X1 U12272 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  AND2_X1 U12273 ( .A1(n9883), .A2(n9739), .ZN(n9746) );
  INV_X1 U12274 ( .A(n9740), .ZN(n9742) );
  NAND2_X1 U12275 ( .A1(n9742), .A2(n9741), .ZN(n9743) );
  INV_X1 U12276 ( .A(n9885), .ZN(n9888) );
  OAI211_X1 U12277 ( .C1(n9746), .C2(n9745), .A(n9888), .B(n13133), .ZN(n9760)
         );
  INV_X1 U12278 ( .A(n13514), .ZN(n9758) );
  NAND2_X1 U12279 ( .A1(n13149), .A2(n13120), .ZN(n9755) );
  NAND2_X1 U12280 ( .A1(n11277), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9753) );
  OR2_X1 U12281 ( .A1(n11317), .A2(n9656), .ZN(n9752) );
  NOR2_X1 U12282 ( .A1(n9747), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9748) );
  OR2_X1 U12283 ( .A1(n9892), .A2(n9748), .ZN(n10361) );
  OR2_X1 U12284 ( .A1(n6847), .A2(n10361), .ZN(n9751) );
  INV_X1 U12285 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9749) );
  OR2_X1 U12286 ( .A1(n11318), .A2(n9749), .ZN(n9750) );
  NAND4_X1 U12287 ( .A1(n9753), .A2(n9752), .A3(n9751), .A4(n9750), .ZN(n13147) );
  NAND2_X1 U12288 ( .A1(n13147), .A2(n13237), .ZN(n9754) );
  AND2_X1 U12289 ( .A1(n9755), .A2(n9754), .ZN(n10237) );
  OAI22_X1 U12290 ( .A1(n10237), .A2(n14554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9756), .ZN(n9757) );
  AOI21_X1 U12291 ( .B1(n13121), .B2(n9758), .A(n9757), .ZN(n9759) );
  OAI211_X1 U12292 ( .C1(n7107), .C2(n14550), .A(n9760), .B(n9759), .ZN(
        P2_U3189) );
  INV_X1 U12293 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9761) );
  INV_X1 U12294 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9763) );
  INV_X1 U12295 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9765) );
  INV_X1 U12296 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U12297 ( .A1(n12058), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9769) );
  NAND2_X1 U12298 ( .A1(n12620), .A2(n9769), .ZN(n12643) );
  INV_X1 U12299 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12300 ( .A1(n6639), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U12301 ( .A1(n12222), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9770) );
  OAI211_X1 U12302 ( .C1(n9772), .C2(n12062), .A(n9771), .B(n9770), .ZN(n9773)
         );
  AOI21_X1 U12303 ( .B1(n12643), .B2(n12024), .A(n9773), .ZN(n12653) );
  INV_X1 U12304 ( .A(P3_U3897), .ZN(n12449) );
  NAND2_X1 U12305 ( .A1(n12449), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n9774) );
  OAI21_X1 U12306 ( .B1(n12653), .B2(n12449), .A(n9774), .ZN(P3_U3519) );
  NAND2_X1 U12307 ( .A1(n9776), .A2(n9775), .ZN(n9778) );
  XNOR2_X1 U12308 ( .A(n9778), .B(n9777), .ZN(n11527) );
  INV_X1 U12309 ( .A(n11527), .ZN(n11462) );
  OAI222_X1 U12310 ( .A1(n13891), .A2(P1_U3086), .B1(n14373), .B2(n11462), 
        .C1(n9779), .C2(n14370), .ZN(P1_U3336) );
  INV_X1 U12311 ( .A(n12620), .ZN(n9780) );
  NAND2_X1 U12312 ( .A1(n9780), .A2(n12024), .ZN(n12228) );
  INV_X1 U12313 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U12314 ( .A1(n12222), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U12315 ( .A1(n6639), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9781) );
  OAI211_X1 U12316 ( .C1(n12062), .C2(n12624), .A(n9782), .B(n9781), .ZN(n9783) );
  INV_X1 U12317 ( .A(n9783), .ZN(n9784) );
  NAND2_X1 U12318 ( .A1(n12449), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n9785) );
  OAI21_X1 U12319 ( .B1(n12241), .B2(n12449), .A(n9785), .ZN(P3_U3521) );
  INV_X1 U12320 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n15392) );
  NAND2_X1 U12321 ( .A1(n6639), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U12322 ( .A1(n6638), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9786) );
  OAI211_X1 U12323 ( .C1(n10977), .C2(n15392), .A(n9787), .B(n9786), .ZN(n9788) );
  INV_X1 U12324 ( .A(n9788), .ZN(n9789) );
  NAND2_X1 U12325 ( .A1(n12449), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n9790) );
  OAI21_X1 U12326 ( .B1(n12636), .B2(n12449), .A(n9790), .ZN(P3_U3520) );
  OR2_X1 U12327 ( .A1(n9791), .A2(n11612), .ZN(n9794) );
  AOI22_X1 U12328 ( .A1(n11529), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11528), 
        .B2(n9792), .ZN(n9793) );
  NAND2_X1 U12329 ( .A1(n9794), .A2(n9793), .ZN(n11765) );
  AOI22_X1 U12330 ( .A1(n11765), .A2(n11699), .B1(n11698), .B2(n13827), .ZN(
        n9795) );
  XNOR2_X1 U12331 ( .A(n9795), .B(n11678), .ZN(n10519) );
  AOI22_X1 U12332 ( .A1(n11765), .A2(n11698), .B1(n11680), .B2(n13827), .ZN(
        n10520) );
  XNOR2_X1 U12333 ( .A(n10519), .B(n10520), .ZN(n9800) );
  OAI21_X1 U12334 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(n9799) );
  AOI21_X1 U12335 ( .B1(n9800), .B2(n9799), .A(n10518), .ZN(n9814) );
  NAND2_X1 U12336 ( .A1(n6644), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9808) );
  OR2_X1 U12337 ( .A1(n11881), .A2(n9801), .ZN(n9807) );
  INV_X1 U12338 ( .A(n10007), .ZN(n9804) );
  NAND2_X1 U12339 ( .A1(n9802), .A2(n10523), .ZN(n9803) );
  NAND2_X1 U12340 ( .A1(n9804), .A2(n9803), .ZN(n10524) );
  OR2_X1 U12341 ( .A1(n11704), .A2(n10524), .ZN(n9806) );
  OR2_X1 U12342 ( .A1(n11656), .A2(n8464), .ZN(n9805) );
  OR2_X1 U12343 ( .A1(n11775), .A2(n14141), .ZN(n9810) );
  NAND2_X1 U12344 ( .A1(n13828), .A2(n14262), .ZN(n9809) );
  NAND2_X1 U12345 ( .A1(n9810), .A2(n9809), .ZN(n10043) );
  AOI22_X1 U12346 ( .A1(n13818), .A2(n10043), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9811) );
  OAI21_X1 U12347 ( .B1(n10047), .B2(n14588), .A(n9811), .ZN(n9812) );
  AOI21_X1 U12348 ( .B1(n11765), .B2(n13798), .A(n9812), .ZN(n9813) );
  OAI21_X1 U12349 ( .B1(n9814), .B2(n14574), .A(n9813), .ZN(P1_U3221) );
  XNOR2_X1 U12350 ( .A(n9816), .B(n9815), .ZN(n14707) );
  NAND2_X1 U12351 ( .A1(n14686), .A2(n14725), .ZN(n14153) );
  XNOR2_X1 U12352 ( .A(n9818), .B(n9817), .ZN(n9819) );
  NAND2_X1 U12353 ( .A1(n9819), .A2(n14504), .ZN(n14702) );
  NOR2_X1 U12354 ( .A1(n14683), .A2(n9820), .ZN(n9821) );
  AOI21_X1 U12355 ( .B1(n14201), .B2(n11751), .A(n9821), .ZN(n9824) );
  INV_X1 U12356 ( .A(n14700), .ZN(n9822) );
  MUX2_X1 U12357 ( .A(n9822), .B(n15340), .S(n14689), .Z(n9823) );
  OAI211_X1 U12358 ( .C1(n14702), .C2(n14130), .A(n9824), .B(n9823), .ZN(n9827) );
  XNOR2_X1 U12359 ( .A(n9825), .B(n11920), .ZN(n14705) );
  NOR2_X1 U12360 ( .A1(n14177), .A2(n14704), .ZN(n14510) );
  INV_X1 U12361 ( .A(n14510), .ZN(n14188) );
  NOR2_X1 U12362 ( .A1(n14705), .A2(n14188), .ZN(n9826) );
  AOI211_X1 U12363 ( .C1(n14707), .C2(n14605), .A(n9827), .B(n9826), .ZN(n9828) );
  INV_X1 U12364 ( .A(n9828), .ZN(P1_U3288) );
  OR2_X1 U12365 ( .A1(n12236), .A2(SI_9_), .ZN(n9831) );
  OR2_X1 U12366 ( .A1(n11984), .A2(n9829), .ZN(n9830) );
  OAI211_X1 U12367 ( .C1(n10145), .C2(n10270), .A(n9831), .B(n9830), .ZN(
        n10533) );
  XNOR2_X1 U12368 ( .A(n10289), .B(n10533), .ZN(n9943) );
  NAND2_X1 U12369 ( .A1(n6639), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U12370 ( .A1(n9832), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U12371 ( .A1(n9859), .A2(n9833), .ZN(n10484) );
  NAND2_X1 U12372 ( .A1(n12024), .A2(n10484), .ZN(n9836) );
  NAND2_X1 U12373 ( .A1(n12222), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U12374 ( .A1(n6638), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9834) );
  NAND4_X1 U12375 ( .A1(n9837), .A2(n9836), .A3(n9835), .A4(n9834), .ZN(n12444) );
  XNOR2_X1 U12376 ( .A(n9943), .B(n12444), .ZN(n9857) );
  OR2_X1 U12377 ( .A1(n11984), .A2(n9838), .ZN(n9840) );
  NAND2_X1 U12378 ( .A1(n10875), .A2(n10114), .ZN(n9839) );
  OAI211_X1 U12379 ( .C1(n12236), .C2(n9841), .A(n9840), .B(n9839), .ZN(n10223) );
  XNOR2_X1 U12380 ( .A(n12117), .B(n10223), .ZN(n9851) );
  XNOR2_X1 U12381 ( .A(n9851), .B(n10479), .ZN(n10165) );
  NAND2_X1 U12382 ( .A1(n10195), .A2(n9842), .ZN(n9844) );
  AND4_X1 U12383 ( .A1(n10163), .A2(n10165), .A3(n9844), .A4(n9843), .ZN(n9845) );
  NAND2_X1 U12384 ( .A1(n9846), .A2(n9845), .ZN(n9855) );
  INV_X1 U12385 ( .A(n10165), .ZN(n9850) );
  OAI21_X1 U12386 ( .B1(n9850), .B2(n9847), .A(n10163), .ZN(n9853) );
  INV_X1 U12387 ( .A(n10163), .ZN(n9848) );
  OAI21_X1 U12388 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9852) );
  AOI22_X1 U12389 ( .A1(n9853), .A2(n9852), .B1(n9851), .B2(n12445), .ZN(n9854) );
  INV_X1 U12390 ( .A(n9952), .ZN(n9948) );
  AOI21_X1 U12391 ( .B1(n9857), .B2(n9856), .A(n9948), .ZN(n9869) );
  NOR2_X1 U12392 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9858), .ZN(n15091) );
  NAND2_X1 U12393 ( .A1(n6639), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U12394 ( .A1(n9859), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12395 ( .A1(n9861), .A2(n9860), .ZN(n9942) );
  NAND2_X1 U12396 ( .A1(n12024), .A2(n9942), .ZN(n9864) );
  NAND2_X1 U12397 ( .A1(n6638), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U12398 ( .A1(n9240), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9862) );
  NAND4_X1 U12399 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(n12443) );
  INV_X1 U12400 ( .A(n12443), .ZN(n12324) );
  OAI22_X1 U12401 ( .A1(n12324), .A2(n12202), .B1(n12174), .B2(n10533), .ZN(
        n9866) );
  AOI211_X1 U12402 ( .C1(n12199), .C2(n12445), .A(n15091), .B(n9866), .ZN(
        n9868) );
  NAND2_X1 U12403 ( .A1(n12207), .A2(n10484), .ZN(n9867) );
  OAI211_X1 U12404 ( .C1(n9869), .C2(n12214), .A(n9868), .B(n9867), .ZN(
        P3_U3171) );
  MUX2_X1 U12405 ( .A(n9870), .B(P1_REG2_REG_4__SCAN_IN), .S(n14689), .Z(n9877) );
  INV_X1 U12406 ( .A(n9871), .ZN(n9875) );
  NAND2_X1 U12407 ( .A1(n14201), .A2(n11743), .ZN(n9874) );
  NAND2_X1 U12408 ( .A1(n14199), .A2(n9872), .ZN(n9873) );
  OAI211_X1 U12409 ( .C1(n9875), .C2(n14130), .A(n9874), .B(n9873), .ZN(n9876)
         );
  AOI211_X1 U12410 ( .C1(n9878), .C2(n14510), .A(n9877), .B(n9876), .ZN(n9879)
         );
  OAI21_X1 U12411 ( .B1(n14153), .B2(n9880), .A(n9879), .ZN(P1_U3289) );
  NAND2_X1 U12412 ( .A1(n10245), .A2(n11362), .ZN(n9882) );
  AOI22_X1 U12413 ( .A1(n11358), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11169), 
        .B2(n14815), .ZN(n9881) );
  NAND2_X2 U12414 ( .A1(n9882), .A2(n9881), .ZN(n11107) );
  NAND2_X1 U12415 ( .A1(n13147), .A2(n13066), .ZN(n9904) );
  XNOR2_X1 U12416 ( .A(n9922), .B(n9904), .ZN(n9889) );
  INV_X1 U12417 ( .A(n9883), .ZN(n9884) );
  NAND3_X1 U12418 ( .A1(n9886), .A2(n13111), .A3(n13148), .ZN(n9887) );
  OAI21_X1 U12419 ( .B1(n9888), .B2(n14552), .A(n9887), .ZN(n9890) );
  NAND2_X1 U12420 ( .A1(n9890), .A2(n9889), .ZN(n9903) );
  NOR2_X1 U12421 ( .A1(n14558), .A2(n10361), .ZN(n9901) );
  NAND2_X1 U12422 ( .A1(n13148), .A2(n13120), .ZN(n9899) );
  NAND2_X1 U12423 ( .A1(n11372), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9897) );
  OR2_X1 U12424 ( .A1(n6658), .A2(n9891), .ZN(n9896) );
  OR2_X1 U12425 ( .A1(n11317), .A2(n9657), .ZN(n9895) );
  NOR2_X1 U12426 ( .A1(n9892), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9893) );
  OR2_X1 U12427 ( .A1(n9909), .A2(n9893), .ZN(n10374) );
  OR2_X1 U12428 ( .A1(n6847), .A2(n10374), .ZN(n9894) );
  NAND4_X1 U12429 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n13146) );
  NAND2_X1 U12430 ( .A1(n13146), .A2(n13237), .ZN(n9898) );
  AND2_X1 U12431 ( .A1(n9899), .A2(n9898), .ZN(n10357) );
  INV_X1 U12432 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n14809) );
  OAI22_X1 U12433 ( .A1(n10357), .A2(n14554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14809), .ZN(n9900) );
  OAI211_X1 U12434 ( .C1(n14552), .C2(n9924), .A(n9903), .B(n9902), .ZN(
        P2_U3208) );
  NAND2_X1 U12435 ( .A1(n9922), .A2(n9904), .ZN(n9905) );
  NAND2_X1 U12436 ( .A1(n10408), .A2(n11362), .ZN(n9907) );
  AOI22_X1 U12437 ( .A1(n11358), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11169), 
        .B2(n13169), .ZN(n9906) );
  XNOR2_X1 U12438 ( .A(n11116), .B(n13067), .ZN(n10326) );
  NAND2_X1 U12439 ( .A1(n13146), .A2(n13066), .ZN(n10327) );
  XNOR2_X1 U12440 ( .A(n10326), .B(n10327), .ZN(n9921) );
  NAND2_X1 U12441 ( .A1(n13147), .A2(n13120), .ZN(n9917) );
  NAND2_X1 U12442 ( .A1(n11277), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9915) );
  OR2_X1 U12443 ( .A1(n9909), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U12444 ( .A1(n10633), .A2(n9910), .ZN(n10338) );
  OR2_X1 U12445 ( .A1(n6847), .A2(n10338), .ZN(n9914) );
  INV_X1 U12446 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9911) );
  OR2_X1 U12447 ( .A1(n11318), .A2(n9911), .ZN(n9913) );
  INV_X1 U12448 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13162) );
  OR2_X1 U12449 ( .A1(n11317), .A2(n13162), .ZN(n9912) );
  NAND4_X1 U12450 ( .A1(n9915), .A2(n9914), .A3(n9913), .A4(n9912), .ZN(n13145) );
  NAND2_X1 U12451 ( .A1(n13145), .A2(n13237), .ZN(n9916) );
  NAND2_X1 U12452 ( .A1(n9917), .A2(n9916), .ZN(n10372) );
  NAND2_X1 U12453 ( .A1(n13137), .A2(n10372), .ZN(n9918) );
  OAI211_X1 U12454 ( .C1(n14558), .C2(n10374), .A(n9919), .B(n9918), .ZN(n9920) );
  AOI21_X1 U12455 ( .B1(n11116), .B2(n13128), .A(n9920), .ZN(n9926) );
  INV_X1 U12456 ( .A(n13147), .ZN(n11109) );
  OAI22_X1 U12457 ( .A1(n9922), .A2(n14552), .B1(n11109), .B2(n13048), .ZN(
        n9923) );
  NAND3_X1 U12458 ( .A1(n9924), .A2(n6935), .A3(n9923), .ZN(n9925) );
  OAI211_X1 U12459 ( .C1(n10330), .C2(n14552), .A(n9926), .B(n9925), .ZN(
        P2_U3196) );
  NOR2_X1 U12460 ( .A1(n13411), .A2(n9927), .ZN(n9930) );
  OAI22_X1 U12461 ( .A1(n13471), .A2(n8394), .B1(n9928), .B2(n13515), .ZN(
        n9929) );
  AOI211_X1 U12462 ( .C1(n13517), .C2(n6820), .A(n9930), .B(n9929), .ZN(n9933)
         );
  NAND2_X1 U12463 ( .A1(n9931), .A2(n14872), .ZN(n9932) );
  OAI211_X1 U12464 ( .C1(n13512), .C2(n9934), .A(n9933), .B(n9932), .ZN(
        P2_U3264) );
  MUX2_X1 U12465 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6641), .Z(n9937) );
  NAND2_X1 U12466 ( .A1(n9937), .A2(SI_21_), .ZN(n10313) );
  OAI21_X1 U12467 ( .B1(n9937), .B2(SI_21_), .A(n10313), .ZN(n9938) );
  INV_X1 U12468 ( .A(n9938), .ZN(n9939) );
  OR2_X1 U12469 ( .A1(n9940), .A2(n9939), .ZN(n9941) );
  NAND2_X1 U12470 ( .A1(n10314), .A2(n9941), .ZN(n11560) );
  OAI222_X1 U12471 ( .A1(n11464), .A2(n11009), .B1(P2_U3088), .B2(n11425), 
        .C1(n13675), .C2(n11560), .ZN(P2_U3306) );
  INV_X1 U12472 ( .A(n9942), .ZN(n10540) );
  NOR2_X1 U12473 ( .A1(n9943), .A2(n12444), .ZN(n9949) );
  NAND2_X1 U12474 ( .A1(n9944), .A2(n12235), .ZN(n9947) );
  NAND2_X1 U12475 ( .A1(n12069), .A2(n9945), .ZN(n9946) );
  OAI211_X1 U12476 ( .C1(n10178), .C2(n10270), .A(n9947), .B(n9946), .ZN(
        n15210) );
  XNOR2_X1 U12477 ( .A(n15210), .B(n10289), .ZN(n10267) );
  XNOR2_X1 U12478 ( .A(n10267), .B(n12443), .ZN(n9950) );
  OAI21_X1 U12479 ( .B1(n9948), .B2(n9949), .A(n9950), .ZN(n9953) );
  NOR2_X1 U12480 ( .A1(n9950), .A2(n9949), .ZN(n9951) );
  NAND3_X1 U12481 ( .A1(n9953), .A2(n12168), .A3(n10269), .ZN(n9957) );
  INV_X1 U12482 ( .A(n15210), .ZN(n10727) );
  NAND2_X1 U12483 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n10151)
         );
  NAND2_X1 U12484 ( .A1(n12444), .A2(n12199), .ZN(n9954) );
  OAI211_X1 U12485 ( .C1(n10757), .C2(n12202), .A(n10151), .B(n9954), .ZN(
        n9955) );
  AOI21_X1 U12486 ( .B1(n10727), .B2(n12212), .A(n9955), .ZN(n9956) );
  OAI211_X1 U12487 ( .C1(n10540), .C2(n9958), .A(n9957), .B(n9956), .ZN(
        P3_U3157) );
  INV_X1 U12488 ( .A(SI_23_), .ZN(n9963) );
  NAND2_X1 U12489 ( .A1(n10320), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9961) );
  XNOR2_X1 U12490 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n10465) );
  XNOR2_X1 U12491 ( .A(n10466), .B(n10465), .ZN(n12008) );
  NAND2_X1 U12492 ( .A1(n12008), .A2(n12979), .ZN(n9962) );
  OAI211_X1 U12493 ( .C1(n9963), .C2(n12985), .A(n9962), .B(n12432), .ZN(
        P3_U3272) );
  OR2_X1 U12494 ( .A1(n9964), .A2(n11612), .ZN(n9967) );
  AOI22_X1 U12495 ( .A1(n11529), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9965), 
        .B2(n11528), .ZN(n9966) );
  AND2_X2 U12496 ( .A1(n9967), .A2(n9966), .ZN(n11774) );
  INV_X1 U12497 ( .A(n11774), .ZN(n14730) );
  XNOR2_X1 U12498 ( .A(n14730), .B(n11775), .ZN(n11927) );
  NAND2_X1 U12499 ( .A1(n14712), .A2(n9969), .ZN(n9970) );
  AND2_X1 U12500 ( .A1(n14715), .A2(n9986), .ZN(n9971) );
  INV_X1 U12501 ( .A(n13827), .ZN(n9972) );
  XNOR2_X1 U12502 ( .A(n11765), .B(n9972), .ZN(n11925) );
  OR2_X1 U12503 ( .A1(n11765), .A2(n9972), .ZN(n9973) );
  NAND2_X1 U12504 ( .A1(n9974), .A2(n9973), .ZN(n9976) );
  INV_X1 U12505 ( .A(n10020), .ZN(n9975) );
  AOI21_X1 U12506 ( .B1(n11927), .B2(n9976), .A(n9975), .ZN(n9992) );
  NAND2_X1 U12507 ( .A1(n11885), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9982) );
  INV_X1 U12508 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9977) );
  OR2_X1 U12509 ( .A1(n11888), .A2(n9977), .ZN(n9981) );
  XNOR2_X1 U12510 ( .A(n10007), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n10651) );
  OR2_X1 U12511 ( .A1(n11671), .A2(n10651), .ZN(n9980) );
  OR2_X1 U12512 ( .A1(n11656), .A2(n9978), .ZN(n9979) );
  NAND4_X1 U12513 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n14576) );
  AOI22_X1 U12514 ( .A1(n14262), .A2(n13827), .B1(n14576), .B2(n14591), .ZN(
        n9991) );
  NAND2_X1 U12515 ( .A1(n9983), .A2(n7517), .ZN(n9985) );
  OR2_X1 U12516 ( .A1(n14712), .A2(n13829), .ZN(n9984) );
  OR2_X1 U12517 ( .A1(n14715), .A2(n13828), .ZN(n9987) );
  OR2_X1 U12518 ( .A1(n11765), .A2(n13827), .ZN(n9988) );
  XNOR2_X1 U12519 ( .A(n10016), .B(n11927), .ZN(n9989) );
  NAND2_X1 U12520 ( .A1(n9989), .A2(n14725), .ZN(n9990) );
  OAI211_X1 U12521 ( .C1(n9992), .C2(n14704), .A(n9991), .B(n9990), .ZN(n14727) );
  INV_X1 U12522 ( .A(n14727), .ZN(n9998) );
  INV_X1 U12523 ( .A(n10045), .ZN(n9994) );
  NAND2_X1 U12524 ( .A1(n11774), .A2(n10045), .ZN(n10002) );
  INV_X1 U12525 ( .A(n10002), .ZN(n9993) );
  AOI211_X1 U12526 ( .C1(n14730), .C2(n9994), .A(n14719), .B(n9993), .ZN(
        n14728) );
  NOR2_X1 U12527 ( .A1(n11774), .A2(n14180), .ZN(n9996) );
  OAI22_X1 U12528 ( .A1(n14686), .A2(n8464), .B1(n10524), .B2(n14683), .ZN(
        n9995) );
  AOI211_X1 U12529 ( .C1(n14728), .C2(n14606), .A(n9996), .B(n9995), .ZN(n9997) );
  OAI21_X1 U12530 ( .B1(n9998), .B2(n14689), .A(n9997), .ZN(P1_U3284) );
  AOI22_X1 U12531 ( .A1(n10000), .A2(n11528), .B1(n11529), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U12532 ( .A1(n11778), .A2(n10002), .ZN(n10003) );
  NAND3_X1 U12533 ( .A1(n10261), .A2(n14504), .A3(n10003), .ZN(n10015) );
  NAND2_X1 U12534 ( .A1(n6645), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U12535 ( .A1(n10007), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10005) );
  INV_X1 U12536 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U12537 ( .A1(n10005), .A2(n10004), .ZN(n10008) );
  AND2_X1 U12538 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n10006) );
  NAND2_X1 U12539 ( .A1(n10007), .A2(n10006), .ZN(n10251) );
  NAND2_X1 U12540 ( .A1(n10008), .A2(n10251), .ZN(n14587) );
  OR2_X1 U12541 ( .A1(n11704), .A2(n14587), .ZN(n10012) );
  OR2_X1 U12542 ( .A1(n11656), .A2(n8996), .ZN(n10011) );
  OR2_X1 U12543 ( .A1(n11881), .A2(n10009), .ZN(n10010) );
  NAND4_X1 U12544 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n13825) );
  NAND2_X1 U12545 ( .A1(n13825), .A2(n14591), .ZN(n10014) );
  NAND2_X1 U12546 ( .A1(n10015), .A2(n10014), .ZN(n10157) );
  INV_X1 U12547 ( .A(n10157), .ZN(n10029) );
  NAND2_X1 U12548 ( .A1(n10016), .A2(n11927), .ZN(n10018) );
  NAND2_X1 U12549 ( .A1(n11774), .A2(n11775), .ZN(n10017) );
  XNOR2_X1 U12550 ( .A(n10244), .B(n7600), .ZN(n10024) );
  INV_X1 U12551 ( .A(n11775), .ZN(n13826) );
  OR2_X1 U12552 ( .A1(n11774), .A2(n13826), .ZN(n10019) );
  AOI21_X1 U12553 ( .B1(n10021), .B2(n10243), .A(n14704), .ZN(n10022) );
  AOI22_X1 U12554 ( .A1(n10022), .A2(n10258), .B1(n14262), .B2(n13826), .ZN(
        n10023) );
  OAI21_X1 U12555 ( .B1(n14289), .B2(n10024), .A(n10023), .ZN(n10158) );
  NAND2_X1 U12556 ( .A1(n10158), .A2(n14686), .ZN(n10028) );
  NAND2_X1 U12557 ( .A1(n14177), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10025) );
  OAI21_X1 U12558 ( .B1(n14683), .B2(n10651), .A(n10025), .ZN(n10026) );
  AOI21_X1 U12559 ( .B1(n11778), .B2(n14201), .A(n10026), .ZN(n10027) );
  OAI211_X1 U12560 ( .C1(n10029), .C2(n14130), .A(n10028), .B(n10027), .ZN(
        P1_U3283) );
  INV_X1 U12561 ( .A(n10046), .ZN(n10030) );
  AOI211_X1 U12562 ( .C1(n14715), .C2(n10031), .A(n14719), .B(n10030), .ZN(
        n14714) );
  OAI22_X1 U12563 ( .A1(n14180), .A2(n7525), .B1(n10032), .B2(n14683), .ZN(
        n10040) );
  XNOR2_X1 U12564 ( .A(n10033), .B(n11924), .ZN(n10038) );
  AOI22_X1 U12565 ( .A1(n14262), .A2(n13829), .B1(n13827), .B2(n14591), .ZN(
        n10037) );
  XNOR2_X1 U12566 ( .A(n10034), .B(n11924), .ZN(n10035) );
  NAND2_X1 U12567 ( .A1(n10035), .A2(n14725), .ZN(n10036) );
  OAI211_X1 U12568 ( .C1(n10038), .C2(n14704), .A(n10037), .B(n10036), .ZN(
        n14713) );
  MUX2_X1 U12569 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n14713), .S(n14686), .Z(
        n10039) );
  AOI211_X1 U12570 ( .C1(n14606), .C2(n14714), .A(n10040), .B(n10039), .ZN(
        n10041) );
  INV_X1 U12571 ( .A(n10041), .ZN(P1_U3286) );
  XNOR2_X1 U12572 ( .A(n10042), .B(n11925), .ZN(n10044) );
  AOI21_X1 U12573 ( .B1(n10044), .B2(n14592), .A(n10043), .ZN(n14721) );
  AOI21_X1 U12574 ( .B1(n11765), .B2(n10046), .A(n10045), .ZN(n14716) );
  NOR2_X1 U12575 ( .A1(n14130), .A2(n14719), .ZN(n14105) );
  INV_X1 U12576 ( .A(n11765), .ZN(n14718) );
  NOR2_X1 U12577 ( .A1(n14718), .A2(n14180), .ZN(n10050) );
  OAI22_X1 U12578 ( .A1(n14686), .A2(n10048), .B1(n10047), .B2(n14683), .ZN(
        n10049) );
  AOI211_X1 U12579 ( .C1(n14716), .C2(n14105), .A(n10050), .B(n10049), .ZN(
        n10053) );
  XNOR2_X1 U12580 ( .A(n10051), .B(n11925), .ZN(n14724) );
  NAND2_X1 U12581 ( .A1(n14724), .A2(n14605), .ZN(n10052) );
  OAI211_X1 U12582 ( .C1(n14721), .C2(n14177), .A(n10053), .B(n10052), .ZN(
        P1_U3285) );
  INV_X1 U12583 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10061) );
  NAND3_X1 U12584 ( .A1(n10055), .A2(n11400), .A3(n10054), .ZN(n10056) );
  AOI21_X1 U12585 ( .B1(n10057), .B2(n10056), .A(n13435), .ZN(n10059) );
  NOR2_X1 U12586 ( .A1(n10059), .A2(n10058), .ZN(n14920) );
  INV_X1 U12587 ( .A(n14920), .ZN(n10060) );
  AOI21_X1 U12588 ( .B1(n14864), .B2(n10061), .A(n10060), .ZN(n10069) );
  XNOR2_X1 U12589 ( .A(n11400), .B(n10062), .ZN(n14923) );
  OAI211_X1 U12590 ( .C1(n10064), .C2(n14921), .A(n13488), .B(n10063), .ZN(
        n14919) );
  NOR2_X1 U12591 ( .A1(n14919), .A2(n13411), .ZN(n10067) );
  OAI22_X1 U12592 ( .A1(n14921), .A2(n14868), .B1(n13471), .B2(n10065), .ZN(
        n10066) );
  AOI211_X1 U12593 ( .C1(n14923), .C2(n14872), .A(n10067), .B(n10066), .ZN(
        n10068) );
  OAI21_X1 U12594 ( .B1(n10069), .B2(n13512), .A(n10068), .ZN(P2_U3262) );
  INV_X1 U12595 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15451) );
  MUX2_X1 U12596 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n15451), .S(n10178), .Z(
        n10085) );
  NAND2_X1 U12597 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n15068), .ZN(n10081) );
  INV_X1 U12598 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U12599 ( .A1(n10114), .A2(n15228), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15068), .ZN(n15072) );
  NAND2_X1 U12600 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n15033), .ZN(n10078) );
  INV_X1 U12601 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15224) );
  AOI22_X1 U12602 ( .A1(n10105), .A2(n15224), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15033), .ZN(n15037) );
  NAND2_X1 U12603 ( .A1(n14997), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10075) );
  INV_X1 U12604 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10093) );
  MUX2_X1 U12605 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10093), .S(n14997), .Z(
        n15001) );
  NAND2_X1 U12606 ( .A1(n14979), .A2(n10073), .ZN(n10074) );
  NAND2_X1 U12607 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14983), .ZN(n14982) );
  NAND2_X1 U12608 ( .A1(n10074), .A2(n14982), .ZN(n15002) );
  NAND2_X1 U12609 ( .A1(n15016), .A2(n10076), .ZN(n10077) );
  XNOR2_X1 U12610 ( .A(n10076), .B(n10137), .ZN(n15020) );
  NAND2_X1 U12611 ( .A1(n15020), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U12612 ( .A1(n10077), .A2(n15019), .ZN(n15038) );
  NAND2_X1 U12613 ( .A1(n15051), .A2(n10079), .ZN(n10080) );
  INV_X1 U12614 ( .A(n15051), .ZN(n10141) );
  NAND2_X1 U12615 ( .A1(n15055), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n15054) );
  NAND2_X1 U12616 ( .A1(n10080), .A2(n15054), .ZN(n15073) );
  NAND2_X1 U12617 ( .A1(n15088), .A2(n10082), .ZN(n10083) );
  XNOR2_X1 U12618 ( .A(n10082), .B(n10145), .ZN(n15094) );
  AOI21_X1 U12619 ( .B1(n10085), .B2(n10084), .A(n10176), .ZN(n10156) );
  INV_X1 U12620 ( .A(n10086), .ZN(n14974) );
  INV_X1 U12621 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10088) );
  INV_X1 U12622 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10087) );
  MUX2_X1 U12623 ( .A(n10088), .B(n10087), .S(n6648), .Z(n10090) );
  NAND2_X1 U12624 ( .A1(n10090), .A2(n10089), .ZN(n14993) );
  INV_X1 U12625 ( .A(n10090), .ZN(n10091) );
  NAND2_X1 U12626 ( .A1(n10091), .A2(n14979), .ZN(n10092) );
  AND2_X1 U12627 ( .A1(n14993), .A2(n10092), .ZN(n14973) );
  OAI21_X1 U12628 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n14994) );
  MUX2_X1 U12629 ( .A(n10094), .B(n10093), .S(n6648), .Z(n10096) );
  NAND2_X1 U12630 ( .A1(n10096), .A2(n10095), .ZN(n10099) );
  INV_X1 U12631 ( .A(n10096), .ZN(n10097) );
  NAND2_X1 U12632 ( .A1(n10097), .A2(n14997), .ZN(n10098) );
  NAND2_X1 U12633 ( .A1(n10099), .A2(n10098), .ZN(n14992) );
  AOI21_X1 U12634 ( .B1(n14994), .B2(n14993), .A(n14992), .ZN(n15012) );
  INV_X1 U12635 ( .A(n10099), .ZN(n15011) );
  INV_X1 U12636 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10100) );
  MUX2_X1 U12637 ( .A(n15009), .B(n10100), .S(n6648), .Z(n10101) );
  NAND2_X1 U12638 ( .A1(n10101), .A2(n10137), .ZN(n15029) );
  INV_X1 U12639 ( .A(n10101), .ZN(n10102) );
  NAND2_X1 U12640 ( .A1(n10102), .A2(n15016), .ZN(n10103) );
  AND2_X1 U12641 ( .A1(n15029), .A2(n10103), .ZN(n15010) );
  OAI21_X1 U12642 ( .B1(n15012), .B2(n15011), .A(n15010), .ZN(n15030) );
  INV_X1 U12643 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10104) );
  MUX2_X1 U12644 ( .A(n10104), .B(n15224), .S(n6648), .Z(n10106) );
  NAND2_X1 U12645 ( .A1(n10106), .A2(n10105), .ZN(n10109) );
  INV_X1 U12646 ( .A(n10106), .ZN(n10107) );
  NAND2_X1 U12647 ( .A1(n10107), .A2(n15033), .ZN(n10108) );
  NAND2_X1 U12648 ( .A1(n10109), .A2(n10108), .ZN(n15028) );
  AOI21_X1 U12649 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(n15047) );
  INV_X1 U12650 ( .A(n10109), .ZN(n15046) );
  INV_X1 U12651 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10207) );
  INV_X1 U12652 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10110) );
  MUX2_X1 U12653 ( .A(n10207), .B(n10110), .S(n6648), .Z(n10111) );
  NAND2_X1 U12654 ( .A1(n10111), .A2(n10141), .ZN(n15064) );
  INV_X1 U12655 ( .A(n10111), .ZN(n10112) );
  NAND2_X1 U12656 ( .A1(n10112), .A2(n15051), .ZN(n10113) );
  AND2_X1 U12657 ( .A1(n15064), .A2(n10113), .ZN(n15045) );
  OAI21_X1 U12658 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15065) );
  INV_X1 U12659 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U12660 ( .A(n10226), .B(n15228), .S(n6648), .Z(n10115) );
  NAND2_X1 U12661 ( .A1(n10115), .A2(n10114), .ZN(n10118) );
  INV_X1 U12662 ( .A(n10115), .ZN(n10116) );
  NAND2_X1 U12663 ( .A1(n10116), .A2(n15068), .ZN(n10117) );
  NAND2_X1 U12664 ( .A1(n10118), .A2(n10117), .ZN(n15063) );
  AOI21_X1 U12665 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n15083) );
  INV_X1 U12666 ( .A(n10118), .ZN(n15082) );
  INV_X1 U12667 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10486) );
  INV_X1 U12668 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U12669 ( .A(n10486), .B(n10119), .S(n6648), .Z(n10120) );
  NAND2_X1 U12670 ( .A1(n10120), .A2(n10145), .ZN(n10127) );
  INV_X1 U12671 ( .A(n10120), .ZN(n10121) );
  NAND2_X1 U12672 ( .A1(n10121), .A2(n15088), .ZN(n10122) );
  AND2_X1 U12673 ( .A1(n10127), .A2(n10122), .ZN(n15081) );
  OAI21_X1 U12674 ( .B1(n15083), .B2(n15082), .A(n15081), .ZN(n15080) );
  INV_X1 U12675 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10541) );
  MUX2_X1 U12676 ( .A(n10541), .B(n15451), .S(n6648), .Z(n10123) );
  NAND2_X1 U12677 ( .A1(n10123), .A2(n10178), .ZN(n10182) );
  INV_X1 U12678 ( .A(n10123), .ZN(n10124) );
  NAND2_X1 U12679 ( .A1(n10124), .A2(n10173), .ZN(n10125) );
  NAND2_X1 U12680 ( .A1(n10182), .A2(n10125), .ZN(n10126) );
  AOI21_X1 U12681 ( .B1(n15080), .B2(n10127), .A(n10126), .ZN(n10184) );
  AND3_X1 U12682 ( .A1(n15080), .A2(n10127), .A3(n10126), .ZN(n10128) );
  OAI21_X1 U12683 ( .B1(n10184), .B2(n10128), .A(n15084), .ZN(n10155) );
  NAND2_X1 U12684 ( .A1(n6651), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U12685 ( .A1(n10131), .A2(n10130), .ZN(n10133) );
  INV_X1 U12686 ( .A(n10134), .ZN(n10132) );
  NAND2_X1 U12687 ( .A1(n14997), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10136) );
  OR2_X1 U12688 ( .A1(n14997), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U12689 ( .A1(n10136), .A2(n10135), .ZN(n14990) );
  NOR2_X1 U12690 ( .A1(n10137), .A2(n10138), .ZN(n10139) );
  NAND2_X1 U12691 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n15033), .ZN(n10140) );
  OAI21_X1 U12692 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n15033), .A(n10140), .ZN(
        n15026) );
  NOR2_X1 U12693 ( .A1(n10141), .A2(n10142), .ZN(n10143) );
  NAND2_X1 U12694 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15068), .ZN(n10144) );
  OAI21_X1 U12695 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15068), .A(n10144), .ZN(
        n15061) );
  MUX2_X1 U12696 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n10541), .S(n10178), .Z(
        n10148) );
  AOI21_X1 U12697 ( .B1(n10149), .B2(n10148), .A(n10172), .ZN(n10150) );
  NOR2_X1 U12698 ( .A1(n15099), .A2(n10150), .ZN(n10153) );
  INV_X1 U12699 ( .A(n15092), .ZN(n12611) );
  INV_X1 U12700 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14399) );
  OAI21_X1 U12701 ( .B1(n12611), .B2(n14399), .A(n10151), .ZN(n10152) );
  AOI211_X1 U12702 ( .C1(n12613), .C2(n10178), .A(n10153), .B(n10152), .ZN(
        n10154) );
  OAI211_X1 U12703 ( .C1(n10156), .C2(n12616), .A(n10155), .B(n10154), .ZN(
        P3_U3192) );
  NOR2_X1 U12704 ( .A1(n10158), .A2(n10157), .ZN(n10162) );
  INV_X1 U12705 ( .A(n14354), .ZN(n10513) );
  NOR2_X1 U12706 ( .A1(n14733), .A2(n9977), .ZN(n10159) );
  AOI21_X1 U12707 ( .B1(n11778), .B2(n10513), .A(n10159), .ZN(n10160) );
  OAI21_X1 U12708 ( .B1(n10162), .B2(n14731), .A(n10160), .ZN(P1_U3489) );
  AOI22_X1 U12709 ( .A1(n11778), .A2(n10515), .B1(n14739), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n10161) );
  OAI21_X1 U12710 ( .B1(n10162), .B2(n14739), .A(n10161), .ZN(P1_U3538) );
  OAI222_X1 U12711 ( .A1(P1_U3086), .A2(n11908), .B1(n14373), .B2(n11560), 
        .C1(n11561), .C2(n14370), .ZN(P1_U3334) );
  MUX2_X1 U12712 ( .A(n15105), .B(n10164), .S(n10163), .Z(n10166) );
  XNOR2_X1 U12713 ( .A(n10166), .B(n10165), .ZN(n10171) );
  AND2_X1 U12714 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n15070) );
  INV_X1 U12715 ( .A(n12444), .ZN(n10167) );
  INV_X1 U12716 ( .A(n10223), .ZN(n10478) );
  OAI22_X1 U12717 ( .A1(n10167), .A2(n12202), .B1(n10478), .B2(n12174), .ZN(
        n10168) );
  AOI211_X1 U12718 ( .C1(n12199), .C2(n15105), .A(n15070), .B(n10168), .ZN(
        n10170) );
  NAND2_X1 U12719 ( .A1(n12207), .A2(n10224), .ZN(n10169) );
  OAI211_X1 U12720 ( .C1(n10171), .C2(n12214), .A(n10170), .B(n10169), .ZN(
        P3_U3161) );
  INV_X1 U12721 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n10175) );
  INV_X1 U12722 ( .A(n10451), .ZN(n10435) );
  AOI21_X1 U12723 ( .B1(n10175), .B2(n10174), .A(n10436), .ZN(n10192) );
  INV_X1 U12724 ( .A(n10176), .ZN(n10177) );
  NAND2_X1 U12725 ( .A1(n10179), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n10447) );
  OAI21_X1 U12726 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n10179), .A(n10447), 
        .ZN(n10190) );
  INV_X1 U12727 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n10180) );
  NOR2_X1 U12728 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10180), .ZN(n10279) );
  AOI21_X1 U12729 ( .B1(n15092), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n10279), 
        .ZN(n10181) );
  OAI21_X1 U12730 ( .B1(n15089), .B2(n10451), .A(n10181), .ZN(n10189) );
  INV_X1 U12731 ( .A(n10182), .ZN(n10183) );
  NOR2_X1 U12732 ( .A1(n10184), .A2(n10183), .ZN(n10186) );
  MUX2_X1 U12733 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6648), .Z(n10452) );
  XNOR2_X1 U12734 ( .A(n10452), .B(n10451), .ZN(n10185) );
  AOI21_X1 U12735 ( .B1(n10186), .B2(n10185), .A(n10455), .ZN(n10187) );
  INV_X1 U12736 ( .A(n15084), .ZN(n12592) );
  NOR2_X1 U12737 ( .A1(n10187), .A2(n12592), .ZN(n10188) );
  AOI211_X1 U12738 ( .C1(n15095), .C2(n10190), .A(n10189), .B(n10188), .ZN(
        n10191) );
  OAI21_X1 U12739 ( .B1(n10192), .B2(n15099), .A(n10191), .ZN(P3_U3193) );
  NAND2_X1 U12740 ( .A1(n10193), .A2(n12297), .ZN(n10194) );
  NAND2_X1 U12741 ( .A1(n10195), .A2(n15109), .ZN(n12300) );
  NAND2_X1 U12742 ( .A1(n12446), .A2(n10196), .ZN(n12302) );
  NAND2_X1 U12743 ( .A1(n15102), .A2(n15101), .ZN(n10197) );
  XNOR2_X1 U12744 ( .A(n10213), .B(n12310), .ZN(n15194) );
  NAND2_X1 U12745 ( .A1(n10198), .A2(n15184), .ZN(n10199) );
  NAND2_X1 U12746 ( .A1(n12446), .A2(n15109), .ZN(n10203) );
  OAI211_X1 U12747 ( .C1(n10204), .C2(n12310), .A(n10217), .B(n15133), .ZN(
        n10206) );
  AOI22_X1 U12748 ( .A1(n15148), .A2(n12446), .B1(n12445), .B2(n15149), .ZN(
        n10205) );
  OAI211_X1 U12749 ( .C1(n15146), .C2(n15194), .A(n10206), .B(n10205), .ZN(
        n15195) );
  INV_X1 U12750 ( .A(n15195), .ZN(n10208) );
  MUX2_X1 U12751 ( .A(n10208), .B(n10207), .S(n12846), .Z(n10212) );
  NOR2_X1 U12752 ( .A1(n10209), .A2(n15209), .ZN(n15196) );
  AOI22_X1 U12753 ( .A1(n15196), .A2(n15122), .B1(n15157), .B2(n10210), .ZN(
        n10211) );
  OAI211_X1 U12754 ( .C1(n15194), .C2(n12723), .A(n10212), .B(n10211), .ZN(
        P3_U3226) );
  INV_X1 U12755 ( .A(n12310), .ZN(n12249) );
  NAND2_X1 U12756 ( .A1(n10213), .A2(n12249), .ZN(n10214) );
  NAND2_X1 U12757 ( .A1(n10479), .A2(n10223), .ZN(n12313) );
  NAND2_X1 U12758 ( .A1(n12445), .A2(n10478), .ZN(n12314) );
  NAND2_X1 U12759 ( .A1(n12313), .A2(n12314), .ZN(n10475) );
  XNOR2_X1 U12760 ( .A(n10476), .B(n10475), .ZN(n10222) );
  NAND2_X1 U12761 ( .A1(n15105), .A2(n10215), .ZN(n10216) );
  OAI21_X1 U12762 ( .B1(n10218), .B2(n10475), .A(n10480), .ZN(n10219) );
  NAND2_X1 U12763 ( .A1(n10219), .A2(n15133), .ZN(n10221) );
  AOI22_X1 U12764 ( .A1(n15105), .A2(n15148), .B1(n15149), .B2(n12444), .ZN(
        n10220) );
  OAI211_X1 U12765 ( .C1(n15146), .C2(n10222), .A(n10221), .B(n10220), .ZN(
        n15199) );
  INV_X1 U12766 ( .A(n15199), .ZN(n10229) );
  INV_X1 U12767 ( .A(n10222), .ZN(n15201) );
  AND2_X1 U12768 ( .A1(n10223), .A2(n15155), .ZN(n15200) );
  AOI22_X1 U12769 ( .A1(n15122), .A2(n15200), .B1(n15157), .B2(n10224), .ZN(
        n10225) );
  OAI21_X1 U12770 ( .B1(n10226), .B2(n15162), .A(n10225), .ZN(n10227) );
  AOI21_X1 U12771 ( .B1(n15201), .B2(n12704), .A(n10227), .ZN(n10228) );
  OAI21_X1 U12772 ( .B1(n10229), .B2(n12846), .A(n10228), .ZN(P3_U3225) );
  INV_X1 U12773 ( .A(n13148), .ZN(n10353) );
  XNOR2_X1 U12774 ( .A(n13518), .B(n10353), .ZN(n11410) );
  INV_X1 U12775 ( .A(n11410), .ZN(n10235) );
  XNOR2_X1 U12776 ( .A(n10350), .B(n10235), .ZN(n13519) );
  AOI21_X1 U12777 ( .B1(n13518), .B2(n10231), .A(n13030), .ZN(n10232) );
  AND2_X1 U12778 ( .A1(n10232), .A2(n10360), .ZN(n13520) );
  OR2_X1 U12779 ( .A1(n11094), .A2(n11096), .ZN(n10233) );
  OAI211_X1 U12780 ( .C1(n10236), .C2(n10235), .A(n10355), .B(n13499), .ZN(
        n10238) );
  NAND2_X1 U12781 ( .A1(n10238), .A2(n10237), .ZN(n13511) );
  AOI211_X1 U12782 ( .C1(n14938), .C2(n13519), .A(n13520), .B(n13511), .ZN(
        n10242) );
  NOR2_X1 U12783 ( .A1(n14960), .A2(n9387), .ZN(n10239) );
  AOI21_X1 U12784 ( .B1(n13518), .B2(n6902), .A(n10239), .ZN(n10240) );
  OAI21_X1 U12785 ( .B1(n10242), .B2(n14959), .A(n10240), .ZN(P2_U3460) );
  AOI22_X1 U12786 ( .A1(n13518), .A2(n10558), .B1(n14968), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n10241) );
  OAI21_X1 U12787 ( .B1(n10242), .B2(n14968), .A(n10241), .ZN(P2_U3509) );
  NAND2_X1 U12788 ( .A1(n10245), .A2(n11897), .ZN(n10248) );
  AOI22_X1 U12789 ( .A1(n11528), .A2(n10246), .B1(n11529), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n10247) );
  OR2_X1 U12790 ( .A1(n11787), .A2(n13825), .ZN(n10404) );
  NAND2_X1 U12791 ( .A1(n11787), .A2(n13825), .ZN(n10406) );
  NAND2_X1 U12792 ( .A1(n10404), .A2(n10406), .ZN(n11930) );
  INV_X1 U12793 ( .A(n11930), .ZN(n10249) );
  XNOR2_X1 U12794 ( .A(n10405), .B(n10249), .ZN(n10492) );
  INV_X1 U12795 ( .A(n10492), .ZN(n10266) );
  NAND2_X1 U12796 ( .A1(n6645), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10256) );
  OR2_X1 U12797 ( .A1(n11881), .A2(n9000), .ZN(n10255) );
  INV_X1 U12798 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12799 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NAND2_X1 U12800 ( .A1(n10414), .A2(n10252), .ZN(n10870) );
  OR2_X1 U12801 ( .A1(n11671), .A2(n10870), .ZN(n10254) );
  OR2_X1 U12802 ( .A1(n11656), .A2(n8991), .ZN(n10253) );
  INV_X1 U12803 ( .A(n14576), .ZN(n10654) );
  OR2_X1 U12804 ( .A1(n11778), .A2(n10654), .ZN(n10257) );
  XNOR2_X1 U12805 ( .A(n10412), .B(n11930), .ZN(n10259) );
  OAI222_X1 U12806 ( .A1(n14141), .A2(n13773), .B1(n10259), .B2(n14704), .C1(
        n14609), .C2(n10654), .ZN(n10490) );
  NAND2_X1 U12807 ( .A1(n10490), .A2(n14686), .ZN(n10265) );
  INV_X1 U12808 ( .A(n10426), .ZN(n10260) );
  AOI211_X1 U12809 ( .C1(n11787), .C2(n10261), .A(n14719), .B(n10260), .ZN(
        n10491) );
  NOR2_X1 U12810 ( .A1(n14582), .A2(n14180), .ZN(n10263) );
  OAI22_X1 U12811 ( .A1(n14686), .A2(n8996), .B1(n14587), .B2(n14683), .ZN(
        n10262) );
  AOI211_X1 U12812 ( .C1(n10491), .C2(n14606), .A(n10263), .B(n10262), .ZN(
        n10264) );
  OAI211_X1 U12813 ( .C1(n10266), .C2(n14153), .A(n10265), .B(n10264), .ZN(
        P1_U3282) );
  NAND2_X1 U12814 ( .A1(n10267), .A2(n12443), .ZN(n10268) );
  OAI22_X1 U12815 ( .A1(n12236), .A2(SI_11_), .B1(n10435), .B2(n10270), .ZN(
        n10271) );
  AOI21_X1 U12816 ( .B1(n10272), .B2(n12235), .A(n10271), .ZN(n10736) );
  XNOR2_X1 U12817 ( .A(n10736), .B(n10289), .ZN(n10615) );
  XNOR2_X1 U12818 ( .A(n10617), .B(n10615), .ZN(n10618) );
  XNOR2_X1 U12819 ( .A(n10618), .B(n10761), .ZN(n10285) );
  INV_X1 U12820 ( .A(n10736), .ZN(n10756) );
  NOR2_X1 U12821 ( .A1(n10756), .A2(n12174), .ZN(n10283) );
  NAND2_X1 U12822 ( .A1(n6639), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U12823 ( .A1(n10273), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12824 ( .A1(n10297), .A2(n10274), .ZN(n10764) );
  NAND2_X1 U12825 ( .A1(n12024), .A2(n10764), .ZN(n10277) );
  NAND2_X1 U12826 ( .A1(n9240), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n10276) );
  NAND2_X1 U12827 ( .A1(n6638), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n10275) );
  INV_X1 U12828 ( .A(n10279), .ZN(n10281) );
  NAND2_X1 U12829 ( .A1(n12443), .A2(n12199), .ZN(n10280) );
  OAI211_X1 U12830 ( .C1(n10922), .C2(n12202), .A(n10281), .B(n10280), .ZN(
        n10282) );
  AOI211_X1 U12831 ( .C1(n10737), .C2(n12207), .A(n10283), .B(n10282), .ZN(
        n10284) );
  OAI21_X1 U12832 ( .B1(n10285), .B2(n12214), .A(n10284), .ZN(P3_U3176) );
  AOI22_X1 U12833 ( .A1(n12069), .A2(SI_12_), .B1(n10875), .B2(n12460), .ZN(
        n10287) );
  NAND2_X1 U12834 ( .A1(n10288), .A2(n10287), .ZN(n14533) );
  INV_X2 U12835 ( .A(n10289), .ZN(n12155) );
  INV_X1 U12836 ( .A(n10922), .ZN(n12442) );
  NAND2_X1 U12837 ( .A1(n10290), .A2(n12442), .ZN(n10620) );
  OAI21_X1 U12838 ( .B1(n10757), .B2(n10615), .A(n10620), .ZN(n10293) );
  INV_X1 U12839 ( .A(n10290), .ZN(n10291) );
  NAND2_X1 U12840 ( .A1(n10291), .A2(n10922), .ZN(n10619) );
  NAND3_X1 U12841 ( .A1(n10620), .A2(n10757), .A3(n10615), .ZN(n10292) );
  OR2_X1 U12842 ( .A1(n10294), .A2(n11984), .ZN(n10296) );
  AOI22_X1 U12843 ( .A1(n12069), .A2(SI_13_), .B1(n10875), .B2(n12484), .ZN(
        n10295) );
  XNOR2_X1 U12844 ( .A(n12076), .B(n12155), .ZN(n10304) );
  NAND2_X1 U12845 ( .A1(n6639), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U12846 ( .A1(n10297), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U12847 ( .A1(n10299), .A2(n10298), .ZN(n10926) );
  NAND2_X1 U12848 ( .A1(n12024), .A2(n10926), .ZN(n10302) );
  NAND2_X1 U12849 ( .A1(n6638), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U12850 ( .A1(n12222), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n10300) );
  NAND4_X1 U12851 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n12441) );
  NOR2_X1 U12852 ( .A1(n10304), .A2(n12441), .ZN(n10503) );
  INV_X1 U12853 ( .A(n10503), .ZN(n10305) );
  NAND2_X1 U12854 ( .A1(n10304), .A2(n12441), .ZN(n10502) );
  NAND2_X1 U12855 ( .A1(n10305), .A2(n10502), .ZN(n10306) );
  XNOR2_X1 U12856 ( .A(n10504), .B(n10306), .ZN(n10312) );
  NAND2_X1 U12857 ( .A1(n12207), .A2(n10926), .ZN(n10309) );
  INV_X1 U12858 ( .A(n12202), .ZN(n12189) );
  NOR2_X1 U12859 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10307), .ZN(n12457) );
  AOI21_X1 U12860 ( .B1(n11974), .B2(n12189), .A(n12457), .ZN(n10308) );
  OAI211_X1 U12861 ( .C1(n10922), .C2(n12209), .A(n10309), .B(n10308), .ZN(
        n10310) );
  AOI21_X1 U12862 ( .B1(n12076), .B2(n12212), .A(n10310), .ZN(n10311) );
  OAI21_X1 U12863 ( .B1(n10312), .B2(n12214), .A(n10311), .ZN(P3_U3174) );
  INV_X1 U12864 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U12865 ( .A(n10317), .B(n10320), .S(n6641), .Z(n10318) );
  NAND2_X1 U12866 ( .A1(n11576), .A2(n10318), .ZN(n10319) );
  NAND2_X1 U12867 ( .A1(n10546), .A2(n10319), .ZN(n11199) );
  OAI222_X1 U12868 ( .A1(n11464), .A2(n10320), .B1(P2_U3088), .B2(n11315), 
        .C1(n13675), .C2(n11199), .ZN(P2_U3305) );
  NAND2_X1 U12869 ( .A1(n10778), .A2(n11362), .ZN(n10325) );
  OAI22_X1 U12870 ( .A1(n11363), .A2(n10322), .B1(n14833), .B2(n10321), .ZN(
        n10323) );
  INV_X1 U12871 ( .A(n10323), .ZN(n10324) );
  INV_X1 U12872 ( .A(n13618), .ZN(n10716) );
  INV_X1 U12873 ( .A(n10326), .ZN(n10328) );
  NAND2_X1 U12874 ( .A1(n10328), .A2(n10327), .ZN(n10329) );
  XNOR2_X1 U12875 ( .A(n13618), .B(n13067), .ZN(n10331) );
  AND2_X1 U12876 ( .A1(n13145), .A2(n13030), .ZN(n10332) );
  NAND2_X1 U12877 ( .A1(n10331), .A2(n10332), .ZN(n10686) );
  INV_X1 U12878 ( .A(n10331), .ZN(n10334) );
  INV_X1 U12879 ( .A(n10332), .ZN(n10333) );
  NAND2_X1 U12880 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  AND2_X1 U12881 ( .A1(n10686), .A2(n10335), .ZN(n10336) );
  OAI211_X1 U12882 ( .C1(n10337), .C2(n10336), .A(n10687), .B(n13133), .ZN(
        n10349) );
  INV_X1 U12883 ( .A(n10338), .ZN(n10714) );
  NAND2_X1 U12884 ( .A1(n13146), .A2(n13120), .ZN(n10345) );
  NAND2_X1 U12885 ( .A1(n11372), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10343) );
  INV_X1 U12886 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10631) );
  XNOR2_X1 U12887 ( .A(n10633), .B(n10631), .ZN(n14557) );
  OR2_X1 U12888 ( .A1(n6847), .A2(n14557), .ZN(n10342) );
  INV_X1 U12889 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10339) );
  OR2_X1 U12890 ( .A1(n6658), .A2(n10339), .ZN(n10341) );
  INV_X1 U12891 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10644) );
  OR2_X1 U12892 ( .A1(n11317), .A2(n10644), .ZN(n10340) );
  NAND4_X1 U12893 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n13144) );
  NAND2_X1 U12894 ( .A1(n13144), .A2(n13237), .ZN(n10344) );
  NAND2_X1 U12895 ( .A1(n10345), .A2(n10344), .ZN(n10721) );
  INV_X1 U12896 ( .A(n10721), .ZN(n10346) );
  INV_X1 U12897 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14822) );
  OAI22_X1 U12898 ( .A1(n10346), .A2(n14554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14822), .ZN(n10347) );
  AOI21_X1 U12899 ( .B1(n10714), .B2(n13121), .A(n10347), .ZN(n10348) );
  OAI211_X1 U12900 ( .C1(n10716), .C2(n14550), .A(n10349), .B(n10348), .ZN(
        P2_U3206) );
  NAND2_X1 U12901 ( .A1(n13518), .A2(n13148), .ZN(n10351) );
  NAND2_X1 U12902 ( .A1(n10352), .A2(n10351), .ZN(n10380) );
  XNOR2_X1 U12903 ( .A(n11107), .B(n13147), .ZN(n11413) );
  XNOR2_X1 U12904 ( .A(n10380), .B(n11413), .ZN(n10555) );
  INV_X1 U12905 ( .A(n10555), .ZN(n10366) );
  OR2_X1 U12906 ( .A1(n13518), .A2(n10353), .ZN(n10354) );
  AOI21_X1 U12907 ( .B1(n10379), .B2(n10356), .A(n6905), .ZN(n10358) );
  OAI21_X1 U12908 ( .B1(n10358), .B2(n13435), .A(n10357), .ZN(n10553) );
  NAND2_X1 U12909 ( .A1(n10553), .A2(n13471), .ZN(n10365) );
  INV_X1 U12910 ( .A(n10375), .ZN(n10359) );
  AOI211_X1 U12911 ( .C1(n11107), .C2(n10360), .A(n13030), .B(n10359), .ZN(
        n10554) );
  NOR2_X1 U12912 ( .A1(n7105), .A2(n14868), .ZN(n10363) );
  OAI22_X1 U12913 ( .A1(n13471), .A2(n9656), .B1(n10361), .B2(n13515), .ZN(
        n10362) );
  AOI211_X1 U12914 ( .C1(n10554), .C2(n14862), .A(n10363), .B(n10362), .ZN(
        n10364) );
  OAI211_X1 U12915 ( .C1(n10366), .C2(n13507), .A(n10365), .B(n10364), .ZN(
        P2_U3254) );
  NAND2_X1 U12916 ( .A1(n11107), .A2(n11109), .ZN(n10367) );
  INV_X1 U12917 ( .A(n13146), .ZN(n10369) );
  NAND2_X1 U12918 ( .A1(n11116), .A2(n10369), .ZN(n10370) );
  NAND2_X1 U12919 ( .A1(n10717), .A2(n10370), .ZN(n11411) );
  AOI21_X1 U12920 ( .B1(n10371), .B2(n11411), .A(n13435), .ZN(n10373) );
  AOI21_X1 U12921 ( .B1(n10373), .B2(n10720), .A(n10372), .ZN(n10589) );
  OAI22_X1 U12922 ( .A1(n13471), .A2(n9657), .B1(n10374), .B2(n13515), .ZN(
        n10378) );
  AOI21_X1 U12923 ( .B1(n10375), .B2(n11116), .A(n13030), .ZN(n10376) );
  NAND2_X1 U12924 ( .A1(n10376), .A2(n10713), .ZN(n10588) );
  NOR2_X1 U12925 ( .A1(n10588), .A2(n13411), .ZN(n10377) );
  AOI211_X1 U12926 ( .C1(n13517), .C2(n11116), .A(n10378), .B(n10377), .ZN(
        n10384) );
  NAND2_X1 U12927 ( .A1(n10380), .A2(n10379), .ZN(n10382) );
  NAND2_X1 U12928 ( .A1(n11107), .A2(n13147), .ZN(n10381) );
  XOR2_X1 U12929 ( .A(n10641), .B(n11411), .Z(n10592) );
  NAND2_X1 U12930 ( .A1(n10592), .A2(n14872), .ZN(n10383) );
  OAI211_X1 U12931 ( .C1(n10589), .C2(n13512), .A(n10384), .B(n10383), .ZN(
        P2_U3253) );
  INV_X1 U12932 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10812) );
  NOR2_X1 U12933 ( .A1(n11488), .A2(n10812), .ZN(n10389) );
  NAND2_X1 U12934 ( .A1(n10786), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10386) );
  NAND2_X1 U12935 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  NOR2_X1 U12936 ( .A1(n14666), .A2(n10387), .ZN(n10388) );
  XOR2_X1 U12937 ( .A(n10394), .B(n10387), .Z(n14661) );
  NOR2_X1 U12938 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14661), .ZN(n14660) );
  NOR2_X1 U12939 ( .A1(n10388), .A2(n14660), .ZN(n10391) );
  AOI211_X1 U12940 ( .C1(n11488), .C2(n10812), .A(n10389), .B(n10391), .ZN(
        n10392) );
  NAND2_X1 U12941 ( .A1(n10400), .A2(n10812), .ZN(n10390) );
  NAND2_X1 U12942 ( .A1(n11488), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10603) );
  NAND3_X1 U12943 ( .A1(n10391), .A2(n10390), .A3(n10603), .ZN(n10604) );
  INV_X1 U12944 ( .A(n10604), .ZN(n10609) );
  NOR3_X1 U12945 ( .A1(n10392), .A2(n10609), .A3(n13867), .ZN(n10403) );
  OAI21_X1 U12946 ( .B1(n10786), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10393), 
        .ZN(n10395) );
  NAND2_X1 U12947 ( .A1(n10394), .A2(n10395), .ZN(n10396) );
  XNOR2_X1 U12948 ( .A(n14666), .B(n10395), .ZN(n14664) );
  NAND2_X1 U12949 ( .A1(n14664), .A2(n10801), .ZN(n14663) );
  NAND2_X1 U12950 ( .A1(n10396), .A2(n14663), .ZN(n10398) );
  XNOR2_X1 U12951 ( .A(n11488), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U12952 ( .A1(n10398), .A2(n10397), .ZN(n10597) );
  AOI211_X1 U12953 ( .C1(n10398), .C2(n10397), .A(n13886), .B(n10597), .ZN(
        n10402) );
  AND2_X1 U12954 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13740) );
  AOI21_X1 U12955 ( .B1(n14656), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n13740), 
        .ZN(n10399) );
  OAI21_X1 U12956 ( .B1(n13885), .B2(n10400), .A(n10399), .ZN(n10401) );
  OR3_X1 U12957 ( .A1(n10403), .A2(n10402), .A3(n10401), .ZN(P1_U3259) );
  NAND2_X1 U12958 ( .A1(n10407), .A2(n10406), .ZN(n10823) );
  NAND2_X1 U12959 ( .A1(n10408), .A2(n11897), .ZN(n10411) );
  AOI22_X1 U12960 ( .A1(n10409), .A2(n11528), .B1(n11529), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10410) );
  XNOR2_X1 U12961 ( .A(n11792), .B(n14578), .ZN(n11928) );
  INV_X1 U12962 ( .A(n11928), .ZN(n10413) );
  XNOR2_X1 U12963 ( .A(n10823), .B(n10413), .ZN(n10425) );
  INV_X1 U12964 ( .A(n13825), .ZN(n10859) );
  OAI211_X1 U12965 ( .C1(n6783), .C2(n11928), .A(n14592), .B(n10777), .ZN(
        n10424) );
  NAND2_X1 U12966 ( .A1(n6644), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10422) );
  INV_X1 U12967 ( .A(n10789), .ZN(n10416) );
  NAND2_X1 U12968 ( .A1(n10414), .A2(n15476), .ZN(n10415) );
  NAND2_X1 U12969 ( .A1(n10416), .A2(n10415), .ZN(n14514) );
  OR2_X1 U12970 ( .A1(n11704), .A2(n14514), .ZN(n10421) );
  OR2_X1 U12971 ( .A1(n11656), .A2(n10417), .ZN(n10420) );
  OR2_X1 U12972 ( .A1(n11881), .A2(n10418), .ZN(n10419) );
  NAND4_X1 U12973 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n14564) );
  AOI22_X1 U12974 ( .A1(n14262), .A2(n13825), .B1(n14564), .B2(n14591), .ZN(
        n10423) );
  OAI211_X1 U12975 ( .C1(n10425), .C2(n14289), .A(n10424), .B(n10423), .ZN(
        n10512) );
  INV_X1 U12976 ( .A(n10512), .ZN(n10433) );
  NAND2_X1 U12977 ( .A1(n10426), .A2(n11792), .ZN(n10427) );
  NAND2_X1 U12978 ( .A1(n10427), .A2(n14504), .ZN(n10428) );
  NOR2_X1 U12979 ( .A1(n14505), .A2(n10428), .ZN(n10511) );
  NOR2_X1 U12980 ( .A1(n14683), .A2(n10870), .ZN(n10429) );
  AOI21_X1 U12981 ( .B1(n14689), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10429), 
        .ZN(n10430) );
  OAI21_X1 U12982 ( .B1(n11791), .B2(n14180), .A(n10430), .ZN(n10431) );
  AOI21_X1 U12983 ( .B1(n10511), .B2(n14606), .A(n10431), .ZN(n10432) );
  OAI21_X1 U12984 ( .B1(n10433), .B2(n14689), .A(n10432), .ZN(P1_U3281) );
  NOR2_X1 U12985 ( .A1(n10435), .A2(n10434), .ZN(n10437) );
  INV_X1 U12986 ( .A(n10441), .ZN(n10443) );
  INV_X1 U12987 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U12988 ( .A1(n12450), .A2(n10766), .ZN(n10439) );
  NAND2_X1 U12989 ( .A1(n12460), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n10438) );
  AND2_X1 U12990 ( .A1(n10439), .A2(n10438), .ZN(n10440) );
  INV_X1 U12991 ( .A(n10440), .ZN(n10442) );
  OAI21_X1 U12992 ( .B1(n10443), .B2(n10442), .A(n12452), .ZN(n10463) );
  INV_X1 U12993 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U12994 ( .A1(n12460), .A2(n10445), .ZN(n10444) );
  OAI21_X1 U12995 ( .B1(n12460), .B2(n10445), .A(n10444), .ZN(n10450) );
  NAND2_X1 U12996 ( .A1(n10451), .A2(n10446), .ZN(n10448) );
  AOI21_X1 U12997 ( .B1(n10450), .B2(n10449), .A(n12454), .ZN(n10461) );
  NOR2_X1 U12998 ( .A1(n10452), .A2(n10451), .ZN(n10454) );
  MUX2_X1 U12999 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6648), .Z(n12459) );
  XOR2_X1 U13000 ( .A(n12460), .B(n12459), .Z(n10453) );
  INV_X1 U13001 ( .A(n12464), .ZN(n10457) );
  OAI21_X1 U13002 ( .B1(n10455), .B2(n10454), .A(n10453), .ZN(n10456) );
  NAND3_X1 U13003 ( .A1(n10457), .A2(n15084), .A3(n10456), .ZN(n10460) );
  AND2_X1 U13004 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n10612) );
  INV_X1 U13005 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14403) );
  NOR2_X1 U13006 ( .A1(n12611), .A2(n14403), .ZN(n10458) );
  AOI211_X1 U13007 ( .C1(n12613), .C2(n12460), .A(n10612), .B(n10458), .ZN(
        n10459) );
  OAI211_X1 U13008 ( .C1(n10461), .C2(n12616), .A(n10460), .B(n10459), .ZN(
        n10462) );
  AOI21_X1 U13009 ( .B1(n12588), .B2(n10463), .A(n10462), .ZN(n10464) );
  INV_X1 U13010 ( .A(n10464), .ZN(P3_U3194) );
  INV_X1 U13011 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10467) );
  NAND2_X1 U13012 ( .A1(n10467), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10468) );
  INV_X1 U13013 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U13014 ( .A1(n10470), .A2(n11237), .ZN(n10471) );
  INV_X1 U13015 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11614) );
  XNOR2_X1 U13016 ( .A(n10561), .B(n11614), .ZN(n12019) );
  INV_X1 U13017 ( .A(n12019), .ZN(n10473) );
  INV_X1 U13018 ( .A(SI_24_), .ZN(n10472) );
  OAI222_X1 U13019 ( .A1(P3_U3151), .A2(n10474), .B1(n12997), .B2(n10473), 
        .C1(n10472), .C2(n12985), .ZN(P3_U3271) );
  INV_X1 U13020 ( .A(n10475), .ZN(n12309) );
  NAND2_X1 U13021 ( .A1(n10476), .A2(n12309), .ZN(n10477) );
  XNOR2_X1 U13022 ( .A(n12444), .B(n10533), .ZN(n12312) );
  XNOR2_X1 U13023 ( .A(n10531), .B(n12312), .ZN(n15203) );
  NAND2_X1 U13024 ( .A1(n10481), .A2(n12312), .ZN(n10536) );
  OAI211_X1 U13025 ( .C1(n10481), .C2(n12312), .A(n10536), .B(n15133), .ZN(
        n10483) );
  AOI22_X1 U13026 ( .A1(n12445), .A2(n15148), .B1(n15149), .B2(n12443), .ZN(
        n10482) );
  OAI211_X1 U13027 ( .C1(n15146), .C2(n15203), .A(n10483), .B(n10482), .ZN(
        n15204) );
  NAND2_X1 U13028 ( .A1(n15204), .A2(n15162), .ZN(n10489) );
  NOR2_X1 U13029 ( .A1(n10533), .A2(n15209), .ZN(n15205) );
  INV_X1 U13030 ( .A(n10484), .ZN(n10485) );
  OAI22_X1 U13031 ( .A1(n15162), .A2(n10486), .B1(n10485), .B2(n12782), .ZN(
        n10487) );
  AOI21_X1 U13032 ( .B1(n15122), .B2(n15205), .A(n10487), .ZN(n10488) );
  OAI211_X1 U13033 ( .C1(n15203), .C2(n12723), .A(n10489), .B(n10488), .ZN(
        P3_U3224) );
  AOI211_X1 U13034 ( .C1(n14725), .C2(n10492), .A(n10491), .B(n10490), .ZN(
        n10497) );
  AOI22_X1 U13035 ( .A1(n11787), .A2(n10515), .B1(n14739), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n10493) );
  OAI21_X1 U13036 ( .B1(n10497), .B2(n14739), .A(n10493), .ZN(P1_U3539) );
  INV_X1 U13037 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10494) );
  OAI22_X1 U13038 ( .A1(n14582), .A2(n14354), .B1(n14733), .B2(n10494), .ZN(
        n10495) );
  INV_X1 U13039 ( .A(n10495), .ZN(n10496) );
  OAI21_X1 U13040 ( .B1(n10497), .B2(n14731), .A(n10496), .ZN(P1_U3492) );
  NAND2_X1 U13041 ( .A1(n10498), .A2(n12235), .ZN(n10501) );
  AOI22_X1 U13042 ( .A1(n12069), .A2(n10499), .B1(n10875), .B2(n12507), .ZN(
        n10500) );
  XNOR2_X1 U13043 ( .A(n12977), .B(n12155), .ZN(n10569) );
  XNOR2_X1 U13044 ( .A(n10569), .B(n11974), .ZN(n10505) );
  OAI211_X1 U13045 ( .C1(n10506), .C2(n10505), .A(n10568), .B(n12168), .ZN(
        n10510) );
  NAND2_X1 U13046 ( .A1(n12441), .A2(n12199), .ZN(n10507) );
  NAND2_X1 U13047 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12490)
         );
  OAI211_X1 U13048 ( .C1(n12836), .C2(n12202), .A(n10507), .B(n12490), .ZN(
        n10508) );
  AOI21_X1 U13049 ( .B1(n12840), .B2(n12207), .A(n10508), .ZN(n10509) );
  OAI211_X1 U13050 ( .C1(n12174), .C2(n12977), .A(n10510), .B(n10509), .ZN(
        P3_U3155) );
  NOR2_X1 U13051 ( .A1(n10512), .A2(n10511), .ZN(n10517) );
  AOI22_X1 U13052 ( .A1(n11792), .A2(n10513), .B1(n14731), .B2(
        P1_REG0_REG_12__SCAN_IN), .ZN(n10514) );
  OAI21_X1 U13053 ( .B1(n10517), .B2(n14731), .A(n10514), .ZN(P1_U3495) );
  AOI22_X1 U13054 ( .A1(n11792), .A2(n10515), .B1(n14739), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n10516) );
  OAI21_X1 U13055 ( .B1(n10517), .B2(n14739), .A(n10516), .ZN(P1_U3540) );
  OAI22_X1 U13056 ( .A1(n11774), .A2(n6646), .B1(n11775), .B2(n11696), .ZN(
        n10659) );
  OAI22_X1 U13057 ( .A1(n11774), .A2(n7432), .B1(n11775), .B2(n6646), .ZN(
        n10522) );
  XNOR2_X1 U13058 ( .A(n10522), .B(n11678), .ZN(n10660) );
  XNOR2_X1 U13059 ( .A(n10661), .B(n10660), .ZN(n10529) );
  OAI22_X1 U13060 ( .A1(n14588), .A2(n10524), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10523), .ZN(n10525) );
  AOI21_X1 U13061 ( .B1(n14579), .B2(n14576), .A(n10525), .ZN(n10527) );
  NAND2_X1 U13062 ( .A1(n14577), .A2(n13827), .ZN(n10526) );
  OAI211_X1 U13063 ( .C1(n11774), .C2(n14581), .A(n10527), .B(n10526), .ZN(
        n10528) );
  AOI21_X1 U13064 ( .B1(n10529), .B2(n14567), .A(n10528), .ZN(n10530) );
  INV_X1 U13065 ( .A(n10530), .ZN(P1_U3231) );
  NOR2_X1 U13066 ( .A1(n12444), .A2(n10533), .ZN(n12318) );
  NAND2_X1 U13067 ( .A1(n12444), .A2(n10533), .ZN(n12320) );
  XNOR2_X1 U13068 ( .A(n12443), .B(n15210), .ZN(n12321) );
  XNOR2_X1 U13069 ( .A(n10734), .B(n12255), .ZN(n15212) );
  OR2_X1 U13070 ( .A1(n12697), .A2(n15136), .ZN(n10532) );
  NAND2_X1 U13071 ( .A1(n15162), .A2(n10532), .ZN(n12787) );
  INV_X1 U13072 ( .A(n10533), .ZN(n10534) );
  NAND2_X1 U13073 ( .A1(n12444), .A2(n10534), .ZN(n10535) );
  NAND2_X1 U13074 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  OAI211_X1 U13075 ( .C1(n10537), .C2(n12321), .A(n10729), .B(n15133), .ZN(
        n10539) );
  AOI22_X1 U13076 ( .A1(n10761), .A2(n15149), .B1(n15148), .B2(n12444), .ZN(
        n10538) );
  NAND2_X1 U13077 ( .A1(n10539), .A2(n10538), .ZN(n15214) );
  NAND2_X1 U13078 ( .A1(n15214), .A2(n15162), .ZN(n10544) );
  OAI22_X1 U13079 ( .A1(n15162), .A2(n10541), .B1(n10540), .B2(n12782), .ZN(
        n10542) );
  AOI21_X1 U13080 ( .B1(n12792), .B2(n10727), .A(n10542), .ZN(n10543) );
  OAI211_X1 U13081 ( .C1(n15212), .C2(n12787), .A(n10544), .B(n10543), .ZN(
        P3_U3223) );
  MUX2_X1 U13082 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6641), .Z(n10547) );
  NAND2_X1 U13083 ( .A1(n10547), .A2(SI_23_), .ZN(n10746) );
  OAI21_X1 U13084 ( .B1(n10547), .B2(SI_23_), .A(n10746), .ZN(n10743) );
  INV_X1 U13085 ( .A(n11595), .ZN(n10550) );
  NAND2_X1 U13086 ( .A1(n13677), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n10549) );
  OR2_X1 U13087 ( .A1(n10548), .A2(P2_U3088), .ZN(n11460) );
  OAI211_X1 U13088 ( .C1(n10550), .C2(n13675), .A(n10549), .B(n11460), .ZN(
        P2_U3304) );
  INV_X1 U13089 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11596) );
  NAND2_X1 U13090 ( .A1(n11595), .A2(n10551), .ZN(n10552) );
  OAI211_X1 U13091 ( .C1(n11596), .C2(n14370), .A(n10552), .B(n11959), .ZN(
        P1_U3332) );
  AOI211_X1 U13092 ( .C1(n14938), .C2(n10555), .A(n10554), .B(n10553), .ZN(
        n10560) );
  NOR2_X1 U13093 ( .A1(n14960), .A2(n9749), .ZN(n10556) );
  AOI21_X1 U13094 ( .B1(n11107), .B2(n6902), .A(n10556), .ZN(n10557) );
  OAI21_X1 U13095 ( .B1(n10560), .B2(n14959), .A(n10557), .ZN(P2_U3463) );
  AOI22_X1 U13096 ( .A1(n11107), .A2(n10558), .B1(n14968), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n10559) );
  OAI21_X1 U13097 ( .B1(n10560), .B2(n14968), .A(n10559), .ZN(P2_U3510) );
  INV_X1 U13098 ( .A(SI_25_), .ZN(n10989) );
  INV_X1 U13099 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11249) );
  XNOR2_X1 U13100 ( .A(n11249), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n10562) );
  XNOR2_X1 U13101 ( .A(n10582), .B(n10562), .ZN(n12031) );
  INV_X1 U13102 ( .A(n12031), .ZN(n10563) );
  OAI222_X1 U13103 ( .A1(n12985), .A2(n10989), .B1(P3_U3151), .B2(n10564), 
        .C1(n12997), .C2(n10563), .ZN(P3_U3270) );
  AOI22_X1 U13104 ( .A1(n12069), .A2(SI_15_), .B1(n10875), .B2(n12536), .ZN(
        n10566) );
  NAND2_X1 U13105 ( .A1(n10567), .A2(n10566), .ZN(n12077) );
  INV_X1 U13106 ( .A(n12077), .ZN(n12973) );
  INV_X1 U13107 ( .A(n11974), .ZN(n12824) );
  OAI21_X1 U13108 ( .B1(n12824), .B2(n10569), .A(n10568), .ZN(n10571) );
  XNOR2_X1 U13109 ( .A(n12077), .B(n12155), .ZN(n10670) );
  XNOR2_X1 U13110 ( .A(n10670), .B(n12836), .ZN(n10570) );
  NAND2_X1 U13111 ( .A1(n10571), .A2(n10570), .ZN(n10671) );
  OAI211_X1 U13112 ( .C1(n10571), .C2(n10570), .A(n10671), .B(n12168), .ZN(
        n10580) );
  NAND2_X1 U13113 ( .A1(n6639), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13114 ( .A1(n6638), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n10575) );
  XNOR2_X1 U13115 ( .A(n10572), .B(P3_REG3_REG_16__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U13116 ( .A1(n12024), .A2(n12812), .ZN(n10574) );
  NAND2_X1 U13117 ( .A1(n12222), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n10573) );
  NAND2_X1 U13118 ( .A1(n11974), .A2(n12199), .ZN(n10577) );
  NAND2_X1 U13119 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12505)
         );
  OAI211_X1 U13120 ( .C1(n12825), .C2(n12202), .A(n10577), .B(n12505), .ZN(
        n10578) );
  AOI21_X1 U13121 ( .B1(n12828), .B2(n12207), .A(n10578), .ZN(n10579) );
  OAI211_X1 U13122 ( .C1(n12973), .C2(n12174), .A(n10580), .B(n10579), .ZN(
        P3_U3181) );
  NAND2_X1 U13123 ( .A1(n11249), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10581) );
  INV_X1 U13124 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11635) );
  NAND2_X1 U13125 ( .A1(n11635), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10583) );
  INV_X1 U13126 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13682) );
  XNOR2_X1 U13127 ( .A(n13682), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n10585) );
  XNOR2_X1 U13128 ( .A(n10771), .B(n10585), .ZN(n12042) );
  INV_X1 U13129 ( .A(n12042), .ZN(n10587) );
  INV_X1 U13130 ( .A(SI_26_), .ZN(n10996) );
  OAI222_X1 U13131 ( .A1(n12997), .A2(n10587), .B1(n12985), .B2(n10996), .C1(
        P3_U3151), .C2(n10586), .ZN(P3_U3269) );
  INV_X1 U13132 ( .A(n11116), .ZN(n10590) );
  OAI211_X1 U13133 ( .C1(n10590), .C2(n14953), .A(n10589), .B(n10588), .ZN(
        n10591) );
  AOI21_X1 U13134 ( .B1(n10592), .B2(n14938), .A(n10591), .ZN(n10595) );
  NAND2_X1 U13135 ( .A1(n14968), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10593) );
  OAI21_X1 U13136 ( .B1(n10595), .B2(n14968), .A(n10593), .ZN(P2_U3511) );
  NAND2_X1 U13137 ( .A1(n14959), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10594) );
  OAI21_X1 U13138 ( .B1(n10595), .B2(n14959), .A(n10594), .ZN(P2_U3466) );
  INV_X1 U13139 ( .A(n10939), .ZN(n11499) );
  INV_X1 U13140 ( .A(n14656), .ZN(n14673) );
  INV_X1 U13141 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13142 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13749)
         );
  OAI21_X1 U13143 ( .B1(n14673), .B2(n10596), .A(n13749), .ZN(n10601) );
  AOI21_X1 U13144 ( .B1(n11488), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10597), 
        .ZN(n10599) );
  XNOR2_X1 U13145 ( .A(n11499), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10598) );
  NOR2_X1 U13146 ( .A1(n10599), .A2(n10598), .ZN(n10940) );
  AOI211_X1 U13147 ( .C1(n10599), .C2(n10598), .A(n13886), .B(n10940), .ZN(
        n10600) );
  AOI211_X1 U13148 ( .C1(n14665), .C2(n11499), .A(n10601), .B(n10600), .ZN(
        n10611) );
  NAND2_X1 U13149 ( .A1(n10939), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10602) );
  OAI211_X1 U13150 ( .C1(n10939), .C2(P1_REG2_REG_17__SCAN_IN), .A(n10602), 
        .B(n10603), .ZN(n10608) );
  INV_X1 U13151 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13152 ( .A1(n10604), .A2(n10603), .ZN(n10606) );
  NAND2_X1 U13153 ( .A1(n10939), .A2(n10607), .ZN(n10605) );
  OAI211_X1 U13154 ( .C1(n10939), .C2(n10607), .A(n10606), .B(n10605), .ZN(
        n10938) );
  OAI211_X1 U13155 ( .C1(n10609), .C2(n10608), .A(n10938), .B(n14669), .ZN(
        n10610) );
  NAND2_X1 U13156 ( .A1(n10611), .A2(n10610), .ZN(P1_U3260) );
  NAND2_X1 U13157 ( .A1(n12207), .A2(n10764), .ZN(n10614) );
  AOI21_X1 U13158 ( .B1(n12441), .B2(n12189), .A(n10612), .ZN(n10613) );
  OAI211_X1 U13159 ( .C1(n10757), .C2(n12209), .A(n10614), .B(n10613), .ZN(
        n10625) );
  INV_X1 U13160 ( .A(n10615), .ZN(n10616) );
  AOI22_X1 U13161 ( .A1(n10618), .A2(n10761), .B1(n10617), .B2(n10616), .ZN(
        n10622) );
  NAND2_X1 U13162 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  XNOR2_X1 U13163 ( .A(n10622), .B(n10621), .ZN(n10623) );
  NOR2_X1 U13164 ( .A1(n10623), .A2(n12214), .ZN(n10624) );
  AOI211_X1 U13165 ( .C1(n12212), .C2(n14533), .A(n10625), .B(n10624), .ZN(
        n10626) );
  INV_X1 U13166 ( .A(n10626), .ZN(P3_U3164) );
  XNOR2_X1 U13167 ( .A(n13618), .B(n13145), .ZN(n11412) );
  INV_X1 U13168 ( .A(n13145), .ZN(n10627) );
  OR2_X1 U13169 ( .A1(n13618), .A2(n10627), .ZN(n10628) );
  NAND2_X1 U13170 ( .A1(n10785), .A2(n11362), .ZN(n10630) );
  AOI22_X1 U13171 ( .A1(n11169), .A2(n13171), .B1(n11358), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n10629) );
  OR2_X1 U13172 ( .A1(n11125), .A2(n13144), .ZN(n10829) );
  NAND2_X1 U13173 ( .A1(n11125), .A2(n13144), .ZN(n10831) );
  NAND2_X1 U13174 ( .A1(n10829), .A2(n10831), .ZN(n11415) );
  XNOR2_X1 U13175 ( .A(n10834), .B(n11415), .ZN(n10639) );
  NAND2_X1 U13176 ( .A1(n11372), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10638) );
  INV_X1 U13177 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13614) );
  OR2_X1 U13178 ( .A1(n6658), .A2(n13614), .ZN(n10637) );
  INV_X1 U13179 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10841) );
  OR2_X1 U13180 ( .A1(n11317), .A2(n10841), .ZN(n10636) );
  INV_X1 U13181 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13166) );
  OAI21_X1 U13182 ( .B1(n10633), .B2(n10631), .A(n13166), .ZN(n10634) );
  NAND2_X1 U13183 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n10632) );
  NAND2_X1 U13184 ( .A1(n10634), .A2(n10696), .ZN(n10840) );
  OR2_X1 U13185 ( .A1(n6847), .A2(n10840), .ZN(n10635) );
  NAND4_X1 U13186 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n13143) );
  AOI22_X1 U13187 ( .A1(n13237), .A2(n13143), .B1(n13145), .B2(n13120), .ZN(
        n14553) );
  OAI21_X1 U13188 ( .B1(n10639), .B2(n13435), .A(n14553), .ZN(n10847) );
  INV_X1 U13189 ( .A(n10847), .ZN(n10649) );
  AND2_X1 U13190 ( .A1(n11116), .A2(n13146), .ZN(n10640) );
  NOR2_X1 U13191 ( .A1(n13618), .A2(n13145), .ZN(n10642) );
  NAND2_X1 U13192 ( .A1(n13618), .A2(n13145), .ZN(n10643) );
  XNOR2_X1 U13193 ( .A(n10830), .B(n11415), .ZN(n10849) );
  INV_X1 U13194 ( .A(n11125), .ZN(n14549) );
  NAND2_X1 U13195 ( .A1(n14549), .A2(n10712), .ZN(n10839) );
  OAI211_X1 U13196 ( .C1(n14549), .C2(n10712), .A(n13488), .B(n10839), .ZN(
        n10846) );
  OAI22_X1 U13197 ( .A1(n13471), .A2(n10644), .B1(n14557), .B2(n13515), .ZN(
        n10645) );
  AOI21_X1 U13198 ( .B1(n11125), .B2(n13517), .A(n10645), .ZN(n10646) );
  OAI21_X1 U13199 ( .B1(n10846), .B2(n13411), .A(n10646), .ZN(n10647) );
  AOI21_X1 U13200 ( .B1(n10849), .B2(n14872), .A(n10647), .ZN(n10648) );
  OAI21_X1 U13201 ( .B1(n10649), .B2(n13512), .A(n10648), .ZN(P2_U3251) );
  OAI21_X1 U13202 ( .B1(n14588), .B2(n10651), .A(n10650), .ZN(n10652) );
  AOI21_X1 U13203 ( .B1(n14577), .B2(n13826), .A(n10652), .ZN(n10653) );
  OAI21_X1 U13204 ( .B1(n10859), .B2(n13806), .A(n10653), .ZN(n10665) );
  NOR2_X1 U13205 ( .A1(n10654), .A2(n11696), .ZN(n10655) );
  AOI21_X1 U13206 ( .B1(n11778), .B2(n10521), .A(n10655), .ZN(n10854) );
  NAND2_X1 U13207 ( .A1(n11778), .A2(n11699), .ZN(n10657) );
  NAND2_X1 U13208 ( .A1(n14576), .A2(n11698), .ZN(n10656) );
  NAND2_X1 U13209 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  XNOR2_X1 U13210 ( .A(n10658), .B(n11678), .ZN(n10853) );
  XOR2_X1 U13211 ( .A(n10854), .B(n10853), .Z(n10663) );
  AOI211_X1 U13212 ( .C1(n10663), .C2(n10662), .A(n14574), .B(n10861), .ZN(
        n10664) );
  AOI211_X1 U13213 ( .C1(n13798), .C2(n11778), .A(n10665), .B(n10664), .ZN(
        n10666) );
  INV_X1 U13214 ( .A(n10666), .ZN(P1_U3217) );
  AOI22_X1 U13215 ( .A1(n12069), .A2(SI_16_), .B1(n10875), .B2(n12541), .ZN(
        n10668) );
  INV_X1 U13216 ( .A(n12906), .ZN(n12814) );
  INV_X1 U13217 ( .A(n10670), .ZN(n10672) );
  XNOR2_X1 U13218 ( .A(n12906), .B(n12155), .ZN(n10878) );
  XNOR2_X1 U13219 ( .A(n10878), .B(n12825), .ZN(n10673) );
  OAI211_X1 U13220 ( .C1(n10674), .C2(n10673), .A(n10879), .B(n12168), .ZN(
        n10685) );
  NAND2_X1 U13221 ( .A1(n6639), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U13222 ( .A1(n12222), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n10680) );
  INV_X1 U13223 ( .A(n10675), .ZN(n10676) );
  NAND2_X1 U13224 ( .A1(n10676), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13225 ( .A1(n10882), .A2(n10677), .ZN(n12800) );
  NAND2_X1 U13226 ( .A1(n12024), .A2(n12800), .ZN(n10679) );
  NAND2_X1 U13227 ( .A1(n6638), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13228 ( .A1(n12806), .A2(n12199), .ZN(n10682) );
  NAND2_X1 U13229 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12532)
         );
  OAI211_X1 U13230 ( .C1(n12779), .C2(n12202), .A(n10682), .B(n12532), .ZN(
        n10683) );
  AOI21_X1 U13231 ( .B1(n12812), .B2(n12207), .A(n10683), .ZN(n10684) );
  OAI211_X1 U13232 ( .C1(n12814), .C2(n12174), .A(n10685), .B(n10684), .ZN(
        P3_U3166) );
  XNOR2_X1 U13233 ( .A(n11125), .B(n13001), .ZN(n10690) );
  NAND2_X1 U13234 ( .A1(n13144), .A2(n13030), .ZN(n10689) );
  XNOR2_X1 U13235 ( .A(n10690), .B(n10689), .ZN(n14548) );
  NAND2_X1 U13236 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NAND2_X1 U13237 ( .A1(n10797), .A2(n11362), .ZN(n10693) );
  AOI22_X1 U13238 ( .A1(n11358), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n11169), 
        .B2(n13185), .ZN(n10692) );
  XNOR2_X1 U13239 ( .A(n11133), .B(n13035), .ZN(n10950) );
  INV_X1 U13240 ( .A(n10954), .ZN(n10710) );
  AOI22_X1 U13241 ( .A1(n10694), .A2(n13133), .B1(n13111), .B2(n13143), .ZN(
        n10709) );
  INV_X1 U13242 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13192) );
  NAND2_X1 U13243 ( .A1(n10696), .A2(n13192), .ZN(n10697) );
  NAND2_X1 U13244 ( .A1(n11159), .A2(n10697), .ZN(n10957) );
  OR2_X1 U13245 ( .A1(n6847), .A2(n10957), .ZN(n10703) );
  INV_X1 U13246 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13188) );
  OR2_X1 U13247 ( .A1(n11317), .A2(n13188), .ZN(n10702) );
  INV_X1 U13248 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10698) );
  OR2_X1 U13249 ( .A1(n6658), .A2(n10698), .ZN(n10701) );
  INV_X1 U13250 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10699) );
  OR2_X1 U13251 ( .A1(n11318), .A2(n10699), .ZN(n10700) );
  NAND4_X1 U13252 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n13248) );
  NAND2_X1 U13253 ( .A1(n13248), .A2(n13237), .ZN(n10705) );
  NAND2_X1 U13254 ( .A1(n13144), .A2(n13120), .ZN(n10704) );
  NAND2_X1 U13255 ( .A1(n10705), .A2(n10704), .ZN(n13610) );
  AOI22_X1 U13256 ( .A1(n13137), .A2(n13610), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10706) );
  OAI21_X1 U13257 ( .B1(n10840), .B2(n14558), .A(n10706), .ZN(n10707) );
  AOI21_X1 U13258 ( .B1(n11133), .B2(n13128), .A(n10707), .ZN(n10708) );
  OAI21_X1 U13259 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(P2_U3213) );
  XNOR2_X1 U13260 ( .A(n10711), .B(n11412), .ZN(n13621) );
  AOI211_X1 U13261 ( .C1(n13618), .C2(n10713), .A(n13066), .B(n10712), .ZN(
        n13617) );
  AOI22_X1 U13262 ( .A1(n13512), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10714), 
        .B2(n14864), .ZN(n10715) );
  OAI21_X1 U13263 ( .B1(n10716), .B2(n14868), .A(n10715), .ZN(n10725) );
  INV_X1 U13264 ( .A(n10717), .ZN(n10718) );
  NOR2_X1 U13265 ( .A1(n11412), .A2(n10718), .ZN(n10719) );
  AOI21_X1 U13266 ( .B1(n10720), .B2(n10719), .A(n13435), .ZN(n10722) );
  AOI21_X1 U13267 ( .B1(n10723), .B2(n10722), .A(n10721), .ZN(n13620) );
  NOR2_X1 U13268 ( .A1(n13620), .A2(n13512), .ZN(n10724) );
  AOI211_X1 U13269 ( .C1(n13617), .C2(n14862), .A(n10725), .B(n10724), .ZN(
        n10726) );
  OAI21_X1 U13270 ( .B1(n13507), .B2(n13621), .A(n10726), .ZN(P2_U3252) );
  NAND2_X1 U13271 ( .A1(n10757), .A2(n10736), .ZN(n12328) );
  NAND2_X1 U13272 ( .A1(n10761), .A2(n10756), .ZN(n12332) );
  NAND2_X1 U13273 ( .A1(n12443), .A2(n10727), .ZN(n10728) );
  INV_X1 U13274 ( .A(n10759), .ZN(n10731) );
  AOI21_X1 U13275 ( .B1(n12254), .B2(n10732), .A(n10731), .ZN(n10733) );
  OAI222_X1 U13276 ( .A1(n15130), .A2(n12324), .B1(n15128), .B2(n10922), .C1(
        n15154), .C2(n10733), .ZN(n14534) );
  INV_X1 U13277 ( .A(n14534), .ZN(n10742) );
  NAND2_X1 U13278 ( .A1(n12443), .A2(n15210), .ZN(n10735) );
  OAI21_X1 U13279 ( .B1(n6782), .B2(n12254), .A(n10755), .ZN(n14536) );
  AND2_X1 U13280 ( .A1(n10736), .A2(n15155), .ZN(n14535) );
  INV_X1 U13281 ( .A(n14535), .ZN(n10739) );
  AOI22_X1 U13282 ( .A1(n12846), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15157), 
        .B2(n10737), .ZN(n10738) );
  OAI21_X1 U13283 ( .B1(n10739), .B2(n10928), .A(n10738), .ZN(n10740) );
  AOI21_X1 U13284 ( .B1(n14536), .B2(n12844), .A(n10740), .ZN(n10741) );
  OAI21_X1 U13285 ( .B1(n10742), .B2(n12846), .A(n10741), .ZN(P3_U3222) );
  INV_X1 U13286 ( .A(n10743), .ZN(n10744) );
  MUX2_X1 U13287 ( .A(n11614), .B(n11237), .S(n6641), .Z(n10750) );
  NAND2_X1 U13288 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  OAI222_X1 U13289 ( .A1(n10753), .A2(P2_U3088), .B1(n13675), .B2(n11613), 
        .C1(n11237), .C2(n11464), .ZN(P2_U3303) );
  OAI222_X1 U13290 ( .A1(P1_U3086), .A2(n10754), .B1(n14373), .B2(n11613), 
        .C1(n11614), .C2(n14370), .ZN(P1_U3331) );
  OR2_X1 U13291 ( .A1(n14533), .A2(n10922), .ZN(n12331) );
  NAND2_X1 U13292 ( .A1(n14533), .A2(n10922), .ZN(n12335) );
  NAND2_X1 U13293 ( .A1(n12331), .A2(n12335), .ZN(n10923) );
  XNOR2_X1 U13294 ( .A(n10924), .B(n10923), .ZN(n14530) );
  NAND2_X1 U13295 ( .A1(n10757), .A2(n10756), .ZN(n10758) );
  NAND2_X1 U13296 ( .A1(n10760), .A2(n10923), .ZN(n10920) );
  OAI211_X1 U13297 ( .C1(n10760), .C2(n10923), .A(n10920), .B(n15133), .ZN(
        n10763) );
  AOI22_X1 U13298 ( .A1(n10761), .A2(n15148), .B1(n15149), .B2(n12441), .ZN(
        n10762) );
  NAND2_X1 U13299 ( .A1(n10763), .A2(n10762), .ZN(n14531) );
  NAND2_X1 U13300 ( .A1(n14531), .A2(n15162), .ZN(n10769) );
  INV_X1 U13301 ( .A(n10764), .ZN(n10765) );
  OAI22_X1 U13302 ( .A1(n15162), .A2(n10766), .B1(n10765), .B2(n12782), .ZN(
        n10767) );
  AOI21_X1 U13303 ( .B1(n14533), .B2(n12792), .A(n10767), .ZN(n10768) );
  OAI211_X1 U13304 ( .C1(n12787), .C2(n14530), .A(n10769), .B(n10768), .ZN(
        P3_U3221) );
  INV_X1 U13305 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14371) );
  AND2_X1 U13306 ( .A1(n14371), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U13307 ( .A1(n13682), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n10772) );
  XNOR2_X1 U13308 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n10773) );
  XNOR2_X1 U13309 ( .A(n11963), .B(n10773), .ZN(n12053) );
  INV_X1 U13310 ( .A(n12053), .ZN(n10774) );
  INV_X1 U13311 ( .A(SI_27_), .ZN(n11003) );
  OAI222_X1 U13312 ( .A1(P3_U3151), .A2(n6648), .B1(n12997), .B2(n10774), .C1(
        n11003), .C2(n12985), .ZN(P3_U3268) );
  OR2_X1 U13313 ( .A1(n10791), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10775) );
  NAND2_X1 U13314 ( .A1(n10808), .A2(n10775), .ZN(n13814) );
  INV_X1 U13315 ( .A(n13814), .ZN(n10820) );
  NAND2_X1 U13316 ( .A1(n11791), .A2(n14578), .ZN(n10776) );
  NAND2_X1 U13317 ( .A1(n10777), .A2(n10776), .ZN(n14508) );
  NAND2_X1 U13318 ( .A1(n10778), .A2(n11897), .ZN(n10783) );
  NOR2_X1 U13319 ( .A1(n8839), .A2(n10779), .ZN(n10780) );
  AOI21_X1 U13320 ( .B1(n10781), .B2(n11528), .A(n10780), .ZN(n10782) );
  XNOR2_X1 U13321 ( .A(n11798), .B(n14610), .ZN(n14502) );
  INV_X1 U13322 ( .A(n14502), .ZN(n14507) );
  NAND2_X1 U13323 ( .A1(n14508), .A2(n14507), .ZN(n14506) );
  OR2_X1 U13324 ( .A1(n11798), .A2(n14610), .ZN(n10784) );
  NAND2_X1 U13325 ( .A1(n10785), .A2(n11897), .ZN(n10788) );
  AOI22_X1 U13326 ( .A1(n10786), .A2(n11528), .B1(n11529), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13327 ( .A1(n6644), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10796) );
  NOR2_X1 U13328 ( .A1(n10789), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10790) );
  OR2_X1 U13329 ( .A1(n10791), .A2(n10790), .ZN(n14595) );
  OR2_X1 U13330 ( .A1(n11704), .A2(n14595), .ZN(n10795) );
  OR2_X1 U13331 ( .A1(n11656), .A2(n14596), .ZN(n10794) );
  OR2_X1 U13332 ( .A1(n11881), .A2(n10792), .ZN(n10793) );
  NAND2_X1 U13333 ( .A1(n14602), .A2(n13772), .ZN(n11801) );
  OR2_X1 U13334 ( .A1(n14602), .A2(n13772), .ZN(n11804) );
  NAND2_X1 U13335 ( .A1(n10797), .A2(n11897), .ZN(n10799) );
  AOI22_X1 U13336 ( .A1(n14666), .A2(n11528), .B1(n11529), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U13337 ( .A1(n6644), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n10805) );
  OR2_X1 U13338 ( .A1(n13814), .A2(n11671), .ZN(n10804) );
  INV_X1 U13339 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10800) );
  OR2_X1 U13340 ( .A1(n11656), .A2(n10800), .ZN(n10803) );
  INV_X1 U13341 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10801) );
  OR2_X1 U13342 ( .A1(n11881), .A2(n10801), .ZN(n10802) );
  NAND2_X1 U13343 ( .A1(n13910), .A2(n10806), .ZN(n11809) );
  XNOR2_X1 U13344 ( .A(n13935), .B(n13934), .ZN(n10819) );
  INV_X1 U13345 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U13346 ( .A1(n10808), .A2(n10807), .ZN(n10809) );
  AND2_X1 U13347 ( .A1(n11503), .A2(n10809), .ZN(n14176) );
  INV_X1 U13348 ( .A(n11704), .ZN(n10810) );
  NAND2_X1 U13349 ( .A1(n14176), .A2(n10810), .ZN(n10816) );
  NAND2_X1 U13350 ( .A1(n11885), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10815) );
  INV_X1 U13351 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10811) );
  OR2_X1 U13352 ( .A1(n11888), .A2(n10811), .ZN(n10814) );
  OR2_X1 U13353 ( .A1(n11656), .A2(n10812), .ZN(n10813) );
  OR2_X1 U13354 ( .A1(n13912), .A2(n14141), .ZN(n10817) );
  OAI21_X1 U13355 ( .B1(n13772), .B2(n14609), .A(n10817), .ZN(n13817) );
  INV_X1 U13356 ( .A(n13817), .ZN(n10818) );
  OAI21_X1 U13357 ( .B1(n10819), .B2(n14704), .A(n10818), .ZN(n14305) );
  AOI21_X1 U13358 ( .B1(n10820), .B2(n14199), .A(n14305), .ZN(n10828) );
  INV_X1 U13359 ( .A(n14172), .ZN(n10821) );
  AOI211_X1 U13360 ( .C1(n13910), .C2(n14600), .A(n14719), .B(n10821), .ZN(
        n14306) );
  OAI22_X1 U13361 ( .A1(n14355), .A2(n14180), .B1(n10800), .B2(n14686), .ZN(
        n10822) );
  AOI21_X1 U13362 ( .B1(n14306), .B2(n14606), .A(n10822), .ZN(n10827) );
  NAND2_X1 U13363 ( .A1(n11791), .A2(n13773), .ZN(n10824) );
  INV_X1 U13364 ( .A(n13772), .ZN(n13824) );
  NAND2_X1 U13365 ( .A1(n14602), .A2(n13824), .ZN(n10825) );
  XNOR2_X1 U13366 ( .A(n13909), .B(n13934), .ZN(n14307) );
  NAND2_X1 U13367 ( .A1(n14307), .A2(n14605), .ZN(n10826) );
  OAI211_X1 U13368 ( .C1(n10828), .C2(n14177), .A(n10827), .B(n10826), .ZN(
        P1_U3278) );
  XNOR2_X1 U13369 ( .A(n11133), .B(n13143), .ZN(n11418) );
  NAND2_X1 U13370 ( .A1(n10830), .A2(n10829), .ZN(n10832) );
  NAND2_X1 U13371 ( .A1(n10832), .A2(n10831), .ZN(n10893) );
  XOR2_X1 U13372 ( .A(n10893), .B(n11418), .Z(n13609) );
  INV_X1 U13373 ( .A(n13144), .ZN(n11127) );
  NAND2_X1 U13374 ( .A1(n11125), .A2(n11127), .ZN(n10833) );
  OR2_X1 U13375 ( .A1(n11125), .A2(n11127), .ZN(n10835) );
  XNOR2_X1 U13376 ( .A(n10901), .B(n11418), .ZN(n10837) );
  NOR2_X1 U13377 ( .A1(n10837), .A2(n13435), .ZN(n13612) );
  OAI21_X1 U13378 ( .B1(n13612), .B2(n13610), .A(n13471), .ZN(n10845) );
  OR2_X2 U13379 ( .A1(n10839), .A2(n11133), .ZN(n10913) );
  INV_X1 U13380 ( .A(n10913), .ZN(n10838) );
  AOI211_X1 U13381 ( .C1(n11133), .C2(n10839), .A(n13066), .B(n10838), .ZN(
        n13611) );
  INV_X1 U13382 ( .A(n11133), .ZN(n13663) );
  NOR2_X1 U13383 ( .A1(n13663), .A2(n14868), .ZN(n10843) );
  OAI22_X1 U13384 ( .A1(n13471), .A2(n10841), .B1(n10840), .B2(n13515), .ZN(
        n10842) );
  AOI211_X1 U13385 ( .C1(n13611), .C2(n14862), .A(n10843), .B(n10842), .ZN(
        n10844) );
  OAI211_X1 U13386 ( .C1(n13609), .C2(n13507), .A(n10845), .B(n10844), .ZN(
        P2_U3250) );
  OAI21_X1 U13387 ( .B1(n14549), .B2(n14953), .A(n10846), .ZN(n10848) );
  AOI211_X1 U13388 ( .C1(n14938), .C2(n10849), .A(n10848), .B(n10847), .ZN(
        n10852) );
  NAND2_X1 U13389 ( .A1(n14968), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10850) );
  OAI21_X1 U13390 ( .B1(n10852), .B2(n14968), .A(n10850), .ZN(P2_U3513) );
  NAND2_X1 U13391 ( .A1(n14959), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10851) );
  OAI21_X1 U13392 ( .B1(n10852), .B2(n14959), .A(n10851), .ZN(P2_U3472) );
  INV_X1 U13393 ( .A(n10853), .ZN(n10855) );
  NOR2_X1 U13394 ( .A1(n10855), .A2(n10854), .ZN(n14573) );
  NAND2_X1 U13395 ( .A1(n11787), .A2(n11699), .ZN(n10857) );
  NAND2_X1 U13396 ( .A1(n13825), .A2(n11698), .ZN(n10856) );
  NAND2_X1 U13397 ( .A1(n10857), .A2(n10856), .ZN(n10858) );
  XNOR2_X1 U13398 ( .A(n10858), .B(n9192), .ZN(n10863) );
  NOR2_X1 U13399 ( .A1(n10859), .A2(n11696), .ZN(n10860) );
  AOI21_X1 U13400 ( .B1(n11787), .B2(n11698), .A(n10860), .ZN(n10862) );
  XNOR2_X1 U13401 ( .A(n10863), .B(n10862), .ZN(n14572) );
  AND2_X1 U13402 ( .A1(n10863), .A2(n10862), .ZN(n10864) );
  OAI22_X1 U13403 ( .A1(n11791), .A2(n6646), .B1(n13773), .B2(n11696), .ZN(
        n11469) );
  OAI22_X1 U13404 ( .A1(n11791), .A2(n7432), .B1(n13773), .B2(n6646), .ZN(
        n10865) );
  XNOR2_X1 U13405 ( .A(n10865), .B(n11678), .ZN(n11470) );
  XOR2_X1 U13406 ( .A(n11469), .B(n11470), .Z(n10866) );
  OAI211_X1 U13407 ( .C1(n10867), .C2(n10866), .A(n11472), .B(n14567), .ZN(
        n10873) );
  NAND2_X1 U13408 ( .A1(n14577), .A2(n13825), .ZN(n10869) );
  OAI211_X1 U13409 ( .C1(n14588), .C2(n10870), .A(n10869), .B(n10868), .ZN(
        n10871) );
  AOI21_X1 U13410 ( .B1(n14579), .B2(n14564), .A(n10871), .ZN(n10872) );
  OAI211_X1 U13411 ( .C1(n11791), .C2(n14581), .A(n10873), .B(n10872), .ZN(
        P1_U3224) );
  NAND2_X1 U13412 ( .A1(n10874), .A2(n12235), .ZN(n10877) );
  AOI22_X1 U13413 ( .A1(n12069), .A2(SI_17_), .B1(n10875), .B2(n12577), .ZN(
        n10876) );
  INV_X1 U13414 ( .A(n12902), .ZN(n12802) );
  XNOR2_X1 U13415 ( .A(n12902), .B(n12155), .ZN(n10966) );
  XNOR2_X1 U13416 ( .A(n10966), .B(n12779), .ZN(n10880) );
  OAI211_X1 U13417 ( .C1(n10881), .C2(n10880), .A(n10967), .B(n12168), .ZN(
        n10892) );
  NAND2_X1 U13418 ( .A1(n10882), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U13419 ( .A1(n10972), .A2(n10883), .ZN(n12781) );
  NAND2_X1 U13420 ( .A1(n12781), .A2(n12024), .ZN(n10888) );
  NAND2_X1 U13421 ( .A1(n6638), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U13422 ( .A1(n6639), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U13423 ( .A1(n12222), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13424 ( .A1(n6815), .A2(n12199), .ZN(n10889) );
  NAND2_X1 U13425 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12555)
         );
  OAI211_X1 U13426 ( .C1(n12091), .C2(n12202), .A(n10889), .B(n12555), .ZN(
        n10890) );
  AOI21_X1 U13427 ( .B1(n12800), .B2(n12207), .A(n10890), .ZN(n10891) );
  OAI211_X1 U13428 ( .C1(n12802), .C2(n12174), .A(n10892), .B(n10891), .ZN(
        P3_U3168) );
  OR2_X1 U13429 ( .A1(n11133), .A2(n13143), .ZN(n10894) );
  NAND2_X1 U13430 ( .A1(n11487), .A2(n11362), .ZN(n10897) );
  AOI22_X1 U13431 ( .A1(n11358), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n13207), 
        .B2(n11169), .ZN(n10896) );
  INV_X1 U13432 ( .A(n13248), .ZN(n13283) );
  XNOR2_X1 U13433 ( .A(n13603), .B(n13283), .ZN(n11416) );
  NAND2_X1 U13434 ( .A1(n10898), .A2(n10904), .ZN(n10899) );
  NAND2_X1 U13435 ( .A1(n13250), .A2(n10899), .ZN(n13606) );
  INV_X1 U13436 ( .A(n13143), .ZN(n10902) );
  NOR2_X1 U13437 ( .A1(n11133), .A2(n10902), .ZN(n10900) );
  NAND2_X1 U13438 ( .A1(n11133), .A2(n10902), .ZN(n10903) );
  XNOR2_X1 U13439 ( .A(n13281), .B(n10904), .ZN(n10905) );
  NAND2_X1 U13440 ( .A1(n10905), .A2(n13499), .ZN(n10912) );
  XNOR2_X1 U13441 ( .A(n11159), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U13442 ( .A1(n13503), .A2(n11370), .ZN(n10909) );
  INV_X1 U13443 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13198) );
  OR2_X1 U13444 ( .A1(n11317), .A2(n13198), .ZN(n10908) );
  NAND2_X1 U13445 ( .A1(n11277), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U13446 ( .A1(n11372), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n10906) );
  NAND4_X1 U13447 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n13286) );
  NAND2_X1 U13448 ( .A1(n13286), .A2(n13237), .ZN(n10911) );
  NAND2_X1 U13449 ( .A1(n13143), .A2(n13120), .ZN(n10910) );
  AND2_X1 U13450 ( .A1(n10911), .A2(n10910), .ZN(n10958) );
  NAND2_X1 U13451 ( .A1(n10912), .A2(n10958), .ZN(n13608) );
  NAND2_X1 U13452 ( .A1(n13608), .A2(n13471), .ZN(n10918) );
  OAI22_X1 U13453 ( .A1(n13471), .A2(n13188), .B1(n10957), .B2(n13515), .ZN(
        n10916) );
  AOI21_X1 U13454 ( .B1(n10913), .B2(n13603), .A(n13066), .ZN(n10914) );
  NAND2_X1 U13455 ( .A1(n10914), .A2(n13501), .ZN(n13605) );
  NOR2_X1 U13456 ( .A1(n13605), .A2(n13411), .ZN(n10915) );
  AOI211_X1 U13457 ( .C1(n13517), .C2(n13603), .A(n10916), .B(n10915), .ZN(
        n10917) );
  OAI211_X1 U13458 ( .C1(n13507), .C2(n13606), .A(n10918), .B(n10917), .ZN(
        P2_U3249) );
  NAND2_X1 U13459 ( .A1(n14533), .A2(n12442), .ZN(n10919) );
  NAND2_X1 U13460 ( .A1(n10920), .A2(n10919), .ZN(n12075) );
  INV_X1 U13461 ( .A(n12441), .ZN(n12837) );
  OR2_X1 U13462 ( .A1(n12076), .A2(n12837), .ZN(n12340) );
  AND2_X1 U13463 ( .A1(n12076), .A2(n12837), .ZN(n12339) );
  XNOR2_X1 U13464 ( .A(n12075), .B(n12342), .ZN(n10921) );
  OAI222_X1 U13465 ( .A1(n15128), .A2(n12824), .B1(n15130), .B2(n10922), .C1(
        n10921), .C2(n15154), .ZN(n14527) );
  INV_X1 U13466 ( .A(n14527), .ZN(n10932) );
  INV_X1 U13467 ( .A(n10923), .ZN(n12253) );
  NAND2_X1 U13468 ( .A1(n10924), .A2(n12253), .ZN(n10925) );
  XOR2_X1 U13469 ( .A(n12342), .B(n11973), .Z(n14529) );
  AND2_X1 U13470 ( .A1(n12076), .A2(n15155), .ZN(n14528) );
  INV_X1 U13471 ( .A(n14528), .ZN(n10929) );
  AOI22_X1 U13472 ( .A1(n12846), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15157), 
        .B2(n10926), .ZN(n10927) );
  OAI21_X1 U13473 ( .B1(n10929), .B2(n10928), .A(n10927), .ZN(n10930) );
  AOI21_X1 U13474 ( .B1(n14529), .B2(n12844), .A(n10930), .ZN(n10931) );
  OAI21_X1 U13475 ( .B1(n10932), .B2(n12846), .A(n10931), .ZN(P3_U3220) );
  MUX2_X1 U13476 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6641), .Z(n10988) );
  XNOR2_X1 U13477 ( .A(n10988), .B(SI_25_), .ZN(n10992) );
  XNOR2_X1 U13478 ( .A(n10993), .B(n10992), .ZN(n11634) );
  INV_X1 U13479 ( .A(n11634), .ZN(n10936) );
  OAI222_X1 U13480 ( .A1(n11464), .A2(n11249), .B1(n13675), .B2(n10936), .C1(
        P2_U3088), .C2(n10935), .ZN(P2_U3302) );
  OAI222_X1 U13481 ( .A1(n10937), .A2(P1_U3086), .B1(n14373), .B2(n10936), 
        .C1(n11635), .C2(n14370), .ZN(P1_U3330) );
  OAI21_X1 U13482 ( .B1(n10607), .B2(n10939), .A(n10938), .ZN(n13876) );
  XNOR2_X1 U13483 ( .A(n13876), .B(n13875), .ZN(n13877) );
  XOR2_X1 U13484 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n13877), .Z(n10949) );
  AOI21_X1 U13485 ( .B1(n11499), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10940), 
        .ZN(n10941) );
  NOR2_X1 U13486 ( .A1(n10941), .A2(n10945), .ZN(n13882) );
  AOI21_X1 U13487 ( .B1(n10941), .B2(n10945), .A(n13882), .ZN(n10943) );
  AND2_X1 U13488 ( .A1(n10943), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n13883) );
  INV_X1 U13489 ( .A(n13883), .ZN(n10942) );
  OAI211_X1 U13490 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n10943), .A(n10942), 
        .B(n14668), .ZN(n10948) );
  NAND2_X1 U13491 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13794)
         );
  NAND2_X1 U13492 ( .A1(n14656), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n10944) );
  OAI211_X1 U13493 ( .C1(n13885), .C2(n10945), .A(n13794), .B(n10944), .ZN(
        n10946) );
  INV_X1 U13494 ( .A(n10946), .ZN(n10947) );
  OAI211_X1 U13495 ( .C1(n10949), .C2(n13867), .A(n10948), .B(n10947), .ZN(
        P1_U3261) );
  NAND2_X1 U13496 ( .A1(n13248), .A2(n13066), .ZN(n13002) );
  XNOR2_X1 U13497 ( .A(n13603), .B(n13035), .ZN(n13087) );
  XOR2_X1 U13498 ( .A(n13002), .B(n13087), .Z(n10956) );
  INV_X1 U13499 ( .A(n10950), .ZN(n10951) );
  OR2_X1 U13500 ( .A1(n10952), .A2(n10951), .ZN(n10953) );
  AOI21_X1 U13501 ( .B1(n10956), .B2(n10955), .A(n13090), .ZN(n10962) );
  NOR2_X1 U13502 ( .A1(n14558), .A2(n10957), .ZN(n10960) );
  OAI22_X1 U13503 ( .A1(n10958), .A2(n14554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13192), .ZN(n10959) );
  AOI211_X1 U13504 ( .C1(n13603), .C2(n13128), .A(n10960), .B(n10959), .ZN(
        n10961) );
  OAI21_X1 U13505 ( .B1(n10962), .B2(n14552), .A(n10961), .ZN(P2_U3198) );
  AOI22_X1 U13506 ( .A1(n12069), .A2(SI_18_), .B1(n10875), .B2(n12599), .ZN(
        n10964) );
  INV_X1 U13507 ( .A(n12791), .ZN(n12967) );
  XNOR2_X1 U13508 ( .A(n12791), .B(n12155), .ZN(n12119) );
  XNOR2_X1 U13509 ( .A(n12119), .B(n12091), .ZN(n10971) );
  INV_X1 U13510 ( .A(n10966), .ZN(n10968) );
  INV_X1 U13511 ( .A(n12118), .ZN(n10969) );
  OAI211_X1 U13512 ( .C1(n10971), .C2(n10970), .A(n10969), .B(n12168), .ZN(
        n10981) );
  INV_X1 U13513 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U13514 ( .A1(n10972), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U13515 ( .A1(n10974), .A2(n10973), .ZN(n12769) );
  NAND2_X1 U13516 ( .A1(n12769), .A2(n12024), .ZN(n10976) );
  AOI22_X1 U13517 ( .A1(n6638), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n6639), .B2(
        P3_REG1_REG_19__SCAN_IN), .ZN(n10975) );
  OAI211_X1 U13518 ( .C1(n10977), .C2(n12961), .A(n10976), .B(n10975), .ZN(
        n12440) );
  NAND2_X1 U13519 ( .A1(n12440), .A2(n12189), .ZN(n10978) );
  NAND2_X1 U13520 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12580)
         );
  OAI211_X1 U13521 ( .C1(n12779), .C2(n12209), .A(n10978), .B(n12580), .ZN(
        n10979) );
  AOI21_X1 U13522 ( .B1(n12781), .B2(n12207), .A(n10979), .ZN(n10980) );
  OAI211_X1 U13523 ( .C1(n12967), .C2(n12174), .A(n10981), .B(n10980), .ZN(
        P3_U3178) );
  MUX2_X1 U13524 ( .A(n10982), .B(P1_REG2_REG_2__SCAN_IN), .S(n14689), .Z(
        n10987) );
  NAND2_X1 U13525 ( .A1(n14201), .A2(n11730), .ZN(n10984) );
  NAND2_X1 U13526 ( .A1(n14199), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10983) );
  OAI211_X1 U13527 ( .C1(n14130), .C2(n10985), .A(n10984), .B(n10983), .ZN(
        n10986) );
  OR2_X1 U13528 ( .A1(n10987), .A2(n10986), .ZN(P1_U3291) );
  INV_X1 U13529 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11962) );
  INV_X1 U13530 ( .A(n10988), .ZN(n10990) );
  NAND2_X1 U13531 ( .A1(n10990), .A2(n10989), .ZN(n10991) );
  MUX2_X1 U13532 ( .A(n14371), .B(n13682), .S(n6641), .Z(n11269) );
  INV_X1 U13533 ( .A(n11269), .ZN(n10994) );
  NAND2_X1 U13534 ( .A1(n10995), .A2(n10994), .ZN(n10997) );
  INV_X1 U13535 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14368) );
  MUX2_X1 U13536 ( .A(n14368), .B(n11962), .S(n6641), .Z(n11004) );
  INV_X1 U13537 ( .A(n11004), .ZN(n10998) );
  XNOR2_X1 U13538 ( .A(n10998), .B(SI_27_), .ZN(n10999) );
  INV_X1 U13539 ( .A(n11666), .ZN(n14369) );
  OAI222_X1 U13540 ( .A1(n11464), .A2(n11962), .B1(n13675), .B2(n14369), .C1(
        n11000), .C2(P2_U3088), .ZN(P2_U3300) );
  NOR2_X1 U13541 ( .A1(n11004), .A2(n11003), .ZN(n11001) );
  NAND2_X1 U13542 ( .A1(n11004), .A2(n11003), .ZN(n11005) );
  INV_X1 U13543 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11966) );
  INV_X1 U13544 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12066) );
  MUX2_X1 U13545 ( .A(n11966), .B(n12066), .S(n6641), .Z(n11302) );
  XNOR2_X1 U13546 ( .A(n11302), .B(SI_28_), .ZN(n11006) );
  INV_X1 U13547 ( .A(n11684), .ZN(n13679) );
  OAI222_X1 U13548 ( .A1(n11008), .A2(P1_U3086), .B1(n14373), .B2(n13679), 
        .C1(n11966), .C2(n14370), .ZN(P1_U3327) );
  OR2_X1 U13549 ( .A1(n11363), .A2(n11009), .ZN(n11010) );
  NAND2_X1 U13550 ( .A1(n13442), .A2(n11067), .ZN(n11023) );
  NAND2_X1 U13551 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n11012) );
  INV_X1 U13552 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13105) );
  INV_X1 U13553 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n15400) );
  NAND2_X1 U13554 ( .A1(n11189), .A2(n15400), .ZN(n11015) );
  NAND2_X1 U13555 ( .A1(n11202), .A2(n11015), .ZN(n13443) );
  OR2_X1 U13556 ( .A1(n13443), .A2(n6847), .ZN(n11021) );
  INV_X1 U13557 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U13558 ( .A1(n11371), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U13559 ( .A1(n11277), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n11017) );
  OAI211_X1 U13560 ( .C1(n13646), .C2(n11318), .A(n11018), .B(n11017), .ZN(
        n11019) );
  INV_X1 U13561 ( .A(n11019), .ZN(n11020) );
  NAND2_X1 U13562 ( .A1(n11021), .A2(n11020), .ZN(n13261) );
  NAND2_X1 U13563 ( .A1(n13261), .A2(n11262), .ZN(n11022) );
  NAND2_X1 U13564 ( .A1(n11315), .A2(n11168), .ZN(n11025) );
  AND2_X1 U13565 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  AOI21_X1 U13566 ( .B1(n11027), .B2(n11142), .A(n11026), .ZN(n11031) );
  NAND2_X1 U13567 ( .A1(n11027), .A2(n11026), .ZN(n11030) );
  NAND3_X1 U13568 ( .A1(n6917), .A2(n11340), .A3(n11028), .ZN(n11029) );
  OAI211_X1 U13569 ( .C1(n6917), .C2(n11031), .A(n11030), .B(n11029), .ZN(
        n11043) );
  INV_X2 U13570 ( .A(n11142), .ZN(n11262) );
  NAND2_X1 U13571 ( .A1(n13157), .A2(n11262), .ZN(n11033) );
  NAND2_X1 U13572 ( .A1(n6820), .A2(n11067), .ZN(n11032) );
  NAND2_X1 U13573 ( .A1(n11033), .A2(n11032), .ZN(n11042) );
  NAND2_X1 U13574 ( .A1(n13156), .A2(n11067), .ZN(n11036) );
  INV_X2 U13575 ( .A(n11142), .ZN(n11340) );
  NAND2_X1 U13576 ( .A1(n11034), .A2(n11340), .ZN(n11035) );
  NAND2_X1 U13577 ( .A1(n11036), .A2(n11035), .ZN(n11044) );
  AND2_X1 U13578 ( .A1(n11034), .A2(n11067), .ZN(n11038) );
  AOI21_X1 U13579 ( .B1(n13156), .B2(n11340), .A(n11038), .ZN(n11045) );
  NAND2_X1 U13580 ( .A1(n11044), .A2(n11045), .ZN(n11039) );
  OAI21_X1 U13581 ( .B1(n11043), .B2(n11042), .A(n11039), .ZN(n11050) );
  AOI22_X1 U13582 ( .A1(n13157), .A2(n11067), .B1(n11340), .B2(n6820), .ZN(
        n11041) );
  AOI21_X1 U13583 ( .B1(n11043), .B2(n11042), .A(n11041), .ZN(n11049) );
  INV_X1 U13584 ( .A(n11044), .ZN(n11047) );
  INV_X1 U13585 ( .A(n11045), .ZN(n11046) );
  NAND2_X1 U13586 ( .A1(n11047), .A2(n11046), .ZN(n11048) );
  NAND2_X1 U13587 ( .A1(n13155), .A2(n11262), .ZN(n11052) );
  NAND2_X1 U13588 ( .A1(n11056), .A2(n11338), .ZN(n11051) );
  NAND2_X1 U13589 ( .A1(n11052), .A2(n11051), .ZN(n11058) );
  AOI22_X1 U13590 ( .A1(n14926), .A2(n11340), .B1(n13154), .B2(n11338), .ZN(
        n11061) );
  NAND2_X1 U13591 ( .A1(n14926), .A2(n11338), .ZN(n11055) );
  NAND2_X1 U13592 ( .A1(n13154), .A2(n11262), .ZN(n11054) );
  NAND2_X1 U13593 ( .A1(n11055), .A2(n11054), .ZN(n11060) );
  OAI22_X1 U13594 ( .A1(n11059), .A2(n11058), .B1(n11061), .B2(n11060), .ZN(
        n11064) );
  AOI22_X1 U13595 ( .A1(n13155), .A2(n11338), .B1(n11340), .B2(n11056), .ZN(
        n11057) );
  AOI21_X1 U13596 ( .B1(n11059), .B2(n11058), .A(n11057), .ZN(n11063) );
  NAND2_X1 U13597 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U13598 ( .A1(n11068), .A2(n11338), .ZN(n11066) );
  NAND2_X1 U13599 ( .A1(n13153), .A2(n11262), .ZN(n11065) );
  NAND2_X1 U13600 ( .A1(n11068), .A2(n11262), .ZN(n11069) );
  OAI21_X1 U13601 ( .B1(n11070), .B2(n11053), .A(n11069), .ZN(n11071) );
  NAND2_X1 U13602 ( .A1(n11075), .A2(n11262), .ZN(n11074) );
  NAND2_X1 U13603 ( .A1(n13152), .A2(n11338), .ZN(n11073) );
  NAND2_X1 U13604 ( .A1(n11074), .A2(n11073), .ZN(n11078) );
  AOI22_X1 U13605 ( .A1(n11075), .A2(n11338), .B1(n11340), .B2(n13152), .ZN(
        n11076) );
  INV_X1 U13606 ( .A(n11077), .ZN(n11080) );
  NAND2_X1 U13607 ( .A1(n11083), .A2(n11338), .ZN(n11082) );
  NAND2_X1 U13608 ( .A1(n13151), .A2(n11262), .ZN(n11081) );
  NAND2_X1 U13609 ( .A1(n11083), .A2(n11262), .ZN(n11084) );
  OAI21_X1 U13610 ( .B1(n11085), .B2(n11053), .A(n11084), .ZN(n11086) );
  NAND2_X1 U13611 ( .A1(n11089), .A2(n11262), .ZN(n11088) );
  NAND2_X1 U13612 ( .A1(n13150), .A2(n11338), .ZN(n11087) );
  AOI22_X1 U13613 ( .A1(n11089), .A2(n11338), .B1(n11340), .B2(n13150), .ZN(
        n11090) );
  NAND2_X1 U13614 ( .A1(n11094), .A2(n11338), .ZN(n11093) );
  NAND2_X1 U13615 ( .A1(n13149), .A2(n11262), .ZN(n11092) );
  NAND2_X1 U13616 ( .A1(n11094), .A2(n11262), .ZN(n11095) );
  OAI21_X1 U13617 ( .B1(n11096), .B2(n11053), .A(n11095), .ZN(n11097) );
  NAND2_X1 U13618 ( .A1(n13518), .A2(n11262), .ZN(n11099) );
  NAND2_X1 U13619 ( .A1(n13148), .A2(n11338), .ZN(n11098) );
  NAND2_X1 U13620 ( .A1(n11099), .A2(n11098), .ZN(n11102) );
  AOI22_X1 U13621 ( .A1(n13518), .A2(n11338), .B1(n11340), .B2(n13148), .ZN(
        n11100) );
  AOI21_X1 U13622 ( .B1(n11103), .B2(n11102), .A(n11100), .ZN(n11101) );
  NOR2_X1 U13623 ( .A1(n11103), .A2(n11102), .ZN(n11104) );
  NAND2_X1 U13624 ( .A1(n11107), .A2(n11338), .ZN(n11106) );
  NAND2_X1 U13625 ( .A1(n13147), .A2(n11262), .ZN(n11105) );
  NAND2_X1 U13626 ( .A1(n11106), .A2(n11105), .ZN(n11113) );
  NAND2_X1 U13627 ( .A1(n11112), .A2(n11113), .ZN(n11111) );
  NAND2_X1 U13628 ( .A1(n11107), .A2(n11262), .ZN(n11108) );
  OAI21_X1 U13629 ( .B1(n11109), .B2(n11053), .A(n11108), .ZN(n11110) );
  NAND2_X1 U13630 ( .A1(n11116), .A2(n11262), .ZN(n11115) );
  NAND2_X1 U13631 ( .A1(n13146), .A2(n11338), .ZN(n11114) );
  AOI22_X1 U13632 ( .A1(n11116), .A2(n11338), .B1(n11340), .B2(n13146), .ZN(
        n11117) );
  NAND2_X1 U13633 ( .A1(n13618), .A2(n11338), .ZN(n11119) );
  NAND2_X1 U13634 ( .A1(n13145), .A2(n11262), .ZN(n11118) );
  NAND2_X1 U13635 ( .A1(n11119), .A2(n11118), .ZN(n11121) );
  AOI22_X1 U13636 ( .A1(n13618), .A2(n11262), .B1(n13145), .B2(n11338), .ZN(
        n11120) );
  NAND2_X1 U13637 ( .A1(n11125), .A2(n11262), .ZN(n11124) );
  NAND2_X1 U13638 ( .A1(n13144), .A2(n11338), .ZN(n11123) );
  NAND2_X1 U13639 ( .A1(n11124), .A2(n11123), .ZN(n11129) );
  NAND2_X1 U13640 ( .A1(n11125), .A2(n11338), .ZN(n11126) );
  OAI21_X1 U13641 ( .B1(n11127), .B2(n11142), .A(n11126), .ZN(n11128) );
  INV_X1 U13642 ( .A(n11129), .ZN(n11130) );
  NAND2_X1 U13643 ( .A1(n11133), .A2(n11338), .ZN(n11132) );
  NAND2_X1 U13644 ( .A1(n13143), .A2(n11262), .ZN(n11131) );
  NAND2_X1 U13645 ( .A1(n11132), .A2(n11131), .ZN(n11135) );
  AOI22_X1 U13646 ( .A1(n11133), .A2(n11262), .B1(n13143), .B2(n11338), .ZN(
        n11134) );
  AOI21_X1 U13647 ( .B1(n11136), .B2(n11135), .A(n11134), .ZN(n11138) );
  NOR2_X1 U13648 ( .A1(n11136), .A2(n11135), .ZN(n11137) );
  NAND2_X1 U13649 ( .A1(n13603), .A2(n11340), .ZN(n11140) );
  NAND2_X1 U13650 ( .A1(n13248), .A2(n11067), .ZN(n11139) );
  NAND2_X1 U13651 ( .A1(n11140), .A2(n11139), .ZN(n11144) );
  NAND2_X1 U13652 ( .A1(n13603), .A2(n11338), .ZN(n11141) );
  OAI21_X1 U13653 ( .B1(n13283), .B2(n11142), .A(n11141), .ZN(n11143) );
  NAND2_X1 U13654 ( .A1(n11498), .A2(n11362), .ZN(n11147) );
  AOI22_X1 U13655 ( .A1(n11358), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n14853), 
        .B2(n11169), .ZN(n11146) );
  NAND2_X1 U13656 ( .A1(n13599), .A2(n11338), .ZN(n11149) );
  NAND2_X1 U13657 ( .A1(n13286), .A2(n11262), .ZN(n11148) );
  NAND2_X1 U13658 ( .A1(n11149), .A2(n11148), .ZN(n11151) );
  AOI22_X1 U13659 ( .A1(n13599), .A2(n11340), .B1(n13286), .B2(n11338), .ZN(
        n11150) );
  AOI22_X1 U13660 ( .A1(n13218), .A2(n11169), .B1(n11358), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U13661 ( .A1(n13289), .A2(n11340), .ZN(n11164) );
  INV_X1 U13662 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n15516) );
  INV_X1 U13663 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n11154) );
  OR2_X1 U13664 ( .A1(n11317), .A2(n11154), .ZN(n11156) );
  INV_X1 U13665 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13596) );
  OR2_X1 U13666 ( .A1(n6658), .A2(n13596), .ZN(n11155) );
  AND2_X1 U13667 ( .A1(n11156), .A2(n11155), .ZN(n11162) );
  INV_X1 U13668 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11158) );
  INV_X1 U13669 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11157) );
  OAI21_X1 U13670 ( .B1(n11159), .B2(n11158), .A(n11157), .ZN(n11160) );
  AND2_X1 U13671 ( .A1(n11160), .A2(n11173), .ZN(n13492) );
  NAND2_X1 U13672 ( .A1(n13492), .A2(n11370), .ZN(n11161) );
  OAI211_X1 U13673 ( .C1(n11318), .C2(n15516), .A(n11162), .B(n11161), .ZN(
        n13254) );
  NAND2_X1 U13674 ( .A1(n13254), .A2(n11067), .ZN(n11163) );
  NAND2_X1 U13675 ( .A1(n11164), .A2(n11163), .ZN(n11165) );
  NAND2_X1 U13676 ( .A1(n13289), .A2(n11067), .ZN(n11167) );
  NAND2_X1 U13677 ( .A1(n13254), .A2(n11262), .ZN(n11166) );
  NAND2_X1 U13678 ( .A1(n11527), .A2(n11362), .ZN(n11171) );
  AOI22_X1 U13679 ( .A1(n11358), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11169), 
        .B2(n11168), .ZN(n11170) );
  NAND2_X1 U13680 ( .A1(n13588), .A2(n11067), .ZN(n11179) );
  INV_X1 U13681 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n11177) );
  INV_X1 U13682 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U13683 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  NAND2_X1 U13684 ( .A1(n11187), .A2(n11174), .ZN(n13476) );
  OR2_X1 U13685 ( .A1(n13476), .A2(n6847), .ZN(n11176) );
  AOI22_X1 U13686 ( .A1(n11371), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n11277), 
        .B2(P2_REG1_REG_19__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U13687 ( .C1(n11318), .C2(n11177), .A(n11176), .B(n11175), .ZN(
        n13292) );
  NAND2_X1 U13688 ( .A1(n13292), .A2(n11262), .ZN(n11178) );
  NAND2_X1 U13689 ( .A1(n11179), .A2(n11178), .ZN(n11181) );
  AOI22_X1 U13690 ( .A1(n13588), .A2(n11340), .B1(n13292), .B2(n11338), .ZN(
        n11180) );
  NOR2_X1 U13691 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  NAND2_X1 U13692 ( .A1(n11358), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U13693 ( .A1(n13457), .A2(n11262), .ZN(n11193) );
  NAND2_X1 U13694 ( .A1(n11187), .A2(n13105), .ZN(n11188) );
  NAND2_X1 U13695 ( .A1(n11189), .A2(n11188), .ZN(n13461) );
  AOI22_X1 U13696 ( .A1(n11371), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n11277), 
        .B2(P2_REG1_REG_20__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U13697 ( .A1(n11372), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n11190) );
  OAI211_X1 U13698 ( .C1(n13461), .C2(n6847), .A(n11191), .B(n11190), .ZN(
        n13258) );
  NAND2_X1 U13699 ( .A1(n13258), .A2(n11338), .ZN(n11192) );
  NAND2_X1 U13700 ( .A1(n11193), .A2(n11192), .ZN(n11195) );
  AOI22_X1 U13701 ( .A1(n13457), .A2(n11067), .B1(n11340), .B2(n13258), .ZN(
        n11194) );
  INV_X1 U13702 ( .A(n13261), .ZN(n13298) );
  NAND2_X1 U13703 ( .A1(n13442), .A2(n11262), .ZN(n11197) );
  OAI21_X1 U13704 ( .B1(n13298), .B2(n11053), .A(n11197), .ZN(n11198) );
  NAND2_X1 U13705 ( .A1(n11358), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U13706 ( .A1(n13423), .A2(n11262), .ZN(n11210) );
  INV_X1 U13707 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U13708 ( .A1(n11202), .A2(n13115), .ZN(n11203) );
  NAND2_X1 U13709 ( .A1(n11217), .A2(n11203), .ZN(n13424) );
  OR2_X1 U13710 ( .A1(n13424), .A2(n6847), .ZN(n11208) );
  INV_X1 U13711 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13642) );
  NAND2_X1 U13712 ( .A1(n11277), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U13713 ( .A1(n11371), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11204) );
  OAI211_X1 U13714 ( .C1(n13642), .C2(n11333), .A(n11205), .B(n11204), .ZN(
        n11206) );
  INV_X1 U13715 ( .A(n11206), .ZN(n11207) );
  NAND2_X1 U13716 ( .A1(n11208), .A2(n11207), .ZN(n13264) );
  NAND2_X1 U13717 ( .A1(n13264), .A2(n11338), .ZN(n11209) );
  NAND2_X1 U13718 ( .A1(n11210), .A2(n11209), .ZN(n11213) );
  AOI22_X1 U13719 ( .A1(n13423), .A2(n11067), .B1(n11340), .B2(n13264), .ZN(
        n11211) );
  INV_X1 U13720 ( .A(n11212), .ZN(n11214) );
  NAND2_X1 U13721 ( .A1(n11595), .A2(n11362), .ZN(n11216) );
  NAND2_X1 U13722 ( .A1(n11358), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U13723 ( .A1(n13568), .A2(n11067), .ZN(n11225) );
  INV_X1 U13724 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U13725 ( .A1(n11217), .A2(n13044), .ZN(n11218) );
  NAND2_X1 U13726 ( .A1(n11255), .A2(n11218), .ZN(n13408) );
  INV_X1 U13727 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n11221) );
  NAND2_X1 U13728 ( .A1(n11277), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n11220) );
  NAND2_X1 U13729 ( .A1(n11371), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11219) );
  OAI211_X1 U13730 ( .C1(n11333), .C2(n11221), .A(n11220), .B(n11219), .ZN(
        n11222) );
  INV_X1 U13731 ( .A(n11222), .ZN(n11223) );
  OAI21_X1 U13732 ( .B1(n13408), .B2(n6847), .A(n11223), .ZN(n13268) );
  NAND2_X1 U13733 ( .A1(n13268), .A2(n11262), .ZN(n11224) );
  NAND2_X1 U13734 ( .A1(n11225), .A2(n11224), .ZN(n11231) );
  NAND2_X1 U13735 ( .A1(n11230), .A2(n11231), .ZN(n11229) );
  NAND2_X1 U13736 ( .A1(n13568), .A2(n11262), .ZN(n11227) );
  NAND2_X1 U13737 ( .A1(n13268), .A2(n11338), .ZN(n11226) );
  NAND2_X1 U13738 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  NAND2_X1 U13739 ( .A1(n11229), .A2(n11228), .ZN(n11235) );
  NAND2_X1 U13740 ( .A1(n11233), .A2(n11232), .ZN(n11234) );
  OR2_X1 U13741 ( .A1(n11363), .A2(n11237), .ZN(n11238) );
  NAND2_X2 U13742 ( .A1(n11239), .A2(n11238), .ZN(n13558) );
  NAND2_X1 U13743 ( .A1(n13558), .A2(n11262), .ZN(n11246) );
  XNOR2_X1 U13744 ( .A(n11255), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U13745 ( .A1(n13395), .A2(n11370), .ZN(n11244) );
  INV_X1 U13746 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13638) );
  NAND2_X1 U13747 ( .A1(n11277), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11241) );
  NAND2_X1 U13748 ( .A1(n11371), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n11240) );
  OAI211_X1 U13749 ( .C1(n13638), .C2(n11333), .A(n11241), .B(n11240), .ZN(
        n11242) );
  INV_X1 U13750 ( .A(n11242), .ZN(n11243) );
  NAND2_X1 U13751 ( .A1(n11244), .A2(n11243), .ZN(n13271) );
  NAND2_X1 U13752 ( .A1(n13271), .A2(n11338), .ZN(n11245) );
  NAND2_X1 U13753 ( .A1(n11246), .A2(n11245), .ZN(n11248) );
  AOI22_X1 U13754 ( .A1(n13558), .A2(n11067), .B1(n11340), .B2(n13271), .ZN(
        n11247) );
  NAND2_X1 U13755 ( .A1(n11634), .A2(n11362), .ZN(n11251) );
  OR2_X1 U13756 ( .A1(n11363), .A2(n11249), .ZN(n11250) );
  NAND2_X1 U13757 ( .A1(n13379), .A2(n11338), .ZN(n11264) );
  NAND2_X1 U13758 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n11252) );
  INV_X1 U13759 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n11254) );
  INV_X1 U13760 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n11253) );
  OAI21_X1 U13761 ( .B1(n11255), .B2(n11254), .A(n11253), .ZN(n11256) );
  AND2_X1 U13762 ( .A1(n11275), .A2(n11256), .ZN(n13380) );
  NAND2_X1 U13763 ( .A1(n13380), .A2(n11370), .ZN(n11261) );
  INV_X1 U13764 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13635) );
  NAND2_X1 U13765 ( .A1(n11371), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U13766 ( .A1(n9136), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11257) );
  OAI211_X1 U13767 ( .C1(n13635), .C2(n11318), .A(n11258), .B(n11257), .ZN(
        n11259) );
  INV_X1 U13768 ( .A(n11259), .ZN(n11260) );
  NAND2_X1 U13769 ( .A1(n11261), .A2(n11260), .ZN(n13274) );
  NAND2_X1 U13770 ( .A1(n13274), .A2(n11262), .ZN(n11263) );
  NAND2_X1 U13771 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  NAND2_X1 U13772 ( .A1(n13379), .A2(n11262), .ZN(n11267) );
  NAND2_X1 U13773 ( .A1(n13274), .A2(n11067), .ZN(n11266) );
  NAND2_X1 U13774 ( .A1(n11267), .A2(n11266), .ZN(n11268) );
  XNOR2_X1 U13775 ( .A(n11269), .B(SI_26_), .ZN(n11270) );
  XNOR2_X2 U13776 ( .A(n11271), .B(n11270), .ZN(n13680) );
  NAND2_X1 U13777 ( .A1(n13680), .A2(n11362), .ZN(n11273) );
  OR2_X1 U13778 ( .A1(n11363), .A2(n13682), .ZN(n11272) );
  NAND2_X1 U13779 ( .A1(n13547), .A2(n11262), .ZN(n11284) );
  INV_X1 U13780 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15298) );
  NAND2_X1 U13781 ( .A1(n11275), .A2(n15298), .ZN(n11276) );
  NAND2_X1 U13782 ( .A1(n11368), .A2(n11276), .ZN(n13362) );
  OR2_X1 U13783 ( .A1(n13362), .A2(n6847), .ZN(n11282) );
  INV_X1 U13784 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n15432) );
  NAND2_X1 U13785 ( .A1(n11371), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U13786 ( .A1(n11277), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11278) );
  OAI211_X1 U13787 ( .C1(n15432), .C2(n11333), .A(n11279), .B(n11278), .ZN(
        n11280) );
  INV_X1 U13788 ( .A(n11280), .ZN(n11281) );
  NAND2_X1 U13789 ( .A1(n11282), .A2(n11281), .ZN(n13278) );
  NAND2_X1 U13790 ( .A1(n13278), .A2(n11338), .ZN(n11283) );
  NAND2_X1 U13791 ( .A1(n11284), .A2(n11283), .ZN(n11288) );
  AOI22_X1 U13792 ( .A1(n13547), .A2(n11338), .B1(n11340), .B2(n13278), .ZN(
        n11285) );
  NAND2_X1 U13793 ( .A1(n11666), .A2(n11362), .ZN(n11293) );
  OR2_X1 U13794 ( .A1(n11363), .A2(n11962), .ZN(n11292) );
  NAND2_X2 U13795 ( .A1(n11293), .A2(n11292), .ZN(n13541) );
  NAND2_X1 U13796 ( .A1(n13541), .A2(n11338), .ZN(n11301) );
  XNOR2_X1 U13797 ( .A(n11368), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U13798 ( .A1(n13350), .A2(n11370), .ZN(n11299) );
  INV_X1 U13799 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U13800 ( .A1(n11371), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U13801 ( .A1(n9136), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11294) );
  OAI211_X1 U13802 ( .C1(n11296), .C2(n11333), .A(n11295), .B(n11294), .ZN(
        n11297) );
  INV_X1 U13803 ( .A(n11297), .ZN(n11298) );
  NAND2_X1 U13804 ( .A1(n11299), .A2(n11298), .ZN(n13279) );
  NAND2_X1 U13805 ( .A1(n13279), .A2(n11262), .ZN(n11300) );
  NAND2_X1 U13806 ( .A1(n11301), .A2(n11300), .ZN(n11383) );
  INV_X1 U13807 ( .A(SI_28_), .ZN(n13000) );
  NAND2_X1 U13808 ( .A1(n11302), .A2(n13000), .ZN(n11303) );
  INV_X1 U13809 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14366) );
  INV_X1 U13810 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13673) );
  MUX2_X1 U13811 ( .A(n14366), .B(n13673), .S(n6641), .Z(n11305) );
  XNOR2_X1 U13812 ( .A(n11305), .B(SI_29_), .ZN(n11326) );
  INV_X1 U13813 ( .A(SI_29_), .ZN(n12994) );
  NAND2_X1 U13814 ( .A1(n11305), .A2(n12994), .ZN(n11343) );
  MUX2_X1 U13815 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6641), .Z(n11306) );
  NAND2_X1 U13816 ( .A1(n11306), .A2(SI_30_), .ZN(n11348) );
  INV_X1 U13817 ( .A(n11306), .ZN(n11307) );
  INV_X1 U13818 ( .A(SI_30_), .ZN(n12989) );
  NAND2_X1 U13819 ( .A1(n11307), .A2(n12989), .ZN(n11344) );
  AND2_X1 U13820 ( .A1(n11348), .A2(n11344), .ZN(n11308) );
  NAND2_X1 U13821 ( .A1(n13669), .A2(n11362), .ZN(n11311) );
  NAND2_X1 U13822 ( .A1(n11358), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11310) );
  INV_X1 U13823 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U13824 ( .A1(n11371), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U13825 ( .A1(n11277), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n11312) );
  OAI211_X1 U13826 ( .C1(n11333), .C2(n13623), .A(n11313), .B(n11312), .ZN(
        n13239) );
  OAI211_X1 U13827 ( .C1(n11315), .C2(n11396), .A(n6640), .B(n11314), .ZN(
        n11316) );
  AOI21_X1 U13828 ( .B1(n13239), .B2(n11338), .A(n11316), .ZN(n11322) );
  INV_X1 U13829 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13530) );
  OR2_X1 U13830 ( .A1(n6658), .A2(n13530), .ZN(n11321) );
  INV_X1 U13831 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13243) );
  OR2_X1 U13832 ( .A1(n11317), .A2(n13243), .ZN(n11320) );
  INV_X1 U13833 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15423) );
  OR2_X1 U13834 ( .A1(n11318), .A2(n15423), .ZN(n11319) );
  AND3_X1 U13835 ( .A1(n11321), .A2(n11320), .A3(n11319), .ZN(n13313) );
  NOR2_X1 U13836 ( .A1(n11322), .A2(n13313), .ZN(n11323) );
  AOI21_X1 U13837 ( .B1(n13246), .B2(n11340), .A(n11323), .ZN(n11442) );
  NAND2_X1 U13838 ( .A1(n13246), .A2(n11067), .ZN(n11325) );
  INV_X1 U13839 ( .A(n13313), .ZN(n13140) );
  NAND2_X1 U13840 ( .A1(n13140), .A2(n11262), .ZN(n11324) );
  NAND2_X1 U13841 ( .A1(n11325), .A2(n11324), .ZN(n11441) );
  NAND2_X1 U13842 ( .A1(n13672), .A2(n11362), .ZN(n11329) );
  OR2_X1 U13843 ( .A1(n11363), .A2(n13673), .ZN(n11328) );
  NAND2_X1 U13844 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n11330) );
  INV_X1 U13845 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U13846 ( .A1(n11371), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U13847 ( .A1(n9136), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11331) );
  OAI211_X1 U13848 ( .C1(n11334), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        n11335) );
  INV_X1 U13849 ( .A(n11335), .ZN(n11336) );
  OAI21_X1 U13850 ( .B1(n13318), .B2(n6847), .A(n11336), .ZN(n13141) );
  AND2_X1 U13851 ( .A1(n13141), .A2(n11338), .ZN(n11339) );
  AOI21_X1 U13852 ( .B1(n13534), .B2(n11340), .A(n11339), .ZN(n11431) );
  NAND2_X1 U13853 ( .A1(n13534), .A2(n11338), .ZN(n11342) );
  NAND2_X1 U13854 ( .A1(n13141), .A2(n11262), .ZN(n11341) );
  NAND2_X1 U13855 ( .A1(n11342), .A2(n11341), .ZN(n11430) );
  OAI22_X1 U13856 ( .A1(n11442), .A2(n11441), .B1(n11431), .B2(n11430), .ZN(
        n11361) );
  NAND2_X1 U13857 ( .A1(n11344), .A2(n11343), .ZN(n11351) );
  MUX2_X1 U13858 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6641), .Z(n11346) );
  INV_X1 U13859 ( .A(SI_31_), .ZN(n12986) );
  XNOR2_X1 U13860 ( .A(n11346), .B(n12986), .ZN(n11350) );
  INV_X1 U13861 ( .A(n11350), .ZN(n11347) );
  NOR2_X1 U13862 ( .A1(n11351), .A2(n11347), .ZN(n11357) );
  XNOR2_X1 U13863 ( .A(n11347), .B(n11348), .ZN(n11356) );
  INV_X1 U13864 ( .A(n11353), .ZN(n11349) );
  NOR2_X1 U13865 ( .A1(n11351), .A2(n11350), .ZN(n11352) );
  NAND2_X1 U13866 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  NAND2_X1 U13867 ( .A1(n13665), .A2(n11362), .ZN(n11360) );
  NAND2_X1 U13868 ( .A1(n11358), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U13869 ( .A1(n11361), .A2(n11438), .ZN(n11440) );
  NAND2_X1 U13870 ( .A1(n11684), .A2(n11362), .ZN(n11365) );
  OR2_X1 U13871 ( .A1(n11363), .A2(n12066), .ZN(n11364) );
  INV_X1 U13872 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n11367) );
  INV_X1 U13873 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11366) );
  OAI21_X1 U13874 ( .B1(n11368), .B2(n11367), .A(n11366), .ZN(n11369) );
  NAND2_X1 U13875 ( .A1(n13331), .A2(n11370), .ZN(n11377) );
  INV_X1 U13876 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U13877 ( .A1(n11371), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U13878 ( .A1(n11372), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11373) );
  OAI211_X1 U13879 ( .C1(n6658), .C2(n15444), .A(n11374), .B(n11373), .ZN(
        n11375) );
  INV_X1 U13880 ( .A(n11375), .ZN(n11376) );
  NAND2_X1 U13881 ( .A1(n11377), .A2(n11376), .ZN(n13142) );
  AND2_X1 U13882 ( .A1(n13142), .A2(n11340), .ZN(n11378) );
  AOI21_X1 U13883 ( .B1(n13336), .B2(n11067), .A(n11378), .ZN(n11433) );
  NAND2_X1 U13884 ( .A1(n13336), .A2(n11262), .ZN(n11380) );
  NAND2_X1 U13885 ( .A1(n13142), .A2(n11338), .ZN(n11379) );
  NAND2_X1 U13886 ( .A1(n11380), .A2(n11379), .ZN(n11432) );
  NAND2_X1 U13887 ( .A1(n11433), .A2(n11432), .ZN(n11381) );
  OAI211_X1 U13888 ( .C1(n11384), .C2(n11383), .A(n11440), .B(n11381), .ZN(
        n11386) );
  AOI22_X1 U13889 ( .A1(n13541), .A2(n11262), .B1(n13279), .B2(n11338), .ZN(
        n11382) );
  AOI21_X1 U13890 ( .B1(n11384), .B2(n11383), .A(n11382), .ZN(n11385) );
  AND2_X1 U13891 ( .A1(n13239), .A2(n11053), .ZN(n11388) );
  NOR2_X1 U13892 ( .A1(n13239), .A2(n11340), .ZN(n11387) );
  MUX2_X1 U13893 ( .A(n11388), .B(n11387), .S(n13233), .Z(n11452) );
  INV_X1 U13894 ( .A(n11452), .ZN(n11392) );
  OAI21_X1 U13895 ( .B1(n6640), .B2(n11427), .A(n13227), .ZN(n11389) );
  OAI21_X1 U13896 ( .B1(n11458), .B2(n11390), .A(n11389), .ZN(n11391) );
  NAND2_X1 U13897 ( .A1(n11392), .A2(n11391), .ZN(n11454) );
  INV_X1 U13898 ( .A(n11454), .ZN(n11393) );
  XNOR2_X1 U13899 ( .A(n13246), .B(n13140), .ZN(n11424) );
  NAND2_X1 U13900 ( .A1(n13336), .A2(n13315), .ZN(n11394) );
  INV_X1 U13901 ( .A(n13279), .ZN(n13310) );
  XNOR2_X1 U13902 ( .A(n13541), .B(n13310), .ZN(n13354) );
  INV_X1 U13903 ( .A(n13274), .ZN(n13306) );
  XNOR2_X1 U13904 ( .A(n13379), .B(n13306), .ZN(n13371) );
  INV_X1 U13905 ( .A(n13278), .ZN(n11395) );
  NAND2_X1 U13906 ( .A1(n13547), .A2(n11395), .ZN(n13309) );
  INV_X1 U13907 ( .A(n13264), .ZN(n13300) );
  XNOR2_X1 U13908 ( .A(n13423), .B(n13300), .ZN(n13420) );
  XNOR2_X1 U13909 ( .A(n13442), .B(n13298), .ZN(n13438) );
  INV_X1 U13910 ( .A(n13292), .ZN(n13291) );
  XNOR2_X1 U13911 ( .A(n13588), .B(n13291), .ZN(n13431) );
  INV_X1 U13912 ( .A(n13258), .ZN(n13259) );
  OR2_X1 U13913 ( .A1(n13457), .A2(n13259), .ZN(n13293) );
  NAND2_X1 U13914 ( .A1(n13457), .A2(n13259), .ZN(n13432) );
  NAND4_X1 U13915 ( .A1(n11397), .A2(n11398), .A3(n11399), .A4(n11396), .ZN(
        n11401) );
  NOR4_X1 U13916 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11406) );
  NAND4_X1 U13917 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11408) );
  NOR4_X1 U13918 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11414) );
  NAND4_X1 U13919 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11417) );
  INV_X1 U13920 ( .A(n13286), .ZN(n13285) );
  XNOR2_X1 U13921 ( .A(n13599), .B(n13285), .ZN(n13505) );
  NOR3_X1 U13922 ( .A1(n11417), .A2(n13505), .A3(n11416), .ZN(n11419) );
  XNOR2_X1 U13923 ( .A(n13289), .B(n13254), .ZN(n13484) );
  NAND4_X1 U13924 ( .A1(n13452), .A2(n11419), .A3(n13484), .A4(n11418), .ZN(
        n11420) );
  NOR4_X1 U13925 ( .A1(n13420), .A2(n13438), .A3(n13431), .A4(n11420), .ZN(
        n11421) );
  XNOR2_X1 U13926 ( .A(n13568), .B(n13268), .ZN(n13405) );
  NAND4_X1 U13927 ( .A1(n13367), .A2(n11421), .A3(n13405), .A4(n13398), .ZN(
        n11422) );
  NOR4_X1 U13928 ( .A1(n13332), .A2(n13354), .A3(n13371), .A4(n11422), .ZN(
        n11423) );
  NAND2_X1 U13929 ( .A1(n11426), .A2(n11425), .ZN(n11448) );
  NOR2_X1 U13930 ( .A1(n11427), .A2(n13227), .ZN(n11428) );
  AOI22_X1 U13931 ( .A1(n11458), .A2(n11429), .B1(n11428), .B2(n6640), .ZN(
        n11450) );
  NAND2_X1 U13932 ( .A1(n11431), .A2(n11430), .ZN(n11437) );
  INV_X1 U13933 ( .A(n11432), .ZN(n11435) );
  INV_X1 U13934 ( .A(n11433), .ZN(n11434) );
  NAND2_X1 U13935 ( .A1(n11435), .A2(n11434), .ZN(n11436) );
  NAND3_X1 U13936 ( .A1(n11438), .A2(n11437), .A3(n11436), .ZN(n11439) );
  NAND2_X1 U13937 ( .A1(n11440), .A2(n11439), .ZN(n11444) );
  NAND2_X1 U13938 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  INV_X1 U13939 ( .A(n11450), .ZN(n11451) );
  NAND2_X1 U13940 ( .A1(n11452), .A2(n11451), .ZN(n11453) );
  NAND4_X1 U13941 ( .A1(n11456), .A2(n13235), .A3(n11455), .A4(n13120), .ZN(
        n11457) );
  OAI211_X1 U13942 ( .C1(n11458), .C2(n11460), .A(n11457), .B(P2_B_REG_SCAN_IN), .ZN(n11459) );
  OAI21_X1 U13943 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(P2_U3328) );
  OAI222_X1 U13944 ( .A1(n11464), .A2(n11463), .B1(n13675), .B2(n11462), .C1(
        n13227), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U13945 ( .A1(n14602), .A2(n11699), .ZN(n11466) );
  NAND2_X1 U13946 ( .A1(n13824), .A2(n10521), .ZN(n11465) );
  NAND2_X1 U13947 ( .A1(n11466), .A2(n11465), .ZN(n11467) );
  XNOR2_X1 U13948 ( .A(n11467), .B(n11678), .ZN(n11479) );
  NOR2_X1 U13949 ( .A1(n13772), .A2(n11696), .ZN(n11468) );
  AOI21_X1 U13950 ( .B1(n14602), .B2(n10521), .A(n11468), .ZN(n11475) );
  INV_X1 U13951 ( .A(n11475), .ZN(n11478) );
  NAND2_X1 U13952 ( .A1(n11470), .A2(n11469), .ZN(n11471) );
  NOR2_X1 U13953 ( .A1(n14610), .A2(n11696), .ZN(n11473) );
  AOI21_X1 U13954 ( .B1(n11798), .B2(n10521), .A(n11473), .ZN(n11476) );
  AOI22_X1 U13955 ( .A1(n11798), .A2(n11699), .B1(n10521), .B2(n14564), .ZN(
        n11474) );
  XNOR2_X1 U13956 ( .A(n11474), .B(n11678), .ZN(n11477) );
  XOR2_X1 U13957 ( .A(n11476), .B(n11477), .Z(n13771) );
  XNOR2_X1 U13958 ( .A(n11479), .B(n11475), .ZN(n14562) );
  OR2_X1 U13959 ( .A1(n11477), .A2(n11476), .ZN(n14559) );
  NAND2_X1 U13960 ( .A1(n13910), .A2(n11699), .ZN(n11481) );
  NAND2_X1 U13961 ( .A1(n14590), .A2(n10521), .ZN(n11480) );
  NAND2_X1 U13962 ( .A1(n11481), .A2(n11480), .ZN(n11482) );
  XNOR2_X1 U13963 ( .A(n11482), .B(n11678), .ZN(n11483) );
  AOI22_X1 U13964 ( .A1(n13910), .A2(n11698), .B1(n11680), .B2(n14590), .ZN(
        n13812) );
  INV_X1 U13965 ( .A(n11483), .ZN(n11484) );
  NAND2_X1 U13966 ( .A1(n11485), .A2(n11484), .ZN(n11486) );
  NAND2_X1 U13967 ( .A1(n13810), .A2(n11486), .ZN(n13738) );
  NAND2_X1 U13968 ( .A1(n11487), .A2(n11897), .ZN(n11490) );
  AOI22_X1 U13969 ( .A1(n11529), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11528), 
        .B2(n11488), .ZN(n11489) );
  OAI22_X1 U13970 ( .A1(n14181), .A2(n6646), .B1(n13912), .B2(n11696), .ZN(
        n11493) );
  OAI22_X1 U13971 ( .A1(n14181), .A2(n7432), .B1(n13912), .B2(n6646), .ZN(
        n11491) );
  XNOR2_X1 U13972 ( .A(n11491), .B(n11678), .ZN(n11492) );
  XOR2_X1 U13973 ( .A(n11493), .B(n11492), .Z(n13739) );
  NAND2_X1 U13974 ( .A1(n13738), .A2(n13739), .ZN(n11497) );
  INV_X1 U13975 ( .A(n11492), .ZN(n11495) );
  INV_X1 U13976 ( .A(n11493), .ZN(n11494) );
  NAND2_X1 U13977 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  NAND2_X1 U13978 ( .A1(n11498), .A2(n11897), .ZN(n11501) );
  AOI22_X1 U13979 ( .A1(n11529), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11528), 
        .B2(n11499), .ZN(n11500) );
  NAND2_X1 U13980 ( .A1(n14158), .A2(n11699), .ZN(n11508) );
  INV_X1 U13981 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11502) );
  AND2_X1 U13982 ( .A1(n11503), .A2(n11502), .ZN(n11504) );
  OR2_X1 U13983 ( .A1(n11504), .A2(n11517), .ZN(n14161) );
  AOI22_X1 U13984 ( .A1(n11885), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6645), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U13985 ( .A1(n11884), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11505) );
  OAI211_X1 U13986 ( .C1(n14161), .C2(n11704), .A(n11506), .B(n11505), .ZN(
        n14173) );
  NAND2_X1 U13987 ( .A1(n14173), .A2(n10521), .ZN(n11507) );
  NAND2_X1 U13988 ( .A1(n11508), .A2(n11507), .ZN(n11509) );
  XNOR2_X1 U13989 ( .A(n11509), .B(n11678), .ZN(n11512) );
  AOI22_X1 U13990 ( .A1(n14158), .A2(n10521), .B1(n11680), .B2(n14173), .ZN(
        n11510) );
  XNOR2_X1 U13991 ( .A(n11512), .B(n11510), .ZN(n13746) );
  INV_X1 U13992 ( .A(n11510), .ZN(n11511) );
  NOR2_X1 U13993 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  AOI22_X1 U13994 ( .A1(n11529), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11528), 
        .B2(n13875), .ZN(n11515) );
  NAND2_X1 U13995 ( .A1(n11517), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11532) );
  OR2_X1 U13996 ( .A1(n11517), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U13997 ( .A1(n11532), .A2(n11518), .ZN(n14143) );
  AOI22_X1 U13998 ( .A1(n11885), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6645), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U13999 ( .A1(n11884), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11519) );
  OAI211_X1 U14000 ( .C1(n14143), .C2(n11671), .A(n11520), .B(n11519), .ZN(
        n14160) );
  INV_X1 U14001 ( .A(n14160), .ZN(n13915) );
  OAI22_X1 U14002 ( .A1(n14147), .A2(n7432), .B1(n13915), .B2(n6646), .ZN(
        n11521) );
  XNOR2_X1 U14003 ( .A(n11521), .B(n11678), .ZN(n11522) );
  OAI22_X1 U14004 ( .A1(n14147), .A2(n6646), .B1(n13915), .B2(n11696), .ZN(
        n11523) );
  XNOR2_X1 U14005 ( .A(n11522), .B(n11523), .ZN(n13793) );
  INV_X1 U14006 ( .A(n11522), .ZN(n11525) );
  INV_X1 U14007 ( .A(n11523), .ZN(n11524) );
  NAND2_X1 U14008 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  NAND2_X1 U14009 ( .A1(n11527), .A2(n11897), .ZN(n11531) );
  AOI22_X1 U14010 ( .A1(n11529), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14677), 
        .B2(n11528), .ZN(n11530) );
  INV_X1 U14011 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14127) );
  INV_X1 U14012 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U14013 ( .A1(n11532), .A2(n13716), .ZN(n11533) );
  NAND2_X1 U14014 ( .A1(n11548), .A2(n11533), .ZN(n14126) );
  OR2_X1 U14015 ( .A1(n14126), .A2(n11704), .ZN(n11535) );
  AOI22_X1 U14016 ( .A1(n11885), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6645), 
        .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n11534) );
  OAI211_X1 U14017 ( .C1(n11656), .C2(n14127), .A(n11535), .B(n11534), .ZN(
        n13823) );
  AND2_X1 U14018 ( .A1(n13823), .A2(n11680), .ZN(n11536) );
  AOI21_X1 U14019 ( .B1(n14133), .B2(n10521), .A(n11536), .ZN(n11540) );
  NAND2_X1 U14020 ( .A1(n14133), .A2(n11699), .ZN(n11538) );
  NAND2_X1 U14021 ( .A1(n13823), .A2(n10521), .ZN(n11537) );
  NAND2_X1 U14022 ( .A1(n11538), .A2(n11537), .ZN(n11539) );
  XNOR2_X1 U14023 ( .A(n11539), .B(n11678), .ZN(n11542) );
  XOR2_X1 U14024 ( .A(n11540), .B(n11542), .Z(n13712) );
  INV_X1 U14025 ( .A(n11540), .ZN(n11541) );
  NAND2_X1 U14026 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  OR2_X1 U14027 ( .A1(n11544), .A2(n11612), .ZN(n11547) );
  OR2_X1 U14028 ( .A1(n8839), .A2(n11545), .ZN(n11546) );
  INV_X1 U14029 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13765) );
  NAND2_X1 U14030 ( .A1(n11548), .A2(n13765), .ZN(n11550) );
  INV_X1 U14031 ( .A(n11564), .ZN(n11549) );
  NAND2_X1 U14032 ( .A1(n11550), .A2(n11549), .ZN(n14115) );
  OR2_X1 U14033 ( .A1(n14115), .A2(n11671), .ZN(n11556) );
  INV_X1 U14034 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14035 ( .A1(n11884), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U14036 ( .A1(n6644), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11551) );
  OAI211_X1 U14037 ( .C1(n11881), .C2(n11553), .A(n11552), .B(n11551), .ZN(
        n11554) );
  INV_X1 U14038 ( .A(n11554), .ZN(n11555) );
  OAI22_X1 U14039 ( .A1(n14272), .A2(n6646), .B1(n13920), .B2(n11696), .ZN(
        n11558) );
  OAI22_X1 U14040 ( .A1(n14272), .A2(n7432), .B1(n13920), .B2(n6646), .ZN(
        n11557) );
  XNOR2_X1 U14041 ( .A(n11557), .B(n11678), .ZN(n11559) );
  XOR2_X1 U14042 ( .A(n11558), .B(n11559), .Z(n13763) );
  OR2_X1 U14043 ( .A1(n11560), .A2(n11612), .ZN(n11563) );
  OR2_X1 U14044 ( .A1(n8839), .A2(n11561), .ZN(n11562) );
  NAND2_X1 U14045 ( .A1(n6645), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11568) );
  INV_X1 U14046 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15517) );
  OR2_X1 U14047 ( .A1(n11881), .A2(n15517), .ZN(n11567) );
  NAND2_X1 U14048 ( .A1(n11564), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11580) );
  OAI21_X1 U14049 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n11564), .A(n11580), 
        .ZN(n14101) );
  OR2_X1 U14050 ( .A1(n11671), .A2(n14101), .ZN(n11566) );
  INV_X1 U14051 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14102) );
  OR2_X1 U14052 ( .A1(n11656), .A2(n14102), .ZN(n11565) );
  OAI22_X1 U14053 ( .A1(n14342), .A2(n6646), .B1(n14080), .B2(n11696), .ZN(
        n11572) );
  AOI22_X1 U14054 ( .A1(n14100), .A2(n11699), .B1(n10521), .B2(n14261), .ZN(
        n11569) );
  XNOR2_X1 U14055 ( .A(n11569), .B(n11678), .ZN(n11574) );
  XOR2_X1 U14056 ( .A(n11572), .B(n11574), .Z(n13723) );
  INV_X1 U14057 ( .A(n13723), .ZN(n11570) );
  INV_X1 U14058 ( .A(n11572), .ZN(n11573) );
  NAND2_X1 U14059 ( .A1(n11574), .A2(n11573), .ZN(n11575) );
  OR2_X1 U14060 ( .A1(n11576), .A2(n6641), .ZN(n11577) );
  XNOR2_X1 U14061 ( .A(n11577), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U14062 ( .A1(n11885), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11586) );
  INV_X1 U14063 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11579) );
  OR2_X1 U14064 ( .A1(n11888), .A2(n11579), .ZN(n11585) );
  INV_X1 U14065 ( .A(n11599), .ZN(n11601) );
  OAI21_X1 U14066 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11581), .A(n11601), 
        .ZN(n14077) );
  OR2_X1 U14067 ( .A1(n11704), .A2(n14077), .ZN(n11584) );
  INV_X1 U14068 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11582) );
  OR2_X1 U14069 ( .A1(n11656), .A2(n11582), .ZN(n11583) );
  NAND4_X1 U14070 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n14087) );
  INV_X1 U14071 ( .A(n14087), .ZN(n13945) );
  OAI22_X1 U14072 ( .A1(n13791), .A2(n6646), .B1(n13945), .B2(n11696), .ZN(
        n11591) );
  NAND2_X1 U14073 ( .A1(n14263), .A2(n11699), .ZN(n11588) );
  NAND2_X1 U14074 ( .A1(n14087), .A2(n10521), .ZN(n11587) );
  NAND2_X1 U14075 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  XNOR2_X1 U14076 ( .A(n11589), .B(n11678), .ZN(n11590) );
  XOR2_X1 U14077 ( .A(n11591), .B(n11590), .Z(n13784) );
  INV_X1 U14078 ( .A(n11590), .ZN(n11593) );
  INV_X1 U14079 ( .A(n11591), .ZN(n11592) );
  NAND2_X1 U14080 ( .A1(n11593), .A2(n11592), .ZN(n11594) );
  NAND2_X1 U14081 ( .A1(n11595), .A2(n11897), .ZN(n11598) );
  OR2_X1 U14082 ( .A1(n8839), .A2(n11596), .ZN(n11597) );
  NAND2_X1 U14083 ( .A1(n6644), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11606) );
  INV_X1 U14084 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14055) );
  OR2_X1 U14085 ( .A1(n11656), .A2(n14055), .ZN(n11605) );
  INV_X1 U14086 ( .A(n11618), .ZN(n11620) );
  INV_X1 U14087 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14088 ( .A1(n11601), .A2(n11600), .ZN(n11602) );
  NAND2_X1 U14089 ( .A1(n11620), .A2(n11602), .ZN(n14054) );
  OR2_X1 U14090 ( .A1(n11704), .A2(n14054), .ZN(n11604) );
  INV_X1 U14091 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n14259) );
  OR2_X1 U14092 ( .A1(n11881), .A2(n14259), .ZN(n11603) );
  OAI22_X1 U14093 ( .A1(n14337), .A2(n6646), .B1(n13924), .B2(n11696), .ZN(
        n11609) );
  OAI22_X1 U14094 ( .A1(n14337), .A2(n7432), .B1(n13924), .B2(n6646), .ZN(
        n11607) );
  XNOR2_X1 U14095 ( .A(n11607), .B(n11678), .ZN(n11608) );
  XOR2_X1 U14096 ( .A(n11609), .B(n11608), .Z(n13695) );
  INV_X1 U14097 ( .A(n11608), .ZN(n11611) );
  INV_X1 U14098 ( .A(n11609), .ZN(n11610) );
  OR2_X1 U14099 ( .A1(n8839), .A2(n11614), .ZN(n11615) );
  NAND2_X2 U14100 ( .A1(n11616), .A2(n11615), .ZN(n14045) );
  NAND2_X1 U14101 ( .A1(n14045), .A2(n11699), .ZN(n11628) );
  NAND2_X1 U14102 ( .A1(n6645), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11626) );
  INV_X1 U14103 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11617) );
  OR2_X1 U14104 ( .A1(n11881), .A2(n11617), .ZN(n11625) );
  INV_X1 U14105 ( .A(n11638), .ZN(n11622) );
  INV_X1 U14106 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14107 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U14108 ( .A1(n11622), .A2(n11621), .ZN(n14040) );
  INV_X1 U14109 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14041) );
  OR2_X1 U14110 ( .A1(n11656), .A2(n14041), .ZN(n11623) );
  NAND4_X1 U14111 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n14020) );
  NAND2_X1 U14112 ( .A1(n14020), .A2(n10521), .ZN(n11627) );
  NAND2_X1 U14113 ( .A1(n11628), .A2(n11627), .ZN(n11629) );
  XNOR2_X1 U14114 ( .A(n11629), .B(n11678), .ZN(n11630) );
  AOI22_X1 U14115 ( .A1(n14045), .A2(n11698), .B1(n11680), .B2(n14020), .ZN(
        n11631) );
  XNOR2_X1 U14116 ( .A(n11630), .B(n11631), .ZN(n13755) );
  INV_X1 U14117 ( .A(n11630), .ZN(n11632) );
  NAND2_X1 U14118 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  NAND2_X1 U14119 ( .A1(n11634), .A2(n11897), .ZN(n11637) );
  OR2_X1 U14120 ( .A1(n8839), .A2(n11635), .ZN(n11636) );
  NAND2_X1 U14121 ( .A1(n14030), .A2(n11699), .ZN(n11645) );
  NAND2_X1 U14122 ( .A1(n11885), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11643) );
  INV_X1 U14123 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n14330) );
  OR2_X1 U14124 ( .A1(n11888), .A2(n14330), .ZN(n11642) );
  NAND2_X1 U14125 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n11638), .ZN(n11654) );
  OAI21_X1 U14126 ( .B1(n11638), .B2(P1_REG3_REG_25__SCAN_IN), .A(n11654), 
        .ZN(n14022) );
  OR2_X1 U14127 ( .A1(n11704), .A2(n14022), .ZN(n11641) );
  INV_X1 U14128 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11639) );
  OR2_X1 U14129 ( .A1(n11656), .A2(n11639), .ZN(n11640) );
  NAND4_X1 U14130 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n13999) );
  NAND2_X1 U14131 ( .A1(n13999), .A2(n10521), .ZN(n11644) );
  NAND2_X1 U14132 ( .A1(n11645), .A2(n11644), .ZN(n11646) );
  XNOR2_X1 U14133 ( .A(n11646), .B(n11678), .ZN(n11647) );
  AOI22_X1 U14134 ( .A1(n14030), .A2(n10521), .B1(n11680), .B2(n13999), .ZN(
        n11648) );
  XNOR2_X1 U14135 ( .A(n11647), .B(n11648), .ZN(n13730) );
  INV_X1 U14136 ( .A(n11647), .ZN(n11649) );
  NAND2_X1 U14137 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  NAND2_X1 U14138 ( .A1(n13680), .A2(n11897), .ZN(n11652) );
  OR2_X1 U14139 ( .A1(n8839), .A2(n14371), .ZN(n11651) );
  NAND2_X1 U14140 ( .A1(n11885), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11660) );
  INV_X1 U14141 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11653) );
  OR2_X1 U14142 ( .A1(n11888), .A2(n11653), .ZN(n11659) );
  INV_X1 U14143 ( .A(n11654), .ZN(n11655) );
  NAND2_X1 U14144 ( .A1(n11655), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11670) );
  OAI21_X1 U14145 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n11655), .A(n11670), 
        .ZN(n14008) );
  OR2_X1 U14146 ( .A1(n11704), .A2(n14008), .ZN(n11658) );
  INV_X1 U14147 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14009) );
  OR2_X1 U14148 ( .A1(n11656), .A2(n14009), .ZN(n11657) );
  OAI22_X1 U14149 ( .A1(n14007), .A2(n6646), .B1(n14021), .B2(n11696), .ZN(
        n11663) );
  OAI22_X1 U14150 ( .A1(n14007), .A2(n7432), .B1(n14021), .B2(n6646), .ZN(
        n11661) );
  XNOR2_X1 U14151 ( .A(n11661), .B(n11678), .ZN(n11662) );
  XOR2_X1 U14152 ( .A(n11663), .B(n11662), .Z(n13801) );
  INV_X1 U14153 ( .A(n11662), .ZN(n11665) );
  INV_X1 U14154 ( .A(n11663), .ZN(n11664) );
  NAND2_X1 U14155 ( .A1(n11666), .A2(n11897), .ZN(n11668) );
  OR2_X1 U14156 ( .A1(n8839), .A2(n14368), .ZN(n11667) );
  NAND2_X1 U14157 ( .A1(n13991), .A2(n11699), .ZN(n11677) );
  NAND2_X1 U14158 ( .A1(n6644), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11675) );
  INV_X1 U14159 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n11669) );
  OR2_X1 U14160 ( .A1(n11656), .A2(n11669), .ZN(n11674) );
  XNOR2_X1 U14161 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n11687), .ZN(n13989) );
  OR2_X1 U14162 ( .A1(n11671), .A2(n13989), .ZN(n11673) );
  INV_X1 U14163 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15350) );
  OR2_X1 U14164 ( .A1(n11881), .A2(n15350), .ZN(n11672) );
  NAND4_X1 U14165 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(
        n14000) );
  NAND2_X1 U14166 ( .A1(n14000), .A2(n10521), .ZN(n11676) );
  NAND2_X1 U14167 ( .A1(n11677), .A2(n11676), .ZN(n11679) );
  XNOR2_X1 U14168 ( .A(n11679), .B(n11678), .ZN(n11681) );
  AOI22_X1 U14169 ( .A1(n13991), .A2(n10521), .B1(n11680), .B2(n14000), .ZN(
        n11682) );
  XNOR2_X1 U14170 ( .A(n11681), .B(n11682), .ZN(n13686) );
  INV_X1 U14171 ( .A(n11681), .ZN(n11683) );
  AOI22_X1 U14172 ( .A1(n13687), .A2(n13686), .B1(n11683), .B2(n11682), .ZN(
        n11703) );
  NAND2_X1 U14173 ( .A1(n11684), .A2(n11897), .ZN(n11686) );
  OR2_X1 U14174 ( .A1(n8839), .A2(n11966), .ZN(n11685) );
  NAND2_X1 U14175 ( .A1(n11885), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11695) );
  INV_X1 U14176 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15326) );
  OR2_X1 U14177 ( .A1(n11888), .A2(n15326), .ZN(n11694) );
  NAND2_X1 U14178 ( .A1(n11688), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13953) );
  INV_X1 U14179 ( .A(n11688), .ZN(n11690) );
  INV_X1 U14180 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11689) );
  NAND2_X1 U14181 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  NAND2_X1 U14182 ( .A1(n13953), .A2(n11691), .ZN(n13967) );
  OR2_X1 U14183 ( .A1(n11704), .A2(n13967), .ZN(n11693) );
  INV_X1 U14184 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13970) );
  OR2_X1 U14185 ( .A1(n11656), .A2(n13970), .ZN(n11692) );
  OAI22_X1 U14186 ( .A1(n14323), .A2(n6646), .B1(n14219), .B2(n11696), .ZN(
        n11697) );
  XNOR2_X1 U14187 ( .A(n11697), .B(n11678), .ZN(n11701) );
  INV_X2 U14188 ( .A(n14323), .ZN(n13974) );
  INV_X1 U14189 ( .A(n14219), .ZN(n13948) );
  AOI22_X1 U14190 ( .A1(n13974), .A2(n11699), .B1(n11698), .B2(n13948), .ZN(
        n11700) );
  XNOR2_X1 U14191 ( .A(n11701), .B(n11700), .ZN(n11702) );
  XNOR2_X1 U14192 ( .A(n11703), .B(n11702), .ZN(n11712) );
  NAND2_X1 U14193 ( .A1(n6644), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14194 ( .A1(n11884), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11707) );
  INV_X1 U14195 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15495) );
  OR2_X1 U14196 ( .A1(n11881), .A2(n15495), .ZN(n11706) );
  OR2_X1 U14197 ( .A1(n11704), .A2(n13953), .ZN(n11705) );
  NAND4_X1 U14198 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n13821) );
  INV_X1 U14199 ( .A(n13821), .ZN(n11872) );
  INV_X1 U14200 ( .A(n14000), .ZN(n13805) );
  OAI22_X1 U14201 ( .A1(n11872), .A2(n14141), .B1(n13805), .B2(n14609), .ZN(
        n14224) );
  AOI22_X1 U14202 ( .A1(n13818), .A2(n14224), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11709) );
  OAI21_X1 U14203 ( .B1(n13967), .B2(n14588), .A(n11709), .ZN(n11710) );
  AOI21_X1 U14204 ( .B1(n13974), .B2(n13798), .A(n11710), .ZN(n11711) );
  OAI21_X1 U14205 ( .B1(n11712), .B2(n14574), .A(n11711), .ZN(P1_U3220) );
  NAND2_X1 U14206 ( .A1(n11883), .A2(n11714), .ZN(n11891) );
  XNOR2_X1 U14207 ( .A(n14376), .B(n13891), .ZN(n11715) );
  NAND2_X1 U14208 ( .A1(n11715), .A2(n11907), .ZN(n11716) );
  NAND2_X1 U14209 ( .A1(n11891), .A2(n11716), .ZN(n11737) );
  MUX2_X1 U14210 ( .A(n14219), .B(n14323), .S(n6808), .Z(n11867) );
  MUX2_X1 U14211 ( .A(n14021), .B(n14007), .S(n6808), .Z(n11857) );
  MUX2_X1 U14212 ( .A(n14337), .B(n13924), .S(n6808), .Z(n11841) );
  MUX2_X1 U14213 ( .A(n14342), .B(n14080), .S(n6808), .Z(n11833) );
  NAND2_X1 U14214 ( .A1(n11721), .A2(n11717), .ZN(n11718) );
  MUX2_X1 U14215 ( .A(n11721), .B(n11720), .S(n11737), .Z(n11722) );
  NAND2_X1 U14216 ( .A1(n11737), .A2(n11728), .ZN(n11726) );
  AND2_X1 U14217 ( .A1(n11726), .A2(n11725), .ZN(n11731) );
  MUX2_X1 U14218 ( .A(n11728), .B(n11727), .S(n11737), .Z(n11729) );
  OAI21_X1 U14219 ( .B1(n11732), .B2(n11731), .A(n11729), .ZN(n11734) );
  NAND3_X1 U14220 ( .A1(n11732), .A2(n11731), .A3(n11730), .ZN(n11733) );
  NAND3_X1 U14221 ( .A1(n11734), .A2(n11733), .A3(n11918), .ZN(n11742) );
  INV_X1 U14222 ( .A(n11735), .ZN(n11739) );
  INV_X1 U14223 ( .A(n11736), .ZN(n11738) );
  MUX2_X1 U14224 ( .A(n11739), .B(n11738), .S(n11737), .Z(n11740) );
  INV_X1 U14225 ( .A(n11740), .ZN(n11741) );
  NAND2_X1 U14226 ( .A1(n11742), .A2(n11741), .ZN(n11746) );
  MUX2_X1 U14227 ( .A(n13831), .B(n11743), .S(n11737), .Z(n11747) );
  NAND2_X1 U14228 ( .A1(n11746), .A2(n11747), .ZN(n11745) );
  MUX2_X1 U14229 ( .A(n11743), .B(n13831), .S(n11737), .Z(n11744) );
  INV_X1 U14230 ( .A(n11746), .ZN(n11749) );
  INV_X1 U14231 ( .A(n11747), .ZN(n11748) );
  NAND2_X1 U14232 ( .A1(n11749), .A2(n11748), .ZN(n11750) );
  MUX2_X1 U14233 ( .A(n11751), .B(n13830), .S(n11737), .Z(n11753) );
  MUX2_X1 U14234 ( .A(n13830), .B(n11751), .S(n11737), .Z(n11752) );
  MUX2_X1 U14235 ( .A(n13829), .B(n14712), .S(n6808), .Z(n11757) );
  NAND2_X1 U14236 ( .A1(n11756), .A2(n11757), .ZN(n11755) );
  MUX2_X1 U14237 ( .A(n14712), .B(n13829), .S(n6808), .Z(n11754) );
  NAND2_X1 U14238 ( .A1(n11755), .A2(n11754), .ZN(n11761) );
  INV_X1 U14239 ( .A(n11756), .ZN(n11759) );
  INV_X1 U14240 ( .A(n11757), .ZN(n11758) );
  NAND2_X1 U14241 ( .A1(n11759), .A2(n11758), .ZN(n11760) );
  MUX2_X1 U14242 ( .A(n13828), .B(n14715), .S(n11898), .Z(n11763) );
  MUX2_X1 U14243 ( .A(n14715), .B(n13828), .S(n11898), .Z(n11762) );
  INV_X1 U14244 ( .A(n11763), .ZN(n11764) );
  MUX2_X1 U14245 ( .A(n13827), .B(n11765), .S(n6808), .Z(n11769) );
  NAND2_X1 U14246 ( .A1(n11768), .A2(n11769), .ZN(n11767) );
  MUX2_X1 U14247 ( .A(n13827), .B(n11765), .S(n11898), .Z(n11766) );
  NAND2_X1 U14248 ( .A1(n11767), .A2(n11766), .ZN(n11773) );
  INV_X1 U14249 ( .A(n11768), .ZN(n11771) );
  INV_X1 U14250 ( .A(n11769), .ZN(n11770) );
  NAND2_X1 U14251 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  MUX2_X1 U14252 ( .A(n11775), .B(n11774), .S(n6808), .Z(n11777) );
  MUX2_X1 U14253 ( .A(n11775), .B(n11774), .S(n11898), .Z(n11776) );
  MUX2_X1 U14254 ( .A(n14576), .B(n11778), .S(n6808), .Z(n11782) );
  NAND2_X1 U14255 ( .A1(n11781), .A2(n11782), .ZN(n11780) );
  MUX2_X1 U14256 ( .A(n14576), .B(n11778), .S(n11898), .Z(n11779) );
  NAND2_X1 U14257 ( .A1(n11780), .A2(n11779), .ZN(n11786) );
  INV_X1 U14258 ( .A(n11781), .ZN(n11784) );
  INV_X1 U14259 ( .A(n11782), .ZN(n11783) );
  NAND2_X1 U14260 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  MUX2_X1 U14261 ( .A(n13825), .B(n11787), .S(n11898), .Z(n11789) );
  MUX2_X1 U14262 ( .A(n13825), .B(n11787), .S(n6808), .Z(n11788) );
  INV_X1 U14263 ( .A(n11789), .ZN(n11790) );
  MUX2_X1 U14264 ( .A(n13773), .B(n11791), .S(n6808), .Z(n11794) );
  MUX2_X1 U14265 ( .A(n11792), .B(n14578), .S(n6808), .Z(n11793) );
  INV_X1 U14266 ( .A(n11794), .ZN(n11795) );
  NOR2_X1 U14267 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  MUX2_X1 U14268 ( .A(n11798), .B(n14564), .S(n6808), .Z(n11799) );
  MUX2_X1 U14269 ( .A(n14564), .B(n11798), .S(n6808), .Z(n11800) );
  AOI21_X1 U14270 ( .B1(n11809), .B2(n11801), .A(n6808), .ZN(n11802) );
  AOI21_X1 U14271 ( .B1(n11803), .B2(n11915), .A(n11802), .ZN(n11808) );
  INV_X1 U14272 ( .A(n11804), .ZN(n11805) );
  OAI21_X1 U14273 ( .B1(n11807), .B2(n11805), .A(n6808), .ZN(n11806) );
  OAI21_X1 U14274 ( .B1(n11808), .B2(n11807), .A(n11806), .ZN(n11810) );
  NAND2_X1 U14275 ( .A1(n14158), .A2(n14173), .ZN(n13913) );
  OR2_X1 U14276 ( .A1(n14158), .A2(n14173), .ZN(n13914) );
  INV_X1 U14277 ( .A(n13912), .ZN(n14159) );
  MUX2_X1 U14278 ( .A(n14159), .B(n14300), .S(n6808), .Z(n11818) );
  INV_X1 U14279 ( .A(n11818), .ZN(n11812) );
  MUX2_X1 U14280 ( .A(n14181), .B(n13912), .S(n6808), .Z(n11819) );
  NAND2_X1 U14281 ( .A1(n11812), .A2(n11811), .ZN(n11813) );
  INV_X1 U14282 ( .A(n14158), .ZN(n14292) );
  NAND4_X1 U14283 ( .A1(n11914), .A2(n11898), .A3(n14292), .A4(n14173), .ZN(
        n11815) );
  OAI21_X1 U14284 ( .B1(n11898), .B2(n11914), .A(n11815), .ZN(n11817) );
  NOR4_X1 U14285 ( .A1(n11913), .A2(n11898), .A3(n14292), .A4(n14173), .ZN(
        n11816) );
  AOI211_X1 U14286 ( .C1(n11913), .C2(n11898), .A(n11817), .B(n11816), .ZN(
        n11823) );
  NAND3_X1 U14287 ( .A1(n11820), .A2(n11819), .A3(n11818), .ZN(n11822) );
  NAND2_X1 U14288 ( .A1(n14133), .A2(n13823), .ZN(n11821) );
  NAND2_X1 U14289 ( .A1(n13917), .A2(n11821), .ZN(n13941) );
  MUX2_X1 U14290 ( .A(n13823), .B(n14133), .S(n6808), .Z(n11824) );
  INV_X1 U14291 ( .A(n11824), .ZN(n11825) );
  MUX2_X1 U14292 ( .A(n14272), .B(n13920), .S(n6808), .Z(n11827) );
  INV_X1 U14293 ( .A(n13920), .ZN(n14088) );
  INV_X1 U14294 ( .A(n14272), .ZN(n11912) );
  MUX2_X1 U14295 ( .A(n14088), .B(n11912), .S(n6808), .Z(n11826) );
  NAND2_X1 U14296 ( .A1(n11827), .A2(n11826), .ZN(n11830) );
  INV_X1 U14297 ( .A(n11826), .ZN(n11829) );
  INV_X1 U14298 ( .A(n11827), .ZN(n11828) );
  MUX2_X1 U14299 ( .A(n14261), .B(n14100), .S(n6808), .Z(n11832) );
  MUX2_X1 U14300 ( .A(n14087), .B(n14263), .S(n6808), .Z(n11838) );
  MUX2_X1 U14301 ( .A(n13791), .B(n13945), .S(n6808), .Z(n11836) );
  INV_X1 U14302 ( .A(n11838), .ZN(n11839) );
  INV_X1 U14303 ( .A(n13924), .ZN(n14076) );
  MUX2_X1 U14304 ( .A(n14076), .B(n13700), .S(n6808), .Z(n11840) );
  MUX2_X1 U14305 ( .A(n14020), .B(n14045), .S(n6808), .Z(n11843) );
  MUX2_X1 U14306 ( .A(n14045), .B(n14020), .S(n6808), .Z(n11846) );
  INV_X1 U14307 ( .A(n11843), .ZN(n11844) );
  MUX2_X1 U14308 ( .A(n14030), .B(n13999), .S(n6808), .Z(n11851) );
  NAND2_X1 U14309 ( .A1(n11848), .A2(n11851), .ZN(n11850) );
  MUX2_X1 U14310 ( .A(n13999), .B(n14030), .S(n6808), .Z(n11849) );
  NAND2_X1 U14311 ( .A1(n11850), .A2(n11849), .ZN(n11855) );
  INV_X1 U14312 ( .A(n11851), .ZN(n11852) );
  NAND2_X1 U14313 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  INV_X2 U14314 ( .A(n14007), .ZN(n14236) );
  INV_X1 U14315 ( .A(n14021), .ZN(n13822) );
  MUX2_X1 U14316 ( .A(n14236), .B(n13822), .S(n6808), .Z(n11856) );
  MUX2_X1 U14317 ( .A(n13991), .B(n14000), .S(n6808), .Z(n11861) );
  NAND2_X1 U14318 ( .A1(n11860), .A2(n11861), .ZN(n11865) );
  MUX2_X1 U14319 ( .A(n14000), .B(n13991), .S(n6808), .Z(n11864) );
  INV_X1 U14320 ( .A(n11861), .ZN(n11862) );
  MUX2_X1 U14321 ( .A(n13974), .B(n13948), .S(n6808), .Z(n11866) );
  OAI21_X1 U14322 ( .B1(n11868), .B2(n11867), .A(n11866), .ZN(n11869) );
  NAND2_X1 U14323 ( .A1(n13672), .A2(n11897), .ZN(n11871) );
  OR2_X1 U14324 ( .A1(n8839), .A2(n14366), .ZN(n11870) );
  MUX2_X1 U14325 ( .A(n13961), .B(n13821), .S(n6808), .Z(n11874) );
  MUX2_X1 U14326 ( .A(n11872), .B(n14321), .S(n6808), .Z(n11873) );
  NAND2_X1 U14327 ( .A1(n13669), .A2(n11897), .ZN(n11877) );
  INV_X1 U14328 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14364) );
  OR2_X1 U14329 ( .A1(n8839), .A2(n14364), .ZN(n11876) );
  INV_X1 U14330 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U14331 ( .A1(n11884), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U14332 ( .A1(n6645), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11879) );
  OAI211_X1 U14333 ( .C1(n11881), .C2(n15450), .A(n11880), .B(n11879), .ZN(
        n13900) );
  INV_X1 U14334 ( .A(n13900), .ZN(n11882) );
  NOR2_X1 U14335 ( .A1(n6808), .A2(n11882), .ZN(n11899) );
  INV_X1 U14336 ( .A(n11883), .ZN(n11889) );
  INV_X1 U14337 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U14338 ( .A1(n11884), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11887) );
  NAND2_X1 U14339 ( .A1(n11885), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11886) );
  OAI211_X1 U14340 ( .C1(n11888), .C2(n14316), .A(n11887), .B(n11886), .ZN(
        n13951) );
  OAI21_X1 U14341 ( .B1(n11899), .B2(n11889), .A(n13951), .ZN(n11890) );
  OAI21_X1 U14342 ( .B1(n14318), .B2(n11898), .A(n11890), .ZN(n11894) );
  INV_X1 U14343 ( .A(n11891), .ZN(n11892) );
  OAI21_X1 U14344 ( .B1(n11892), .B2(n13900), .A(n13951), .ZN(n11893) );
  MUX2_X1 U14345 ( .A(n14318), .B(n11893), .S(n6808), .Z(n11895) );
  NAND2_X1 U14346 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  INV_X1 U14347 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14358) );
  INV_X1 U14348 ( .A(n14314), .ZN(n13901) );
  INV_X1 U14349 ( .A(n11899), .ZN(n11900) );
  NAND2_X1 U14350 ( .A1(n11901), .A2(n14677), .ZN(n11906) );
  NAND2_X1 U14351 ( .A1(n8275), .A2(n11902), .ZN(n11903) );
  NAND2_X1 U14352 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  AND2_X1 U14353 ( .A1(n11906), .A2(n11905), .ZN(n11946) );
  INV_X1 U14354 ( .A(n11946), .ZN(n11909) );
  NAND2_X1 U14355 ( .A1(n11908), .A2(n11907), .ZN(n11941) );
  NAND2_X1 U14356 ( .A1(n11909), .A2(n11941), .ZN(n11942) );
  INV_X1 U14357 ( .A(n11942), .ZN(n11910) );
  NAND2_X1 U14358 ( .A1(n11944), .A2(n11910), .ZN(n11952) );
  XNOR2_X1 U14359 ( .A(n13991), .B(n13805), .ZN(n13983) );
  XNOR2_X1 U14360 ( .A(n13974), .B(n14219), .ZN(n13933) );
  XNOR2_X2 U14361 ( .A(n14236), .B(n13822), .ZN(n13996) );
  XNOR2_X1 U14362 ( .A(n13700), .B(n13924), .ZN(n13923) );
  XNOR2_X1 U14363 ( .A(n13791), .B(n14087), .ZN(n14070) );
  NAND2_X1 U14364 ( .A1(n14100), .A2(n14261), .ZN(n11911) );
  XNOR2_X1 U14365 ( .A(n11912), .B(n13920), .ZN(n13919) );
  NAND2_X1 U14366 ( .A1(n13940), .A2(n11914), .ZN(n14149) );
  XNOR2_X1 U14367 ( .A(n14300), .B(n13912), .ZN(n14184) );
  AND4_X1 U14368 ( .A1(n11918), .A2(n11917), .A3(n14193), .A4(n11916), .ZN(
        n11921) );
  NAND4_X1 U14369 ( .A1(n11922), .A2(n11921), .A3(n11920), .A4(n11919), .ZN(
        n11923) );
  OR3_X1 U14370 ( .A1(n11925), .A2(n11924), .A3(n11923), .ZN(n11926) );
  NOR2_X1 U14371 ( .A1(n11927), .A2(n11926), .ZN(n11929) );
  NAND4_X1 U14372 ( .A1(n11930), .A2(n11929), .A3(n7600), .A4(n11928), .ZN(
        n11931) );
  OR4_X1 U14373 ( .A1(n14603), .A2(n14502), .A3(n14184), .A4(n11931), .ZN(
        n11932) );
  NOR2_X1 U14374 ( .A1(n14149), .A2(n11932), .ZN(n11933) );
  XNOR2_X1 U14375 ( .A(n14158), .B(n14173), .ZN(n14156) );
  NAND4_X1 U14376 ( .A1(n13941), .A2(n11933), .A3(n13934), .A4(n14156), .ZN(
        n11934) );
  OR4_X1 U14377 ( .A1(n14070), .A2(n14090), .A3(n13919), .A4(n11934), .ZN(
        n11935) );
  NOR2_X1 U14378 ( .A1(n13923), .A2(n11935), .ZN(n11936) );
  XNOR2_X1 U14379 ( .A(n14030), .B(n13999), .ZN(n14018) );
  XNOR2_X1 U14380 ( .A(n14045), .B(n14020), .ZN(n13947) );
  NAND4_X1 U14381 ( .A1(n13996), .A2(n11936), .A3(n14018), .A4(n13947), .ZN(
        n11937) );
  XNOR2_X1 U14382 ( .A(n7129), .B(n13951), .ZN(n11938) );
  XNOR2_X1 U14383 ( .A(n13961), .B(n13821), .ZN(n13950) );
  NAND3_X1 U14384 ( .A1(n11939), .A2(n11938), .A3(n13950), .ZN(n11940) );
  XNOR2_X1 U14385 ( .A(n11940), .B(n14677), .ZN(n11949) );
  INV_X1 U14386 ( .A(n11941), .ZN(n11948) );
  NOR2_X1 U14387 ( .A1(n11943), .A2(n11942), .ZN(n11945) );
  MUX2_X1 U14388 ( .A(n11946), .B(n11945), .S(n11944), .Z(n11947) );
  OAI211_X1 U14389 ( .C1(n11953), .C2(n11952), .A(n11951), .B(n11950), .ZN(
        n11955) );
  NAND2_X1 U14390 ( .A1(n11955), .A2(n11954), .ZN(n11961) );
  NAND3_X1 U14391 ( .A1(n11957), .A2(n11956), .A3(n14262), .ZN(n11958) );
  OAI211_X1 U14392 ( .C1(n14376), .C2(n11959), .A(n11958), .B(P1_B_REG_SCAN_IN), .ZN(n11960) );
  NAND2_X1 U14393 ( .A1(n11961), .A2(n11960), .ZN(P1_U3242) );
  NAND2_X1 U14394 ( .A1(n14368), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11964) );
  AND2_X1 U14395 ( .A1(n11966), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U14396 ( .A1(n12066), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11968) );
  XNOR2_X1 U14397 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12216) );
  XNOR2_X1 U14398 ( .A(n12218), .B(n12216), .ZN(n12991) );
  NAND2_X1 U14399 ( .A1(n12991), .A2(n12235), .ZN(n11970) );
  NAND2_X1 U14400 ( .A1(n12069), .A2(SI_29_), .ZN(n11969) );
  NAND2_X1 U14401 ( .A1(n11972), .A2(n12636), .ZN(n12410) );
  NAND2_X1 U14402 ( .A1(n12977), .A2(n11974), .ZN(n12345) );
  NAND2_X1 U14403 ( .A1(n12344), .A2(n12345), .ZN(n12833) );
  OR2_X1 U14404 ( .A1(n12077), .A2(n12836), .ZN(n12348) );
  NAND2_X1 U14405 ( .A1(n12077), .A2(n12836), .ZN(n12354) );
  NAND2_X1 U14406 ( .A1(n12348), .A2(n12354), .ZN(n12821) );
  NAND2_X1 U14407 ( .A1(n12827), .A2(n12826), .ZN(n11975) );
  NAND2_X1 U14408 ( .A1(n11975), .A2(n12354), .ZN(n12810) );
  OR2_X1 U14409 ( .A1(n12906), .A2(n12825), .ZN(n12356) );
  NAND2_X1 U14410 ( .A1(n12906), .A2(n12825), .ZN(n12355) );
  NAND2_X1 U14411 ( .A1(n12356), .A2(n12355), .ZN(n12086) );
  OR2_X1 U14412 ( .A1(n12902), .A2(n12779), .ZN(n12363) );
  NAND2_X1 U14413 ( .A1(n12902), .A2(n12779), .ZN(n12360) );
  NAND2_X1 U14414 ( .A1(n12363), .A2(n12360), .ZN(n12260) );
  NAND2_X1 U14415 ( .A1(n12791), .A2(n12091), .ZN(n12364) );
  NAND2_X1 U14416 ( .A1(n11976), .A2(n12235), .ZN(n11979) );
  AOI22_X1 U14417 ( .A1(n12069), .A2(n11977), .B1(n10875), .B2(n12601), .ZN(
        n11978) );
  NAND2_X1 U14418 ( .A1(n12963), .A2(n12440), .ZN(n12371) );
  OR2_X1 U14419 ( .A1(n12963), .A2(n12440), .ZN(n12370) );
  NAND2_X1 U14420 ( .A1(n11981), .A2(n12235), .ZN(n11983) );
  NAND2_X1 U14421 ( .A1(n12069), .A2(SI_20_), .ZN(n11982) );
  XNOR2_X1 U14422 ( .A(n12753), .B(n12741), .ZN(n12754) );
  OR2_X1 U14423 ( .A1(n12753), .A2(n12741), .ZN(n12375) );
  NAND2_X1 U14424 ( .A1(n12069), .A2(SI_21_), .ZN(n11986) );
  NAND2_X1 U14425 ( .A1(n11988), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U14426 ( .A1(n11999), .A2(n11989), .ZN(n12745) );
  NAND2_X1 U14427 ( .A1(n12745), .A2(n12024), .ZN(n11995) );
  INV_X1 U14428 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U14429 ( .A1(n12222), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U14430 ( .A1(n6639), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n11990) );
  OAI211_X1 U14431 ( .C1(n12062), .C2(n11992), .A(n11991), .B(n11990), .ZN(
        n11993) );
  INV_X1 U14432 ( .A(n11993), .ZN(n11994) );
  NAND2_X1 U14433 ( .A1(n11995), .A2(n11994), .ZN(n12439) );
  NAND2_X1 U14434 ( .A1(n12164), .A2(n12752), .ZN(n12380) );
  OR2_X1 U14435 ( .A1(n12164), .A2(n12752), .ZN(n12379) );
  NAND2_X1 U14436 ( .A1(n11996), .A2(n12235), .ZN(n11998) );
  NAND2_X1 U14437 ( .A1(n12069), .A2(SI_22_), .ZN(n11997) );
  NAND2_X1 U14438 ( .A1(n11999), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n12000) );
  NAND2_X1 U14439 ( .A1(n12011), .A2(n12000), .ZN(n12734) );
  NAND2_X1 U14440 ( .A1(n12734), .A2(n12024), .ZN(n12006) );
  INV_X1 U14441 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U14442 ( .A1(n6639), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n12002) );
  NAND2_X1 U14443 ( .A1(n12222), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n12001) );
  OAI211_X1 U14444 ( .C1(n12003), .C2(n12062), .A(n12002), .B(n12001), .ZN(
        n12004) );
  INV_X1 U14445 ( .A(n12004), .ZN(n12005) );
  NAND2_X1 U14446 ( .A1(n12006), .A2(n12005), .ZN(n12714) );
  NAND2_X1 U14447 ( .A1(n12733), .A2(n12742), .ZN(n12383) );
  NAND2_X1 U14448 ( .A1(n12731), .A2(n12383), .ZN(n12007) );
  NAND2_X1 U14449 ( .A1(n12007), .A2(n12382), .ZN(n12711) );
  NAND2_X1 U14450 ( .A1(n12008), .A2(n12235), .ZN(n12010) );
  NAND2_X1 U14451 ( .A1(n12069), .A2(SI_23_), .ZN(n12009) );
  NAND2_X1 U14452 ( .A1(n12011), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U14453 ( .A1(n12022), .A2(n12012), .ZN(n12719) );
  NAND2_X1 U14454 ( .A1(n12719), .A2(n12024), .ZN(n12017) );
  INV_X1 U14455 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12721) );
  NAND2_X1 U14456 ( .A1(n6639), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U14457 ( .A1(n12222), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n12013) );
  OAI211_X1 U14458 ( .C1(n12721), .C2(n12062), .A(n12014), .B(n12013), .ZN(
        n12015) );
  INV_X1 U14459 ( .A(n12015), .ZN(n12016) );
  NAND2_X1 U14460 ( .A1(n12945), .A2(n12730), .ZN(n12018) );
  NAND2_X1 U14461 ( .A1(n12392), .A2(n12018), .ZN(n12097) );
  NAND2_X1 U14462 ( .A1(n12019), .A2(n12235), .ZN(n12021) );
  NAND2_X1 U14463 ( .A1(n12069), .A2(SI_24_), .ZN(n12020) );
  NAND2_X1 U14464 ( .A1(n12022), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n12023) );
  NAND2_X1 U14465 ( .A1(n12034), .A2(n12023), .ZN(n12701) );
  NAND2_X1 U14466 ( .A1(n12701), .A2(n12024), .ZN(n12030) );
  INV_X1 U14467 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U14468 ( .A1(n6639), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U14469 ( .A1(n12222), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U14470 ( .C1(n12027), .C2(n12062), .A(n12026), .B(n12025), .ZN(
        n12028) );
  INV_X1 U14471 ( .A(n12028), .ZN(n12029) );
  NAND2_X1 U14472 ( .A1(n12030), .A2(n12029), .ZN(n12715) );
  OR2_X1 U14473 ( .A1(n12700), .A2(n12679), .ZN(n12391) );
  NAND2_X1 U14474 ( .A1(n12700), .A2(n12679), .ZN(n12390) );
  NAND2_X1 U14475 ( .A1(n12391), .A2(n12390), .ZN(n12693) );
  NAND2_X1 U14476 ( .A1(n12031), .A2(n12235), .ZN(n12033) );
  NAND2_X1 U14477 ( .A1(n12069), .A2(SI_25_), .ZN(n12032) );
  NAND2_X1 U14478 ( .A1(n12034), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n12035) );
  NAND2_X1 U14479 ( .A1(n12045), .A2(n12035), .ZN(n12687) );
  NAND2_X1 U14480 ( .A1(n12687), .A2(n12024), .ZN(n12041) );
  INV_X1 U14481 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12038) );
  NAND2_X1 U14482 ( .A1(n6639), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n12037) );
  NAND2_X1 U14483 ( .A1(n12222), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n12036) );
  OAI211_X1 U14484 ( .C1(n12038), .C2(n12062), .A(n12037), .B(n12036), .ZN(
        n12039) );
  INV_X1 U14485 ( .A(n12039), .ZN(n12040) );
  OR2_X1 U14486 ( .A1(n12866), .A2(n12695), .ZN(n12398) );
  NAND2_X1 U14487 ( .A1(n12866), .A2(n12695), .ZN(n12399) );
  NAND2_X1 U14488 ( .A1(n12042), .A2(n12235), .ZN(n12044) );
  NAND2_X1 U14489 ( .A1(n12069), .A2(SI_26_), .ZN(n12043) );
  NAND2_X1 U14490 ( .A1(n12045), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U14491 ( .A1(n12056), .A2(n12046), .ZN(n12671) );
  NAND2_X1 U14492 ( .A1(n12671), .A2(n12024), .ZN(n12051) );
  INV_X1 U14493 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U14494 ( .A1(n12222), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U14495 ( .A1(n6639), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n12047) );
  OAI211_X1 U14496 ( .C1(n12062), .C2(n12673), .A(n12048), .B(n12047), .ZN(
        n12049) );
  INV_X1 U14497 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U14498 ( .A1(n12051), .A2(n12050), .ZN(n12436) );
  NAND2_X1 U14499 ( .A1(n12664), .A2(n12402), .ZN(n12052) );
  NAND2_X1 U14500 ( .A1(n12861), .A2(n12680), .ZN(n12403) );
  NAND2_X1 U14501 ( .A1(n12053), .A2(n12235), .ZN(n12055) );
  NAND2_X1 U14502 ( .A1(n12069), .A2(SI_27_), .ZN(n12054) );
  NAND2_X1 U14503 ( .A1(n12056), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U14504 ( .A1(n12058), .A2(n12057), .ZN(n12658) );
  NAND2_X1 U14505 ( .A1(n12658), .A2(n12024), .ZN(n12065) );
  INV_X1 U14506 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12061) );
  NAND2_X1 U14507 ( .A1(n12222), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U14508 ( .A1(n6639), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n12059) );
  OAI211_X1 U14509 ( .C1(n12062), .C2(n12061), .A(n12060), .B(n12059), .ZN(
        n12063) );
  INV_X1 U14510 ( .A(n12063), .ZN(n12064) );
  NAND2_X1 U14511 ( .A1(n12657), .A2(n12667), .ZN(n12640) );
  XNOR2_X1 U14512 ( .A(n12066), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n12067) );
  XNOR2_X1 U14513 ( .A(n12068), .B(n12067), .ZN(n12995) );
  NAND2_X1 U14514 ( .A1(n12995), .A2(n12235), .ZN(n12071) );
  NAND2_X1 U14515 ( .A1(n12069), .A2(SI_28_), .ZN(n12070) );
  NAND2_X1 U14516 ( .A1(n12161), .A2(n12653), .ZN(n12106) );
  INV_X1 U14517 ( .A(n12106), .ZN(n12073) );
  INV_X1 U14518 ( .A(n12640), .ZN(n12072) );
  NOR2_X1 U14519 ( .A1(n12073), .A2(n12072), .ZN(n12408) );
  INV_X1 U14520 ( .A(n12107), .ZN(n12407) );
  OR2_X1 U14521 ( .A1(n12076), .A2(n12441), .ZN(n12074) );
  NAND2_X1 U14522 ( .A1(n12075), .A2(n12074), .ZN(n12818) );
  NAND2_X1 U14523 ( .A1(n12076), .A2(n12441), .ZN(n12817) );
  OR2_X1 U14524 ( .A1(n12977), .A2(n12824), .ZN(n12819) );
  NAND2_X1 U14525 ( .A1(n12077), .A2(n12806), .ZN(n12078) );
  AND2_X1 U14526 ( .A1(n12819), .A2(n12078), .ZN(n12080) );
  AND2_X1 U14527 ( .A1(n12817), .A2(n12080), .ZN(n12085) );
  INV_X1 U14528 ( .A(n12078), .ZN(n12079) );
  OR2_X1 U14529 ( .A1(n12079), .A2(n12821), .ZN(n12083) );
  INV_X1 U14530 ( .A(n12080), .ZN(n12081) );
  OR2_X1 U14531 ( .A1(n12081), .A2(n12833), .ZN(n12082) );
  NAND2_X1 U14532 ( .A1(n12805), .A2(n12086), .ZN(n12088) );
  NAND2_X1 U14533 ( .A1(n12906), .A2(n6815), .ZN(n12087) );
  NAND2_X1 U14534 ( .A1(n12795), .A2(n12260), .ZN(n12090) );
  INV_X1 U14535 ( .A(n12779), .ZN(n12807) );
  NAND2_X1 U14536 ( .A1(n12902), .A2(n12807), .ZN(n12089) );
  OR2_X1 U14537 ( .A1(n12791), .A2(n12796), .ZN(n12092) );
  INV_X1 U14538 ( .A(n12440), .ZN(n12780) );
  OR2_X1 U14539 ( .A1(n12963), .A2(n12780), .ZN(n12093) );
  NAND2_X1 U14540 ( .A1(n12753), .A2(n12764), .ZN(n12094) );
  OR2_X1 U14541 ( .A1(n12164), .A2(n12439), .ZN(n12726) );
  AND2_X1 U14542 ( .A1(n7650), .A2(n12726), .ZN(n12095) );
  NAND2_X1 U14543 ( .A1(n12727), .A2(n12095), .ZN(n12708) );
  NAND2_X1 U14544 ( .A1(n12733), .A2(n12714), .ZN(n12707) );
  NAND2_X1 U14545 ( .A1(n12945), .A2(n12438), .ZN(n12096) );
  AND2_X1 U14546 ( .A1(n12707), .A2(n12096), .ZN(n12099) );
  INV_X1 U14547 ( .A(n12096), .ZN(n12098) );
  AND2_X1 U14548 ( .A1(n12700), .A2(n12715), .ZN(n12100) );
  OAI22_X1 U14549 ( .A1(n12692), .A2(n12100), .B1(n12715), .B2(n12700), .ZN(
        n12683) );
  NAND2_X1 U14550 ( .A1(n12866), .A2(n12437), .ZN(n12101) );
  OR2_X1 U14551 ( .A1(n12436), .A2(n12861), .ZN(n12102) );
  NAND2_X1 U14552 ( .A1(n12861), .A2(n12436), .ZN(n12103) );
  OR2_X1 U14553 ( .A1(n12657), .A2(n12435), .ZN(n12105) );
  XNOR2_X1 U14554 ( .A(n12108), .B(n12266), .ZN(n12114) );
  NAND2_X1 U14555 ( .A1(n12109), .A2(P3_B_REG_SCAN_IN), .ZN(n12110) );
  NAND2_X1 U14556 ( .A1(n15149), .A2(n12110), .ZN(n12618) );
  NOR2_X1 U14557 ( .A1(n12241), .A2(n12618), .ZN(n12112) );
  NOR2_X1 U14558 ( .A1(n12653), .A2(n15130), .ZN(n12111) );
  OAI21_X1 U14559 ( .B1(n12627), .B2(n12918), .A(n12115), .ZN(P3_U3488) );
  OAI21_X1 U14560 ( .B1(n12627), .B2(n12978), .A(n12116), .ZN(P3_U3456) );
  XNOR2_X1 U14561 ( .A(n6832), .B(n12117), .ZN(n12152) );
  XNOR2_X1 U14562 ( .A(n12152), .B(n12435), .ZN(n12153) );
  XNOR2_X1 U14563 ( .A(n12733), .B(n12117), .ZN(n12125) );
  XNOR2_X1 U14564 ( .A(n12164), .B(n12117), .ZN(n12123) );
  XNOR2_X1 U14565 ( .A(n12753), .B(n12117), .ZN(n12122) );
  XNOR2_X1 U14566 ( .A(n12963), .B(n12155), .ZN(n12120) );
  INV_X1 U14567 ( .A(n12120), .ZN(n12121) );
  XNOR2_X1 U14568 ( .A(n12120), .B(n12780), .ZN(n12145) );
  XNOR2_X1 U14569 ( .A(n12122), .B(n12764), .ZN(n12194) );
  XNOR2_X1 U14570 ( .A(n12123), .B(n12752), .ZN(n12166) );
  INV_X1 U14571 ( .A(n12124), .ZN(n12126) );
  XNOR2_X1 U14572 ( .A(n12700), .B(n12155), .ZN(n12128) );
  XNOR2_X1 U14573 ( .A(n12128), .B(n12679), .ZN(n12183) );
  INV_X1 U14574 ( .A(n12128), .ZN(n12129) );
  XNOR2_X1 U14575 ( .A(n12866), .B(n12155), .ZN(n12130) );
  XNOR2_X1 U14576 ( .A(n12130), .B(n12437), .ZN(n12176) );
  XNOR2_X1 U14577 ( .A(n12861), .B(n12155), .ZN(n12131) );
  XNOR2_X1 U14578 ( .A(n12131), .B(n12680), .ZN(n12206) );
  INV_X1 U14579 ( .A(n12131), .ZN(n12132) );
  XOR2_X1 U14580 ( .A(n12153), .B(n12154), .Z(n12137) );
  NOR2_X1 U14581 ( .A1(n12653), .A2(n12202), .ZN(n12135) );
  AOI22_X1 U14582 ( .A1(n12658), .A2(n12207), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12133) );
  OAI21_X1 U14583 ( .B1(n12680), .B2(n12209), .A(n12133), .ZN(n12134) );
  AOI211_X1 U14584 ( .C1(n12657), .C2(n12212), .A(n12135), .B(n12134), .ZN(
        n12136) );
  OAI21_X1 U14585 ( .B1(n12137), .B2(n12214), .A(n12136), .ZN(P3_U3154) );
  XNOR2_X1 U14586 ( .A(n12138), .B(n12730), .ZN(n12143) );
  AOI22_X1 U14587 ( .A1(n12714), .A2(n12199), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12140) );
  NAND2_X1 U14588 ( .A1(n12719), .A2(n12207), .ZN(n12139) );
  OAI211_X1 U14589 ( .C1(n12679), .C2(n12202), .A(n12140), .B(n12139), .ZN(
        n12141) );
  AOI21_X1 U14590 ( .B1(n12945), .B2(n12212), .A(n12141), .ZN(n12142) );
  OAI21_X1 U14591 ( .B1(n12143), .B2(n12214), .A(n12142), .ZN(P3_U3156) );
  AOI211_X1 U14592 ( .C1(n12146), .C2(n12145), .A(n12214), .B(n12144), .ZN(
        n12147) );
  INV_X1 U14593 ( .A(n12147), .ZN(n12151) );
  NAND2_X1 U14594 ( .A1(n12796), .A2(n12199), .ZN(n12148) );
  NAND2_X1 U14595 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12610)
         );
  OAI211_X1 U14596 ( .C1(n12741), .C2(n12202), .A(n12148), .B(n12610), .ZN(
        n12149) );
  AOI21_X1 U14597 ( .B1(n12769), .B2(n12207), .A(n12149), .ZN(n12150) );
  OAI211_X1 U14598 ( .C1(n12174), .C2(n12963), .A(n12151), .B(n12150), .ZN(
        P3_U3159) );
  XNOR2_X1 U14599 ( .A(n12641), .B(n12155), .ZN(n12156) );
  XNOR2_X1 U14600 ( .A(n12157), .B(n12156), .ZN(n12163) );
  NOR2_X1 U14601 ( .A1(n12636), .A2(n12202), .ZN(n12160) );
  AOI22_X1 U14602 ( .A1(n12643), .A2(n12207), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12158) );
  OAI21_X1 U14603 ( .B1(n12667), .B2(n12209), .A(n12158), .ZN(n12159) );
  AOI211_X1 U14604 ( .C1(n12161), .C2(n12212), .A(n12160), .B(n12159), .ZN(
        n12162) );
  OAI21_X1 U14605 ( .B1(n12163), .B2(n12214), .A(n12162), .ZN(P3_U3160) );
  INV_X1 U14606 ( .A(n12164), .ZN(n12955) );
  OAI21_X1 U14607 ( .B1(n12167), .B2(n12166), .A(n12165), .ZN(n12169) );
  NAND2_X1 U14608 ( .A1(n12169), .A2(n12168), .ZN(n12173) );
  AOI22_X1 U14609 ( .A1(n12764), .A2(n12199), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12170) );
  OAI21_X1 U14610 ( .B1(n12742), .B2(n12202), .A(n12170), .ZN(n12171) );
  AOI21_X1 U14611 ( .B1(n12745), .B2(n12207), .A(n12171), .ZN(n12172) );
  OAI211_X1 U14612 ( .C1(n12955), .C2(n12174), .A(n12173), .B(n12172), .ZN(
        P3_U3163) );
  XOR2_X1 U14613 ( .A(n12176), .B(n12175), .Z(n12181) );
  AOI22_X1 U14614 ( .A1(n12715), .A2(n12199), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12178) );
  NAND2_X1 U14615 ( .A1(n12687), .A2(n12207), .ZN(n12177) );
  OAI211_X1 U14616 ( .C1(n12680), .C2(n12202), .A(n12178), .B(n12177), .ZN(
        n12179) );
  AOI21_X1 U14617 ( .B1(n12866), .B2(n12212), .A(n12179), .ZN(n12180) );
  OAI21_X1 U14618 ( .B1(n12181), .B2(n12214), .A(n12180), .ZN(P3_U3165) );
  XOR2_X1 U14619 ( .A(n12183), .B(n12182), .Z(n12188) );
  AOI22_X1 U14620 ( .A1(n12438), .A2(n12199), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12185) );
  NAND2_X1 U14621 ( .A1(n12701), .A2(n12207), .ZN(n12184) );
  OAI211_X1 U14622 ( .C1(n12695), .C2(n12202), .A(n12185), .B(n12184), .ZN(
        n12186) );
  AOI21_X1 U14623 ( .B1(n12700), .B2(n12212), .A(n12186), .ZN(n12187) );
  OAI21_X1 U14624 ( .B1(n12188), .B2(n12214), .A(n12187), .ZN(P3_U3169) );
  AOI22_X1 U14625 ( .A1(n12439), .A2(n12189), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12191) );
  NAND2_X1 U14626 ( .A1(n12207), .A2(n12758), .ZN(n12190) );
  OAI211_X1 U14627 ( .C1(n12780), .C2(n12209), .A(n12191), .B(n12190), .ZN(
        n12196) );
  AOI211_X1 U14628 ( .C1(n12194), .C2(n12193), .A(n12214), .B(n12192), .ZN(
        n12195) );
  AOI211_X1 U14629 ( .C1(n12212), .C2(n12753), .A(n12196), .B(n12195), .ZN(
        n12197) );
  INV_X1 U14630 ( .A(n12197), .ZN(P3_U3173) );
  XNOR2_X1 U14631 ( .A(n12198), .B(n12742), .ZN(n12205) );
  AOI22_X1 U14632 ( .A1(n12439), .A2(n12199), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12201) );
  NAND2_X1 U14633 ( .A1(n12734), .A2(n12207), .ZN(n12200) );
  OAI211_X1 U14634 ( .C1(n12730), .C2(n12202), .A(n12201), .B(n12200), .ZN(
        n12203) );
  AOI21_X1 U14635 ( .B1(n12733), .B2(n12212), .A(n12203), .ZN(n12204) );
  OAI21_X1 U14636 ( .B1(n12205), .B2(n12214), .A(n12204), .ZN(P3_U3175) );
  NOR2_X1 U14637 ( .A1(n12667), .A2(n12202), .ZN(n12211) );
  AOI22_X1 U14638 ( .A1(n12671), .A2(n12207), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12208) );
  OAI21_X1 U14639 ( .B1(n12695), .B2(n12209), .A(n12208), .ZN(n12210) );
  AOI211_X1 U14640 ( .C1(n12861), .C2(n12212), .A(n12211), .B(n12210), .ZN(
        n12213) );
  OAI21_X1 U14641 ( .B1(n12215), .B2(n12214), .A(n12213), .ZN(P3_U3180) );
  INV_X1 U14642 ( .A(n12216), .ZN(n12217) );
  NAND2_X1 U14643 ( .A1(n14366), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12219) );
  INV_X1 U14644 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13671) );
  XNOR2_X1 U14645 ( .A(n13671), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12231) );
  XNOR2_X1 U14646 ( .A(n12232), .B(n12231), .ZN(n12987) );
  NAND2_X1 U14647 ( .A1(n12987), .A2(n12235), .ZN(n12221) );
  OR2_X1 U14648 ( .A1(n12236), .A2(n12989), .ZN(n12220) );
  INV_X1 U14649 ( .A(n12922), .ZN(n12851) );
  NAND2_X1 U14650 ( .A1(n12222), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U14651 ( .A1(n6638), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U14652 ( .A1(n6639), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12224) );
  AND3_X1 U14653 ( .A1(n12226), .A2(n12225), .A3(n12224), .ZN(n12227) );
  INV_X1 U14654 ( .A(n12619), .ZN(n12434) );
  NAND2_X1 U14655 ( .A1(n12229), .A2(n12413), .ZN(n12230) );
  OAI211_X1 U14656 ( .C1(n12851), .C2(n12434), .A(n12230), .B(n12410), .ZN(
        n12243) );
  XNOR2_X1 U14657 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12233) );
  XNOR2_X1 U14658 ( .A(n12234), .B(n12233), .ZN(n12980) );
  NAND2_X1 U14659 ( .A1(n12980), .A2(n12235), .ZN(n12238) );
  OR2_X1 U14660 ( .A1(n12236), .A2(n12986), .ZN(n12237) );
  NAND2_X1 U14661 ( .A1(n12922), .A2(n12241), .ZN(n12239) );
  NAND2_X1 U14662 ( .A1(n12240), .A2(n12619), .ZN(n12416) );
  OR2_X1 U14663 ( .A1(n12922), .A2(n12241), .ZN(n12242) );
  NAND2_X1 U14664 ( .A1(n12416), .A2(n12242), .ZN(n12419) );
  XNOR2_X1 U14665 ( .A(n12244), .B(n12614), .ZN(n12425) );
  INV_X1 U14666 ( .A(n12245), .ZN(n12424) );
  NAND2_X1 U14667 ( .A1(n12402), .A2(n12403), .ZN(n12665) );
  INV_X1 U14668 ( .A(n12684), .ZN(n12263) );
  NOR2_X1 U14669 ( .A1(n15126), .A2(n12246), .ZN(n12248) );
  INV_X1 U14670 ( .A(n15145), .ZN(n12247) );
  NAND4_X1 U14671 ( .A1(n12248), .A2(n15113), .A3(n15101), .A4(n12247), .ZN(
        n12252) );
  NAND4_X1 U14672 ( .A1(n12250), .A2(n12249), .A3(n12309), .A4(n12297), .ZN(
        n12251) );
  NOR3_X1 U14673 ( .A1(n12252), .A2(n12251), .A3(n12312), .ZN(n12256) );
  NAND4_X1 U14674 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12257) );
  NOR3_X1 U14675 ( .A1(n12833), .A2(n12342), .A3(n12257), .ZN(n12258) );
  NAND4_X1 U14676 ( .A1(n12777), .A2(n12826), .A3(n12811), .A4(n12258), .ZN(
        n12259) );
  NOR4_X1 U14677 ( .A1(n12743), .A2(n6680), .A3(n12260), .A4(n12259), .ZN(
        n12261) );
  INV_X1 U14678 ( .A(n12754), .ZN(n12373) );
  NAND4_X1 U14679 ( .A1(n12710), .A2(n12732), .A3(n12261), .A4(n12373), .ZN(
        n12262) );
  NOR4_X1 U14680 ( .A1(n12665), .A2(n12263), .A3(n12693), .A4(n12262), .ZN(
        n12264) );
  NAND3_X1 U14681 ( .A1(n12641), .A2(n12651), .A3(n12264), .ZN(n12265) );
  XNOR2_X1 U14682 ( .A(n12268), .B(n12614), .ZN(n12270) );
  AND2_X1 U14683 ( .A1(n12284), .A2(n12271), .ZN(n12288) );
  INV_X1 U14684 ( .A(n12272), .ZN(n12279) );
  NOR2_X1 U14685 ( .A1(n12279), .A2(n12273), .ZN(n12277) );
  OAI21_X1 U14686 ( .B1(n15144), .B2(n12275), .A(n12274), .ZN(n12276) );
  MUX2_X1 U14687 ( .A(n12277), .B(n12276), .S(n12397), .Z(n12281) );
  INV_X1 U14688 ( .A(n12282), .ZN(n12278) );
  AOI211_X1 U14689 ( .C1(n12282), .C2(n12281), .A(n15126), .B(n12280), .ZN(
        n12286) );
  AOI21_X1 U14690 ( .B1(n12291), .B2(n12283), .A(n12397), .ZN(n12285) );
  OAI21_X1 U14691 ( .B1(n12286), .B2(n12285), .A(n12284), .ZN(n12287) );
  OAI21_X1 U14692 ( .B1(n12409), .B2(n12288), .A(n12287), .ZN(n12290) );
  NAND3_X1 U14693 ( .A1(n12294), .A2(n12293), .A3(n12302), .ZN(n12295) );
  NAND2_X1 U14694 ( .A1(n12295), .A2(n12300), .ZN(n12305) );
  NAND3_X1 U14695 ( .A1(n12298), .A2(n12297), .A3(n12296), .ZN(n12301) );
  NAND3_X1 U14696 ( .A1(n12301), .A2(n12300), .A3(n12299), .ZN(n12303) );
  NAND2_X1 U14697 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  MUX2_X1 U14698 ( .A(n12305), .B(n12304), .S(n12409), .Z(n12311) );
  MUX2_X1 U14699 ( .A(n12307), .B(n12306), .S(n12409), .Z(n12308) );
  OAI211_X1 U14700 ( .C1(n12311), .C2(n12310), .A(n12309), .B(n12308), .ZN(
        n12317) );
  INV_X1 U14701 ( .A(n12312), .ZN(n12316) );
  MUX2_X1 U14702 ( .A(n12314), .B(n12313), .S(n12397), .Z(n12315) );
  NAND3_X1 U14703 ( .A1(n12317), .A2(n12316), .A3(n12315), .ZN(n12323) );
  INV_X1 U14704 ( .A(n12318), .ZN(n12319) );
  MUX2_X1 U14705 ( .A(n12320), .B(n12319), .S(n12409), .Z(n12322) );
  NOR2_X1 U14706 ( .A1(n12443), .A2(n12397), .ZN(n12326) );
  NOR2_X1 U14707 ( .A1(n12324), .A2(n12409), .ZN(n12325) );
  MUX2_X1 U14708 ( .A(n12326), .B(n12325), .S(n15210), .Z(n12327) );
  AOI21_X1 U14709 ( .B1(n12335), .B2(n12328), .A(n12409), .ZN(n12329) );
  OAI21_X1 U14710 ( .B1(n12330), .B2(n12329), .A(n12331), .ZN(n12338) );
  INV_X1 U14711 ( .A(n12331), .ZN(n12334) );
  INV_X1 U14712 ( .A(n12332), .ZN(n12333) );
  OAI21_X1 U14713 ( .B1(n12334), .B2(n12333), .A(n12409), .ZN(n12337) );
  INV_X1 U14714 ( .A(n12335), .ZN(n12336) );
  AOI22_X1 U14715 ( .A1(n12338), .A2(n12337), .B1(n12409), .B2(n12336), .ZN(
        n12343) );
  INV_X1 U14716 ( .A(n12833), .ZN(n12839) );
  MUX2_X1 U14717 ( .A(n12340), .B(n7152), .S(n12409), .Z(n12341) );
  OAI211_X1 U14718 ( .C1(n12343), .C2(n12342), .A(n12839), .B(n12341), .ZN(
        n12347) );
  MUX2_X1 U14719 ( .A(n12345), .B(n12344), .S(n12397), .Z(n12346) );
  INV_X1 U14720 ( .A(n12356), .ZN(n12350) );
  INV_X1 U14721 ( .A(n12348), .ZN(n12349) );
  OAI21_X1 U14722 ( .B1(n12350), .B2(n12349), .A(n12397), .ZN(n12352) );
  INV_X1 U14723 ( .A(n12355), .ZN(n12351) );
  AOI21_X1 U14724 ( .B1(n12353), .B2(n12352), .A(n12351), .ZN(n12358) );
  AOI21_X1 U14725 ( .B1(n12355), .B2(n12354), .A(n12397), .ZN(n12357) );
  OAI22_X1 U14726 ( .A1(n12358), .A2(n12357), .B1(n12397), .B2(n12356), .ZN(
        n12359) );
  NAND3_X1 U14727 ( .A1(n12359), .A2(n12798), .A3(n12777), .ZN(n12369) );
  NOR2_X1 U14728 ( .A1(n12785), .A2(n12360), .ZN(n12362) );
  AND2_X1 U14729 ( .A1(n12364), .A2(n12397), .ZN(n12361) );
  NAND2_X1 U14730 ( .A1(n12370), .A2(n12361), .ZN(n12366) );
  OAI22_X1 U14731 ( .A1(n12397), .A2(n6736), .B1(n12362), .B2(n12366), .ZN(
        n12368) );
  INV_X1 U14732 ( .A(n12363), .ZN(n12365) );
  NAND3_X1 U14733 ( .A1(n12366), .A2(n12365), .A3(n12364), .ZN(n12367) );
  NAND3_X1 U14734 ( .A1(n12369), .A2(n12368), .A3(n12367), .ZN(n12374) );
  MUX2_X1 U14735 ( .A(n12371), .B(n12370), .S(n12409), .Z(n12372) );
  NAND3_X1 U14736 ( .A1(n12374), .A2(n12373), .A3(n12372), .ZN(n12378) );
  NAND2_X1 U14737 ( .A1(n12753), .A2(n12741), .ZN(n12376) );
  MUX2_X1 U14738 ( .A(n12376), .B(n12375), .S(n12409), .Z(n12377) );
  AOI21_X1 U14739 ( .B1(n12378), .B2(n12377), .A(n12743), .ZN(n12386) );
  MUX2_X1 U14740 ( .A(n12380), .B(n12379), .S(n12409), .Z(n12381) );
  NAND2_X1 U14741 ( .A1(n12732), .A2(n12381), .ZN(n12385) );
  MUX2_X1 U14742 ( .A(n12383), .B(n12382), .S(n12397), .Z(n12384) );
  OAI21_X1 U14743 ( .B1(n12386), .B2(n12385), .A(n12384), .ZN(n12388) );
  NOR2_X1 U14744 ( .A1(n12438), .A2(n12397), .ZN(n12387) );
  AOI22_X1 U14745 ( .A1(n12388), .A2(n12710), .B1(n12387), .B2(n12945), .ZN(
        n12389) );
  NOR2_X1 U14746 ( .A1(n12389), .A2(n12693), .ZN(n12396) );
  INV_X1 U14747 ( .A(n12390), .ZN(n12394) );
  OAI21_X1 U14748 ( .B1(n12394), .B2(n12392), .A(n12391), .ZN(n12393) );
  MUX2_X1 U14749 ( .A(n12394), .B(n12393), .S(n12397), .Z(n12395) );
  MUX2_X1 U14750 ( .A(n12399), .B(n12398), .S(n12397), .Z(n12400) );
  NAND3_X1 U14751 ( .A1(n12401), .A2(n12663), .A3(n12400), .ZN(n12405) );
  MUX2_X1 U14752 ( .A(n12403), .B(n12402), .S(n12409), .Z(n12404) );
  NAND3_X1 U14753 ( .A1(n12405), .A2(n12651), .A3(n12404), .ZN(n12412) );
  NAND2_X1 U14754 ( .A1(n12641), .A2(n12409), .ZN(n12411) );
  OAI21_X1 U14755 ( .B1(n12412), .B2(n12411), .A(n12410), .ZN(n12414) );
  OAI21_X1 U14756 ( .B1(n12415), .B2(n12414), .A(n12413), .ZN(n12420) );
  INV_X1 U14757 ( .A(n12416), .ZN(n12417) );
  NOR4_X1 U14758 ( .A1(n12428), .A2(n12427), .A3(n12998), .A4(n12426), .ZN(
        n12431) );
  OAI21_X1 U14759 ( .B1(n12432), .B2(n12429), .A(P3_B_REG_SCAN_IN), .ZN(n12430) );
  MUX2_X1 U14760 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12434), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14761 ( .A(n12435), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12449), .Z(
        P3_U3518) );
  MUX2_X1 U14762 ( .A(n12436), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12449), .Z(
        P3_U3517) );
  MUX2_X1 U14763 ( .A(n12437), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12449), .Z(
        P3_U3516) );
  MUX2_X1 U14764 ( .A(n12715), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12449), .Z(
        P3_U3515) );
  MUX2_X1 U14765 ( .A(n12438), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12449), .Z(
        P3_U3514) );
  MUX2_X1 U14766 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12714), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14767 ( .A(n12439), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12449), .Z(
        P3_U3512) );
  MUX2_X1 U14768 ( .A(n12440), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12449), .Z(
        P3_U3510) );
  MUX2_X1 U14769 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12796), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14770 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12807), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14771 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n6815), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14772 ( .A(n12441), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12449), .Z(
        P3_U3504) );
  MUX2_X1 U14773 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12442), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14774 ( .A(n12443), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12449), .Z(
        P3_U3501) );
  MUX2_X1 U14775 ( .A(n12444), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12449), .Z(
        P3_U3500) );
  MUX2_X1 U14776 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12445), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14777 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n15105), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14778 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12446), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14779 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n15104), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14780 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12447), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14781 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15150), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14782 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12448), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14783 ( .A(n15147), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12449), .Z(
        P3_U3491) );
  INV_X1 U14784 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15443) );
  NAND2_X1 U14785 ( .A1(n12450), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12451) );
  AOI21_X1 U14786 ( .B1(n15443), .B2(n12453), .A(n12473), .ZN(n12471) );
  INV_X1 U14787 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U14788 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12456), .ZN(n12478) );
  OAI21_X1 U14789 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12456), .A(n12478), 
        .ZN(n12469) );
  AOI21_X1 U14790 ( .B1(n15092), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12457), 
        .ZN(n12458) );
  OAI21_X1 U14791 ( .B1(n15089), .B2(n12477), .A(n12458), .ZN(n12468) );
  INV_X1 U14792 ( .A(n12459), .ZN(n12461) );
  NOR2_X1 U14793 ( .A1(n12461), .A2(n12460), .ZN(n12463) );
  MUX2_X1 U14794 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6648), .Z(n12481) );
  XNOR2_X1 U14795 ( .A(n12481), .B(n12477), .ZN(n12462) );
  INV_X1 U14796 ( .A(n12482), .ZN(n12466) );
  OAI21_X1 U14797 ( .B1(n12464), .B2(n12463), .A(n12462), .ZN(n12465) );
  AOI21_X1 U14798 ( .B1(n12466), .B2(n12465), .A(n12592), .ZN(n12467) );
  AOI211_X1 U14799 ( .C1(n12469), .C2(n15095), .A(n12468), .B(n12467), .ZN(
        n12470) );
  OAI21_X1 U14800 ( .B1(n12471), .B2(n15099), .A(n12470), .ZN(P3_U3195) );
  NOR2_X1 U14801 ( .A1(n12484), .A2(n12472), .ZN(n12474) );
  XNOR2_X1 U14802 ( .A(n12507), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12485) );
  AOI21_X1 U14803 ( .B1(n12475), .B2(n12485), .A(n12499), .ZN(n12498) );
  NAND2_X1 U14804 ( .A1(n12477), .A2(n12476), .ZN(n12479) );
  INV_X1 U14805 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12916) );
  XNOR2_X1 U14806 ( .A(n12507), .B(n12916), .ZN(n12486) );
  OAI21_X1 U14807 ( .B1(n12480), .B2(n12486), .A(n12502), .ZN(n12496) );
  INV_X1 U14808 ( .A(n12481), .ZN(n12483) );
  AOI21_X1 U14809 ( .B1(n12484), .B2(n12483), .A(n12482), .ZN(n12489) );
  INV_X1 U14810 ( .A(n12485), .ZN(n12487) );
  MUX2_X1 U14811 ( .A(n12487), .B(n12486), .S(n6648), .Z(n12488) );
  NAND2_X1 U14812 ( .A1(n12489), .A2(n12488), .ZN(n12511) );
  OAI211_X1 U14813 ( .C1(n12489), .C2(n12488), .A(n12511), .B(n15084), .ZN(
        n12494) );
  INV_X1 U14814 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12491) );
  OAI21_X1 U14815 ( .B1(n12611), .B2(n12491), .A(n12490), .ZN(n12492) );
  INV_X1 U14816 ( .A(n12492), .ZN(n12493) );
  OAI211_X1 U14817 ( .C1(n15089), .C2(n12507), .A(n12494), .B(n12493), .ZN(
        n12495) );
  AOI21_X1 U14818 ( .B1(n15095), .B2(n12496), .A(n12495), .ZN(n12497) );
  OAI21_X1 U14819 ( .B1(n12498), .B2(n15099), .A(n12497), .ZN(P3_U3196) );
  INV_X1 U14820 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12501) );
  AOI21_X1 U14821 ( .B1(n12501), .B2(n12500), .A(n12520), .ZN(n12518) );
  INV_X1 U14822 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14410) );
  NAND2_X1 U14823 ( .A1(n12507), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U14824 ( .A1(n12508), .A2(n12502), .ZN(n12526) );
  OAI21_X1 U14825 ( .B1(n12503), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12528), 
        .ZN(n12504) );
  NAND2_X1 U14826 ( .A1(n15095), .A2(n12504), .ZN(n12506) );
  OAI211_X1 U14827 ( .C1(n14410), .C2(n12611), .A(n12506), .B(n12505), .ZN(
        n12516) );
  NAND2_X1 U14828 ( .A1(n12507), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12509) );
  MUX2_X1 U14829 ( .A(n12509), .B(n12508), .S(n6648), .Z(n12510) );
  NAND2_X1 U14830 ( .A1(n12511), .A2(n12510), .ZN(n12534) );
  XNOR2_X1 U14831 ( .A(n12534), .B(n12527), .ZN(n12513) );
  MUX2_X1 U14832 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6648), .Z(n12512) );
  NOR2_X1 U14833 ( .A1(n12513), .A2(n12512), .ZN(n12535) );
  AOI21_X1 U14834 ( .B1(n12513), .B2(n12512), .A(n12535), .ZN(n12514) );
  NOR2_X1 U14835 ( .A1(n12514), .A2(n12592), .ZN(n12515) );
  AOI211_X1 U14836 ( .C1(n12613), .C2(n12536), .A(n12516), .B(n12515), .ZN(
        n12517) );
  OAI21_X1 U14837 ( .B1(n12518), .B2(n15099), .A(n12517), .ZN(P3_U3197) );
  NOR2_X1 U14838 ( .A1(n12536), .A2(n12519), .ZN(n12521) );
  INV_X1 U14839 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12538) );
  NOR2_X1 U14840 ( .A1(n12541), .A2(n12538), .ZN(n12542) );
  INV_X1 U14841 ( .A(n12542), .ZN(n12564) );
  NAND2_X1 U14842 ( .A1(n12541), .A2(n12538), .ZN(n12522) );
  NAND2_X1 U14843 ( .A1(n12564), .A2(n12522), .ZN(n12524) );
  INV_X1 U14844 ( .A(n12565), .ZN(n12523) );
  AOI21_X1 U14845 ( .B1(n12525), .B2(n12524), .A(n12523), .ZN(n12550) );
  NAND2_X1 U14846 ( .A1(n12527), .A2(n12526), .ZN(n12529) );
  NAND2_X1 U14847 ( .A1(n12529), .A2(n12528), .ZN(n12531) );
  XNOR2_X1 U14848 ( .A(n12541), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12530) );
  OAI21_X1 U14849 ( .B1(n12531), .B2(n12530), .A(n12552), .ZN(n12548) );
  INV_X1 U14850 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14473) );
  NAND2_X1 U14851 ( .A1(n12613), .A2(n12541), .ZN(n12533) );
  OAI211_X1 U14852 ( .C1(n14473), .C2(n12611), .A(n12533), .B(n12532), .ZN(
        n12547) );
  INV_X1 U14853 ( .A(n12534), .ZN(n12537) );
  AOI21_X1 U14854 ( .B1(n12537), .B2(n12536), .A(n12535), .ZN(n12559) );
  INV_X1 U14855 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12540) );
  MUX2_X1 U14856 ( .A(n12538), .B(n12540), .S(n6648), .Z(n12539) );
  NAND2_X1 U14857 ( .A1(n12539), .A2(n12541), .ZN(n12557) );
  INV_X1 U14858 ( .A(n12557), .ZN(n12543) );
  NOR2_X1 U14859 ( .A1(n12541), .A2(n12540), .ZN(n12551) );
  MUX2_X1 U14860 ( .A(n12542), .B(n12551), .S(n6648), .Z(n12558) );
  NOR2_X1 U14861 ( .A1(n12543), .A2(n12558), .ZN(n12544) );
  XNOR2_X1 U14862 ( .A(n12559), .B(n12544), .ZN(n12545) );
  NOR2_X1 U14863 ( .A1(n12545), .A2(n12592), .ZN(n12546) );
  AOI211_X1 U14864 ( .C1(n15095), .C2(n12548), .A(n12547), .B(n12546), .ZN(
        n12549) );
  OAI21_X1 U14865 ( .B1(n12550), .B2(n15099), .A(n12549), .ZN(P3_U3198) );
  INV_X1 U14866 ( .A(n12551), .ZN(n12553) );
  XNOR2_X1 U14867 ( .A(n12578), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U14868 ( .A1(n15092), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12554) );
  OAI211_X1 U14869 ( .C1(n12616), .C2(n12556), .A(n12555), .B(n12554), .ZN(
        n12563) );
  MUX2_X1 U14870 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6648), .Z(n12572) );
  XOR2_X1 U14871 ( .A(n12577), .B(n12572), .Z(n12561) );
  OAI21_X1 U14872 ( .B1(n12559), .B2(n12558), .A(n12557), .ZN(n12560) );
  NOR2_X1 U14873 ( .A1(n12560), .A2(n12561), .ZN(n12570) );
  AOI211_X1 U14874 ( .C1(n12561), .C2(n12560), .A(n12592), .B(n12570), .ZN(
        n12562) );
  AOI211_X1 U14875 ( .C1(n12613), .C2(n12577), .A(n12563), .B(n12562), .ZN(
        n12569) );
  OAI21_X1 U14876 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12566), .A(n12587), 
        .ZN(n12567) );
  NAND2_X1 U14877 ( .A1(n12567), .A2(n12588), .ZN(n12568) );
  NAND2_X1 U14878 ( .A1(n12569), .A2(n12568), .ZN(P3_U3199) );
  MUX2_X1 U14879 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6648), .Z(n12574) );
  AOI21_X1 U14880 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(n12600) );
  XNOR2_X1 U14881 ( .A(n12600), .B(n12599), .ZN(n12573) );
  NOR2_X1 U14882 ( .A1(n12573), .A2(n12574), .ZN(n12598) );
  AOI21_X1 U14883 ( .B1(n12574), .B2(n12573), .A(n12598), .ZN(n12593) );
  XNOR2_X1 U14884 ( .A(n12599), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12606) );
  INV_X1 U14885 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n15323) );
  INV_X1 U14886 ( .A(n12575), .ZN(n12576) );
  OAI22_X1 U14887 ( .A1(n12578), .A2(n15323), .B1(n12577), .B2(n12576), .ZN(
        n12607) );
  NAND2_X1 U14888 ( .A1(n15092), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12579) );
  OAI211_X1 U14889 ( .C1(n12581), .C2(n12616), .A(n12580), .B(n12579), .ZN(
        n12582) );
  INV_X1 U14890 ( .A(n12583), .ZN(n12586) );
  NAND2_X1 U14891 ( .A1(n12605), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12594) );
  INV_X1 U14892 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12784) );
  NAND2_X1 U14893 ( .A1(n12599), .A2(n12784), .ZN(n12584) );
  NAND2_X1 U14894 ( .A1(n12594), .A2(n12584), .ZN(n12585) );
  AND3_X1 U14895 ( .A1(n12587), .A2(n12586), .A3(n12585), .ZN(n12589) );
  OAI21_X1 U14896 ( .B1(n12596), .B2(n12589), .A(n12588), .ZN(n12590) );
  OAI211_X1 U14897 ( .C1(n12593), .C2(n12592), .A(n12591), .B(n12590), .ZN(
        P3_U3200) );
  XNOR2_X1 U14898 ( .A(n12601), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12602) );
  INV_X1 U14899 ( .A(n12594), .ZN(n12595) );
  AOI21_X1 U14900 ( .B1(n12600), .B2(n12599), .A(n12598), .ZN(n12604) );
  XNOR2_X1 U14901 ( .A(n12601), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12608) );
  MUX2_X1 U14902 ( .A(n12602), .B(n12608), .S(n6648), .Z(n12603) );
  XNOR2_X1 U14903 ( .A(n12604), .B(n12603), .ZN(n12617) );
  AOI22_X1 U14904 ( .A1(n12607), .A2(n12606), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12605), .ZN(n12609) );
  OAI21_X1 U14905 ( .B1(n12611), .B2(n15447), .A(n12610), .ZN(n12612) );
  AOI21_X1 U14906 ( .B1(n12614), .B2(n12613), .A(n12612), .ZN(n12615) );
  NOR2_X1 U14907 ( .A1(n12619), .A2(n12618), .ZN(n12919) );
  NOR2_X1 U14908 ( .A1(n12620), .A2(n12782), .ZN(n12629) );
  AOI21_X1 U14909 ( .B1(n12919), .B2(n15162), .A(n12629), .ZN(n12622) );
  NAND2_X1 U14910 ( .A1(n12846), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12621) );
  OAI211_X1 U14911 ( .C1(n12921), .C2(n12842), .A(n12622), .B(n12621), .ZN(
        P3_U3202) );
  NAND2_X1 U14912 ( .A1(n12922), .A2(n12792), .ZN(n12623) );
  OAI211_X1 U14913 ( .C1(n15162), .C2(n12624), .A(n12623), .B(n12622), .ZN(
        P3_U3203) );
  INV_X1 U14914 ( .A(n12625), .ZN(n12632) );
  NAND2_X1 U14915 ( .A1(n12626), .A2(n15162), .ZN(n12631) );
  NOR2_X1 U14916 ( .A1(n12627), .A2(n12842), .ZN(n12628) );
  AOI211_X1 U14917 ( .C1(n12846), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12629), 
        .B(n12628), .ZN(n12630) );
  OAI211_X1 U14918 ( .C1(n12632), .C2(n12787), .A(n12631), .B(n12630), .ZN(
        P3_U3204) );
  OAI211_X1 U14919 ( .C1(n12635), .C2(n12634), .A(n12633), .B(n15133), .ZN(
        n12639) );
  OAI22_X1 U14920 ( .A1(n12636), .A2(n15128), .B1(n12667), .B2(n15130), .ZN(
        n12637) );
  INV_X1 U14921 ( .A(n12637), .ZN(n12638) );
  NAND2_X1 U14922 ( .A1(n12650), .A2(n12640), .ZN(n12642) );
  XNOR2_X1 U14923 ( .A(n12642), .B(n12641), .ZN(n12852) );
  AOI22_X1 U14924 ( .A1(n12643), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12644) );
  OAI21_X1 U14925 ( .B1(n12929), .B2(n12842), .A(n12644), .ZN(n12645) );
  AOI21_X1 U14926 ( .B1(n12852), .B2(n12844), .A(n12645), .ZN(n12646) );
  OAI21_X1 U14927 ( .B1(n12854), .B2(n12846), .A(n12646), .ZN(P3_U3205) );
  INV_X1 U14928 ( .A(n12647), .ZN(n12648) );
  AOI21_X1 U14929 ( .B1(n12651), .B2(n12649), .A(n12648), .ZN(n12656) );
  OAI22_X1 U14930 ( .A1(n12653), .A2(n15128), .B1(n12680), .B2(n15130), .ZN(
        n12654) );
  AOI21_X1 U14931 ( .B1(n12858), .B2(n12697), .A(n12654), .ZN(n12655) );
  INV_X1 U14932 ( .A(n12857), .ZN(n12662) );
  INV_X1 U14933 ( .A(n12657), .ZN(n12933) );
  AOI22_X1 U14934 ( .A1(n12658), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12659) );
  OAI21_X1 U14935 ( .B1(n12933), .B2(n12842), .A(n12659), .ZN(n12660) );
  AOI21_X1 U14936 ( .B1(n12858), .B2(n12704), .A(n12660), .ZN(n12661) );
  OAI21_X1 U14937 ( .B1(n12662), .B2(n12846), .A(n12661), .ZN(P3_U3206) );
  XNOR2_X1 U14938 ( .A(n12664), .B(n12663), .ZN(n12863) );
  INV_X1 U14939 ( .A(n12863), .ZN(n12677) );
  XNOR2_X1 U14940 ( .A(n12666), .B(n12665), .ZN(n12670) );
  OAI22_X1 U14941 ( .A1(n12667), .A2(n15128), .B1(n12695), .B2(n15130), .ZN(
        n12668) );
  AOI21_X1 U14942 ( .B1(n12863), .B2(n12697), .A(n12668), .ZN(n12669) );
  OAI21_X1 U14943 ( .B1(n12670), .B2(n15154), .A(n12669), .ZN(n12862) );
  NAND2_X1 U14944 ( .A1(n12862), .A2(n15162), .ZN(n12676) );
  NAND2_X1 U14945 ( .A1(n12671), .A2(n15157), .ZN(n12672) );
  OAI21_X1 U14946 ( .B1(n15162), .B2(n12673), .A(n12672), .ZN(n12674) );
  AOI21_X1 U14947 ( .B1(n12861), .B2(n12792), .A(n12674), .ZN(n12675) );
  OAI211_X1 U14948 ( .C1(n12723), .C2(n12677), .A(n12676), .B(n12675), .ZN(
        P3_U3207) );
  XNOR2_X1 U14949 ( .A(n12678), .B(n12684), .ZN(n12867) );
  OAI22_X1 U14950 ( .A1(n12680), .A2(n15128), .B1(n12679), .B2(n15130), .ZN(
        n12686) );
  INV_X1 U14951 ( .A(n12681), .ZN(n12682) );
  AOI211_X1 U14952 ( .C1(n12684), .C2(n12683), .A(n15154), .B(n12682), .ZN(
        n12685) );
  AOI211_X1 U14953 ( .C1(n12867), .C2(n12697), .A(n12686), .B(n12685), .ZN(
        n12869) );
  INV_X1 U14954 ( .A(n12866), .ZN(n12689) );
  AOI22_X1 U14955 ( .A1(n12687), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12688) );
  OAI21_X1 U14956 ( .B1(n12689), .B2(n12842), .A(n12688), .ZN(n12690) );
  AOI21_X1 U14957 ( .B1(n12867), .B2(n12704), .A(n12690), .ZN(n12691) );
  OAI21_X1 U14958 ( .B1(n12869), .B2(n12846), .A(n12691), .ZN(P3_U3208) );
  XNOR2_X1 U14959 ( .A(n12692), .B(n12693), .ZN(n12699) );
  OAI21_X1 U14960 ( .B1(n6665), .B2(n6833), .A(n12694), .ZN(n12871) );
  OAI22_X1 U14961 ( .A1(n12695), .A2(n15128), .B1(n12730), .B2(n15130), .ZN(
        n12696) );
  AOI21_X1 U14962 ( .B1(n12871), .B2(n12697), .A(n12696), .ZN(n12698) );
  OAI21_X1 U14963 ( .B1(n12699), .B2(n15154), .A(n12698), .ZN(n12870) );
  INV_X1 U14964 ( .A(n12870), .ZN(n12706) );
  INV_X1 U14965 ( .A(n12700), .ZN(n12942) );
  AOI22_X1 U14966 ( .A1(n12701), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12702) );
  OAI21_X1 U14967 ( .B1(n12942), .B2(n12842), .A(n12702), .ZN(n12703) );
  AOI21_X1 U14968 ( .B1(n12871), .B2(n12704), .A(n12703), .ZN(n12705) );
  OAI21_X1 U14969 ( .B1(n12706), .B2(n12846), .A(n12705), .ZN(P3_U3209) );
  NAND2_X1 U14970 ( .A1(n12708), .A2(n12707), .ZN(n12709) );
  XNOR2_X1 U14971 ( .A(n12709), .B(n12710), .ZN(n12718) );
  OR2_X1 U14972 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  NAND2_X1 U14973 ( .A1(n12713), .A2(n12712), .ZN(n12874) );
  AOI22_X1 U14974 ( .A1(n12715), .A2(n15149), .B1(n15148), .B2(n12714), .ZN(
        n12716) );
  OAI21_X1 U14975 ( .B1(n12874), .B2(n15146), .A(n12716), .ZN(n12717) );
  AOI21_X1 U14976 ( .B1(n12718), .B2(n15133), .A(n12717), .ZN(n12876) );
  NAND2_X1 U14977 ( .A1(n12719), .A2(n15157), .ZN(n12720) );
  OAI21_X1 U14978 ( .B1(n15162), .B2(n12721), .A(n12720), .ZN(n12722) );
  AOI21_X1 U14979 ( .B1(n12945), .B2(n12792), .A(n12722), .ZN(n12725) );
  OR2_X1 U14980 ( .A1(n12874), .A2(n12723), .ZN(n12724) );
  OAI211_X1 U14981 ( .C1(n12876), .C2(n12846), .A(n12725), .B(n12724), .ZN(
        P3_U3210) );
  NAND2_X1 U14982 ( .A1(n12727), .A2(n12726), .ZN(n12728) );
  XNOR2_X1 U14983 ( .A(n12728), .B(n12732), .ZN(n12729) );
  OAI222_X1 U14984 ( .A1(n15128), .A2(n12730), .B1(n15130), .B2(n12752), .C1(
        n15154), .C2(n12729), .ZN(n12880) );
  INV_X1 U14985 ( .A(n12880), .ZN(n12738) );
  XOR2_X1 U14986 ( .A(n12731), .B(n12732), .Z(n12881) );
  INV_X1 U14987 ( .A(n12733), .ZN(n12951) );
  AOI22_X1 U14988 ( .A1(n12734), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12735) );
  OAI21_X1 U14989 ( .B1(n12951), .B2(n12842), .A(n12735), .ZN(n12736) );
  AOI21_X1 U14990 ( .B1(n12881), .B2(n12844), .A(n12736), .ZN(n12737) );
  OAI21_X1 U14991 ( .B1(n12738), .B2(n12846), .A(n12737), .ZN(P3_U3211) );
  XNOR2_X1 U14992 ( .A(n12739), .B(n12743), .ZN(n12740) );
  OAI222_X1 U14993 ( .A1(n15128), .A2(n12742), .B1(n15130), .B2(n12741), .C1(
        n15154), .C2(n12740), .ZN(n12884) );
  INV_X1 U14994 ( .A(n12884), .ZN(n12749) );
  XNOR2_X1 U14995 ( .A(n12744), .B(n12743), .ZN(n12885) );
  AOI22_X1 U14996 ( .A1(n12745), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n12746) );
  OAI21_X1 U14997 ( .B1(n12955), .B2(n12842), .A(n12746), .ZN(n12747) );
  AOI21_X1 U14998 ( .B1(n12885), .B2(n12844), .A(n12747), .ZN(n12748) );
  OAI21_X1 U14999 ( .B1(n12749), .B2(n12846), .A(n12748), .ZN(P3_U3212) );
  XNOR2_X1 U15000 ( .A(n12750), .B(n12754), .ZN(n12751) );
  OAI222_X1 U15001 ( .A1(n15128), .A2(n12752), .B1(n15130), .B2(n12780), .C1(
        n15154), .C2(n12751), .ZN(n12888) );
  INV_X1 U15002 ( .A(n12753), .ZN(n12959) );
  NAND2_X1 U15003 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  AND2_X1 U15004 ( .A1(n12757), .A2(n12756), .ZN(n12889) );
  NAND2_X1 U15005 ( .A1(n12889), .A2(n12844), .ZN(n12760) );
  AOI22_X1 U15006 ( .A1(n12758), .A2(n15157), .B1(n12846), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n12759) );
  OAI211_X1 U15007 ( .C1(n12959), .C2(n12842), .A(n12760), .B(n12759), .ZN(
        n12761) );
  AOI21_X1 U15008 ( .B1(n12888), .B2(n15162), .A(n12761), .ZN(n12762) );
  INV_X1 U15009 ( .A(n12762), .ZN(P3_U3213) );
  OAI211_X1 U15010 ( .C1(n6775), .C2(n6680), .A(n15133), .B(n12763), .ZN(
        n12766) );
  AOI22_X1 U15011 ( .A1(n12764), .A2(n15149), .B1(n15148), .B2(n12796), .ZN(
        n12765) );
  NAND2_X1 U15012 ( .A1(n12766), .A2(n12765), .ZN(n12892) );
  INV_X1 U15013 ( .A(n12892), .ZN(n12773) );
  NAND2_X1 U15014 ( .A1(n12898), .A2(n12767), .ZN(n12768) );
  XNOR2_X1 U15015 ( .A(n12768), .B(n6680), .ZN(n12893) );
  AOI22_X1 U15016 ( .A1(n12846), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12769), 
        .B2(n15157), .ZN(n12770) );
  OAI21_X1 U15017 ( .B1(n12963), .B2(n12842), .A(n12770), .ZN(n12771) );
  AOI21_X1 U15018 ( .B1(n12893), .B2(n12844), .A(n12771), .ZN(n12772) );
  OAI21_X1 U15019 ( .B1(n12773), .B2(n12846), .A(n12772), .ZN(P3_U3214) );
  INV_X1 U15020 ( .A(n12774), .ZN(n12775) );
  AOI21_X1 U15021 ( .B1(n12777), .B2(n12776), .A(n12775), .ZN(n12778) );
  OAI222_X1 U15022 ( .A1(n15128), .A2(n12780), .B1(n15130), .B2(n12779), .C1(
        n15154), .C2(n12778), .ZN(n12897) );
  INV_X1 U15023 ( .A(n12897), .ZN(n12794) );
  INV_X1 U15024 ( .A(n12781), .ZN(n12783) );
  OAI22_X1 U15025 ( .A1(n15162), .A2(n12784), .B1(n12783), .B2(n12782), .ZN(
        n12790) );
  INV_X1 U15026 ( .A(n12898), .ZN(n12788) );
  AND2_X1 U15027 ( .A1(n12786), .A2(n12785), .ZN(n12896) );
  NOR3_X1 U15028 ( .A1(n12788), .A2(n12896), .A3(n12787), .ZN(n12789) );
  AOI211_X1 U15029 ( .C1(n12792), .C2(n12791), .A(n12790), .B(n12789), .ZN(
        n12793) );
  OAI21_X1 U15030 ( .B1(n12794), .B2(n12846), .A(n12793), .ZN(P3_U3215) );
  XNOR2_X1 U15031 ( .A(n12795), .B(n12798), .ZN(n12797) );
  AOI222_X1 U15032 ( .A1(n15133), .A2(n12797), .B1(n12796), .B2(n15149), .C1(
        n6815), .C2(n15148), .ZN(n12905) );
  XNOR2_X1 U15033 ( .A(n12799), .B(n12798), .ZN(n12903) );
  AOI22_X1 U15034 ( .A1(n12846), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15157), 
        .B2(n12800), .ZN(n12801) );
  OAI21_X1 U15035 ( .B1(n12802), .B2(n12842), .A(n12801), .ZN(n12803) );
  AOI21_X1 U15036 ( .B1(n12903), .B2(n12844), .A(n12803), .ZN(n12804) );
  OAI21_X1 U15037 ( .B1(n12905), .B2(n12846), .A(n12804), .ZN(P3_U3216) );
  XNOR2_X1 U15038 ( .A(n12805), .B(n12811), .ZN(n12808) );
  AOI222_X1 U15039 ( .A1(n15133), .A2(n12808), .B1(n12807), .B2(n15149), .C1(
        n12806), .C2(n15148), .ZN(n12909) );
  OAI21_X1 U15040 ( .B1(n12811), .B2(n12810), .A(n12809), .ZN(n12907) );
  AOI22_X1 U15041 ( .A1(n12846), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12812), 
        .B2(n15157), .ZN(n12813) );
  OAI21_X1 U15042 ( .B1(n12814), .B2(n12842), .A(n12813), .ZN(n12815) );
  AOI21_X1 U15043 ( .B1(n12907), .B2(n12844), .A(n12815), .ZN(n12816) );
  OAI21_X1 U15044 ( .B1(n12909), .B2(n12846), .A(n12816), .ZN(P3_U3217) );
  NAND2_X1 U15045 ( .A1(n12818), .A2(n12817), .ZN(n12834) );
  NAND2_X1 U15046 ( .A1(n12834), .A2(n12833), .ZN(n12820) );
  NAND2_X1 U15047 ( .A1(n12820), .A2(n12819), .ZN(n12822) );
  XNOR2_X1 U15048 ( .A(n12822), .B(n12821), .ZN(n12823) );
  OAI222_X1 U15049 ( .A1(n15128), .A2(n12825), .B1(n15130), .B2(n12824), .C1(
        n12823), .C2(n15154), .ZN(n12910) );
  INV_X1 U15050 ( .A(n12910), .ZN(n12832) );
  XNOR2_X1 U15051 ( .A(n12827), .B(n12826), .ZN(n12911) );
  AOI22_X1 U15052 ( .A1(n12846), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15157), 
        .B2(n12828), .ZN(n12829) );
  OAI21_X1 U15053 ( .B1(n12973), .B2(n12842), .A(n12829), .ZN(n12830) );
  AOI21_X1 U15054 ( .B1(n12911), .B2(n12844), .A(n12830), .ZN(n12831) );
  OAI21_X1 U15055 ( .B1(n12832), .B2(n12846), .A(n12831), .ZN(P3_U3218) );
  XNOR2_X1 U15056 ( .A(n12834), .B(n12833), .ZN(n12835) );
  OAI222_X1 U15057 ( .A1(n15130), .A2(n12837), .B1(n15128), .B2(n12836), .C1(
        n12835), .C2(n15154), .ZN(n12914) );
  INV_X1 U15058 ( .A(n12914), .ZN(n12847) );
  OAI21_X1 U15059 ( .B1(n6774), .B2(n12839), .A(n12838), .ZN(n12915) );
  AOI22_X1 U15060 ( .A1(n12846), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15157), 
        .B2(n12840), .ZN(n12841) );
  OAI21_X1 U15061 ( .B1(n12977), .B2(n12842), .A(n12841), .ZN(n12843) );
  AOI21_X1 U15062 ( .B1(n12915), .B2(n12844), .A(n12843), .ZN(n12845) );
  OAI21_X1 U15063 ( .B1(n12847), .B2(n12846), .A(n12845), .ZN(P3_U3219) );
  NAND2_X1 U15064 ( .A1(n15231), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U15065 ( .A1(n12919), .A2(n15227), .ZN(n12850) );
  OAI211_X1 U15066 ( .C1(n12921), .C2(n12918), .A(n12848), .B(n12850), .ZN(
        P3_U3490) );
  NAND2_X1 U15067 ( .A1(n15231), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12849) );
  OAI211_X1 U15068 ( .C1(n12851), .C2(n12918), .A(n12850), .B(n12849), .ZN(
        P3_U3489) );
  NAND2_X1 U15069 ( .A1(n12852), .A2(n14537), .ZN(n12853) );
  NAND2_X1 U15070 ( .A1(n12854), .A2(n12853), .ZN(n12926) );
  MUX2_X1 U15071 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12926), .S(n15227), .Z(
        n12855) );
  INV_X1 U15072 ( .A(n12855), .ZN(n12856) );
  OAI21_X1 U15073 ( .B1(n12929), .B2(n12918), .A(n12856), .ZN(P3_U3487) );
  INV_X1 U15074 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12859) );
  MUX2_X1 U15075 ( .A(n12859), .B(n12930), .S(n15227), .Z(n12860) );
  INV_X1 U15076 ( .A(n12861), .ZN(n12937) );
  INV_X1 U15077 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12864) );
  AOI21_X1 U15078 ( .B1(n15206), .B2(n12863), .A(n12862), .ZN(n12934) );
  MUX2_X1 U15079 ( .A(n12864), .B(n12934), .S(n15227), .Z(n12865) );
  OAI21_X1 U15080 ( .B1(n12937), .B2(n12918), .A(n12865), .ZN(P3_U3485) );
  AOI22_X1 U15081 ( .A1(n12867), .A2(n15206), .B1(n15155), .B2(n12866), .ZN(
        n12868) );
  NAND2_X1 U15082 ( .A1(n12869), .A2(n12868), .ZN(n12938) );
  MUX2_X1 U15083 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12938), .S(n15227), .Z(
        P3_U3484) );
  INV_X1 U15084 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12872) );
  AOI21_X1 U15085 ( .B1(n15206), .B2(n12871), .A(n12870), .ZN(n12939) );
  MUX2_X1 U15086 ( .A(n12872), .B(n12939), .S(n15227), .Z(n12873) );
  OAI21_X1 U15087 ( .B1(n12942), .B2(n12918), .A(n12873), .ZN(P3_U3483) );
  INV_X1 U15088 ( .A(n15206), .ZN(n15185) );
  OR2_X1 U15089 ( .A1(n12874), .A2(n15185), .ZN(n12875) );
  NAND2_X1 U15090 ( .A1(n12876), .A2(n12875), .ZN(n12943) );
  MUX2_X1 U15091 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12943), .S(n15227), .Z(
        n12877) );
  AOI21_X1 U15092 ( .B1(n12878), .B2(n12945), .A(n12877), .ZN(n12879) );
  INV_X1 U15093 ( .A(n12879), .ZN(P3_U3482) );
  INV_X1 U15094 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12882) );
  AOI21_X1 U15095 ( .B1(n14537), .B2(n12881), .A(n12880), .ZN(n12948) );
  MUX2_X1 U15096 ( .A(n12882), .B(n12948), .S(n15227), .Z(n12883) );
  OAI21_X1 U15097 ( .B1(n12951), .B2(n12918), .A(n12883), .ZN(P3_U3481) );
  INV_X1 U15098 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12886) );
  AOI21_X1 U15099 ( .B1(n12885), .B2(n14537), .A(n12884), .ZN(n12952) );
  MUX2_X1 U15100 ( .A(n12886), .B(n12952), .S(n15227), .Z(n12887) );
  OAI21_X1 U15101 ( .B1(n12955), .B2(n12918), .A(n12887), .ZN(P3_U3480) );
  INV_X1 U15102 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12890) );
  AOI21_X1 U15103 ( .B1(n12889), .B2(n14537), .A(n12888), .ZN(n12956) );
  MUX2_X1 U15104 ( .A(n12890), .B(n12956), .S(n15227), .Z(n12891) );
  OAI21_X1 U15105 ( .B1(n12959), .B2(n12918), .A(n12891), .ZN(P3_U3479) );
  INV_X1 U15106 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12894) );
  AOI21_X1 U15107 ( .B1(n14537), .B2(n12893), .A(n12892), .ZN(n12960) );
  MUX2_X1 U15108 ( .A(n12894), .B(n12960), .S(n15227), .Z(n12895) );
  OAI21_X1 U15109 ( .B1(n12918), .B2(n12963), .A(n12895), .ZN(P3_U3478) );
  INV_X1 U15110 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12900) );
  INV_X1 U15111 ( .A(n14537), .ZN(n15211) );
  NOR2_X1 U15112 ( .A1(n12896), .A2(n15211), .ZN(n12899) );
  AOI21_X1 U15113 ( .B1(n12899), .B2(n12898), .A(n12897), .ZN(n12964) );
  MUX2_X1 U15114 ( .A(n12900), .B(n12964), .S(n15227), .Z(n12901) );
  OAI21_X1 U15115 ( .B1(n12967), .B2(n12918), .A(n12901), .ZN(P3_U3477) );
  AOI22_X1 U15116 ( .A1(n12903), .A2(n14537), .B1(n15155), .B2(n12902), .ZN(
        n12904) );
  NAND2_X1 U15117 ( .A1(n12905), .A2(n12904), .ZN(n12968) );
  MUX2_X1 U15118 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12968), .S(n15227), .Z(
        P3_U3476) );
  AOI22_X1 U15119 ( .A1(n12907), .A2(n14537), .B1(n15155), .B2(n12906), .ZN(
        n12908) );
  NAND2_X1 U15120 ( .A1(n12909), .A2(n12908), .ZN(n12969) );
  MUX2_X1 U15121 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12969), .S(n15227), .Z(
        P3_U3475) );
  INV_X1 U15122 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12912) );
  AOI21_X1 U15123 ( .B1(n12911), .B2(n14537), .A(n12910), .ZN(n12970) );
  MUX2_X1 U15124 ( .A(n12912), .B(n12970), .S(n15227), .Z(n12913) );
  OAI21_X1 U15125 ( .B1(n12973), .B2(n12918), .A(n12913), .ZN(P3_U3474) );
  AOI21_X1 U15126 ( .B1(n14537), .B2(n12915), .A(n12914), .ZN(n12974) );
  MUX2_X1 U15127 ( .A(n12916), .B(n12974), .S(n15227), .Z(n12917) );
  OAI21_X1 U15128 ( .B1(n12918), .B2(n12977), .A(n12917), .ZN(P3_U3473) );
  NAND2_X1 U15129 ( .A1(n15215), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U15130 ( .A1(n12919), .A2(n15217), .ZN(n12923) );
  OAI211_X1 U15131 ( .C1(n12921), .C2(n12978), .A(n12920), .B(n12923), .ZN(
        P3_U3458) );
  INV_X1 U15132 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12925) );
  INV_X1 U15133 ( .A(n12978), .ZN(n12946) );
  NAND2_X1 U15134 ( .A1(n12922), .A2(n12946), .ZN(n12924) );
  OAI211_X1 U15135 ( .C1(n15217), .C2(n12925), .A(n12924), .B(n12923), .ZN(
        P3_U3457) );
  MUX2_X1 U15136 ( .A(n12926), .B(P3_REG0_REG_28__SCAN_IN), .S(n15215), .Z(
        n12927) );
  INV_X1 U15137 ( .A(n12927), .ZN(n12928) );
  OAI21_X1 U15138 ( .B1(n12929), .B2(n12978), .A(n12928), .ZN(P3_U3455) );
  INV_X1 U15139 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12931) );
  MUX2_X1 U15140 ( .A(n12931), .B(n12930), .S(n15217), .Z(n12932) );
  INV_X1 U15141 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12935) );
  MUX2_X1 U15142 ( .A(n12935), .B(n12934), .S(n15217), .Z(n12936) );
  OAI21_X1 U15143 ( .B1(n12937), .B2(n12978), .A(n12936), .ZN(P3_U3453) );
  MUX2_X1 U15144 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12938), .S(n15217), .Z(
        P3_U3452) );
  INV_X1 U15145 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12940) );
  MUX2_X1 U15146 ( .A(n12940), .B(n12939), .S(n15217), .Z(n12941) );
  OAI21_X1 U15147 ( .B1(n12942), .B2(n12978), .A(n12941), .ZN(P3_U3451) );
  MUX2_X1 U15148 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12943), .S(n15217), .Z(
        n12944) );
  AOI21_X1 U15149 ( .B1(n12946), .B2(n12945), .A(n12944), .ZN(n12947) );
  INV_X1 U15150 ( .A(n12947), .ZN(P3_U3450) );
  INV_X1 U15151 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12949) );
  MUX2_X1 U15152 ( .A(n12949), .B(n12948), .S(n15217), .Z(n12950) );
  OAI21_X1 U15153 ( .B1(n12951), .B2(n12978), .A(n12950), .ZN(P3_U3449) );
  INV_X1 U15154 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12953) );
  MUX2_X1 U15155 ( .A(n12953), .B(n12952), .S(n15217), .Z(n12954) );
  OAI21_X1 U15156 ( .B1(n12955), .B2(n12978), .A(n12954), .ZN(P3_U3448) );
  INV_X1 U15157 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12957) );
  MUX2_X1 U15158 ( .A(n12957), .B(n12956), .S(n15217), .Z(n12958) );
  OAI21_X1 U15159 ( .B1(n12959), .B2(n12978), .A(n12958), .ZN(P3_U3447) );
  MUX2_X1 U15160 ( .A(n12961), .B(n12960), .S(n15217), .Z(n12962) );
  OAI21_X1 U15161 ( .B1(n12978), .B2(n12963), .A(n12962), .ZN(P3_U3446) );
  INV_X1 U15162 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12965) );
  MUX2_X1 U15163 ( .A(n12965), .B(n12964), .S(n15217), .Z(n12966) );
  OAI21_X1 U15164 ( .B1(n12967), .B2(n12978), .A(n12966), .ZN(P3_U3444) );
  MUX2_X1 U15165 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12968), .S(n15217), .Z(
        P3_U3441) );
  MUX2_X1 U15166 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12969), .S(n15217), .Z(
        P3_U3438) );
  INV_X1 U15167 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12971) );
  MUX2_X1 U15168 ( .A(n12971), .B(n12970), .S(n15217), .Z(n12972) );
  OAI21_X1 U15169 ( .B1(n12973), .B2(n12978), .A(n12972), .ZN(P3_U3435) );
  INV_X1 U15170 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12975) );
  MUX2_X1 U15171 ( .A(n12975), .B(n12974), .S(n15217), .Z(n12976) );
  OAI21_X1 U15172 ( .B1(n12978), .B2(n12977), .A(n12976), .ZN(P3_U3432) );
  NAND2_X1 U15173 ( .A1(n12980), .A2(n12979), .ZN(n12984) );
  OR4_X1 U15174 ( .A1(n12982), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12981), .A4(
        P3_U3151), .ZN(n12983) );
  OAI211_X1 U15175 ( .C1(n12986), .C2(n12985), .A(n12984), .B(n12983), .ZN(
        P3_U3264) );
  INV_X1 U15176 ( .A(n12987), .ZN(n12988) );
  OAI222_X1 U15177 ( .A1(n12990), .A2(P3_U3151), .B1(n12985), .B2(n12989), 
        .C1(n12997), .C2(n12988), .ZN(P3_U3265) );
  INV_X1 U15178 ( .A(n12991), .ZN(n12993) );
  OAI222_X1 U15179 ( .A1(n12985), .A2(n12994), .B1(n12997), .B2(n12993), .C1(
        n12992), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15180 ( .A(n12995), .ZN(n12996) );
  XNOR2_X1 U15181 ( .A(n13588), .B(n13001), .ZN(n13012) );
  NAND2_X1 U15182 ( .A1(n13292), .A2(n13030), .ZN(n13011) );
  NAND2_X1 U15183 ( .A1(n13286), .A2(n13066), .ZN(n13004) );
  INV_X1 U15184 ( .A(n13004), .ZN(n13007) );
  XNOR2_X1 U15185 ( .A(n13599), .B(n13035), .ZN(n13006) );
  INV_X1 U15186 ( .A(n13002), .ZN(n13003) );
  NOR2_X1 U15187 ( .A1(n13087), .A2(n13003), .ZN(n13005) );
  XNOR2_X1 U15188 ( .A(n13006), .B(n13004), .ZN(n13088) );
  OAI21_X1 U15189 ( .B1(n13007), .B2(n13006), .A(n13094), .ZN(n13125) );
  XNOR2_X1 U15190 ( .A(n13289), .B(n13035), .ZN(n13049) );
  AND2_X1 U15191 ( .A1(n13254), .A2(n13030), .ZN(n13008) );
  NAND2_X1 U15192 ( .A1(n13049), .A2(n13008), .ZN(n13009) );
  OAI21_X1 U15193 ( .B1(n13049), .B2(n13008), .A(n13009), .ZN(n13124) );
  INV_X1 U15194 ( .A(n13009), .ZN(n13010) );
  XNOR2_X1 U15195 ( .A(n13012), .B(n13011), .ZN(n13051) );
  XNOR2_X1 U15196 ( .A(n13457), .B(n13035), .ZN(n13016) );
  INV_X1 U15197 ( .A(n13016), .ZN(n13014) );
  AND2_X1 U15198 ( .A1(n13258), .A2(n13030), .ZN(n13015) );
  INV_X1 U15199 ( .A(n13015), .ZN(n13013) );
  NAND2_X1 U15200 ( .A1(n13014), .A2(n13013), .ZN(n13101) );
  AND2_X1 U15201 ( .A1(n13016), .A2(n13015), .ZN(n13102) );
  NAND2_X1 U15202 ( .A1(n13261), .A2(n13066), .ZN(n13018) );
  XNOR2_X1 U15203 ( .A(n13442), .B(n13035), .ZN(n13017) );
  XOR2_X1 U15204 ( .A(n13018), .B(n13017), .Z(n13074) );
  INV_X1 U15205 ( .A(n13017), .ZN(n13019) );
  XNOR2_X1 U15206 ( .A(n13423), .B(n13035), .ZN(n13021) );
  NAND2_X1 U15207 ( .A1(n13264), .A2(n13066), .ZN(n13110) );
  INV_X1 U15208 ( .A(n13020), .ZN(n13023) );
  INV_X1 U15209 ( .A(n13021), .ZN(n13022) );
  INV_X1 U15210 ( .A(n13268), .ZN(n13302) );
  NOR2_X1 U15211 ( .A1(n13302), .A2(n13488), .ZN(n13040) );
  NAND2_X1 U15212 ( .A1(n13271), .A2(n13066), .ZN(n13026) );
  XNOR2_X1 U15213 ( .A(n13558), .B(n13035), .ZN(n13025) );
  XOR2_X1 U15214 ( .A(n13026), .B(n13025), .Z(n13095) );
  XNOR2_X1 U15215 ( .A(n13379), .B(n13035), .ZN(n13028) );
  NAND2_X1 U15216 ( .A1(n13274), .A2(n13066), .ZN(n13027) );
  XNOR2_X1 U15217 ( .A(n13028), .B(n13027), .ZN(n13080) );
  INV_X1 U15218 ( .A(n13027), .ZN(n13029) );
  AND2_X1 U15219 ( .A1(n13278), .A2(n13030), .ZN(n13032) );
  XNOR2_X1 U15220 ( .A(n13547), .B(n13035), .ZN(n13031) );
  NOR2_X1 U15221 ( .A1(n13031), .A2(n13032), .ZN(n13033) );
  AOI21_X1 U15222 ( .B1(n13032), .B2(n13031), .A(n13033), .ZN(n13131) );
  INV_X1 U15223 ( .A(n13033), .ZN(n13034) );
  NAND2_X1 U15224 ( .A1(n13279), .A2(n13066), .ZN(n13062) );
  XNOR2_X1 U15225 ( .A(n13541), .B(n13035), .ZN(n13061) );
  XOR2_X1 U15226 ( .A(n13062), .B(n13061), .Z(n13064) );
  XNOR2_X1 U15227 ( .A(n13065), .B(n13064), .ZN(n13039) );
  AOI22_X1 U15228 ( .A1(n13142), .A2(n13237), .B1(n13120), .B2(n13278), .ZN(
        n13344) );
  AOI22_X1 U15229 ( .A1(n13350), .A2(n13121), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13036) );
  OAI21_X1 U15230 ( .B1(n13344), .B2(n14554), .A(n13036), .ZN(n13037) );
  AOI21_X1 U15231 ( .B1(n13541), .B2(n13128), .A(n13037), .ZN(n13038) );
  OAI21_X1 U15232 ( .B1(n13039), .B2(n14552), .A(n13038), .ZN(P2_U3186) );
  NAND2_X1 U15233 ( .A1(n13268), .A2(n13111), .ZN(n13043) );
  OR2_X1 U15234 ( .A1(n13040), .A2(n14552), .ZN(n13042) );
  MUX2_X1 U15235 ( .A(n13043), .B(n13042), .S(n13041), .Z(n13047) );
  INV_X1 U15236 ( .A(n13271), .ZN(n13304) );
  OAI22_X1 U15237 ( .A1(n13304), .A2(n13135), .B1(n13300), .B2(n13316), .ZN(
        n13567) );
  OAI22_X1 U15238 ( .A1(n13408), .A2(n14558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13044), .ZN(n13045) );
  AOI21_X1 U15239 ( .B1(n13567), .B2(n13137), .A(n13045), .ZN(n13046) );
  OAI211_X1 U15240 ( .C1(n7116), .C2(n14550), .A(n13047), .B(n13046), .ZN(
        P2_U3188) );
  INV_X1 U15241 ( .A(n13254), .ZN(n13288) );
  NOR2_X1 U15242 ( .A1(n13048), .A2(n13288), .ZN(n13050) );
  AOI22_X1 U15243 ( .A1(n13123), .A2(n13133), .B1(n13050), .B2(n13049), .ZN(
        n13060) );
  INV_X1 U15244 ( .A(n13051), .ZN(n13059) );
  INV_X1 U15245 ( .A(n13588), .ZN(n13472) );
  NOR2_X1 U15246 ( .A1(n13472), .A2(n14550), .ZN(n13056) );
  NAND2_X1 U15247 ( .A1(n13258), .A2(n13237), .ZN(n13053) );
  NAND2_X1 U15248 ( .A1(n13254), .A2(n13120), .ZN(n13052) );
  NAND2_X1 U15249 ( .A1(n13053), .A2(n13052), .ZN(n13587) );
  NAND2_X1 U15250 ( .A1(n13587), .A2(n13137), .ZN(n13054) );
  NAND2_X1 U15251 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13230)
         );
  OAI211_X1 U15252 ( .C1(n14558), .C2(n13476), .A(n13054), .B(n13230), .ZN(
        n13055) );
  AOI211_X1 U15253 ( .C1(n13057), .C2(n13133), .A(n13056), .B(n13055), .ZN(
        n13058) );
  OAI21_X1 U15254 ( .B1(n13060), .B2(n13059), .A(n13058), .ZN(P2_U3191) );
  INV_X1 U15255 ( .A(n13061), .ZN(n13063) );
  NAND2_X1 U15256 ( .A1(n13142), .A2(n13066), .ZN(n13068) );
  XNOR2_X1 U15257 ( .A(n13068), .B(n13067), .ZN(n13069) );
  XNOR2_X1 U15258 ( .A(n13336), .B(n13069), .ZN(n13070) );
  AOI22_X1 U15259 ( .A1(n13279), .A2(n13120), .B1(n13141), .B2(n13237), .ZN(
        n13328) );
  AOI22_X1 U15260 ( .A1(n13331), .A2(n13121), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13071) );
  OAI21_X1 U15261 ( .B1(n13328), .B2(n14554), .A(n13071), .ZN(n13072) );
  AOI21_X1 U15262 ( .B1(n13336), .B2(n13128), .A(n13072), .ZN(n13073) );
  XNOR2_X1 U15263 ( .A(n13075), .B(n13074), .ZN(n13079) );
  AOI22_X1 U15264 ( .A1(n13264), .A2(n13237), .B1(n13120), .B2(n13258), .ZN(
        n13434) );
  NOR2_X1 U15265 ( .A1(n13434), .A2(n14554), .ZN(n13077) );
  OAI22_X1 U15266 ( .A1(n14558), .A2(n13443), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15400), .ZN(n13076) );
  AOI211_X1 U15267 ( .C1(n13442), .C2(n13128), .A(n13077), .B(n13076), .ZN(
        n13078) );
  OAI21_X1 U15268 ( .B1(n13079), .B2(n14552), .A(n13078), .ZN(P2_U3195) );
  AOI22_X1 U15269 ( .A1(n13278), .A2(n13237), .B1(n13120), .B2(n13271), .ZN(
        n13373) );
  AOI22_X1 U15270 ( .A1(n13380), .A2(n13121), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13081) );
  OAI21_X1 U15271 ( .B1(n13373), .B2(n14554), .A(n13081), .ZN(n13082) );
  AOI21_X1 U15272 ( .B1(n13379), .B2(n13128), .A(n13082), .ZN(n13083) );
  OAI21_X1 U15273 ( .B1(n13084), .B2(n14552), .A(n13083), .ZN(P2_U3197) );
  INV_X1 U15274 ( .A(n13503), .ZN(n13086) );
  OAI22_X1 U15275 ( .A1(n13288), .A2(n13135), .B1(n13283), .B2(n13316), .ZN(
        n13498) );
  AOI22_X1 U15276 ( .A1(n13498), .A2(n13137), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13085) );
  OAI21_X1 U15277 ( .B1(n13086), .B2(n14558), .A(n13085), .ZN(n13092) );
  AOI22_X1 U15278 ( .A1(n13087), .A2(n13133), .B1(n13111), .B2(n13248), .ZN(
        n13089) );
  NOR3_X1 U15279 ( .A1(n13090), .A2(n13089), .A3(n13088), .ZN(n13091) );
  AOI211_X1 U15280 ( .C1(n13599), .C2(n13128), .A(n13092), .B(n13091), .ZN(
        n13093) );
  OAI21_X1 U15281 ( .B1(n13094), .B2(n14552), .A(n13093), .ZN(P2_U3200) );
  XNOR2_X1 U15282 ( .A(n13096), .B(n13095), .ZN(n13100) );
  AOI22_X1 U15283 ( .A1(n13274), .A2(n13237), .B1(n13120), .B2(n13268), .ZN(
        n13391) );
  AOI22_X1 U15284 ( .A1(n13395), .A2(n13121), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13097) );
  OAI21_X1 U15285 ( .B1(n13391), .B2(n14554), .A(n13097), .ZN(n13098) );
  AOI21_X1 U15286 ( .B1(n13558), .B2(n13128), .A(n13098), .ZN(n13099) );
  OAI21_X1 U15287 ( .B1(n13100), .B2(n14552), .A(n13099), .ZN(P2_U3201) );
  INV_X1 U15288 ( .A(n13101), .ZN(n13103) );
  NOR2_X1 U15289 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  XNOR2_X1 U15290 ( .A(n6755), .B(n13104), .ZN(n13109) );
  NOR2_X1 U15291 ( .A1(n14558), .A2(n13461), .ZN(n13107) );
  AOI22_X1 U15292 ( .A1(n13261), .A2(n13237), .B1(n13120), .B2(n13292), .ZN(
        n13455) );
  OAI22_X1 U15293 ( .A1(n13455), .A2(n14554), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13105), .ZN(n13106) );
  AOI211_X1 U15294 ( .C1(n13457), .C2(n13128), .A(n13107), .B(n13106), .ZN(
        n13108) );
  OAI21_X1 U15295 ( .B1(n13109), .B2(n14552), .A(n13108), .ZN(P2_U3205) );
  INV_X1 U15296 ( .A(n13423), .ZN(n13644) );
  NAND2_X1 U15297 ( .A1(n13110), .A2(n13133), .ZN(n13114) );
  NAND2_X1 U15298 ( .A1(n13264), .A2(n13111), .ZN(n13113) );
  MUX2_X1 U15299 ( .A(n13114), .B(n13113), .S(n13112), .Z(n13119) );
  AOI22_X1 U15300 ( .A1(n13268), .A2(n13237), .B1(n13120), .B2(n13261), .ZN(
        n13417) );
  INV_X1 U15301 ( .A(n13417), .ZN(n13117) );
  OAI22_X1 U15302 ( .A1(n14558), .A2(n13424), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13115), .ZN(n13116) );
  AOI21_X1 U15303 ( .B1(n13117), .B2(n13137), .A(n13116), .ZN(n13118) );
  OAI211_X1 U15304 ( .C1(n13644), .C2(n14550), .A(n13119), .B(n13118), .ZN(
        P2_U3207) );
  AOI22_X1 U15305 ( .A1(n13292), .A2(n13237), .B1(n13120), .B2(n13286), .ZN(
        n13490) );
  NAND2_X1 U15306 ( .A1(n13121), .A2(n13492), .ZN(n13122) );
  NAND2_X1 U15307 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13204)
         );
  OAI211_X1 U15308 ( .C1(n13490), .C2(n14554), .A(n13122), .B(n13204), .ZN(
        n13127) );
  AOI211_X1 U15309 ( .C1(n13125), .C2(n13124), .A(n14552), .B(n13123), .ZN(
        n13126) );
  AOI211_X1 U15310 ( .C1(n13289), .C2(n13128), .A(n13127), .B(n13126), .ZN(
        n13129) );
  INV_X1 U15311 ( .A(n13129), .ZN(P2_U3210) );
  INV_X1 U15312 ( .A(n13547), .ZN(n13365) );
  OAI21_X1 U15313 ( .B1(n13132), .B2(n13131), .A(n13130), .ZN(n13134) );
  NAND2_X1 U15314 ( .A1(n13134), .A2(n13133), .ZN(n13139) );
  OAI22_X1 U15315 ( .A1(n13310), .A2(n13135), .B1(n13306), .B2(n13316), .ZN(
        n13359) );
  OAI22_X1 U15316 ( .A1(n13362), .A2(n14558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15298), .ZN(n13136) );
  AOI21_X1 U15317 ( .B1(n13359), .B2(n13137), .A(n13136), .ZN(n13138) );
  OAI211_X1 U15318 ( .C1(n13365), .C2(n14550), .A(n13139), .B(n13138), .ZN(
        P2_U3212) );
  MUX2_X1 U15319 ( .A(n13239), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13158), .Z(
        P2_U3562) );
  MUX2_X1 U15320 ( .A(n13140), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13158), .Z(
        P2_U3561) );
  MUX2_X1 U15321 ( .A(n13141), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13158), .Z(
        P2_U3560) );
  MUX2_X1 U15322 ( .A(n13142), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13158), .Z(
        P2_U3559) );
  MUX2_X1 U15323 ( .A(n13279), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13158), .Z(
        P2_U3558) );
  MUX2_X1 U15324 ( .A(n13278), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13158), .Z(
        P2_U3557) );
  MUX2_X1 U15325 ( .A(n13274), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13158), .Z(
        P2_U3556) );
  MUX2_X1 U15326 ( .A(n13271), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13158), .Z(
        P2_U3555) );
  MUX2_X1 U15327 ( .A(n13268), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13158), .Z(
        P2_U3554) );
  MUX2_X1 U15328 ( .A(n13264), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13158), .Z(
        P2_U3553) );
  MUX2_X1 U15329 ( .A(n13261), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13158), .Z(
        P2_U3552) );
  MUX2_X1 U15330 ( .A(n13258), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13158), .Z(
        P2_U3551) );
  MUX2_X1 U15331 ( .A(n13292), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13158), .Z(
        P2_U3550) );
  MUX2_X1 U15332 ( .A(n13254), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13158), .Z(
        P2_U3549) );
  INV_X2 U15333 ( .A(P2_U3947), .ZN(n13158) );
  MUX2_X1 U15334 ( .A(n13286), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13158), .Z(
        P2_U3548) );
  MUX2_X1 U15335 ( .A(n13248), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13158), .Z(
        P2_U3547) );
  MUX2_X1 U15336 ( .A(n13143), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13158), .Z(
        P2_U3546) );
  MUX2_X1 U15337 ( .A(n13144), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13158), .Z(
        P2_U3545) );
  MUX2_X1 U15338 ( .A(n13145), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13158), .Z(
        P2_U3544) );
  MUX2_X1 U15339 ( .A(n13146), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13158), .Z(
        P2_U3543) );
  MUX2_X1 U15340 ( .A(n13147), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13158), .Z(
        P2_U3542) );
  MUX2_X1 U15341 ( .A(n13148), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13158), .Z(
        P2_U3541) );
  MUX2_X1 U15342 ( .A(n13149), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13158), .Z(
        P2_U3540) );
  MUX2_X1 U15343 ( .A(n13150), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13158), .Z(
        P2_U3539) );
  MUX2_X1 U15344 ( .A(n13151), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13158), .Z(
        P2_U3538) );
  MUX2_X1 U15345 ( .A(n13152), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13158), .Z(
        P2_U3537) );
  MUX2_X1 U15346 ( .A(n13153), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13158), .Z(
        P2_U3536) );
  MUX2_X1 U15347 ( .A(n13154), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13158), .Z(
        P2_U3535) );
  MUX2_X1 U15348 ( .A(n13155), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13158), .Z(
        P2_U3534) );
  MUX2_X1 U15349 ( .A(n13156), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13158), .Z(
        P2_U3533) );
  MUX2_X1 U15350 ( .A(n13157), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13158), .Z(
        P2_U3532) );
  MUX2_X1 U15351 ( .A(n6917), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13158), .Z(
        P2_U3531) );
  AOI21_X1 U15352 ( .B1(n13161), .B2(n9657), .A(n13160), .ZN(n14830) );
  MUX2_X1 U15353 ( .A(n13162), .B(P2_REG2_REG_13__SCAN_IN), .S(n14833), .Z(
        n14829) );
  NAND2_X1 U15354 ( .A1(n14830), .A2(n14829), .ZN(n14828) );
  OAI21_X1 U15355 ( .B1(n13162), .B2(n14833), .A(n14828), .ZN(n13163) );
  NAND2_X1 U15356 ( .A1(n13171), .A2(n13163), .ZN(n13164) );
  XNOR2_X1 U15357 ( .A(n14845), .B(n13163), .ZN(n14842) );
  NAND2_X1 U15358 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14842), .ZN(n14841) );
  NAND2_X1 U15359 ( .A1(n13164), .A2(n14841), .ZN(n13184) );
  XNOR2_X1 U15360 ( .A(n13184), .B(n13178), .ZN(n13165) );
  NAND2_X1 U15361 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13165), .ZN(n13186) );
  OAI211_X1 U15362 ( .C1(n13165), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14856), 
        .B(n13186), .ZN(n13177) );
  NOR2_X1 U15363 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13166), .ZN(n13167) );
  AOI21_X1 U15364 ( .B1(n14840), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n13167), 
        .ZN(n13176) );
  INV_X1 U15365 ( .A(n14833), .ZN(n13170) );
  OAI21_X1 U15366 ( .B1(n13169), .B2(P2_REG1_REG_12__SCAN_IN), .A(n13168), 
        .ZN(n14824) );
  XOR2_X1 U15367 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14833), .Z(n14825) );
  NOR2_X1 U15368 ( .A1(n14824), .A2(n14825), .ZN(n14823) );
  AOI21_X1 U15369 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n13170), .A(n14823), 
        .ZN(n14837) );
  XNOR2_X1 U15370 ( .A(n13171), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14836) );
  NOR2_X1 U15371 ( .A1(n14837), .A2(n14836), .ZN(n14835) );
  AOI21_X1 U15372 ( .B1(n13172), .B2(n13614), .A(n13180), .ZN(n13173) );
  NAND2_X1 U15373 ( .A1(n13225), .A2(n13173), .ZN(n13175) );
  NAND2_X1 U15374 ( .A1(n14854), .A2(n13185), .ZN(n13174) );
  NAND4_X1 U15375 ( .A1(n13177), .A2(n13176), .A3(n13175), .A4(n13174), .ZN(
        P2_U3229) );
  NOR2_X1 U15376 ( .A1(n13179), .A2(n13178), .ZN(n13181) );
  NOR2_X1 U15377 ( .A1(n13181), .A2(n13180), .ZN(n13183) );
  XNOR2_X1 U15378 ( .A(n13207), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13182) );
  AOI211_X1 U15379 ( .C1(n13183), .C2(n13182), .A(n13206), .B(n14847), .ZN(
        n13197) );
  NAND2_X1 U15380 ( .A1(n13185), .A2(n13184), .ZN(n13187) );
  NAND2_X1 U15381 ( .A1(n13187), .A2(n13186), .ZN(n13191) );
  NOR2_X1 U15382 ( .A1(n13201), .A2(n13188), .ZN(n13189) );
  AOI21_X1 U15383 ( .B1(n13188), .B2(n13201), .A(n13189), .ZN(n13190) );
  NAND2_X1 U15384 ( .A1(n13190), .A2(n13191), .ZN(n13200) );
  OAI211_X1 U15385 ( .C1(n13191), .C2(n13190), .A(n14856), .B(n13200), .ZN(
        n13195) );
  NOR2_X1 U15386 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13192), .ZN(n13193) );
  AOI21_X1 U15387 ( .B1(n14840), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n13193), 
        .ZN(n13194) );
  OAI211_X1 U15388 ( .C1(n14846), .C2(n13201), .A(n13195), .B(n13194), .ZN(
        n13196) );
  OR2_X1 U15389 ( .A1(n13197), .A2(n13196), .ZN(P2_U3230) );
  NOR2_X1 U15390 ( .A1(n13202), .A2(n13198), .ZN(n13199) );
  AOI21_X1 U15391 ( .B1(n13198), .B2(n13202), .A(n13199), .ZN(n14858) );
  OAI21_X1 U15392 ( .B1(n13201), .B2(n13188), .A(n13200), .ZN(n14857) );
  NAND2_X1 U15393 ( .A1(n14858), .A2(n14857), .ZN(n14855) );
  OAI21_X1 U15394 ( .B1(n13198), .B2(n13202), .A(n14855), .ZN(n13217) );
  XNOR2_X1 U15395 ( .A(n13217), .B(n13218), .ZN(n13203) );
  NOR2_X1 U15396 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13203), .ZN(n13220) );
  AOI21_X1 U15397 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13203), .A(n13220), 
        .ZN(n13212) );
  INV_X1 U15398 ( .A(n14840), .ZN(n14861) );
  INV_X1 U15399 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13205) );
  OAI21_X1 U15400 ( .B1(n14861), .B2(n13205), .A(n13204), .ZN(n13210) );
  XNOR2_X1 U15401 ( .A(n14853), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14849) );
  XNOR2_X1 U15402 ( .A(n6703), .B(n13213), .ZN(n13208) );
  NOR2_X1 U15403 ( .A1(n13596), .A2(n13208), .ZN(n13215) );
  AOI211_X1 U15404 ( .C1(n13208), .C2(n13596), .A(n13215), .B(n14847), .ZN(
        n13209) );
  AOI211_X1 U15405 ( .C1(n14854), .C2(n13218), .A(n13210), .B(n13209), .ZN(
        n13211) );
  OAI21_X1 U15406 ( .B1(n13212), .B2(n14802), .A(n13211), .ZN(P2_U3232) );
  NOR2_X1 U15407 ( .A1(n6703), .A2(n13213), .ZN(n13214) );
  NOR2_X1 U15408 ( .A1(n13215), .A2(n13214), .ZN(n13216) );
  XNOR2_X1 U15409 ( .A(n13216), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13226) );
  INV_X1 U15410 ( .A(n13226), .ZN(n13223) );
  NOR2_X1 U15411 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  NOR2_X1 U15412 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  XOR2_X1 U15413 ( .A(n13221), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13224) );
  OAI21_X1 U15414 ( .B1(n13224), .B2(n14802), .A(n14846), .ZN(n13222) );
  AOI21_X1 U15415 ( .B1(n13223), .B2(n13225), .A(n13222), .ZN(n13229) );
  AOI22_X1 U15416 ( .A1(n13226), .A2(n13225), .B1(n14856), .B2(n13224), .ZN(
        n13228) );
  MUX2_X1 U15417 ( .A(n13229), .B(n13228), .S(n13227), .Z(n13231) );
  OAI211_X1 U15418 ( .C1(n7735), .C2(n14861), .A(n13231), .B(n13230), .ZN(
        P2_U3233) );
  INV_X1 U15419 ( .A(n13541), .ZN(n13232) );
  INV_X1 U15420 ( .A(n13442), .ZN(n13648) );
  NAND2_X1 U15421 ( .A1(n13232), .A2(n13361), .ZN(n13348) );
  NAND2_X1 U15422 ( .A1(n13628), .A2(n13317), .ZN(n13242) );
  XNOR2_X1 U15423 ( .A(n13242), .B(n13625), .ZN(n13234) );
  NAND2_X1 U15424 ( .A1(n13234), .A2(n13488), .ZN(n13525) );
  NAND2_X1 U15425 ( .A1(n13235), .A2(P2_B_REG_SCAN_IN), .ZN(n13236) );
  NAND2_X1 U15426 ( .A1(n13237), .A2(n13236), .ZN(n13314) );
  INV_X1 U15427 ( .A(n13314), .ZN(n13238) );
  NAND2_X1 U15428 ( .A1(n13239), .A2(n13238), .ZN(n13528) );
  NOR2_X1 U15429 ( .A1(n13512), .A2(n13528), .ZN(n13244) );
  NOR2_X1 U15430 ( .A1(n13625), .A2(n14868), .ZN(n13240) );
  AOI211_X1 U15431 ( .C1(n13512), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13244), 
        .B(n13240), .ZN(n13241) );
  OAI21_X1 U15432 ( .B1(n13525), .B2(n13411), .A(n13241), .ZN(P2_U3234) );
  OAI211_X1 U15433 ( .C1(n13628), .C2(n13317), .A(n13488), .B(n13242), .ZN(
        n13529) );
  NOR2_X1 U15434 ( .A1(n13471), .A2(n13243), .ZN(n13245) );
  AOI211_X1 U15435 ( .C1(n13246), .C2(n13517), .A(n13245), .B(n13244), .ZN(
        n13247) );
  OAI21_X1 U15436 ( .B1(n13529), .B2(n13411), .A(n13247), .ZN(P2_U3235) );
  NAND2_X1 U15437 ( .A1(n13603), .A2(n13248), .ZN(n13249) );
  OR2_X1 U15438 ( .A1(n13599), .A2(n13286), .ZN(n13251) );
  NAND2_X1 U15439 ( .A1(n13599), .A2(n13286), .ZN(n13252) );
  NAND2_X1 U15440 ( .A1(n13253), .A2(n13252), .ZN(n13485) );
  OR2_X1 U15441 ( .A1(n13289), .A2(n13254), .ZN(n13255) );
  NAND2_X1 U15442 ( .A1(n13588), .A2(n13292), .ZN(n13256) );
  OR2_X1 U15443 ( .A1(n13588), .A2(n13292), .ZN(n13257) );
  NOR2_X1 U15444 ( .A1(n13457), .A2(n13258), .ZN(n13260) );
  INV_X1 U15445 ( .A(n13457), .ZN(n13652) );
  NAND2_X1 U15446 ( .A1(n13442), .A2(n13261), .ZN(n13262) );
  NAND2_X1 U15447 ( .A1(n13263), .A2(n13262), .ZN(n13419) );
  NAND2_X1 U15448 ( .A1(n13419), .A2(n13420), .ZN(n13266) );
  NAND2_X1 U15449 ( .A1(n13423), .A2(n13264), .ZN(n13265) );
  AND2_X1 U15450 ( .A1(n13568), .A2(n13268), .ZN(n13267) );
  OR2_X1 U15451 ( .A1(n13568), .A2(n13268), .ZN(n13269) );
  NAND2_X1 U15452 ( .A1(n13558), .A2(n13271), .ZN(n13272) );
  OR2_X1 U15453 ( .A1(n13379), .A2(n13274), .ZN(n13273) );
  NAND2_X1 U15454 ( .A1(n13379), .A2(n13274), .ZN(n13275) );
  AND2_X1 U15455 ( .A1(n13547), .A2(n13278), .ZN(n13277) );
  NAND2_X1 U15456 ( .A1(n13541), .A2(n13279), .ZN(n13280) );
  NAND2_X1 U15457 ( .A1(n13539), .A2(n13280), .ZN(n13333) );
  NAND2_X1 U15458 ( .A1(n13333), .A2(n13332), .ZN(n13334) );
  AND2_X1 U15459 ( .A1(n13603), .A2(n13283), .ZN(n13282) );
  OR2_X1 U15460 ( .A1(n13603), .A2(n13283), .ZN(n13284) );
  AND2_X1 U15461 ( .A1(n13289), .A2(n13288), .ZN(n13287) );
  OR2_X1 U15462 ( .A1(n13289), .A2(n13288), .ZN(n13290) );
  NAND2_X1 U15463 ( .A1(n13294), .A2(n13293), .ZN(n13295) );
  NAND2_X1 U15464 ( .A1(n13295), .A2(n13432), .ZN(n13297) );
  OR2_X1 U15465 ( .A1(n13442), .A2(n13298), .ZN(n13296) );
  NAND2_X1 U15466 ( .A1(n13442), .A2(n13298), .ZN(n13299) );
  OR2_X1 U15467 ( .A1(n13423), .A2(n13300), .ZN(n13301) );
  OR2_X1 U15468 ( .A1(n13568), .A2(n13302), .ZN(n13303) );
  INV_X1 U15469 ( .A(n13398), .ZN(n13386) );
  NAND2_X1 U15470 ( .A1(n13558), .A2(n13304), .ZN(n13305) );
  INV_X1 U15471 ( .A(n13371), .ZN(n13375) );
  NAND2_X1 U15472 ( .A1(n13379), .A2(n13306), .ZN(n13307) );
  INV_X1 U15473 ( .A(n13354), .ZN(n13342) );
  NAND2_X1 U15474 ( .A1(n13532), .A2(n13471), .ZN(n13324) );
  AOI211_X1 U15475 ( .C1(n13534), .C2(n6664), .A(n13066), .B(n13317), .ZN(
        n13533) );
  INV_X1 U15476 ( .A(n13534), .ZN(n13321) );
  INV_X1 U15477 ( .A(n13318), .ZN(n13319) );
  AOI22_X1 U15478 ( .A1(n13319), .A2(n14864), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13512), .ZN(n13320) );
  OAI21_X1 U15479 ( .B1(n13321), .B2(n14868), .A(n13320), .ZN(n13322) );
  AOI21_X1 U15480 ( .B1(n13533), .B2(n14862), .A(n13322), .ZN(n13323) );
  OAI211_X1 U15481 ( .C1(n13535), .C2(n13507), .A(n13324), .B(n13323), .ZN(
        P2_U3236) );
  NAND2_X1 U15482 ( .A1(n13325), .A2(n13332), .ZN(n13326) );
  NAND3_X1 U15483 ( .A1(n13327), .A2(n13499), .A3(n13326), .ZN(n13329) );
  INV_X1 U15484 ( .A(n13537), .ZN(n13330) );
  AOI21_X1 U15485 ( .B1(n13331), .B2(n14864), .A(n13330), .ZN(n13341) );
  INV_X1 U15486 ( .A(n13538), .ZN(n13339) );
  NAND2_X1 U15487 ( .A1(n13348), .A2(n13336), .ZN(n13335) );
  NAND3_X1 U15488 ( .A1(n6664), .A2(n13488), .A3(n13335), .ZN(n13536) );
  AOI22_X1 U15489 ( .A1(n13336), .A2(n13517), .B1(n13512), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13337) );
  OAI21_X1 U15490 ( .B1(n13536), .B2(n13411), .A(n13337), .ZN(n13338) );
  AOI21_X1 U15491 ( .B1(n13339), .B2(n14872), .A(n13338), .ZN(n13340) );
  OAI21_X1 U15492 ( .B1(n13341), .B2(n13512), .A(n13340), .ZN(P2_U3237) );
  XNOR2_X1 U15493 ( .A(n13343), .B(n13342), .ZN(n13346) );
  INV_X1 U15494 ( .A(n13344), .ZN(n13345) );
  AOI21_X1 U15495 ( .B1(n13346), .B2(n13499), .A(n13345), .ZN(n13544) );
  INV_X1 U15496 ( .A(n13361), .ZN(n13347) );
  AOI21_X1 U15497 ( .B1(n13347), .B2(n13541), .A(n13030), .ZN(n13349) );
  NAND2_X1 U15498 ( .A1(n13349), .A2(n13348), .ZN(n13542) );
  AOI22_X1 U15499 ( .A1(n13350), .A2(n14864), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13512), .ZN(n13352) );
  NAND2_X1 U15500 ( .A1(n13541), .A2(n13517), .ZN(n13351) );
  OAI211_X1 U15501 ( .C1(n13542), .C2(n13411), .A(n13352), .B(n13351), .ZN(
        n13353) );
  INV_X1 U15502 ( .A(n13353), .ZN(n13357) );
  OR2_X1 U15503 ( .A1(n13355), .A2(n13354), .ZN(n13540) );
  NAND3_X1 U15504 ( .A1(n13540), .A2(n14872), .A3(n13539), .ZN(n13356) );
  OAI211_X1 U15505 ( .C1(n13544), .C2(n13512), .A(n13357), .B(n13356), .ZN(
        P2_U3238) );
  XNOR2_X1 U15506 ( .A(n13358), .B(n13367), .ZN(n13360) );
  AOI21_X1 U15507 ( .B1(n13360), .B2(n13499), .A(n13359), .ZN(n13549) );
  AOI211_X1 U15508 ( .C1(n13547), .C2(n13377), .A(n13066), .B(n13361), .ZN(
        n13546) );
  INV_X1 U15509 ( .A(n13362), .ZN(n13363) );
  AOI22_X1 U15510 ( .A1(n13363), .A2(n14864), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13512), .ZN(n13364) );
  OAI21_X1 U15511 ( .B1(n13365), .B2(n14868), .A(n13364), .ZN(n13369) );
  XOR2_X1 U15512 ( .A(n13367), .B(n13366), .Z(n13550) );
  NOR2_X1 U15513 ( .A1(n13550), .A2(n13507), .ZN(n13368) );
  AOI211_X1 U15514 ( .C1(n13546), .C2(n14862), .A(n13369), .B(n13368), .ZN(
        n13370) );
  OAI21_X1 U15515 ( .B1(n13512), .B2(n13549), .A(n13370), .ZN(P2_U3239) );
  XNOR2_X1 U15516 ( .A(n13372), .B(n13371), .ZN(n13374) );
  INV_X1 U15517 ( .A(n13551), .ZN(n13385) );
  XNOR2_X1 U15518 ( .A(n13376), .B(n13375), .ZN(n13553) );
  INV_X1 U15519 ( .A(n13377), .ZN(n13378) );
  AOI211_X1 U15520 ( .C1(n13379), .C2(n13393), .A(n13066), .B(n13378), .ZN(
        n13552) );
  NAND2_X1 U15521 ( .A1(n13552), .A2(n14862), .ZN(n13382) );
  AOI22_X1 U15522 ( .A1(n13380), .A2(n14864), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13512), .ZN(n13381) );
  OAI211_X1 U15523 ( .C1(n7112), .C2(n14868), .A(n13382), .B(n13381), .ZN(
        n13383) );
  AOI21_X1 U15524 ( .B1(n14872), .B2(n13553), .A(n13383), .ZN(n13384) );
  OAI21_X1 U15525 ( .B1(n13385), .B2(n13512), .A(n13384), .ZN(P2_U3240) );
  NAND2_X1 U15526 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  NAND2_X1 U15527 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  NAND2_X1 U15528 ( .A1(n13390), .A2(n13499), .ZN(n13392) );
  NAND2_X1 U15529 ( .A1(n13392), .A2(n13391), .ZN(n13563) );
  AOI21_X1 U15530 ( .B1(n13558), .B2(n13409), .A(n13066), .ZN(n13394) );
  NAND2_X1 U15531 ( .A1(n13394), .A2(n13393), .ZN(n13559) );
  AOI22_X1 U15532 ( .A1(n13395), .A2(n14864), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13512), .ZN(n13397) );
  NAND2_X1 U15533 ( .A1(n13558), .A2(n13517), .ZN(n13396) );
  OAI211_X1 U15534 ( .C1(n13559), .C2(n13411), .A(n13397), .B(n13396), .ZN(
        n13401) );
  NAND2_X1 U15535 ( .A1(n13399), .A2(n13398), .ZN(n13556) );
  AND3_X1 U15536 ( .A1(n13557), .A2(n14872), .A3(n13556), .ZN(n13400) );
  AOI211_X1 U15537 ( .C1(n13563), .C2(n13471), .A(n13401), .B(n13400), .ZN(
        n13402) );
  INV_X1 U15538 ( .A(n13402), .ZN(P2_U3241) );
  XOR2_X1 U15539 ( .A(n13405), .B(n13403), .Z(n13571) );
  OAI211_X1 U15540 ( .C1(n13406), .C2(n13405), .A(n13499), .B(n6836), .ZN(
        n13569) );
  INV_X1 U15541 ( .A(n13567), .ZN(n13407) );
  OAI211_X1 U15542 ( .C1(n13515), .C2(n13408), .A(n13569), .B(n13407), .ZN(
        n13414) );
  AOI211_X1 U15543 ( .C1(n13568), .C2(n13421), .A(n13066), .B(n7115), .ZN(
        n13566) );
  INV_X1 U15544 ( .A(n13566), .ZN(n13412) );
  AOI22_X1 U15545 ( .A1(n13568), .A2(n13517), .B1(n13512), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13410) );
  OAI21_X1 U15546 ( .B1(n13412), .B2(n13411), .A(n13410), .ZN(n13413) );
  AOI21_X1 U15547 ( .B1(n13414), .B2(n13471), .A(n13413), .ZN(n13415) );
  OAI21_X1 U15548 ( .B1(n13571), .B2(n13507), .A(n13415), .ZN(P2_U3242) );
  XNOR2_X1 U15549 ( .A(n13416), .B(n13420), .ZN(n13418) );
  OAI21_X1 U15550 ( .B1(n13418), .B2(n13435), .A(n13417), .ZN(n13572) );
  INV_X1 U15551 ( .A(n13572), .ZN(n13430) );
  XOR2_X1 U15552 ( .A(n13419), .B(n13420), .Z(n13574) );
  INV_X1 U15553 ( .A(n13421), .ZN(n13422) );
  AOI211_X1 U15554 ( .C1(n13423), .C2(n13439), .A(n13066), .B(n13422), .ZN(
        n13573) );
  NAND2_X1 U15555 ( .A1(n13573), .A2(n14862), .ZN(n13427) );
  INV_X1 U15556 ( .A(n13424), .ZN(n13425) );
  AOI22_X1 U15557 ( .A1(n13425), .A2(n14864), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13512), .ZN(n13426) );
  OAI211_X1 U15558 ( .C1(n13644), .C2(n14868), .A(n13427), .B(n13426), .ZN(
        n13428) );
  AOI21_X1 U15559 ( .B1(n13574), .B2(n14872), .A(n13428), .ZN(n13429) );
  OAI21_X1 U15560 ( .B1(n13430), .B2(n13512), .A(n13429), .ZN(P2_U3243) );
  NAND2_X1 U15561 ( .A1(n13475), .A2(n13474), .ZN(n13473) );
  NAND3_X1 U15562 ( .A1(n13473), .A2(n13452), .A3(n6769), .ZN(n13451) );
  NAND2_X1 U15563 ( .A1(n13451), .A2(n13432), .ZN(n13433) );
  XNOR2_X1 U15564 ( .A(n13433), .B(n13438), .ZN(n13436) );
  OAI21_X1 U15565 ( .B1(n13436), .B2(n13435), .A(n13434), .ZN(n13577) );
  INV_X1 U15566 ( .A(n13577), .ZN(n13449) );
  XOR2_X1 U15567 ( .A(n13438), .B(n13437), .Z(n13579) );
  INV_X1 U15568 ( .A(n13460), .ZN(n13441) );
  INV_X1 U15569 ( .A(n13439), .ZN(n13440) );
  AOI211_X1 U15570 ( .C1(n13442), .C2(n13441), .A(n13066), .B(n13440), .ZN(
        n13578) );
  NAND2_X1 U15571 ( .A1(n13578), .A2(n14862), .ZN(n13446) );
  INV_X1 U15572 ( .A(n13443), .ZN(n13444) );
  AOI22_X1 U15573 ( .A1(n13444), .A2(n14864), .B1(n13512), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13445) );
  OAI211_X1 U15574 ( .C1(n13648), .C2(n14868), .A(n13446), .B(n13445), .ZN(
        n13447) );
  AOI21_X1 U15575 ( .B1(n13579), .B2(n14872), .A(n13447), .ZN(n13448) );
  OAI21_X1 U15576 ( .B1(n13449), .B2(n13512), .A(n13448), .ZN(P2_U3244) );
  XOR2_X1 U15577 ( .A(n13450), .B(n13452), .Z(n13584) );
  INV_X1 U15578 ( .A(n13584), .ZN(n13467) );
  INV_X1 U15579 ( .A(n13451), .ZN(n13454) );
  AOI21_X1 U15580 ( .B1(n13473), .B2(n6769), .A(n13452), .ZN(n13453) );
  OAI21_X1 U15581 ( .B1(n13454), .B2(n13453), .A(n13499), .ZN(n13456) );
  NAND2_X1 U15582 ( .A1(n13456), .A2(n13455), .ZN(n13582) );
  NAND2_X1 U15583 ( .A1(n6773), .A2(n13457), .ZN(n13458) );
  NAND2_X1 U15584 ( .A1(n13458), .A2(n13488), .ZN(n13459) );
  NOR2_X1 U15585 ( .A1(n13460), .A2(n13459), .ZN(n13583) );
  NAND2_X1 U15586 ( .A1(n13583), .A2(n14862), .ZN(n13464) );
  INV_X1 U15587 ( .A(n13461), .ZN(n13462) );
  AOI22_X1 U15588 ( .A1(n13512), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13462), 
        .B2(n14864), .ZN(n13463) );
  OAI211_X1 U15589 ( .C1(n13652), .C2(n14868), .A(n13464), .B(n13463), .ZN(
        n13465) );
  AOI21_X1 U15590 ( .B1(n13582), .B2(n13471), .A(n13465), .ZN(n13466) );
  OAI21_X1 U15591 ( .B1(n13467), .B2(n13507), .A(n13466), .ZN(P2_U3245) );
  XNOR2_X1 U15592 ( .A(n13468), .B(n13474), .ZN(n13591) );
  AOI21_X1 U15593 ( .B1(n6682), .B2(n13588), .A(n13066), .ZN(n13469) );
  AND2_X1 U15594 ( .A1(n13469), .A2(n6773), .ZN(n13586) );
  INV_X1 U15595 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13470) );
  OAI22_X1 U15596 ( .A1(n13472), .A2(n14868), .B1(n13471), .B2(n13470), .ZN(
        n13480) );
  OAI211_X1 U15597 ( .C1(n13475), .C2(n13474), .A(n13499), .B(n13473), .ZN(
        n13590) );
  INV_X1 U15598 ( .A(n13476), .ZN(n13477) );
  AOI21_X1 U15599 ( .B1(n13477), .B2(n14864), .A(n13587), .ZN(n13478) );
  AOI21_X1 U15600 ( .B1(n13590), .B2(n13478), .A(n13512), .ZN(n13479) );
  AOI211_X1 U15601 ( .C1(n13586), .C2(n14862), .A(n13480), .B(n13479), .ZN(
        n13481) );
  OAI21_X1 U15602 ( .B1(n13507), .B2(n13591), .A(n13481), .ZN(P2_U3246) );
  XNOR2_X1 U15603 ( .A(n13482), .B(n13484), .ZN(n13483) );
  NAND2_X1 U15604 ( .A1(n13483), .A2(n13499), .ZN(n13595) );
  NAND2_X1 U15605 ( .A1(n13485), .A2(n13484), .ZN(n13486) );
  NAND2_X1 U15606 ( .A1(n13487), .A2(n13486), .ZN(n13593) );
  OAI211_X1 U15607 ( .C1(n13489), .C2(n13656), .A(n6682), .B(n13488), .ZN(
        n13491) );
  NAND2_X1 U15608 ( .A1(n13491), .A2(n13490), .ZN(n13592) );
  NAND2_X1 U15609 ( .A1(n13592), .A2(n14862), .ZN(n13494) );
  AOI22_X1 U15610 ( .A1(n13512), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13492), 
        .B2(n14864), .ZN(n13493) );
  OAI211_X1 U15611 ( .C1(n13656), .C2(n14868), .A(n13494), .B(n13493), .ZN(
        n13495) );
  AOI21_X1 U15612 ( .B1(n13593), .B2(n14872), .A(n13495), .ZN(n13496) );
  OAI21_X1 U15613 ( .B1(n13595), .B2(n13512), .A(n13496), .ZN(P2_U3247) );
  XNOR2_X1 U15614 ( .A(n6916), .B(n13505), .ZN(n13500) );
  AOI21_X1 U15615 ( .B1(n13500), .B2(n13499), .A(n13498), .ZN(n13601) );
  XNOR2_X1 U15616 ( .A(n13501), .B(n13599), .ZN(n13502) );
  NOR2_X1 U15617 ( .A1(n13502), .A2(n13030), .ZN(n13598) );
  AOI22_X1 U15618 ( .A1(n13512), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13503), 
        .B2(n14864), .ZN(n13504) );
  OAI21_X1 U15619 ( .B1(n7111), .B2(n14868), .A(n13504), .ZN(n13509) );
  XNOR2_X1 U15620 ( .A(n13506), .B(n13505), .ZN(n13602) );
  NOR2_X1 U15621 ( .A1(n13602), .A2(n13507), .ZN(n13508) );
  AOI211_X1 U15622 ( .C1(n13598), .C2(n14862), .A(n13509), .B(n13508), .ZN(
        n13510) );
  OAI21_X1 U15623 ( .B1(n13512), .B2(n13601), .A(n13510), .ZN(P2_U3248) );
  NAND2_X1 U15624 ( .A1(n13511), .A2(n13471), .ZN(n13524) );
  NAND2_X1 U15625 ( .A1(n13512), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n13513) );
  OAI21_X1 U15626 ( .B1(n13515), .B2(n13514), .A(n13513), .ZN(n13516) );
  AOI21_X1 U15627 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(n13523) );
  NAND2_X1 U15628 ( .A1(n13519), .A2(n14872), .ZN(n13522) );
  NAND2_X1 U15629 ( .A1(n13520), .A2(n14862), .ZN(n13521) );
  NAND4_X1 U15630 ( .A1(n13524), .A2(n13523), .A3(n13522), .A4(n13521), .ZN(
        P2_U3255) );
  INV_X1 U15631 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13526) );
  AND2_X1 U15632 ( .A1(n13525), .A2(n13528), .ZN(n13622) );
  MUX2_X1 U15633 ( .A(n13526), .B(n13622), .S(n14970), .Z(n13527) );
  AND2_X1 U15634 ( .A1(n13529), .A2(n13528), .ZN(n13626) );
  MUX2_X1 U15635 ( .A(n13530), .B(n13626), .S(n14970), .Z(n13531) );
  OAI21_X1 U15636 ( .B1(n13628), .B2(n13616), .A(n13531), .ZN(P2_U3529) );
  NAND3_X1 U15637 ( .A1(n13540), .A2(n14938), .A3(n13539), .ZN(n13545) );
  NAND2_X1 U15638 ( .A1(n13541), .A2(n14927), .ZN(n13543) );
  NAND4_X1 U15639 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13632) );
  MUX2_X1 U15640 ( .A(n13632), .B(P2_REG1_REG_27__SCAN_IN), .S(n14968), .Z(
        P2_U3526) );
  AOI21_X1 U15641 ( .B1(n14927), .B2(n13547), .A(n13546), .ZN(n13548) );
  OAI211_X1 U15642 ( .C1(n13550), .C2(n14931), .A(n13549), .B(n13548), .ZN(
        n13633) );
  MUX2_X1 U15643 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13633), .S(n14970), .Z(
        P2_U3525) );
  INV_X1 U15644 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13554) );
  MUX2_X1 U15645 ( .A(n13554), .B(n13634), .S(n14970), .Z(n13555) );
  OAI21_X1 U15646 ( .B1(n7112), .B2(n13616), .A(n13555), .ZN(P2_U3524) );
  INV_X1 U15647 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13564) );
  NAND3_X1 U15648 ( .A1(n13557), .A2(n13556), .A3(n14938), .ZN(n13561) );
  NAND2_X1 U15649 ( .A1(n13558), .A2(n14927), .ZN(n13560) );
  NAND3_X1 U15650 ( .A1(n13561), .A2(n13560), .A3(n13559), .ZN(n13562) );
  NOR2_X1 U15651 ( .A1(n13563), .A2(n13562), .ZN(n13637) );
  MUX2_X1 U15652 ( .A(n13564), .B(n13637), .S(n14970), .Z(n13565) );
  INV_X1 U15653 ( .A(n13565), .ZN(P2_U3523) );
  AOI211_X1 U15654 ( .C1(n14927), .C2(n13568), .A(n13567), .B(n13566), .ZN(
        n13570) );
  OAI211_X1 U15655 ( .C1(n13571), .C2(n14931), .A(n13570), .B(n13569), .ZN(
        n13640) );
  MUX2_X1 U15656 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13640), .S(n14970), .Z(
        P2_U3522) );
  INV_X1 U15657 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13575) );
  AOI211_X1 U15658 ( .C1(n14938), .C2(n13574), .A(n13573), .B(n13572), .ZN(
        n13641) );
  MUX2_X1 U15659 ( .A(n13575), .B(n13641), .S(n14970), .Z(n13576) );
  OAI21_X1 U15660 ( .B1(n13644), .B2(n13616), .A(n13576), .ZN(P2_U3521) );
  INV_X1 U15661 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13580) );
  AOI211_X1 U15662 ( .C1(n14938), .C2(n13579), .A(n13578), .B(n13577), .ZN(
        n13645) );
  MUX2_X1 U15663 ( .A(n13580), .B(n13645), .S(n14970), .Z(n13581) );
  OAI21_X1 U15664 ( .B1(n13648), .B2(n13616), .A(n13581), .ZN(P2_U3520) );
  INV_X1 U15665 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n15475) );
  AOI211_X1 U15666 ( .C1(n14938), .C2(n13584), .A(n13583), .B(n13582), .ZN(
        n13649) );
  MUX2_X1 U15667 ( .A(n15475), .B(n13649), .S(n14970), .Z(n13585) );
  OAI21_X1 U15668 ( .B1(n13652), .B2(n13616), .A(n13585), .ZN(P2_U3519) );
  AOI211_X1 U15669 ( .C1(n14927), .C2(n13588), .A(n13587), .B(n13586), .ZN(
        n13589) );
  OAI211_X1 U15670 ( .C1(n14931), .C2(n13591), .A(n13590), .B(n13589), .ZN(
        n13653) );
  MUX2_X1 U15671 ( .A(n13653), .B(P2_REG1_REG_19__SCAN_IN), .S(n14968), .Z(
        P2_U3518) );
  AOI21_X1 U15672 ( .B1(n13593), .B2(n14938), .A(n13592), .ZN(n13594) );
  AND2_X1 U15673 ( .A1(n13595), .A2(n13594), .ZN(n13654) );
  MUX2_X1 U15674 ( .A(n13596), .B(n13654), .S(n14970), .Z(n13597) );
  OAI21_X1 U15675 ( .B1(n13656), .B2(n13616), .A(n13597), .ZN(P2_U3517) );
  AOI21_X1 U15676 ( .B1(n14927), .B2(n13599), .A(n13598), .ZN(n13600) );
  OAI211_X1 U15677 ( .C1(n14931), .C2(n13602), .A(n13601), .B(n13600), .ZN(
        n13657) );
  MUX2_X1 U15678 ( .A(n13657), .B(P2_REG1_REG_17__SCAN_IN), .S(n14968), .Z(
        P2_U3516) );
  NAND2_X1 U15679 ( .A1(n13603), .A2(n14927), .ZN(n13604) );
  OAI211_X1 U15680 ( .C1(n13606), .C2(n14931), .A(n13605), .B(n13604), .ZN(
        n13607) );
  OR2_X1 U15681 ( .A1(n13608), .A2(n13607), .ZN(n13658) );
  MUX2_X1 U15682 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13658), .S(n14970), .Z(
        P2_U3515) );
  NOR2_X1 U15683 ( .A1(n13609), .A2(n14931), .ZN(n13613) );
  NOR4_X1 U15684 ( .A1(n13613), .A2(n13612), .A3(n13611), .A4(n13610), .ZN(
        n13659) );
  MUX2_X1 U15685 ( .A(n13614), .B(n13659), .S(n14970), .Z(n13615) );
  OAI21_X1 U15686 ( .B1(n13663), .B2(n13616), .A(n13615), .ZN(P2_U3514) );
  AOI21_X1 U15687 ( .B1(n14927), .B2(n13618), .A(n13617), .ZN(n13619) );
  OAI211_X1 U15688 ( .C1(n14931), .C2(n13621), .A(n13620), .B(n13619), .ZN(
        n13664) );
  MUX2_X1 U15689 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13664), .S(n14970), .Z(
        P2_U3512) );
  MUX2_X1 U15690 ( .A(n13623), .B(n13622), .S(n14960), .Z(n13624) );
  OAI21_X1 U15691 ( .B1(n13625), .B2(n13662), .A(n13624), .ZN(P2_U3498) );
  MUX2_X1 U15692 ( .A(n15423), .B(n13626), .S(n14960), .Z(n13627) );
  OAI21_X1 U15693 ( .B1(n13628), .B2(n13662), .A(n13627), .ZN(P2_U3497) );
  MUX2_X1 U15694 ( .A(n13632), .B(P2_REG0_REG_27__SCAN_IN), .S(n14959), .Z(
        P2_U3494) );
  MUX2_X1 U15695 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13633), .S(n14960), .Z(
        P2_U3493) );
  MUX2_X1 U15696 ( .A(n13635), .B(n13634), .S(n14960), .Z(n13636) );
  OAI21_X1 U15697 ( .B1(n7112), .B2(n13662), .A(n13636), .ZN(P2_U3492) );
  MUX2_X1 U15698 ( .A(n13638), .B(n13637), .S(n14960), .Z(n13639) );
  INV_X1 U15699 ( .A(n13639), .ZN(P2_U3491) );
  MUX2_X1 U15700 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13640), .S(n14960), .Z(
        P2_U3490) );
  MUX2_X1 U15701 ( .A(n13642), .B(n13641), .S(n14960), .Z(n13643) );
  OAI21_X1 U15702 ( .B1(n13644), .B2(n13662), .A(n13643), .ZN(P2_U3489) );
  MUX2_X1 U15703 ( .A(n13646), .B(n13645), .S(n14960), .Z(n13647) );
  OAI21_X1 U15704 ( .B1(n13648), .B2(n13662), .A(n13647), .ZN(P2_U3488) );
  INV_X1 U15705 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13650) );
  MUX2_X1 U15706 ( .A(n13650), .B(n13649), .S(n14960), .Z(n13651) );
  OAI21_X1 U15707 ( .B1(n13652), .B2(n13662), .A(n13651), .ZN(P2_U3487) );
  MUX2_X1 U15708 ( .A(n13653), .B(P2_REG0_REG_19__SCAN_IN), .S(n14959), .Z(
        P2_U3486) );
  MUX2_X1 U15709 ( .A(n15516), .B(n13654), .S(n14960), .Z(n13655) );
  OAI21_X1 U15710 ( .B1(n13656), .B2(n13662), .A(n13655), .ZN(P2_U3484) );
  MUX2_X1 U15711 ( .A(n13657), .B(P2_REG0_REG_17__SCAN_IN), .S(n14959), .Z(
        P2_U3481) );
  MUX2_X1 U15712 ( .A(n13658), .B(P2_REG0_REG_16__SCAN_IN), .S(n14959), .Z(
        P2_U3478) );
  INV_X1 U15713 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13660) );
  MUX2_X1 U15714 ( .A(n13660), .B(n13659), .S(n14960), .Z(n13661) );
  OAI21_X1 U15715 ( .B1(n13663), .B2(n13662), .A(n13661), .ZN(P2_U3475) );
  MUX2_X1 U15716 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13664), .S(n14960), .Z(
        P2_U3469) );
  INV_X1 U15717 ( .A(n13665), .ZN(n14363) );
  NOR4_X1 U15718 ( .A1(n13666), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8652), .A4(
        P2_U3088), .ZN(n13667) );
  AOI21_X1 U15719 ( .B1(n13677), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13667), 
        .ZN(n13668) );
  OAI21_X1 U15720 ( .B1(n14363), .B2(n13675), .A(n13668), .ZN(P2_U3296) );
  INV_X1 U15721 ( .A(n13669), .ZN(n14365) );
  OAI222_X1 U15722 ( .A1(n13675), .A2(n14365), .B1(P2_U3088), .B2(n13670), 
        .C1(n13671), .C2(n13681), .ZN(P2_U3297) );
  INV_X1 U15723 ( .A(n13672), .ZN(n14367) );
  OAI222_X1 U15724 ( .A1(n13675), .A2(n14367), .B1(P2_U3088), .B2(n13674), 
        .C1(n13673), .C2(n13681), .ZN(P2_U3298) );
  AOI21_X1 U15725 ( .B1(n13677), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13676), 
        .ZN(n13678) );
  OAI21_X1 U15726 ( .B1(n13679), .B2(n13675), .A(n13678), .ZN(P2_U3299) );
  INV_X1 U15727 ( .A(n13680), .ZN(n14372) );
  OAI222_X1 U15728 ( .A1(P2_U3088), .A2(n13683), .B1(n13675), .B2(n14372), 
        .C1(n13682), .C2(n13681), .ZN(P2_U3301) );
  INV_X1 U15729 ( .A(n13684), .ZN(n13685) );
  MUX2_X1 U15730 ( .A(n13685), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U15731 ( .A(n13687), .B(n13686), .ZN(n13688) );
  NAND2_X1 U15732 ( .A1(n13688), .A2(n14567), .ZN(n13693) );
  INV_X1 U15733 ( .A(n13989), .ZN(n13689) );
  AOI22_X1 U15734 ( .A1(n13778), .A2(n13689), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13690) );
  OAI21_X1 U15735 ( .B1(n13806), .B2(n14219), .A(n13690), .ZN(n13691) );
  AOI21_X1 U15736 ( .B1(n14577), .B2(n13822), .A(n13691), .ZN(n13692) );
  OAI211_X1 U15737 ( .C1(n14327), .C2(n14581), .A(n13693), .B(n13692), .ZN(
        P1_U3214) );
  XOR2_X1 U15738 ( .A(n13695), .B(n13694), .Z(n13702) );
  NAND2_X1 U15739 ( .A1(n14087), .A2(n14262), .ZN(n13697) );
  NAND2_X1 U15740 ( .A1(n14020), .A2(n14591), .ZN(n13696) );
  NAND2_X1 U15741 ( .A1(n13697), .A2(n13696), .ZN(n14050) );
  AOI22_X1 U15742 ( .A1(n13818), .A2(n14050), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13698) );
  OAI21_X1 U15743 ( .B1(n14054), .B2(n14588), .A(n13698), .ZN(n13699) );
  AOI21_X1 U15744 ( .B1(n13700), .B2(n13798), .A(n13699), .ZN(n13701) );
  OAI21_X1 U15745 ( .B1(n13702), .B2(n14574), .A(n13701), .ZN(P1_U3216) );
  AND2_X1 U15746 ( .A1(n13704), .A2(n13703), .ZN(n13707) );
  OAI211_X1 U15747 ( .C1(n13707), .C2(n13706), .A(n14567), .B(n13705), .ZN(
        n13711) );
  AOI22_X1 U15748 ( .A1(n14577), .A2(n14196), .B1(n13798), .B2(n7320), .ZN(
        n13710) );
  MUX2_X1 U15749 ( .A(n14588), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13709) );
  NAND2_X1 U15750 ( .A1(n14579), .A2(n13831), .ZN(n13708) );
  NAND4_X1 U15751 ( .A1(n13711), .A2(n13710), .A3(n13709), .A4(n13708), .ZN(
        P1_U3218) );
  AOI21_X1 U15752 ( .B1(n13713), .B2(n13712), .A(n14574), .ZN(n13715) );
  NAND2_X1 U15753 ( .A1(n13715), .A2(n13714), .ZN(n13719) );
  OAI22_X1 U15754 ( .A1(n13920), .A2(n14141), .B1(n13915), .B2(n14609), .ZN(
        n14124) );
  NOR2_X1 U15755 ( .A1(n13716), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13894) );
  NOR2_X1 U15756 ( .A1(n14588), .A2(n14126), .ZN(n13717) );
  AOI211_X1 U15757 ( .C1(n14124), .C2(n13818), .A(n13894), .B(n13717), .ZN(
        n13718) );
  OAI211_X1 U15758 ( .C1(n14347), .C2(n14581), .A(n13719), .B(n13718), .ZN(
        P1_U3219) );
  INV_X1 U15759 ( .A(n13720), .ZN(n13721) );
  AOI21_X1 U15760 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n13729) );
  INV_X1 U15761 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13724) );
  OAI22_X1 U15762 ( .A1(n14588), .A2(n14101), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13724), .ZN(n13725) );
  AOI21_X1 U15763 ( .B1(n14577), .B2(n14088), .A(n13725), .ZN(n13726) );
  OAI21_X1 U15764 ( .B1(n13945), .B2(n13806), .A(n13726), .ZN(n13727) );
  AOI21_X1 U15765 ( .B1(n14100), .B2(n13798), .A(n13727), .ZN(n13728) );
  OAI21_X1 U15766 ( .B1(n13729), .B2(n14574), .A(n13728), .ZN(P1_U3223) );
  XNOR2_X1 U15767 ( .A(n13731), .B(n13730), .ZN(n13732) );
  NAND2_X1 U15768 ( .A1(n13732), .A2(n14567), .ZN(n13737) );
  INV_X1 U15769 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13733) );
  OAI22_X1 U15770 ( .A1(n14588), .A2(n14022), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13733), .ZN(n13735) );
  NOR2_X1 U15771 ( .A1(n13806), .A2(n14021), .ZN(n13734) );
  AOI211_X1 U15772 ( .C1(n14577), .C2(n14020), .A(n13735), .B(n13734), .ZN(
        n13736) );
  OAI211_X1 U15773 ( .C1(n14332), .C2(n14581), .A(n13737), .B(n13736), .ZN(
        P1_U3225) );
  XOR2_X1 U15774 ( .A(n13739), .B(n13738), .Z(n13745) );
  INV_X1 U15775 ( .A(n14173), .ZN(n14140) );
  NAND2_X1 U15776 ( .A1(n14577), .A2(n14590), .ZN(n13742) );
  AOI21_X1 U15777 ( .B1(n13778), .B2(n14176), .A(n13740), .ZN(n13741) );
  OAI211_X1 U15778 ( .C1(n14140), .C2(n13806), .A(n13742), .B(n13741), .ZN(
        n13743) );
  AOI21_X1 U15779 ( .B1(n14300), .B2(n13798), .A(n13743), .ZN(n13744) );
  OAI21_X1 U15780 ( .B1(n13745), .B2(n14574), .A(n13744), .ZN(P1_U3226) );
  XNOR2_X1 U15781 ( .A(n6866), .B(n13746), .ZN(n13748) );
  NAND2_X1 U15782 ( .A1(n13748), .A2(n14567), .ZN(n13753) );
  OAI21_X1 U15783 ( .B1(n14588), .B2(n14161), .A(n13749), .ZN(n13751) );
  NOR2_X1 U15784 ( .A1(n13806), .A2(n13915), .ZN(n13750) );
  AOI211_X1 U15785 ( .C1(n14577), .C2(n14159), .A(n13751), .B(n13750), .ZN(
        n13752) );
  OAI211_X1 U15786 ( .C1(n14292), .C2(n14581), .A(n13753), .B(n13752), .ZN(
        P1_U3228) );
  XOR2_X1 U15787 ( .A(n13755), .B(n13754), .Z(n13761) );
  OR2_X1 U15788 ( .A1(n14609), .A2(n13924), .ZN(n13757) );
  NAND2_X1 U15789 ( .A1(n13999), .A2(n14591), .ZN(n13756) );
  NAND2_X1 U15790 ( .A1(n13757), .A2(n13756), .ZN(n14037) );
  AOI22_X1 U15791 ( .A1(n13818), .A2(n14037), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13758) );
  OAI21_X1 U15792 ( .B1(n14040), .B2(n14588), .A(n13758), .ZN(n13759) );
  AOI21_X1 U15793 ( .B1(n14045), .B2(n13798), .A(n13759), .ZN(n13760) );
  OAI21_X1 U15794 ( .B1(n13761), .B2(n14574), .A(n13760), .ZN(P1_U3229) );
  OAI211_X1 U15795 ( .C1(n13764), .C2(n13763), .A(n13762), .B(n14567), .ZN(
        n13769) );
  INV_X1 U15796 ( .A(n14115), .ZN(n13767) );
  AOI22_X1 U15797 ( .A1(n13823), .A2(n14262), .B1(n14591), .B2(n14261), .ZN(
        n14270) );
  OAI22_X1 U15798 ( .A1(n14270), .A2(n13776), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13765), .ZN(n13766) );
  AOI21_X1 U15799 ( .B1(n13767), .B2(n13778), .A(n13766), .ZN(n13768) );
  OAI211_X1 U15800 ( .C1(n14272), .C2(n14581), .A(n13769), .B(n13768), .ZN(
        P1_U3233) );
  OAI211_X1 U15801 ( .C1(n13771), .C2(n13770), .A(n14560), .B(n14567), .ZN(
        n13781) );
  INV_X1 U15802 ( .A(n14514), .ZN(n13779) );
  OR2_X1 U15803 ( .A1(n13772), .A2(n14141), .ZN(n13775) );
  OR2_X1 U15804 ( .A1(n14609), .A2(n13773), .ZN(n13774) );
  AND2_X1 U15805 ( .A1(n13775), .A2(n13774), .ZN(n14617) );
  OAI22_X1 U15806 ( .A1(n13776), .A2(n14617), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15476), .ZN(n13777) );
  AOI21_X1 U15807 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(n13780) );
  OAI211_X1 U15808 ( .C1(n14619), .C2(n14581), .A(n13781), .B(n13780), .ZN(
        P1_U3234) );
  OAI21_X1 U15809 ( .B1(n13784), .B2(n13783), .A(n13782), .ZN(n13785) );
  NAND2_X1 U15810 ( .A1(n13785), .A2(n14567), .ZN(n13790) );
  INV_X1 U15811 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13786) );
  OAI22_X1 U15812 ( .A1(n14588), .A2(n14077), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13786), .ZN(n13788) );
  NOR2_X1 U15813 ( .A1(n13806), .A2(n13924), .ZN(n13787) );
  AOI211_X1 U15814 ( .C1(n14577), .C2(n14261), .A(n13788), .B(n13787), .ZN(
        n13789) );
  OAI211_X1 U15815 ( .C1(n14581), .C2(n13791), .A(n13790), .B(n13789), .ZN(
        P1_U3235) );
  XOR2_X1 U15816 ( .A(n13793), .B(n13792), .Z(n13800) );
  INV_X1 U15817 ( .A(n13823), .ZN(n14142) );
  OAI21_X1 U15818 ( .B1(n14588), .B2(n14143), .A(n13794), .ZN(n13795) );
  AOI21_X1 U15819 ( .B1(n14577), .B2(n14173), .A(n13795), .ZN(n13796) );
  OAI21_X1 U15820 ( .B1(n14142), .B2(n13806), .A(n13796), .ZN(n13797) );
  AOI21_X1 U15821 ( .B1(n7628), .B2(n13798), .A(n13797), .ZN(n13799) );
  OAI21_X1 U15822 ( .B1(n13800), .B2(n14574), .A(n13799), .ZN(P1_U3238) );
  XNOR2_X1 U15823 ( .A(n13802), .B(n13801), .ZN(n13803) );
  INV_X1 U15824 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13804) );
  OAI22_X1 U15825 ( .A1(n14588), .A2(n14008), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13804), .ZN(n13808) );
  NOR2_X1 U15826 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  AOI211_X1 U15827 ( .C1(n14577), .C2(n13999), .A(n13808), .B(n13807), .ZN(
        n13809) );
  OAI21_X1 U15828 ( .B1(n13812), .B2(n13811), .A(n13810), .ZN(n13813) );
  NAND2_X1 U15829 ( .A1(n13813), .A2(n14567), .ZN(n13820) );
  NAND2_X1 U15830 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14671)
         );
  INV_X1 U15831 ( .A(n14671), .ZN(n13816) );
  NOR2_X1 U15832 ( .A1(n14588), .A2(n13814), .ZN(n13815) );
  AOI211_X1 U15833 ( .C1(n13818), .C2(n13817), .A(n13816), .B(n13815), .ZN(
        n13819) );
  OAI211_X1 U15834 ( .C1(n14355), .C2(n14581), .A(n13820), .B(n13819), .ZN(
        P1_U3241) );
  MUX2_X1 U15835 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13900), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15836 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13951), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15837 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13821), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15838 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13948), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15839 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14000), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15840 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13822), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15841 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13999), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15842 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14020), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14076), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15844 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14087), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15845 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14261), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15846 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14088), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15847 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13823), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15848 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14160), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15849 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14173), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15850 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14159), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15851 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14590), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15852 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13824), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15853 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14564), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15854 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14578), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15855 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13825), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15856 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14576), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15857 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13826), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15858 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13827), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15859 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13828), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13829), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15861 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13830), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15862 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13831), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15863 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13832), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15864 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14196), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15865 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14192), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15866 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14195), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U15867 ( .A1(n14673), .A2(n14379), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13833), .ZN(n13834) );
  AOI21_X1 U15868 ( .B1(n13835), .B2(n14665), .A(n13834), .ZN(n13844) );
  OAI211_X1 U15869 ( .C1(n13838), .C2(n13837), .A(n14668), .B(n13836), .ZN(
        n13843) );
  OAI211_X1 U15870 ( .C1(n13841), .C2(n13840), .A(n14669), .B(n13839), .ZN(
        n13842) );
  NAND3_X1 U15871 ( .A1(n13844), .A2(n13843), .A3(n13842), .ZN(P1_U3244) );
  OAI211_X1 U15872 ( .C1(n13847), .C2(n13846), .A(n14668), .B(n13845), .ZN(
        n13857) );
  INV_X1 U15873 ( .A(n13864), .ZN(n13852) );
  NAND3_X1 U15874 ( .A1(n13850), .A2(n13849), .A3(n13848), .ZN(n13851) );
  NAND3_X1 U15875 ( .A1(n14669), .A2(n13852), .A3(n13851), .ZN(n13856) );
  NAND2_X1 U15876 ( .A1(n14665), .A2(n13853), .ZN(n13855) );
  AOI22_X1 U15877 ( .A1(n14656), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13854) );
  NAND4_X1 U15878 ( .A1(n13857), .A2(n13856), .A3(n13855), .A4(n13854), .ZN(
        P1_U3246) );
  AOI21_X1 U15879 ( .B1(n14656), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n13858), .ZN(
        n13873) );
  XOR2_X1 U15880 ( .A(n13860), .B(n13859), .Z(n13869) );
  INV_X1 U15881 ( .A(n13861), .ZN(n13866) );
  NOR3_X1 U15882 ( .A1(n13864), .A2(n13863), .A3(n13862), .ZN(n13865) );
  NOR3_X1 U15883 ( .A1(n13867), .A2(n13866), .A3(n13865), .ZN(n13868) );
  AOI21_X1 U15884 ( .B1(n14668), .B2(n13869), .A(n13868), .ZN(n13872) );
  NAND2_X1 U15885 ( .A1(n14665), .A2(n13870), .ZN(n13871) );
  NAND4_X1 U15886 ( .A1(n13874), .A2(n13873), .A3(n13872), .A4(n13871), .ZN(
        P1_U3247) );
  NAND2_X1 U15887 ( .A1(n13876), .A2(n13875), .ZN(n13880) );
  INV_X1 U15888 ( .A(n13877), .ZN(n13878) );
  NAND2_X1 U15889 ( .A1(n13878), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U15890 ( .A1(n13880), .A2(n13879), .ZN(n13881) );
  XOR2_X1 U15891 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13881), .Z(n13890) );
  INV_X1 U15892 ( .A(n13890), .ZN(n13888) );
  NOR2_X1 U15893 ( .A1(n13883), .A2(n13882), .ZN(n13884) );
  XNOR2_X1 U15894 ( .A(n13884), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13889) );
  OAI21_X1 U15895 ( .B1(n13889), .B2(n13886), .A(n13885), .ZN(n13887) );
  AOI21_X1 U15896 ( .B1(n13888), .B2(n14669), .A(n13887), .ZN(n13893) );
  AOI22_X1 U15897 ( .A1(n13890), .A2(n14669), .B1(n14668), .B2(n13889), .ZN(
        n13892) );
  MUX2_X1 U15898 ( .A(n13893), .B(n13892), .S(n13891), .Z(n13896) );
  INV_X1 U15899 ( .A(n13894), .ZN(n13895) );
  OAI211_X1 U15900 ( .C1(n7734), .C2(n14673), .A(n13896), .B(n13895), .ZN(
        P1_U3262) );
  NAND2_X1 U15901 ( .A1(n14097), .A2(n14342), .ZN(n14098) );
  NAND2_X1 U15902 ( .A1(n14007), .A2(n14027), .ZN(n14004) );
  XNOR2_X1 U15903 ( .A(n14314), .B(n13904), .ZN(n13897) );
  NAND2_X1 U15904 ( .A1(n13897), .A2(n14504), .ZN(n14210) );
  NOR2_X1 U15905 ( .A1(n14653), .A2(n13898), .ZN(n13899) );
  NOR2_X1 U15906 ( .A1(n14141), .A2(n13899), .ZN(n13952) );
  NAND2_X1 U15907 ( .A1(n13952), .A2(n13900), .ZN(n14212) );
  NOR2_X1 U15908 ( .A1(n14177), .A2(n14212), .ZN(n13907) );
  AOI21_X1 U15909 ( .B1(n14689), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13907), 
        .ZN(n13903) );
  NAND2_X1 U15910 ( .A1(n13901), .A2(n14201), .ZN(n13902) );
  OAI211_X1 U15911 ( .C1(n14210), .C2(n14130), .A(n13903), .B(n13902), .ZN(
        P1_U3263) );
  OAI211_X1 U15912 ( .C1(n14318), .C2(n13905), .A(n14504), .B(n13904), .ZN(
        n14213) );
  NOR2_X1 U15913 ( .A1(n14318), .A2(n14180), .ZN(n13906) );
  AOI211_X1 U15914 ( .C1(n14689), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13907), 
        .B(n13906), .ZN(n13908) );
  OAI21_X1 U15915 ( .B1(n14130), .B2(n14213), .A(n13908), .ZN(P1_U3264) );
  OR2_X1 U15916 ( .A1(n13910), .A2(n14590), .ZN(n13911) );
  AND2_X1 U15917 ( .A1(n14147), .A2(n13915), .ZN(n13916) );
  NAND2_X1 U15918 ( .A1(n13918), .A2(n13917), .ZN(n14112) );
  OR2_X1 U15919 ( .A1(n14272), .A2(n13920), .ZN(n14091) );
  AND2_X1 U15920 ( .A1(n14090), .A2(n14091), .ZN(n13921) );
  OR2_X1 U15921 ( .A1(n14263), .A2(n14087), .ZN(n13922) );
  OR2_X1 U15922 ( .A1(n14337), .A2(n13924), .ZN(n13925) );
  NOR2_X1 U15923 ( .A1(n14045), .A2(n14020), .ZN(n13926) );
  NAND2_X1 U15924 ( .A1(n14014), .A2(n6647), .ZN(n14016) );
  NAND2_X1 U15925 ( .A1(n14030), .A2(n13999), .ZN(n13927) );
  NAND2_X1 U15926 ( .A1(n14016), .A2(n13927), .ZN(n13995) );
  NAND2_X1 U15927 ( .A1(n13995), .A2(n13994), .ZN(n13929) );
  OR2_X1 U15928 ( .A1(n14007), .A2(n14021), .ZN(n13928) );
  INV_X1 U15929 ( .A(n13983), .ZN(n13930) );
  OR2_X1 U15930 ( .A1(n14000), .A2(n13991), .ZN(n13931) );
  NAND2_X1 U15931 ( .A1(n13937), .A2(n13936), .ZN(n14169) );
  OR2_X1 U15932 ( .A1(n14181), .A2(n14159), .ZN(n13938) );
  OR2_X1 U15933 ( .A1(n14158), .A2(n14140), .ZN(n13939) );
  OR2_X2 U15934 ( .A1(n14150), .A2(n14149), .ZN(n14286) );
  NAND2_X1 U15935 ( .A1(n14286), .A2(n13940), .ZN(n14121) );
  OR2_X2 U15936 ( .A1(n14121), .A2(n7627), .ZN(n14123) );
  NAND2_X1 U15937 ( .A1(n14133), .A2(n14142), .ZN(n13942) );
  NAND2_X1 U15938 ( .A1(n14272), .A2(n14088), .ZN(n13943) );
  INV_X1 U15939 ( .A(n14090), .ZN(n14085) );
  NAND2_X1 U15940 ( .A1(n14342), .A2(n14261), .ZN(n13944) );
  NAND2_X1 U15941 ( .A1(n14084), .A2(n13944), .ZN(n14071) );
  OR2_X2 U15942 ( .A1(n14071), .A2(n14070), .ZN(n14073) );
  NAND2_X1 U15943 ( .A1(n14263), .A2(n13945), .ZN(n13946) );
  INV_X1 U15944 ( .A(n14045), .ZN(n14252) );
  NOR2_X1 U15945 ( .A1(n14323), .A2(n13948), .ZN(n13949) );
  NAND2_X1 U15946 ( .A1(n14222), .A2(n14510), .ZN(n13963) );
  NAND2_X1 U15947 ( .A1(n14686), .A2(n14262), .ZN(n14594) );
  NAND2_X1 U15948 ( .A1(n13952), .A2(n13951), .ZN(n14217) );
  OAI22_X1 U15949 ( .A1(n13954), .A2(n14217), .B1(n14683), .B2(n13953), .ZN(
        n13955) );
  AOI21_X1 U15950 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14689), .A(n13955), 
        .ZN(n13956) );
  OAI21_X1 U15951 ( .B1(n14594), .B2(n14219), .A(n13956), .ZN(n13960) );
  INV_X1 U15952 ( .A(n13971), .ZN(n13958) );
  OAI211_X1 U15953 ( .C1(n14321), .C2(n13958), .A(n14504), .B(n13957), .ZN(
        n14218) );
  NOR2_X1 U15954 ( .A1(n14218), .A2(n14130), .ZN(n13959) );
  AOI211_X1 U15955 ( .C1(n14201), .C2(n13961), .A(n13960), .B(n13959), .ZN(
        n13962) );
  OAI211_X1 U15956 ( .C1(n14216), .C2(n14153), .A(n13963), .B(n13962), .ZN(
        P1_U3356) );
  XNOR2_X1 U15957 ( .A(n13966), .B(n13965), .ZN(n14229) );
  NAND2_X1 U15958 ( .A1(n14229), .A2(n14510), .ZN(n13976) );
  INV_X1 U15959 ( .A(n13967), .ZN(n13968) );
  AOI22_X1 U15960 ( .A1(n14686), .A2(n14224), .B1(n13968), .B2(n14199), .ZN(
        n13969) );
  OAI21_X1 U15961 ( .B1(n13970), .B2(n14686), .A(n13969), .ZN(n13973) );
  OAI211_X1 U15962 ( .C1(n14323), .C2(n13978), .A(n14504), .B(n13971), .ZN(
        n14225) );
  NOR2_X1 U15963 ( .A1(n14225), .A2(n14130), .ZN(n13972) );
  AOI211_X1 U15964 ( .C1(n14201), .C2(n13974), .A(n13973), .B(n13972), .ZN(
        n13975) );
  OAI211_X1 U15965 ( .C1(n14153), .C2(n14227), .A(n13976), .B(n13975), .ZN(
        P1_U3265) );
  AND2_X1 U15966 ( .A1(n13991), .A2(n14004), .ZN(n13977) );
  INV_X1 U15967 ( .A(n13981), .ZN(n13979) );
  OAI22_X1 U15968 ( .A1(n13980), .A2(n14704), .B1(n13979), .B2(n14289), .ZN(
        n13985) );
  INV_X1 U15969 ( .A(n13980), .ZN(n13982) );
  OAI22_X1 U15970 ( .A1(n13982), .A2(n14704), .B1(n14289), .B2(n13981), .ZN(
        n13984) );
  MUX2_X1 U15971 ( .A(n13985), .B(n13984), .S(n13983), .Z(n13987) );
  OAI22_X1 U15972 ( .A1(n14021), .A2(n14609), .B1(n14219), .B2(n14141), .ZN(
        n13986) );
  OR2_X1 U15973 ( .A1(n14232), .A2(n14689), .ZN(n13993) );
  NAND2_X1 U15974 ( .A1(n14177), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n13988) );
  OAI21_X1 U15975 ( .B1(n13989), .B2(n14683), .A(n13988), .ZN(n13990) );
  AOI21_X1 U15976 ( .B1(n13991), .B2(n14201), .A(n13990), .ZN(n13992) );
  OAI211_X1 U15977 ( .C1(n14130), .C2(n14231), .A(n13993), .B(n13992), .ZN(
        P1_U3266) );
  XNOR2_X1 U15978 ( .A(n13995), .B(n13994), .ZN(n14239) );
  XNOR2_X1 U15979 ( .A(n13997), .B(n13996), .ZN(n13998) );
  NAND2_X1 U15980 ( .A1(n13998), .A2(n14592), .ZN(n14237) );
  INV_X1 U15981 ( .A(n14237), .ZN(n14003) );
  NAND2_X1 U15982 ( .A1(n13999), .A2(n14262), .ZN(n14002) );
  NAND2_X1 U15983 ( .A1(n14000), .A2(n14591), .ZN(n14001) );
  NAND2_X1 U15984 ( .A1(n14002), .A2(n14001), .ZN(n14235) );
  OAI21_X1 U15985 ( .B1(n14003), .B2(n14235), .A(n14686), .ZN(n14013) );
  INV_X1 U15986 ( .A(n14027), .ZN(n14006) );
  INV_X1 U15987 ( .A(n14004), .ZN(n14005) );
  AOI211_X1 U15988 ( .C1(n14236), .C2(n14006), .A(n14719), .B(n14005), .ZN(
        n14234) );
  NOR2_X1 U15989 ( .A1(n14007), .A2(n14180), .ZN(n14011) );
  OAI22_X1 U15990 ( .A1(n14686), .A2(n14009), .B1(n14008), .B2(n14683), .ZN(
        n14010) );
  AOI211_X1 U15991 ( .C1(n14234), .C2(n14606), .A(n14011), .B(n14010), .ZN(
        n14012) );
  OAI211_X1 U15992 ( .C1(n14239), .C2(n14153), .A(n14013), .B(n14012), .ZN(
        P1_U3267) );
  OR2_X1 U15993 ( .A1(n14014), .A2(n6647), .ZN(n14015) );
  NAND2_X1 U15994 ( .A1(n14016), .A2(n14015), .ZN(n14240) );
  OAI21_X1 U15995 ( .B1(n14019), .B2(n14018), .A(n14017), .ZN(n14246) );
  NAND2_X1 U15996 ( .A1(n14246), .A2(n14510), .ZN(n14032) );
  INV_X1 U15997 ( .A(n14020), .ZN(n14243) );
  OR2_X1 U15998 ( .A1(n14021), .A2(n14141), .ZN(n14241) );
  OAI22_X1 U15999 ( .A1(n14689), .A2(n14241), .B1(n14022), .B2(n14683), .ZN(
        n14023) );
  AOI21_X1 U16000 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14689), .A(n14023), 
        .ZN(n14024) );
  OAI21_X1 U16001 ( .B1(n14243), .B2(n14594), .A(n14024), .ZN(n14029) );
  NAND2_X1 U16002 ( .A1(n14030), .A2(n6685), .ZN(n14025) );
  NAND2_X1 U16003 ( .A1(n14025), .A2(n14504), .ZN(n14026) );
  OR2_X1 U16004 ( .A1(n14027), .A2(n14026), .ZN(n14242) );
  NOR2_X1 U16005 ( .A1(n14242), .A2(n14130), .ZN(n14028) );
  AOI211_X1 U16006 ( .C1(n14201), .C2(n14030), .A(n14029), .B(n14028), .ZN(
        n14031) );
  OAI211_X1 U16007 ( .C1(n14240), .C2(n14153), .A(n14032), .B(n14031), .ZN(
        P1_U3268) );
  XNOR2_X1 U16008 ( .A(n14033), .B(n14034), .ZN(n14249) );
  INV_X1 U16009 ( .A(n14249), .ZN(n14048) );
  XNOR2_X1 U16010 ( .A(n14035), .B(n14034), .ZN(n14036) );
  NAND2_X1 U16011 ( .A1(n14036), .A2(n14592), .ZN(n14039) );
  INV_X1 U16012 ( .A(n14037), .ZN(n14038) );
  NAND2_X1 U16013 ( .A1(n14039), .A2(n14038), .ZN(n14254) );
  NAND2_X1 U16014 ( .A1(n14254), .A2(n14686), .ZN(n14047) );
  OAI22_X1 U16015 ( .A1(n14686), .A2(n14041), .B1(n14040), .B2(n14683), .ZN(
        n14044) );
  AOI21_X1 U16016 ( .B1(n14045), .B2(n14053), .A(n14719), .ZN(n14042) );
  NAND2_X1 U16017 ( .A1(n14042), .A2(n6685), .ZN(n14250) );
  NOR2_X1 U16018 ( .A1(n14250), .A2(n14130), .ZN(n14043) );
  AOI211_X1 U16019 ( .C1(n14201), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n14046) );
  OAI211_X1 U16020 ( .C1(n14048), .C2(n14153), .A(n14047), .B(n14046), .ZN(
        P1_U3269) );
  XNOR2_X1 U16021 ( .A(n14049), .B(n14058), .ZN(n14051) );
  AOI21_X1 U16022 ( .B1(n14051), .B2(n14592), .A(n14050), .ZN(n14258) );
  OR2_X1 U16023 ( .A1(n14337), .A2(n14065), .ZN(n14052) );
  AND3_X1 U16024 ( .A1(n14053), .A2(n14504), .A3(n14052), .ZN(n14255) );
  OAI22_X1 U16025 ( .A1(n14686), .A2(n14055), .B1(n14054), .B2(n14683), .ZN(
        n14057) );
  NOR2_X1 U16026 ( .A1(n14337), .A2(n14180), .ZN(n14056) );
  AOI211_X1 U16027 ( .C1(n14255), .C2(n14606), .A(n14057), .B(n14056), .ZN(
        n14063) );
  NAND2_X1 U16028 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  NAND2_X1 U16029 ( .A1(n14256), .A2(n14605), .ZN(n14062) );
  OAI211_X1 U16030 ( .C1(n14258), .C2(n14689), .A(n14063), .B(n14062), .ZN(
        P1_U3270) );
  AND2_X1 U16031 ( .A1(n14263), .A2(n14098), .ZN(n14064) );
  OR3_X1 U16032 ( .A1(n14065), .A2(n14064), .A3(n14719), .ZN(n14264) );
  INV_X1 U16033 ( .A(n14070), .ZN(n14067) );
  NAND3_X1 U16034 ( .A1(n14089), .A2(n14067), .A3(n14066), .ZN(n14068) );
  AOI21_X1 U16035 ( .B1(n14069), .B2(n14068), .A(n14289), .ZN(n14075) );
  NAND2_X1 U16036 ( .A1(n14071), .A2(n14070), .ZN(n14072) );
  AOI21_X1 U16037 ( .B1(n14073), .B2(n14072), .A(n14704), .ZN(n14074) );
  AOI211_X1 U16038 ( .C1(n14591), .C2(n14076), .A(n14075), .B(n14074), .ZN(
        n14266) );
  OR2_X1 U16039 ( .A1(n14266), .A2(n14689), .ZN(n14083) );
  NOR2_X1 U16040 ( .A1(n14683), .A2(n14077), .ZN(n14078) );
  AOI21_X1 U16041 ( .B1(n14689), .B2(P1_REG2_REG_22__SCAN_IN), .A(n14078), 
        .ZN(n14079) );
  OAI21_X1 U16042 ( .B1(n14594), .B2(n14080), .A(n14079), .ZN(n14081) );
  AOI21_X1 U16043 ( .B1(n14263), .B2(n14201), .A(n14081), .ZN(n14082) );
  OAI211_X1 U16044 ( .C1(n14264), .C2(n14130), .A(n14083), .B(n14082), .ZN(
        P1_U3271) );
  OAI211_X1 U16045 ( .C1(n14086), .C2(n14085), .A(n14084), .B(n14592), .ZN(
        n14096) );
  AOI22_X1 U16046 ( .A1(n14088), .A2(n14262), .B1(n14591), .B2(n14087), .ZN(
        n14095) );
  INV_X1 U16047 ( .A(n14089), .ZN(n14093) );
  AOI21_X1 U16048 ( .B1(n14110), .B2(n14091), .A(n14090), .ZN(n14092) );
  OAI21_X1 U16049 ( .B1(n14093), .B2(n14092), .A(n14725), .ZN(n14094) );
  NAND3_X1 U16050 ( .A1(n14096), .A2(n14095), .A3(n14094), .ZN(n14267) );
  INV_X1 U16051 ( .A(n14267), .ZN(n14107) );
  INV_X1 U16052 ( .A(n14097), .ZN(n14114) );
  INV_X1 U16053 ( .A(n14098), .ZN(n14099) );
  AOI21_X1 U16054 ( .B1(n14100), .B2(n14114), .A(n14099), .ZN(n14268) );
  NOR2_X1 U16055 ( .A1(n14342), .A2(n14180), .ZN(n14104) );
  OAI22_X1 U16056 ( .A1(n14686), .A2(n14102), .B1(n14101), .B2(n14683), .ZN(
        n14103) );
  AOI211_X1 U16057 ( .C1(n14268), .C2(n14105), .A(n14104), .B(n14103), .ZN(
        n14106) );
  OAI21_X1 U16058 ( .B1(n14107), .B2(n14689), .A(n14106), .ZN(P1_U3272) );
  OAI21_X1 U16059 ( .B1(n14109), .B2(n14113), .A(n14108), .ZN(n14276) );
  INV_X1 U16060 ( .A(n14110), .ZN(n14111) );
  AOI21_X1 U16061 ( .B1(n14113), .B2(n14112), .A(n14111), .ZN(n14274) );
  OAI211_X1 U16062 ( .C1(n14272), .C2(n14129), .A(n14114), .B(n14504), .ZN(
        n14271) );
  OAI22_X1 U16063 ( .A1(n14270), .A2(n14689), .B1(n14115), .B2(n14683), .ZN(
        n14117) );
  NOR2_X1 U16064 ( .A1(n14272), .A2(n14180), .ZN(n14116) );
  AOI211_X1 U16065 ( .C1(n14689), .C2(P1_REG2_REG_20__SCAN_IN), .A(n14117), 
        .B(n14116), .ZN(n14118) );
  OAI21_X1 U16066 ( .B1(n14271), .B2(n14130), .A(n14118), .ZN(n14119) );
  AOI21_X1 U16067 ( .B1(n14274), .B2(n14605), .A(n14119), .ZN(n14120) );
  OAI21_X1 U16068 ( .B1(n14188), .B2(n14276), .A(n14120), .ZN(P1_U3273) );
  NAND2_X1 U16069 ( .A1(n14121), .A2(n7627), .ZN(n14122) );
  NAND2_X1 U16070 ( .A1(n14123), .A2(n14122), .ZN(n14125) );
  AOI21_X1 U16071 ( .B1(n14125), .B2(n14592), .A(n14124), .ZN(n14278) );
  OAI22_X1 U16072 ( .A1(n14686), .A2(n14127), .B1(n14126), .B2(n14683), .ZN(
        n14132) );
  OAI21_X1 U16073 ( .B1(n14347), .B2(n14138), .A(n14504), .ZN(n14128) );
  OR2_X1 U16074 ( .A1(n14129), .A2(n14128), .ZN(n14277) );
  NOR2_X1 U16075 ( .A1(n14277), .A2(n14130), .ZN(n14131) );
  AOI211_X1 U16076 ( .C1(n14201), .C2(n14133), .A(n14132), .B(n14131), .ZN(
        n14136) );
  XNOR2_X1 U16077 ( .A(n14134), .B(n7627), .ZN(n14279) );
  OR2_X1 U16078 ( .A1(n14279), .A2(n14153), .ZN(n14135) );
  OAI211_X1 U16079 ( .C1(n14278), .C2(n14177), .A(n14136), .B(n14135), .ZN(
        P1_U3274) );
  XOR2_X1 U16080 ( .A(n14149), .B(n14137), .Z(n14290) );
  OAI21_X1 U16081 ( .B1(n14157), .B2(n14147), .A(n14504), .ZN(n14139) );
  NOR2_X1 U16082 ( .A1(n14139), .A2(n14138), .ZN(n14282) );
  OAI22_X1 U16083 ( .A1(n14142), .A2(n14141), .B1(n14140), .B2(n14609), .ZN(
        n14283) );
  INV_X1 U16084 ( .A(n14143), .ZN(n14144) );
  AOI22_X1 U16085 ( .A1(n14283), .A2(n14686), .B1(n14144), .B2(n14199), .ZN(
        n14146) );
  NAND2_X1 U16086 ( .A1(n14177), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14145) );
  OAI211_X1 U16087 ( .C1(n14147), .C2(n14180), .A(n14146), .B(n14145), .ZN(
        n14148) );
  AOI21_X1 U16088 ( .B1(n14282), .B2(n14606), .A(n14148), .ZN(n14152) );
  NAND2_X1 U16089 ( .A1(n14150), .A2(n14149), .ZN(n14285) );
  NAND3_X1 U16090 ( .A1(n14286), .A2(n14285), .A3(n14510), .ZN(n14151) );
  OAI211_X1 U16091 ( .C1(n14290), .C2(n14153), .A(n14152), .B(n14151), .ZN(
        P1_U3275) );
  XOR2_X1 U16092 ( .A(n14156), .B(n14154), .Z(n14297) );
  XOR2_X1 U16093 ( .A(n14156), .B(n14155), .Z(n14295) );
  AOI211_X1 U16094 ( .C1(n14158), .C2(n14170), .A(n14719), .B(n14157), .ZN(
        n14294) );
  NAND2_X1 U16095 ( .A1(n14294), .A2(n14606), .ZN(n14164) );
  AOI22_X1 U16096 ( .A1(n14160), .A2(n14591), .B1(n14262), .B2(n14159), .ZN(
        n14291) );
  OAI22_X1 U16097 ( .A1(n14291), .A2(n14689), .B1(n14161), .B2(n14683), .ZN(
        n14162) );
  AOI21_X1 U16098 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14689), .A(n14162), 
        .ZN(n14163) );
  OAI211_X1 U16099 ( .C1(n14292), .C2(n14180), .A(n14164), .B(n14163), .ZN(
        n14165) );
  AOI21_X1 U16100 ( .B1(n14295), .B2(n14605), .A(n14165), .ZN(n14166) );
  OAI21_X1 U16101 ( .B1(n14297), .B2(n14188), .A(n14166), .ZN(P1_U3276) );
  INV_X1 U16102 ( .A(n14167), .ZN(n14168) );
  AOI21_X1 U16103 ( .B1(n14184), .B2(n14169), .A(n14168), .ZN(n14304) );
  INV_X1 U16104 ( .A(n14170), .ZN(n14171) );
  AOI211_X1 U16105 ( .C1(n14300), .C2(n14172), .A(n14719), .B(n14171), .ZN(
        n14298) );
  NAND2_X1 U16106 ( .A1(n14173), .A2(n14591), .ZN(n14175) );
  NAND2_X1 U16107 ( .A1(n14590), .A2(n14262), .ZN(n14174) );
  NAND2_X1 U16108 ( .A1(n14175), .A2(n14174), .ZN(n14299) );
  AOI22_X1 U16109 ( .A1(n14686), .A2(n14299), .B1(n14176), .B2(n14199), .ZN(
        n14179) );
  NAND2_X1 U16110 ( .A1(n14177), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14178) );
  OAI211_X1 U16111 ( .C1(n14181), .C2(n14180), .A(n14179), .B(n14178), .ZN(
        n14182) );
  AOI21_X1 U16112 ( .B1(n14298), .B2(n14606), .A(n14182), .ZN(n14187) );
  OAI21_X1 U16113 ( .B1(n14185), .B2(n14184), .A(n14183), .ZN(n14301) );
  NAND2_X1 U16114 ( .A1(n14301), .A2(n14605), .ZN(n14186) );
  OAI211_X1 U16115 ( .C1(n14304), .C2(n14188), .A(n14187), .B(n14186), .ZN(
        P1_U3277) );
  NOR2_X1 U16116 ( .A1(n14694), .A2(n14189), .ZN(n14190) );
  NOR2_X1 U16117 ( .A1(n14191), .A2(n14190), .ZN(n14205) );
  XOR2_X1 U16118 ( .A(n14192), .B(n14205), .Z(n14194) );
  INV_X1 U16119 ( .A(n14193), .ZN(n14204) );
  MUX2_X1 U16120 ( .A(n14194), .B(n14204), .S(n14195), .Z(n14197) );
  AOI222_X1 U16121 ( .A1(n14592), .A2(n14197), .B1(n14196), .B2(n14591), .C1(
        n14195), .C2(n14262), .ZN(n14695) );
  MUX2_X1 U16122 ( .A(n14198), .B(n14695), .S(n14686), .Z(n14209) );
  AOI22_X1 U16123 ( .A1(n14201), .A2(n14200), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14199), .ZN(n14208) );
  OAI21_X1 U16124 ( .B1(n14204), .B2(n14203), .A(n14202), .ZN(n14698) );
  INV_X1 U16125 ( .A(n14205), .ZN(n14206) );
  NOR2_X1 U16126 ( .A1(n14206), .A2(n14719), .ZN(n14692) );
  AOI22_X1 U16127 ( .A1(n14605), .A2(n14698), .B1(n14606), .B2(n14692), .ZN(
        n14207) );
  NAND3_X1 U16128 ( .A1(n14209), .A2(n14208), .A3(n14207), .ZN(P1_U3292) );
  AND2_X1 U16129 ( .A1(n14210), .A2(n14212), .ZN(n14311) );
  MUX2_X1 U16130 ( .A(n15450), .B(n14311), .S(n14741), .Z(n14211) );
  OAI21_X1 U16131 ( .B1(n14314), .B2(n14309), .A(n14211), .ZN(P1_U3559) );
  INV_X1 U16132 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14214) );
  AND2_X1 U16133 ( .A1(n14213), .A2(n14212), .ZN(n14315) );
  MUX2_X1 U16134 ( .A(n14214), .B(n14315), .S(n14741), .Z(n14215) );
  OAI21_X1 U16135 ( .B1(n14318), .B2(n14309), .A(n14215), .ZN(P1_U3558) );
  NOR2_X1 U16136 ( .A1(n14216), .A2(n14289), .ZN(n14221) );
  OAI211_X1 U16137 ( .C1(n14219), .C2(n14609), .A(n14218), .B(n14217), .ZN(
        n14220) );
  OAI21_X1 U16138 ( .B1(n14321), .B2(n14309), .A(n14223), .ZN(P1_U3557) );
  INV_X1 U16139 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n14230) );
  INV_X1 U16140 ( .A(n14224), .ZN(n14226) );
  OAI211_X1 U16141 ( .C1(n14227), .C2(n14289), .A(n14226), .B(n14225), .ZN(
        n14228) );
  AOI21_X1 U16142 ( .B1(n14229), .B2(n14592), .A(n14228), .ZN(n14322) );
  MUX2_X1 U16143 ( .A(n15350), .B(n14324), .S(n14741), .Z(n14233) );
  OAI21_X1 U16144 ( .B1(n14327), .B2(n14309), .A(n14233), .ZN(P1_U3555) );
  AOI211_X1 U16145 ( .C1(n14236), .C2(n14729), .A(n14235), .B(n14234), .ZN(
        n14238) );
  OAI211_X1 U16146 ( .C1(n14239), .C2(n14289), .A(n14238), .B(n14237), .ZN(
        n14328) );
  MUX2_X1 U16147 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14328), .S(n14741), .Z(
        P1_U3554) );
  INV_X1 U16148 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n14247) );
  NOR2_X1 U16149 ( .A1(n14240), .A2(n14289), .ZN(n14245) );
  OAI211_X1 U16150 ( .C1(n14243), .C2(n14609), .A(n14242), .B(n14241), .ZN(
        n14244) );
  AOI211_X1 U16151 ( .C1(n14246), .C2(n14592), .A(n14245), .B(n14244), .ZN(
        n14329) );
  MUX2_X1 U16152 ( .A(n14247), .B(n14329), .S(n14741), .Z(n14248) );
  OAI21_X1 U16153 ( .B1(n14332), .B2(n14309), .A(n14248), .ZN(P1_U3553) );
  NAND2_X1 U16154 ( .A1(n14249), .A2(n14725), .ZN(n14251) );
  OAI211_X1 U16155 ( .C1(n14252), .C2(n14717), .A(n14251), .B(n14250), .ZN(
        n14253) );
  MUX2_X1 U16156 ( .A(n14333), .B(P1_REG1_REG_24__SCAN_IN), .S(n14739), .Z(
        P1_U3552) );
  AOI21_X1 U16157 ( .B1(n14256), .B2(n14725), .A(n14255), .ZN(n14257) );
  AND2_X1 U16158 ( .A1(n14258), .A2(n14257), .ZN(n14334) );
  MUX2_X1 U16159 ( .A(n14259), .B(n14334), .S(n14741), .Z(n14260) );
  OAI21_X1 U16160 ( .B1(n14337), .B2(n14309), .A(n14260), .ZN(P1_U3551) );
  AOI22_X1 U16161 ( .A1(n14263), .A2(n14729), .B1(n14262), .B2(n14261), .ZN(
        n14265) );
  NAND3_X1 U16162 ( .A1(n14266), .A2(n14265), .A3(n14264), .ZN(n14338) );
  MUX2_X1 U16163 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14338), .S(n14741), .Z(
        P1_U3550) );
  AOI21_X1 U16164 ( .B1(n14504), .B2(n14268), .A(n14267), .ZN(n14339) );
  MUX2_X1 U16165 ( .A(n15517), .B(n14339), .S(n14741), .Z(n14269) );
  OAI21_X1 U16166 ( .B1(n14342), .B2(n14309), .A(n14269), .ZN(P1_U3549) );
  OAI211_X1 U16167 ( .C1(n14272), .C2(n14717), .A(n14271), .B(n14270), .ZN(
        n14273) );
  AOI21_X1 U16168 ( .B1(n14274), .B2(n14725), .A(n14273), .ZN(n14275) );
  OAI21_X1 U16169 ( .B1(n14704), .B2(n14276), .A(n14275), .ZN(n14343) );
  MUX2_X1 U16170 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14343), .S(n14741), .Z(
        P1_U3548) );
  OAI211_X1 U16171 ( .C1(n14279), .C2(n14289), .A(n14278), .B(n14277), .ZN(
        n14344) );
  MUX2_X1 U16172 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14344), .S(n14741), .Z(
        n14280) );
  INV_X1 U16173 ( .A(n14280), .ZN(n14281) );
  OAI21_X1 U16174 ( .B1(n14347), .B2(n14309), .A(n14281), .ZN(P1_U3547) );
  AOI211_X1 U16175 ( .C1(n7628), .C2(n14729), .A(n14283), .B(n14282), .ZN(
        n14288) );
  NAND3_X1 U16176 ( .A1(n14286), .A2(n14592), .A3(n14285), .ZN(n14287) );
  OAI211_X1 U16177 ( .C1(n14290), .C2(n14289), .A(n14288), .B(n14287), .ZN(
        n14348) );
  MUX2_X1 U16178 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14348), .S(n14741), .Z(
        P1_U3546) );
  OAI21_X1 U16179 ( .B1(n14292), .B2(n14717), .A(n14291), .ZN(n14293) );
  AOI211_X1 U16180 ( .C1(n14295), .C2(n14725), .A(n14294), .B(n14293), .ZN(
        n14296) );
  OAI21_X1 U16181 ( .B1(n14297), .B2(n14704), .A(n14296), .ZN(n14349) );
  MUX2_X1 U16182 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14349), .S(n14741), .Z(
        P1_U3545) );
  AOI211_X1 U16183 ( .C1(n14300), .C2(n14729), .A(n14299), .B(n14298), .ZN(
        n14303) );
  NAND2_X1 U16184 ( .A1(n14301), .A2(n14725), .ZN(n14302) );
  OAI211_X1 U16185 ( .C1(n14304), .C2(n14704), .A(n14303), .B(n14302), .ZN(
        n14350) );
  MUX2_X1 U16186 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14350), .S(n14741), .Z(
        P1_U3544) );
  AOI211_X1 U16187 ( .C1(n14725), .C2(n14307), .A(n14306), .B(n14305), .ZN(
        n14351) );
  MUX2_X1 U16188 ( .A(n10801), .B(n14351), .S(n14741), .Z(n14308) );
  OAI21_X1 U16189 ( .B1(n14355), .B2(n14309), .A(n14308), .ZN(P1_U3543) );
  MUX2_X1 U16190 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14310), .S(n14741), .Z(
        P1_U3528) );
  INV_X1 U16191 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14312) );
  MUX2_X1 U16192 ( .A(n14312), .B(n14311), .S(n14733), .Z(n14313) );
  OAI21_X1 U16193 ( .B1(n14314), .B2(n14354), .A(n14313), .ZN(P1_U3527) );
  MUX2_X1 U16194 ( .A(n14316), .B(n14315), .S(n14733), .Z(n14317) );
  OAI21_X1 U16195 ( .B1(n14318), .B2(n14354), .A(n14317), .ZN(P1_U3526) );
  INV_X1 U16196 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n14320) );
  INV_X1 U16197 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14325) );
  MUX2_X1 U16198 ( .A(n14325), .B(n14324), .S(n14733), .Z(n14326) );
  OAI21_X1 U16199 ( .B1(n14327), .B2(n14354), .A(n14326), .ZN(P1_U3523) );
  MUX2_X1 U16200 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14328), .S(n14733), .Z(
        P1_U3522) );
  MUX2_X1 U16201 ( .A(n14330), .B(n14329), .S(n14733), .Z(n14331) );
  OAI21_X1 U16202 ( .B1(n14332), .B2(n14354), .A(n14331), .ZN(P1_U3521) );
  MUX2_X1 U16203 ( .A(n14333), .B(P1_REG0_REG_24__SCAN_IN), .S(n14731), .Z(
        P1_U3520) );
  INV_X1 U16204 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14335) );
  MUX2_X1 U16205 ( .A(n14335), .B(n14334), .S(n14733), .Z(n14336) );
  OAI21_X1 U16206 ( .B1(n14337), .B2(n14354), .A(n14336), .ZN(P1_U3519) );
  MUX2_X1 U16207 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14338), .S(n14733), .Z(
        P1_U3518) );
  INV_X1 U16208 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14340) );
  MUX2_X1 U16209 ( .A(n14340), .B(n14339), .S(n14733), .Z(n14341) );
  OAI21_X1 U16210 ( .B1(n14342), .B2(n14354), .A(n14341), .ZN(P1_U3517) );
  MUX2_X1 U16211 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14343), .S(n14733), .Z(
        P1_U3516) );
  MUX2_X1 U16212 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14344), .S(n14733), .Z(
        n14345) );
  INV_X1 U16213 ( .A(n14345), .ZN(n14346) );
  OAI21_X1 U16214 ( .B1(n14347), .B2(n14354), .A(n14346), .ZN(P1_U3515) );
  MUX2_X1 U16215 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14348), .S(n14733), .Z(
        P1_U3513) );
  MUX2_X1 U16216 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14349), .S(n14733), .Z(
        P1_U3510) );
  MUX2_X1 U16217 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14350), .S(n14733), .Z(
        P1_U3507) );
  INV_X1 U16218 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14352) );
  MUX2_X1 U16219 ( .A(n14352), .B(n14351), .S(n14733), .Z(n14353) );
  OAI21_X1 U16220 ( .B1(n14355), .B2(n14354), .A(n14353), .ZN(P1_U3504) );
  NAND4_X1 U16221 ( .A1(n14357), .A2(n14356), .A3(P1_IR_REG_31__SCAN_IN), .A4(
        P1_STATE_REG_SCAN_IN), .ZN(n14359) );
  OAI22_X1 U16222 ( .A1(n14360), .A2(n14359), .B1(n14358), .B2(n14370), .ZN(
        n14361) );
  INV_X1 U16223 ( .A(n14361), .ZN(n14362) );
  OAI21_X1 U16224 ( .B1(n14363), .B2(n14373), .A(n14362), .ZN(P1_U3324) );
  OAI222_X1 U16225 ( .A1(n14373), .A2(n14365), .B1(n8172), .B2(P1_U3086), .C1(
        n14364), .C2(n14370), .ZN(P1_U3325) );
  OAI222_X1 U16226 ( .A1(n14373), .A2(n14367), .B1(n8173), .B2(P1_U3086), .C1(
        n14366), .C2(n14370), .ZN(P1_U3326) );
  OAI222_X1 U16227 ( .A1(n14653), .A2(P1_U3086), .B1(n14373), .B2(n14369), 
        .C1(n14368), .C2(n14370), .ZN(P1_U3328) );
  OAI222_X1 U16228 ( .A1(P1_U3086), .A2(n14374), .B1(n14373), .B2(n14372), 
        .C1(n14371), .C2(n14370), .ZN(P1_U3329) );
  MUX2_X1 U16229 ( .A(n14376), .B(n14375), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16230 ( .A(n14377), .ZN(n14378) );
  MUX2_X1 U16231 ( .A(n14378), .B(n14654), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  NOR2_X1 U16232 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14473), .ZN(n14472) );
  INV_X1 U16233 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14674) );
  NOR2_X1 U16234 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14674), .ZN(n14409) );
  INV_X1 U16235 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14408) );
  XNOR2_X1 U16236 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14408), .ZN(n14469) );
  INV_X1 U16237 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14406) );
  INV_X1 U16238 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14401) );
  INV_X1 U16239 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14419) );
  INV_X1 U16240 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14396) );
  XNOR2_X1 U16241 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14422) );
  INV_X1 U16242 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14394) );
  INV_X1 U16243 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16244 ( .A1(n14381), .A2(n15343), .ZN(n14383) );
  NOR2_X1 U16245 ( .A1(n14386), .A2(n15435), .ZN(n14388) );
  AND2_X1 U16246 ( .A1(n15486), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14389) );
  NOR2_X1 U16247 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14390), .ZN(n14392) );
  XNOR2_X1 U16248 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14390), .ZN(n14450) );
  INV_X1 U16249 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14449) );
  XNOR2_X1 U16250 ( .A(n14394), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U16251 ( .A1(n14422), .A2(n14421), .ZN(n14395) );
  NAND2_X1 U16252 ( .A1(n14419), .A2(n14418), .ZN(n14398) );
  NOR2_X1 U16253 ( .A1(n14419), .A2(n14418), .ZN(n14397) );
  XNOR2_X1 U16254 ( .A(n14401), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14462) );
  XNOR2_X1 U16255 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n14417) );
  NAND2_X1 U16256 ( .A1(n14416), .A2(n14417), .ZN(n14402) );
  OAI21_X1 U16257 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14403), .A(n14402), 
        .ZN(n14404) );
  INV_X1 U16258 ( .A(n14404), .ZN(n14414) );
  AND2_X1 U16259 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14406), .ZN(n14405) );
  OAI22_X1 U16260 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14410), .B1(n14409), 
        .B2(n14413), .ZN(n14475) );
  NAND2_X1 U16261 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14473), .ZN(n14411) );
  OAI21_X1 U16262 ( .B1(n14472), .B2(n14475), .A(n14411), .ZN(n14476) );
  XOR2_X1 U16263 ( .A(n10596), .B(n14476), .Z(n14477) );
  XNOR2_X1 U16264 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14477), .ZN(n14516) );
  XOR2_X1 U16265 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n14412) );
  XOR2_X1 U16266 ( .A(n14413), .B(n14412), .Z(n14644) );
  XNOR2_X1 U16267 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n14415) );
  XNOR2_X1 U16268 ( .A(n14415), .B(n14414), .ZN(n14636) );
  XOR2_X1 U16269 ( .A(n14417), .B(n14416), .Z(n14464) );
  XNOR2_X1 U16270 ( .A(n14419), .B(n14418), .ZN(n14420) );
  XNOR2_X1 U16271 ( .A(n14420), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14498) );
  XOR2_X1 U16272 ( .A(n14422), .B(n14421), .Z(n14457) );
  INV_X1 U16273 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14780) );
  NOR2_X1 U16274 ( .A1(n14437), .A2(n14780), .ZN(n14438) );
  INV_X1 U16275 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14428) );
  NOR2_X1 U16276 ( .A1(n14427), .A2(n14428), .ZN(n14429) );
  OAI21_X1 U16277 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14426), .A(n14425), .ZN(
        n15615) );
  NAND2_X1 U16278 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15615), .ZN(n15631) );
  XOR2_X1 U16279 ( .A(n14431), .B(n14430), .Z(n14432) );
  NOR2_X1 U16280 ( .A1(n14433), .A2(n14432), .ZN(n14434) );
  XNOR2_X1 U16281 ( .A(n14433), .B(n14432), .ZN(n14487) );
  INV_X1 U16282 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14486) );
  XOR2_X1 U16283 ( .A(n14435), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15626) );
  NAND2_X1 U16284 ( .A1(n15627), .A2(n15626), .ZN(n14436) );
  NOR2_X1 U16285 ( .A1(n15627), .A2(n15626), .ZN(n15625) );
  XNOR2_X1 U16286 ( .A(n14780), .B(n14437), .ZN(n15617) );
  NOR2_X1 U16287 ( .A1(n15618), .A2(n15617), .ZN(n15616) );
  NAND2_X1 U16288 ( .A1(n14440), .A2(n14441), .ZN(n14442) );
  INV_X1 U16289 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15620) );
  INV_X1 U16290 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14793) );
  NOR2_X1 U16291 ( .A1(n14443), .A2(n14793), .ZN(n14446) );
  XNOR2_X1 U16292 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14445) );
  XNOR2_X1 U16293 ( .A(n14445), .B(n14444), .ZN(n14489) );
  INV_X1 U16294 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14448) );
  NOR2_X1 U16295 ( .A1(n6649), .A2(n14448), .ZN(n14451) );
  XNOR2_X1 U16296 ( .A(n14450), .B(n14449), .ZN(n15623) );
  XNOR2_X1 U16297 ( .A(n14453), .B(n14452), .ZN(n14455) );
  NAND2_X1 U16298 ( .A1(n14454), .A2(n14455), .ZN(n14456) );
  INV_X1 U16299 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14808) );
  NOR2_X1 U16300 ( .A1(n14457), .A2(n14458), .ZN(n14459) );
  INV_X1 U16301 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14495) );
  XNOR2_X1 U16302 ( .A(n14458), .B(n14457), .ZN(n14494) );
  NAND2_X1 U16303 ( .A1(n14498), .A2(n14497), .ZN(n14460) );
  XNOR2_X1 U16304 ( .A(n14462), .B(n14461), .ZN(n14629) );
  NAND2_X1 U16305 ( .A1(n14630), .A2(n14629), .ZN(n14463) );
  NOR2_X1 U16306 ( .A1(n14630), .A2(n14629), .ZN(n14628) );
  NAND2_X1 U16307 ( .A1(n14464), .A2(n14465), .ZN(n14466) );
  INV_X1 U16308 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15507) );
  XOR2_X1 U16309 ( .A(n14469), .B(n14468), .Z(n14470) );
  INV_X1 U16310 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14642) );
  AOI21_X1 U16311 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14473), .A(n14472), 
        .ZN(n14474) );
  XOR2_X1 U16312 ( .A(n14475), .B(n14474), .Z(n14648) );
  XNOR2_X1 U16313 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n14481) );
  NOR2_X1 U16314 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14476), .ZN(n14480) );
  INV_X1 U16315 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14478) );
  NOR2_X1 U16316 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  NOR2_X1 U16317 ( .A1(n14480), .A2(n14479), .ZN(n14520) );
  XNOR2_X1 U16318 ( .A(n14481), .B(n14520), .ZN(n14522) );
  NAND2_X1 U16319 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  OAI21_X1 U16320 ( .B1(n14523), .B2(n14522), .A(n14524), .ZN(n14482) );
  XNOR2_X1 U16321 ( .A(n14482), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16322 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14483) );
  OAI21_X1 U16323 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14483), 
        .ZN(U28) );
  AOI21_X1 U16324 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14484) );
  OAI21_X1 U16325 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14484), 
        .ZN(U29) );
  AOI21_X1 U16326 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(SUB_1596_U61) );
  AOI21_X1 U16327 ( .B1(n14490), .B2(n14489), .A(n6650), .ZN(SUB_1596_U57) );
  OAI21_X1 U16328 ( .B1(n14492), .B2(n14808), .A(n14491), .ZN(SUB_1596_U55) );
  AOI21_X1 U16329 ( .B1(n14495), .B2(n14494), .A(n14493), .ZN(SUB_1596_U54) );
  AOI21_X1 U16330 ( .B1(n14498), .B2(n14497), .A(n14496), .ZN(n14499) );
  XOR2_X1 U16331 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14499), .Z(SUB_1596_U70)
         );
  OAI211_X1 U16332 ( .C1(n14619), .C2(n14675), .A(n14617), .B(n14686), .ZN(
        n14500) );
  OAI21_X1 U16333 ( .B1(n14686), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14500), 
        .ZN(n14513) );
  OAI21_X1 U16334 ( .B1(n14503), .B2(n14502), .A(n14501), .ZN(n14623) );
  OAI211_X1 U16335 ( .C1(n14505), .C2(n14619), .A(n14601), .B(n14504), .ZN(
        n14618) );
  INV_X1 U16336 ( .A(n14618), .ZN(n14511) );
  OAI21_X1 U16337 ( .B1(n14508), .B2(n14507), .A(n14506), .ZN(n14620) );
  INV_X1 U16338 ( .A(n14620), .ZN(n14509) );
  AOI222_X1 U16339 ( .A1(n14623), .A2(n14605), .B1(n14606), .B2(n14511), .C1(
        n14510), .C2(n14509), .ZN(n14512) );
  OAI211_X1 U16340 ( .C1(n14514), .C2(n14683), .A(n14513), .B(n14512), .ZN(
        P1_U3280) );
  OAI21_X1 U16341 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14518) );
  XNOR2_X1 U16342 ( .A(n14518), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U16343 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14521) );
  AND2_X1 U16344 ( .A1(n14521), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n14519) );
  OAI22_X1 U16345 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14521), .B1(n14520), 
        .B2(n14519), .ZN(n14526) );
  AOI211_X1 U16346 ( .C1(n14529), .C2(n14537), .A(n14528), .B(n14527), .ZN(
        n14540) );
  INV_X1 U16347 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U16348 ( .A1(n15227), .A2(n14540), .B1(n15431), .B2(n15231), .ZN(
        P3_U3472) );
  NOR2_X1 U16349 ( .A1(n14530), .A2(n15211), .ZN(n14532) );
  AOI211_X1 U16350 ( .C1(n15155), .C2(n14533), .A(n14532), .B(n14531), .ZN(
        n14542) );
  AOI22_X1 U16351 ( .A1(n15227), .A2(n14542), .B1(n10445), .B2(n15231), .ZN(
        P3_U3471) );
  AOI211_X1 U16352 ( .C1(n14537), .C2(n14536), .A(n14535), .B(n14534), .ZN(
        n14544) );
  INV_X1 U16353 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14538) );
  AOI22_X1 U16354 ( .A1(n15227), .A2(n14544), .B1(n14538), .B2(n15231), .ZN(
        P3_U3470) );
  INV_X1 U16355 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U16356 ( .A1(n15217), .A2(n14540), .B1(n14539), .B2(n15215), .ZN(
        P3_U3429) );
  INV_X1 U16357 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14541) );
  AOI22_X1 U16358 ( .A1(n15217), .A2(n14542), .B1(n14541), .B2(n15215), .ZN(
        P3_U3426) );
  INV_X1 U16359 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14543) );
  AOI22_X1 U16360 ( .A1(n15217), .A2(n14544), .B1(n14543), .B2(n15215), .ZN(
        P3_U3423) );
  INV_X1 U16361 ( .A(n14545), .ZN(n14546) );
  AOI21_X1 U16362 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14551) );
  OAI222_X1 U16363 ( .A1(n14554), .A2(n14553), .B1(n14552), .B2(n14551), .C1(
        n14550), .C2(n14549), .ZN(n14555) );
  INV_X1 U16364 ( .A(n14555), .ZN(n14556) );
  NAND2_X1 U16365 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14834)
         );
  OAI211_X1 U16366 ( .C1(n14558), .C2(n14557), .A(n14556), .B(n14834), .ZN(
        P2_U3187) );
  AND2_X1 U16367 ( .A1(n14560), .A2(n14559), .ZN(n14563) );
  OAI21_X1 U16368 ( .B1(n14563), .B2(n14562), .A(n14561), .ZN(n14568) );
  INV_X1 U16369 ( .A(n14602), .ZN(n14611) );
  AOI22_X1 U16370 ( .A1(n14579), .A2(n14590), .B1(n14577), .B2(n14564), .ZN(
        n14565) );
  OAI21_X1 U16371 ( .B1(n14611), .B2(n14581), .A(n14565), .ZN(n14566) );
  AOI21_X1 U16372 ( .B1(n14568), .B2(n14567), .A(n14566), .ZN(n14570) );
  OAI211_X1 U16373 ( .C1(n14588), .C2(n14595), .A(n14570), .B(n14569), .ZN(
        P1_U3215) );
  OAI21_X1 U16374 ( .B1(n10861), .B2(n14573), .A(n14572), .ZN(n14575) );
  AOI21_X1 U16375 ( .B1(n7446), .B2(n14575), .A(n14574), .ZN(n14584) );
  AOI22_X1 U16376 ( .A1(n14579), .A2(n14578), .B1(n14577), .B2(n14576), .ZN(
        n14580) );
  OAI21_X1 U16377 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n14583) );
  NOR2_X1 U16378 ( .A1(n14584), .A2(n14583), .ZN(n14586) );
  OAI211_X1 U16379 ( .C1(n14588), .C2(n14587), .A(n14586), .B(n14585), .ZN(
        P1_U3236) );
  XNOR2_X1 U16380 ( .A(n14589), .B(n14603), .ZN(n14593) );
  AOI22_X1 U16381 ( .A1(n14593), .A2(n14592), .B1(n14591), .B2(n14590), .ZN(
        n14615) );
  OAI21_X1 U16382 ( .B1(n14611), .B2(n14675), .A(n14615), .ZN(n14599) );
  NOR2_X1 U16383 ( .A1(n14594), .A2(n14610), .ZN(n14598) );
  OAI22_X1 U16384 ( .A1(n14686), .A2(n14596), .B1(n14595), .B2(n14683), .ZN(
        n14597) );
  AOI211_X1 U16385 ( .C1(n14599), .C2(n14686), .A(n14598), .B(n14597), .ZN(
        n14608) );
  AOI211_X1 U16386 ( .C1(n14602), .C2(n14601), .A(n14719), .B(n6806), .ZN(
        n14612) );
  XNOR2_X1 U16387 ( .A(n14604), .B(n14603), .ZN(n14614) );
  AOI22_X1 U16388 ( .A1(n14612), .A2(n14606), .B1(n14614), .B2(n14605), .ZN(
        n14607) );
  NAND2_X1 U16389 ( .A1(n14608), .A2(n14607), .ZN(P1_U3279) );
  OAI22_X1 U16390 ( .A1(n14611), .A2(n14717), .B1(n14610), .B2(n14609), .ZN(
        n14613) );
  AOI211_X1 U16391 ( .C1(n14725), .C2(n14614), .A(n14613), .B(n14612), .ZN(
        n14616) );
  AND2_X1 U16392 ( .A1(n14616), .A2(n14615), .ZN(n14625) );
  AOI22_X1 U16393 ( .A1(n14741), .A2(n14625), .B1(n10792), .B2(n14739), .ZN(
        P1_U3542) );
  OAI211_X1 U16394 ( .C1(n14619), .C2(n14717), .A(n14618), .B(n14617), .ZN(
        n14622) );
  NOR2_X1 U16395 ( .A1(n14620), .A2(n14704), .ZN(n14621) );
  AOI211_X1 U16396 ( .C1(n14725), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        n14627) );
  AOI22_X1 U16397 ( .A1(n14741), .A2(n14627), .B1(n10418), .B2(n14739), .ZN(
        P1_U3541) );
  INV_X1 U16398 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U16399 ( .A1(n14733), .A2(n14625), .B1(n14624), .B2(n14731), .ZN(
        P1_U3501) );
  INV_X1 U16400 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U16401 ( .A1(n14733), .A2(n14627), .B1(n14626), .B2(n14731), .ZN(
        P1_U3498) );
  AOI21_X1 U16402 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(n14631) );
  XOR2_X1 U16403 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14631), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16404 ( .B1(n14633), .B2(n15507), .A(n14632), .ZN(SUB_1596_U68) );
  OAI21_X1 U16405 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14637) );
  XNOR2_X1 U16406 ( .A(n14637), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI222_X1 U16407 ( .A1(n14642), .A2(n14641), .B1(n14642), .B2(n14640), .C1(
        n14639), .C2(n14638), .ZN(SUB_1596_U66) );
  OAI21_X1 U16408 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n14646) );
  XNOR2_X1 U16409 ( .A(n14646), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  OAI21_X1 U16410 ( .B1(n14649), .B2(n14648), .A(n14647), .ZN(n14650) );
  XNOR2_X1 U16411 ( .A(n14650), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AOI21_X1 U16412 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n14655) );
  XNOR2_X1 U16413 ( .A(n14655), .B(n14654), .ZN(n14659) );
  AOI22_X1 U16414 ( .A1(n14656), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14657) );
  OAI21_X1 U16415 ( .B1(n14659), .B2(n14658), .A(n14657), .ZN(P1_U3243) );
  AOI21_X1 U16416 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14661), .A(n14660), 
        .ZN(n14662) );
  INV_X1 U16417 ( .A(n14662), .ZN(n14670) );
  OAI21_X1 U16418 ( .B1(n14664), .B2(n10801), .A(n14663), .ZN(n14667) );
  AOI222_X1 U16419 ( .A1(n14670), .A2(n14669), .B1(n14668), .B2(n14667), .C1(
        n14666), .C2(n14665), .ZN(n14672) );
  OAI211_X1 U16420 ( .C1(n14674), .C2(n14673), .A(n14672), .B(n14671), .ZN(
        P1_U3258) );
  OAI21_X1 U16421 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(n14679) );
  NAND2_X1 U16422 ( .A1(n14679), .A2(n14678), .ZN(n14680) );
  OAI211_X1 U16423 ( .C1(n14683), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        n14684) );
  INV_X1 U16424 ( .A(n14684), .ZN(n14688) );
  AND2_X1 U16425 ( .A1(n14686), .A2(n14685), .ZN(n14687) );
  AOI22_X1 U16426 ( .A1(n8203), .A2(n14689), .B1(n14688), .B2(n14687), .ZN(
        P1_U3293) );
  AND2_X1 U16427 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14691), .ZN(P1_U3294) );
  INV_X1 U16428 ( .A(n14691), .ZN(n14690) );
  INV_X1 U16429 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16430 ( .A1(n14690), .A2(n15335), .ZN(P1_U3295) );
  AND2_X1 U16431 ( .A1(n14691), .A2(P1_D_REG_29__SCAN_IN), .ZN(P1_U3296) );
  INV_X1 U16432 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15434) );
  NOR2_X1 U16433 ( .A1(n14690), .A2(n15434), .ZN(P1_U3297) );
  AND2_X1 U16434 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14691), .ZN(P1_U3298) );
  AND2_X1 U16435 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14691), .ZN(P1_U3299) );
  INV_X1 U16436 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15371) );
  NOR2_X1 U16437 ( .A1(n14690), .A2(n15371), .ZN(P1_U3300) );
  AND2_X1 U16438 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14691), .ZN(P1_U3301) );
  AND2_X1 U16439 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14691), .ZN(P1_U3302) );
  AND2_X1 U16440 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14691), .ZN(P1_U3303) );
  AND2_X1 U16441 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14691), .ZN(P1_U3304) );
  AND2_X1 U16442 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14691), .ZN(P1_U3305) );
  AND2_X1 U16443 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14691), .ZN(P1_U3306) );
  AND2_X1 U16444 ( .A1(n14691), .A2(P1_D_REG_18__SCAN_IN), .ZN(P1_U3307) );
  AND2_X1 U16445 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14691), .ZN(P1_U3308) );
  AND2_X1 U16446 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14691), .ZN(P1_U3309) );
  AND2_X1 U16447 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14691), .ZN(P1_U3310) );
  AND2_X1 U16448 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14691), .ZN(P1_U3311) );
  AND2_X1 U16449 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14691), .ZN(P1_U3312) );
  INV_X1 U16450 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15372) );
  NOR2_X1 U16451 ( .A1(n14690), .A2(n15372), .ZN(P1_U3313) );
  AND2_X1 U16452 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14691), .ZN(P1_U3314) );
  INV_X1 U16453 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15465) );
  NOR2_X1 U16454 ( .A1(n14690), .A2(n15465), .ZN(P1_U3315) );
  INV_X1 U16455 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15523) );
  NOR2_X1 U16456 ( .A1(n14690), .A2(n15523), .ZN(P1_U3316) );
  AND2_X1 U16457 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14691), .ZN(P1_U3317) );
  AND2_X1 U16458 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14691), .ZN(P1_U3318) );
  AND2_X1 U16459 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14691), .ZN(P1_U3319) );
  AND2_X1 U16460 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14691), .ZN(P1_U3320) );
  AND2_X1 U16461 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14691), .ZN(P1_U3321) );
  INV_X1 U16462 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15325) );
  NOR2_X1 U16463 ( .A1(n14690), .A2(n15325), .ZN(P1_U3322) );
  AND2_X1 U16464 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14691), .ZN(P1_U3323) );
  INV_X1 U16465 ( .A(n14692), .ZN(n14693) );
  OAI21_X1 U16466 ( .B1(n14694), .B2(n14717), .A(n14693), .ZN(n14697) );
  INV_X1 U16467 ( .A(n14695), .ZN(n14696) );
  AOI211_X1 U16468 ( .C1(n14725), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        n14734) );
  INV_X1 U16469 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14699) );
  AOI22_X1 U16470 ( .A1(n14733), .A2(n14734), .B1(n14699), .B2(n14731), .ZN(
        P1_U3462) );
  NOR2_X1 U16471 ( .A1(n14701), .A2(n14700), .ZN(n14703) );
  OAI211_X1 U16472 ( .C1(n14705), .C2(n14704), .A(n14703), .B(n14702), .ZN(
        n14706) );
  AOI21_X1 U16473 ( .B1(n14725), .B2(n14707), .A(n14706), .ZN(n14735) );
  INV_X1 U16474 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14708) );
  AOI22_X1 U16475 ( .A1(n14733), .A2(n14735), .B1(n14708), .B2(n14731), .ZN(
        P1_U3474) );
  INV_X1 U16476 ( .A(n14709), .ZN(n14711) );
  AOI211_X1 U16477 ( .C1(n14712), .C2(n14729), .A(n14711), .B(n14710), .ZN(
        n14736) );
  AOI22_X1 U16478 ( .A1(n14733), .A2(n14736), .B1(n9198), .B2(n14731), .ZN(
        P1_U3477) );
  AOI211_X1 U16479 ( .C1(n14715), .C2(n14729), .A(n14714), .B(n14713), .ZN(
        n14737) );
  AOI22_X1 U16480 ( .A1(n14733), .A2(n14737), .B1(n9322), .B2(n14731), .ZN(
        P1_U3480) );
  INV_X1 U16481 ( .A(n14716), .ZN(n14720) );
  OAI22_X1 U16482 ( .A1(n14720), .A2(n14719), .B1(n14718), .B2(n14717), .ZN(
        n14723) );
  INV_X1 U16483 ( .A(n14721), .ZN(n14722) );
  AOI211_X1 U16484 ( .C1(n14725), .C2(n14724), .A(n14723), .B(n14722), .ZN(
        n14738) );
  INV_X1 U16485 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14726) );
  AOI22_X1 U16486 ( .A1(n14733), .A2(n14738), .B1(n14726), .B2(n14731), .ZN(
        P1_U3483) );
  AOI211_X1 U16487 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14740) );
  INV_X1 U16488 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16489 ( .A1(n14733), .A2(n14740), .B1(n14732), .B2(n14731), .ZN(
        P1_U3486) );
  AOI22_X1 U16490 ( .A1(n14741), .A2(n14734), .B1(n8174), .B2(n14739), .ZN(
        P1_U3529) );
  AOI22_X1 U16491 ( .A1(n14741), .A2(n14735), .B1(n8938), .B2(n14739), .ZN(
        P1_U3533) );
  AOI22_X1 U16492 ( .A1(n14741), .A2(n14736), .B1(n8058), .B2(n14739), .ZN(
        P1_U3534) );
  AOI22_X1 U16493 ( .A1(n14741), .A2(n14737), .B1(n8059), .B2(n14739), .ZN(
        P1_U3535) );
  AOI22_X1 U16494 ( .A1(n14741), .A2(n14738), .B1(n9526), .B2(n14739), .ZN(
        P1_U3536) );
  AOI22_X1 U16495 ( .A1(n14741), .A2(n14740), .B1(n9801), .B2(n14739), .ZN(
        P1_U3537) );
  NOR2_X1 U16496 ( .A1(n14840), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16497 ( .A1(n14840), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14754) );
  INV_X1 U16498 ( .A(n14742), .ZN(n14745) );
  INV_X1 U16499 ( .A(n14743), .ZN(n14744) );
  AOI211_X1 U16500 ( .C1(n14746), .C2(n14745), .A(n14744), .B(n14847), .ZN(
        n14747) );
  AOI21_X1 U16501 ( .B1(n14854), .B2(n14748), .A(n14747), .ZN(n14753) );
  OAI211_X1 U16502 ( .C1(n14751), .C2(n14750), .A(n14856), .B(n14749), .ZN(
        n14752) );
  NAND3_X1 U16503 ( .A1(n14754), .A2(n14753), .A3(n14752), .ZN(P2_U3215) );
  AOI22_X1 U16504 ( .A1(n14840), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14766) );
  NOR2_X1 U16505 ( .A1(n14756), .A2(n14755), .ZN(n14757) );
  NOR3_X1 U16506 ( .A1(n14847), .A2(n14758), .A3(n14757), .ZN(n14759) );
  AOI21_X1 U16507 ( .B1(n14854), .B2(n14760), .A(n14759), .ZN(n14765) );
  XOR2_X1 U16508 ( .A(n14762), .B(n14761), .Z(n14763) );
  NAND2_X1 U16509 ( .A1(n14856), .A2(n14763), .ZN(n14764) );
  NAND3_X1 U16510 ( .A1(n14766), .A2(n14765), .A3(n14764), .ZN(P2_U3216) );
  INV_X1 U16511 ( .A(n14767), .ZN(n14772) );
  AOI211_X1 U16512 ( .C1(n14770), .C2(n14769), .A(n14768), .B(n14847), .ZN(
        n14771) );
  AOI211_X1 U16513 ( .C1(n14854), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14779) );
  AOI211_X1 U16514 ( .C1(n14776), .C2(n14775), .A(n14774), .B(n14802), .ZN(
        n14777) );
  INV_X1 U16515 ( .A(n14777), .ZN(n14778) );
  OAI211_X1 U16516 ( .C1(n14861), .C2(n14780), .A(n14779), .B(n14778), .ZN(
        P2_U3218) );
  INV_X1 U16517 ( .A(n14781), .ZN(n14786) );
  AOI211_X1 U16518 ( .C1(n14784), .C2(n14783), .A(n14847), .B(n14782), .ZN(
        n14785) );
  AOI211_X1 U16519 ( .C1(n14854), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14792) );
  OAI211_X1 U16520 ( .C1(n14790), .C2(n14789), .A(n14788), .B(n14856), .ZN(
        n14791) );
  OAI211_X1 U16521 ( .C1(n14861), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        P2_U3220) );
  INV_X1 U16522 ( .A(n14794), .ZN(n14799) );
  AOI211_X1 U16523 ( .C1(n14797), .C2(n14796), .A(n14847), .B(n14795), .ZN(
        n14798) );
  AOI211_X1 U16524 ( .C1(n14854), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14807) );
  AOI211_X1 U16525 ( .C1(n14804), .C2(n14803), .A(n14802), .B(n14801), .ZN(
        n14805) );
  INV_X1 U16526 ( .A(n14805), .ZN(n14806) );
  OAI211_X1 U16527 ( .C1(n14861), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        P2_U3222) );
  INV_X1 U16528 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15311) );
  NOR2_X1 U16529 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14809), .ZN(n14814) );
  AOI211_X1 U16530 ( .C1(n14812), .C2(n14811), .A(n14847), .B(n14810), .ZN(
        n14813) );
  AOI211_X1 U16531 ( .C1(n14854), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14821) );
  OAI21_X1 U16532 ( .B1(n14818), .B2(n14817), .A(n14816), .ZN(n14819) );
  NAND2_X1 U16533 ( .A1(n14819), .A2(n14856), .ZN(n14820) );
  OAI211_X1 U16534 ( .C1(n14861), .C2(n15311), .A(n14821), .B(n14820), .ZN(
        P2_U3225) );
  NOR2_X1 U16535 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14822), .ZN(n14827) );
  AOI211_X1 U16536 ( .C1(n14825), .C2(n14824), .A(n14847), .B(n14823), .ZN(
        n14826) );
  AOI211_X1 U16537 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n14840), .A(n14827), 
        .B(n14826), .ZN(n14832) );
  OAI211_X1 U16538 ( .C1(n14830), .C2(n14829), .A(n14828), .B(n14856), .ZN(
        n14831) );
  OAI211_X1 U16539 ( .C1(n14846), .C2(n14833), .A(n14832), .B(n14831), .ZN(
        P2_U3227) );
  INV_X1 U16540 ( .A(n14834), .ZN(n14839) );
  AOI211_X1 U16541 ( .C1(n14837), .C2(n14836), .A(n14835), .B(n14847), .ZN(
        n14838) );
  AOI211_X1 U16542 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n14840), .A(n14839), 
        .B(n14838), .ZN(n14844) );
  OAI211_X1 U16543 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n14842), .A(n14856), 
        .B(n14841), .ZN(n14843) );
  OAI211_X1 U16544 ( .C1(n14846), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        P2_U3228) );
  NOR2_X1 U16545 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11158), .ZN(n14852) );
  AOI211_X1 U16546 ( .C1(n14850), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n14851) );
  AOI211_X1 U16547 ( .C1(n14854), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        n14860) );
  OAI211_X1 U16548 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        n14859) );
  OAI211_X1 U16549 ( .C1(n14861), .C2(n6909), .A(n14860), .B(n14859), .ZN(
        P2_U3231) );
  NAND2_X1 U16550 ( .A1(n14863), .A2(n14862), .ZN(n14867) );
  AOI22_X1 U16551 ( .A1(n13512), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14865), 
        .B2(n14864), .ZN(n14866) );
  OAI211_X1 U16552 ( .C1(n14869), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14870) );
  AOI21_X1 U16553 ( .B1(n14872), .B2(n14871), .A(n14870), .ZN(n14873) );
  OAI21_X1 U16554 ( .B1(n13512), .B2(n14874), .A(n14873), .ZN(P2_U3258) );
  INV_X1 U16555 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n14876) );
  NOR2_X1 U16556 ( .A1(n14904), .A2(n14876), .ZN(P2_U3266) );
  INV_X1 U16557 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U16558 ( .A1(n14904), .A2(n14877), .ZN(P2_U3267) );
  INV_X1 U16559 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14878) );
  NOR2_X1 U16560 ( .A1(n14887), .A2(n14878), .ZN(P2_U3268) );
  INV_X1 U16561 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U16562 ( .A1(n14887), .A2(n14879), .ZN(P2_U3269) );
  INV_X1 U16563 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14880) );
  NOR2_X1 U16564 ( .A1(n14887), .A2(n14880), .ZN(P2_U3270) );
  INV_X1 U16565 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14881) );
  NOR2_X1 U16566 ( .A1(n14887), .A2(n14881), .ZN(P2_U3271) );
  NOR2_X1 U16567 ( .A1(n14887), .A2(n15320), .ZN(P2_U3272) );
  INV_X1 U16568 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14882) );
  NOR2_X1 U16569 ( .A1(n14887), .A2(n14882), .ZN(P2_U3273) );
  INV_X1 U16570 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14883) );
  NOR2_X1 U16571 ( .A1(n14887), .A2(n14883), .ZN(P2_U3274) );
  INV_X1 U16572 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14884) );
  NOR2_X1 U16573 ( .A1(n14887), .A2(n14884), .ZN(P2_U3275) );
  INV_X1 U16574 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14885) );
  NOR2_X1 U16575 ( .A1(n14887), .A2(n14885), .ZN(P2_U3276) );
  INV_X1 U16576 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14886) );
  NOR2_X1 U16577 ( .A1(n14887), .A2(n14886), .ZN(P2_U3277) );
  INV_X1 U16578 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14888) );
  NOR2_X1 U16579 ( .A1(n14904), .A2(n14888), .ZN(P2_U3278) );
  INV_X1 U16580 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15493) );
  NOR2_X1 U16581 ( .A1(n14904), .A2(n15493), .ZN(P2_U3279) );
  INV_X1 U16582 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14889) );
  NOR2_X1 U16583 ( .A1(n14904), .A2(n14889), .ZN(P2_U3280) );
  INV_X1 U16584 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U16585 ( .A1(n14904), .A2(n14890), .ZN(P2_U3281) );
  INV_X1 U16586 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n14891) );
  NOR2_X1 U16587 ( .A1(n14904), .A2(n14891), .ZN(P2_U3282) );
  NOR2_X1 U16588 ( .A1(n14904), .A2(n15478), .ZN(P2_U3283) );
  INV_X1 U16589 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14892) );
  NOR2_X1 U16590 ( .A1(n14904), .A2(n14892), .ZN(P2_U3284) );
  INV_X1 U16591 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14893) );
  NOR2_X1 U16592 ( .A1(n14904), .A2(n14893), .ZN(P2_U3285) );
  NOR2_X1 U16593 ( .A1(n14904), .A2(n14894), .ZN(P2_U3286) );
  INV_X1 U16594 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14895) );
  NOR2_X1 U16595 ( .A1(n14904), .A2(n14895), .ZN(P2_U3287) );
  INV_X1 U16596 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14896) );
  NOR2_X1 U16597 ( .A1(n14904), .A2(n14896), .ZN(P2_U3288) );
  INV_X1 U16598 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14897) );
  NOR2_X1 U16599 ( .A1(n14904), .A2(n14897), .ZN(P2_U3289) );
  INV_X1 U16600 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14898) );
  NOR2_X1 U16601 ( .A1(n14904), .A2(n14898), .ZN(P2_U3290) );
  INV_X1 U16602 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14899) );
  NOR2_X1 U16603 ( .A1(n14904), .A2(n14899), .ZN(P2_U3291) );
  INV_X1 U16604 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U16605 ( .A1(n14904), .A2(n14900), .ZN(P2_U3292) );
  INV_X1 U16606 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14901) );
  NOR2_X1 U16607 ( .A1(n14904), .A2(n14901), .ZN(P2_U3293) );
  NOR2_X1 U16608 ( .A1(n14904), .A2(n15483), .ZN(P2_U3294) );
  INV_X1 U16609 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14902) );
  NOR2_X1 U16610 ( .A1(n14904), .A2(n14902), .ZN(P2_U3295) );
  OAI22_X1 U16611 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n14904), .B1(n14907), .B2(
        n14903), .ZN(n14905) );
  INV_X1 U16612 ( .A(n14905), .ZN(P2_U3416) );
  AOI21_X1 U16613 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(P2_U3417) );
  AOI211_X1 U16614 ( .C1(n14958), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        n14961) );
  AOI22_X1 U16615 ( .A1(n14960), .A2(n14961), .B1(n8334), .B2(n14959), .ZN(
        P2_U3430) );
  AOI22_X1 U16616 ( .A1(n14960), .A2(n14912), .B1(n8348), .B2(n14959), .ZN(
        P2_U3433) );
  NAND2_X1 U16617 ( .A1(n14913), .A2(n14958), .ZN(n14915) );
  OAI211_X1 U16618 ( .C1(n14916), .C2(n14953), .A(n14915), .B(n14914), .ZN(
        n14917) );
  NOR2_X1 U16619 ( .A1(n14918), .A2(n14917), .ZN(n14962) );
  AOI22_X1 U16620 ( .A1(n14960), .A2(n14962), .B1(n8361), .B2(n14959), .ZN(
        P2_U3436) );
  OAI211_X1 U16621 ( .C1(n14921), .C2(n14953), .A(n14920), .B(n14919), .ZN(
        n14922) );
  AOI21_X1 U16622 ( .B1(n14938), .B2(n14923), .A(n14922), .ZN(n14963) );
  INV_X1 U16623 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14924) );
  AOI22_X1 U16624 ( .A1(n14960), .A2(n14963), .B1(n14924), .B2(n14959), .ZN(
        P2_U3439) );
  AOI21_X1 U16625 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14929) );
  OAI211_X1 U16626 ( .C1(n14931), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14932) );
  INV_X1 U16627 ( .A(n14932), .ZN(n14965) );
  AOI22_X1 U16628 ( .A1(n14960), .A2(n14965), .B1(n8787), .B2(n14959), .ZN(
        P2_U3442) );
  INV_X1 U16629 ( .A(n14933), .ZN(n14939) );
  INV_X1 U16630 ( .A(n14934), .ZN(n14935) );
  OAI21_X1 U16631 ( .B1(n14936), .B2(n14953), .A(n14935), .ZN(n14937) );
  AOI21_X1 U16632 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(n14940) );
  AND2_X1 U16633 ( .A1(n14941), .A2(n14940), .ZN(n14966) );
  AOI22_X1 U16634 ( .A1(n14960), .A2(n14966), .B1(n8907), .B2(n14959), .ZN(
        P2_U3445) );
  INV_X1 U16635 ( .A(n14942), .ZN(n14948) );
  INV_X1 U16636 ( .A(n14943), .ZN(n14944) );
  OAI21_X1 U16637 ( .B1(n14945), .B2(n14953), .A(n14944), .ZN(n14947) );
  AOI211_X1 U16638 ( .C1(n14958), .C2(n14948), .A(n14947), .B(n14946), .ZN(
        n14967) );
  AOI22_X1 U16639 ( .A1(n14960), .A2(n14967), .B1(n9137), .B2(n14959), .ZN(
        P2_U3454) );
  NOR2_X1 U16640 ( .A1(n14950), .A2(n14949), .ZN(n14956) );
  OAI211_X1 U16641 ( .C1(n14954), .C2(n14953), .A(n14952), .B(n14951), .ZN(
        n14955) );
  AOI211_X1 U16642 ( .C1(n14958), .C2(n14957), .A(n14956), .B(n14955), .ZN(
        n14969) );
  AOI22_X1 U16643 ( .A1(n14960), .A2(n14969), .B1(n9255), .B2(n14959), .ZN(
        P2_U3457) );
  AOI22_X1 U16644 ( .A1(n14970), .A2(n14961), .B1(n8252), .B2(n14968), .ZN(
        P2_U3499) );
  AOI22_X1 U16645 ( .A1(n14970), .A2(n14962), .B1(n8389), .B2(n14968), .ZN(
        P2_U3501) );
  AOI22_X1 U16646 ( .A1(n14970), .A2(n14963), .B1(n8728), .B2(n14968), .ZN(
        P2_U3502) );
  INV_X1 U16647 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U16648 ( .A1(n14970), .A2(n14965), .B1(n14964), .B2(n14968), .ZN(
        P2_U3503) );
  INV_X1 U16649 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U16650 ( .A1(n14970), .A2(n14966), .B1(n15519), .B2(n14968), .ZN(
        P2_U3504) );
  AOI22_X1 U16651 ( .A1(n14970), .A2(n14967), .B1(n8880), .B2(n14968), .ZN(
        P2_U3507) );
  AOI22_X1 U16652 ( .A1(n14970), .A2(n14969), .B1(n9254), .B2(n14968), .ZN(
        P2_U3508) );
  NOR2_X1 U16653 ( .A1(P3_U3897), .A2(n15092), .ZN(P3_U3150) );
  AOI21_X1 U16654 ( .B1(n10088), .B2(n14972), .A(n14971), .ZN(n14987) );
  INV_X1 U16655 ( .A(n14994), .ZN(n14977) );
  NOR3_X1 U16656 ( .A1(n14975), .A2(n14974), .A3(n14973), .ZN(n14976) );
  OAI21_X1 U16657 ( .B1(n14977), .B2(n14976), .A(n15084), .ZN(n14978) );
  OAI21_X1 U16658 ( .B1(n15089), .B2(n14979), .A(n14978), .ZN(n14980) );
  AOI211_X1 U16659 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n15092), .A(n14981), .B(
        n14980), .ZN(n14986) );
  OAI21_X1 U16660 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14983), .A(n14982), .ZN(
        n14984) );
  NAND2_X1 U16661 ( .A1(n15095), .A2(n14984), .ZN(n14985) );
  OAI211_X1 U16662 ( .C1(n14987), .C2(n15099), .A(n14986), .B(n14985), .ZN(
        P3_U3185) );
  INV_X1 U16663 ( .A(n14988), .ZN(n14989) );
  AOI21_X1 U16664 ( .B1(n14991), .B2(n14990), .A(n14989), .ZN(n15006) );
  AND3_X1 U16665 ( .A1(n14994), .A2(n14993), .A3(n14992), .ZN(n14995) );
  OAI21_X1 U16666 ( .B1(n15012), .B2(n14995), .A(n15084), .ZN(n14996) );
  OAI21_X1 U16667 ( .B1(n15089), .B2(n14997), .A(n14996), .ZN(n14998) );
  AOI211_X1 U16668 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n15092), .A(n14999), .B(
        n14998), .ZN(n15005) );
  OAI21_X1 U16669 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15003) );
  NAND2_X1 U16670 ( .A1(n15095), .A2(n15003), .ZN(n15004) );
  OAI211_X1 U16671 ( .C1(n15006), .C2(n15099), .A(n15005), .B(n15004), .ZN(
        P3_U3186) );
  AOI21_X1 U16672 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15024) );
  INV_X1 U16673 ( .A(n15030), .ZN(n15014) );
  NOR3_X1 U16674 ( .A1(n15012), .A2(n15011), .A3(n15010), .ZN(n15013) );
  OAI21_X1 U16675 ( .B1(n15014), .B2(n15013), .A(n15084), .ZN(n15015) );
  OAI21_X1 U16676 ( .B1(n15089), .B2(n15016), .A(n15015), .ZN(n15017) );
  AOI211_X1 U16677 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15092), .A(n15018), .B(
        n15017), .ZN(n15023) );
  OAI21_X1 U16678 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15020), .A(n15019), .ZN(
        n15021) );
  NAND2_X1 U16679 ( .A1(n15095), .A2(n15021), .ZN(n15022) );
  OAI211_X1 U16680 ( .C1(n15024), .C2(n15099), .A(n15023), .B(n15022), .ZN(
        P3_U3187) );
  AOI21_X1 U16681 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(n15042) );
  AND3_X1 U16682 ( .A1(n15030), .A2(n15029), .A3(n15028), .ZN(n15031) );
  OAI21_X1 U16683 ( .B1(n15047), .B2(n15031), .A(n15084), .ZN(n15032) );
  OAI21_X1 U16684 ( .B1(n15089), .B2(n15033), .A(n15032), .ZN(n15034) );
  AOI211_X1 U16685 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n15092), .A(n15035), .B(
        n15034), .ZN(n15041) );
  OAI21_X1 U16686 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15039) );
  NAND2_X1 U16687 ( .A1(n15039), .A2(n15095), .ZN(n15040) );
  OAI211_X1 U16688 ( .C1(n15042), .C2(n15099), .A(n15041), .B(n15040), .ZN(
        P3_U3188) );
  AOI21_X1 U16689 ( .B1(n10207), .B2(n15044), .A(n15043), .ZN(n15059) );
  INV_X1 U16690 ( .A(n15065), .ZN(n15049) );
  NOR3_X1 U16691 ( .A1(n15047), .A2(n15046), .A3(n15045), .ZN(n15048) );
  OAI21_X1 U16692 ( .B1(n15049), .B2(n15048), .A(n15084), .ZN(n15050) );
  OAI21_X1 U16693 ( .B1(n15089), .B2(n15051), .A(n15050), .ZN(n15052) );
  AOI211_X1 U16694 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15092), .A(n15053), .B(
        n15052), .ZN(n15058) );
  OAI21_X1 U16695 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15055), .A(n15054), .ZN(
        n15056) );
  NAND2_X1 U16696 ( .A1(n15056), .A2(n15095), .ZN(n15057) );
  OAI211_X1 U16697 ( .C1(n15059), .C2(n15099), .A(n15058), .B(n15057), .ZN(
        P3_U3189) );
  AOI21_X1 U16698 ( .B1(n15062), .B2(n15061), .A(n15060), .ZN(n15077) );
  AND3_X1 U16699 ( .A1(n15065), .A2(n15064), .A3(n15063), .ZN(n15066) );
  OAI21_X1 U16700 ( .B1(n15083), .B2(n15066), .A(n15084), .ZN(n15067) );
  OAI21_X1 U16701 ( .B1(n15089), .B2(n15068), .A(n15067), .ZN(n15069) );
  AOI211_X1 U16702 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n15092), .A(n15070), .B(
        n15069), .ZN(n15076) );
  OAI21_X1 U16703 ( .B1(n15073), .B2(n15072), .A(n15071), .ZN(n15074) );
  NAND2_X1 U16704 ( .A1(n15074), .A2(n15095), .ZN(n15075) );
  OAI211_X1 U16705 ( .C1(n15077), .C2(n15099), .A(n15076), .B(n15075), .ZN(
        P3_U3190) );
  AOI21_X1 U16706 ( .B1(n10486), .B2(n15079), .A(n15078), .ZN(n15100) );
  INV_X1 U16707 ( .A(n15080), .ZN(n15086) );
  NOR3_X1 U16708 ( .A1(n15083), .A2(n15082), .A3(n15081), .ZN(n15085) );
  OAI21_X1 U16709 ( .B1(n15086), .B2(n15085), .A(n15084), .ZN(n15087) );
  OAI21_X1 U16710 ( .B1(n15089), .B2(n15088), .A(n15087), .ZN(n15090) );
  AOI211_X1 U16711 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15092), .A(n15091), .B(
        n15090), .ZN(n15098) );
  OAI21_X1 U16712 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15094), .A(n15093), .ZN(
        n15096) );
  NAND2_X1 U16713 ( .A1(n15096), .A2(n15095), .ZN(n15097) );
  OAI211_X1 U16714 ( .C1(n15100), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        P3_U3191) );
  XNOR2_X1 U16715 ( .A(n15102), .B(n10201), .ZN(n15108) );
  INV_X1 U16716 ( .A(n15108), .ZN(n15192) );
  OAI211_X1 U16717 ( .C1(n10202), .C2(n10201), .A(n15133), .B(n15103), .ZN(
        n15107) );
  AOI22_X1 U16718 ( .A1(n15149), .A2(n15105), .B1(n15104), .B2(n15148), .ZN(
        n15106) );
  OAI211_X1 U16719 ( .C1(n15146), .C2(n15108), .A(n15107), .B(n15106), .ZN(
        n15190) );
  AOI21_X1 U16720 ( .B1(n15136), .B2(n15192), .A(n15190), .ZN(n15112) );
  AND2_X1 U16721 ( .A1(n15109), .A2(n15155), .ZN(n15191) );
  AOI22_X1 U16722 ( .A1(n15122), .A2(n15191), .B1(n15157), .B2(n15110), .ZN(
        n15111) );
  OAI221_X1 U16723 ( .B1(n12846), .B2(n15112), .C1(n15162), .C2(n10104), .A(
        n15111), .ZN(P3_U3227) );
  XNOR2_X1 U16724 ( .A(n15114), .B(n9362), .ZN(n15119) );
  INV_X1 U16725 ( .A(n15119), .ZN(n15177) );
  AOI22_X1 U16726 ( .A1(n15148), .A2(n15150), .B1(n15115), .B2(n15149), .ZN(
        n15118) );
  OAI211_X1 U16727 ( .C1(n6780), .C2(n9362), .A(n15133), .B(n15116), .ZN(
        n15117) );
  OAI211_X1 U16728 ( .C1(n15119), .C2(n15146), .A(n15118), .B(n15117), .ZN(
        n15175) );
  AOI21_X1 U16729 ( .B1(n15136), .B2(n15177), .A(n15175), .ZN(n15124) );
  AND2_X1 U16730 ( .A1(n15120), .A2(n15155), .ZN(n15176) );
  AOI22_X1 U16731 ( .A1(n15122), .A2(n15176), .B1(n15157), .B2(n15121), .ZN(
        n15123) );
  OAI221_X1 U16732 ( .B1(n12846), .B2(n15124), .C1(n15162), .C2(n10088), .A(
        n15123), .ZN(P3_U3230) );
  XNOR2_X1 U16733 ( .A(n15125), .B(n15126), .ZN(n15170) );
  XNOR2_X1 U16734 ( .A(n15127), .B(n15126), .ZN(n15134) );
  OAI22_X1 U16735 ( .A1(n15131), .A2(n15130), .B1(n15129), .B2(n15128), .ZN(
        n15132) );
  AOI21_X1 U16736 ( .B1(n15134), .B2(n15133), .A(n15132), .ZN(n15135) );
  OAI21_X1 U16737 ( .B1(n15146), .B2(n15170), .A(n15135), .ZN(n15171) );
  INV_X1 U16738 ( .A(n15136), .ZN(n15160) );
  AND2_X1 U16739 ( .A1(n15137), .A2(n15155), .ZN(n15172) );
  AOI22_X1 U16740 ( .A1(n15172), .A2(n15158), .B1(P3_REG3_REG_2__SCAN_IN), 
        .B2(n15157), .ZN(n15138) );
  OAI21_X1 U16741 ( .B1(n15170), .B2(n15160), .A(n15138), .ZN(n15139) );
  NOR2_X1 U16742 ( .A1(n15171), .A2(n15139), .ZN(n15140) );
  AOI22_X1 U16743 ( .A1(n12846), .A2(n15141), .B1(n15140), .B2(n15162), .ZN(
        P3_U3231) );
  INV_X1 U16744 ( .A(n15142), .ZN(n15143) );
  XNOR2_X1 U16745 ( .A(n15145), .B(n15143), .ZN(n15153) );
  XNOR2_X1 U16746 ( .A(n15145), .B(n15144), .ZN(n15165) );
  OR2_X1 U16747 ( .A1(n15165), .A2(n15146), .ZN(n15152) );
  AOI22_X1 U16748 ( .A1(n15150), .A2(n15149), .B1(n15148), .B2(n15147), .ZN(
        n15151) );
  OAI211_X1 U16749 ( .C1(n15154), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15166) );
  AND2_X1 U16750 ( .A1(n15156), .A2(n15155), .ZN(n15167) );
  AOI22_X1 U16751 ( .A1(n15167), .A2(n15158), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15157), .ZN(n15159) );
  OAI21_X1 U16752 ( .B1(n15165), .B2(n15160), .A(n15159), .ZN(n15161) );
  NOR2_X1 U16753 ( .A1(n15166), .A2(n15161), .ZN(n15163) );
  AOI22_X1 U16754 ( .A1(n12846), .A2(n15164), .B1(n15163), .B2(n15162), .ZN(
        P3_U3232) );
  INV_X1 U16755 ( .A(n15165), .ZN(n15168) );
  AOI211_X1 U16756 ( .C1(n15206), .C2(n15168), .A(n15167), .B(n15166), .ZN(
        n15219) );
  INV_X1 U16757 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U16758 ( .A1(n15217), .A2(n15219), .B1(n15169), .B2(n15215), .ZN(
        P3_U3393) );
  INV_X1 U16759 ( .A(n15170), .ZN(n15173) );
  AOI211_X1 U16760 ( .C1(n15173), .C2(n15206), .A(n15172), .B(n15171), .ZN(
        n15220) );
  INV_X1 U16761 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U16762 ( .A1(n15217), .A2(n15220), .B1(n15174), .B2(n15215), .ZN(
        P3_U3396) );
  AOI211_X1 U16763 ( .C1(n15177), .C2(n15206), .A(n15176), .B(n15175), .ZN(
        n15221) );
  INV_X1 U16764 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U16765 ( .A1(n15217), .A2(n15221), .B1(n15178), .B2(n15215), .ZN(
        P3_U3399) );
  INV_X1 U16766 ( .A(n15179), .ZN(n15182) );
  AOI211_X1 U16767 ( .C1(n15182), .C2(n15206), .A(n15181), .B(n15180), .ZN(
        n15222) );
  INV_X1 U16768 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U16769 ( .A1(n15217), .A2(n15222), .B1(n15183), .B2(n15215), .ZN(
        P3_U3402) );
  OAI22_X1 U16770 ( .A1(n15186), .A2(n15185), .B1(n15184), .B2(n15209), .ZN(
        n15187) );
  NOR2_X1 U16771 ( .A1(n15188), .A2(n15187), .ZN(n15223) );
  INV_X1 U16772 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U16773 ( .A1(n15217), .A2(n15223), .B1(n15189), .B2(n15215), .ZN(
        P3_U3405) );
  AOI211_X1 U16774 ( .C1(n15192), .C2(n15206), .A(n15191), .B(n15190), .ZN(
        n15225) );
  INV_X1 U16775 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U16776 ( .A1(n15217), .A2(n15225), .B1(n15193), .B2(n15215), .ZN(
        P3_U3408) );
  INV_X1 U16777 ( .A(n15194), .ZN(n15197) );
  AOI211_X1 U16778 ( .C1(n15197), .C2(n15206), .A(n15196), .B(n15195), .ZN(
        n15226) );
  INV_X1 U16779 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15198) );
  AOI22_X1 U16780 ( .A1(n15217), .A2(n15226), .B1(n15198), .B2(n15215), .ZN(
        P3_U3411) );
  AOI211_X1 U16781 ( .C1(n15201), .C2(n15206), .A(n15200), .B(n15199), .ZN(
        n15229) );
  INV_X1 U16782 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15202) );
  AOI22_X1 U16783 ( .A1(n15217), .A2(n15229), .B1(n15202), .B2(n15215), .ZN(
        P3_U3414) );
  INV_X1 U16784 ( .A(n15203), .ZN(n15207) );
  AOI211_X1 U16785 ( .C1(n15207), .C2(n15206), .A(n15205), .B(n15204), .ZN(
        n15230) );
  INV_X1 U16786 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15208) );
  AOI22_X1 U16787 ( .A1(n15217), .A2(n15230), .B1(n15208), .B2(n15215), .ZN(
        P3_U3417) );
  OAI22_X1 U16788 ( .A1(n15212), .A2(n15211), .B1(n15210), .B2(n15209), .ZN(
        n15213) );
  NOR2_X1 U16789 ( .A1(n15214), .A2(n15213), .ZN(n15232) );
  INV_X1 U16790 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U16791 ( .A1(n15217), .A2(n15232), .B1(n15216), .B2(n15215), .ZN(
        P3_U3420) );
  AOI22_X1 U16792 ( .A1(n15227), .A2(n15219), .B1(n15218), .B2(n15231), .ZN(
        P3_U3460) );
  AOI22_X1 U16793 ( .A1(n15227), .A2(n15220), .B1(n10071), .B2(n15231), .ZN(
        P3_U3461) );
  AOI22_X1 U16794 ( .A1(n15227), .A2(n15221), .B1(n10087), .B2(n15231), .ZN(
        P3_U3462) );
  AOI22_X1 U16795 ( .A1(n15227), .A2(n15222), .B1(n10093), .B2(n15231), .ZN(
        P3_U3463) );
  AOI22_X1 U16796 ( .A1(n15227), .A2(n15223), .B1(n10100), .B2(n15231), .ZN(
        P3_U3464) );
  AOI22_X1 U16797 ( .A1(n15227), .A2(n15225), .B1(n15224), .B2(n15231), .ZN(
        P3_U3465) );
  AOI22_X1 U16798 ( .A1(n15227), .A2(n15226), .B1(n10110), .B2(n15231), .ZN(
        P3_U3466) );
  AOI22_X1 U16799 ( .A1(n15227), .A2(n15229), .B1(n15228), .B2(n15231), .ZN(
        P3_U3467) );
  AOI22_X1 U16800 ( .A1(n15227), .A2(n15230), .B1(n10119), .B2(n15231), .ZN(
        P3_U3468) );
  AOI22_X1 U16801 ( .A1(n15227), .A2(n15232), .B1(n15451), .B2(n15231), .ZN(
        P3_U3469) );
  NAND2_X1 U16802 ( .A1(n15233), .A2(P3_D_REG_25__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U16803 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput151), .B1(SI_5_), 
        .B2(keyinput179), .ZN(n15234) );
  OAI221_X1 U16804 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput151), .C1(SI_5_), .C2(keyinput179), .A(n15234), .ZN(n15241) );
  AOI22_X1 U16805 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput195), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput244), .ZN(n15235) );
  OAI221_X1 U16806 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput195), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput244), .A(n15235), .ZN(n15240) );
  AOI22_X1 U16807 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput236), .B1(
        P2_REG0_REG_8__SCAN_IN), .B2(keyinput136), .ZN(n15236) );
  OAI221_X1 U16808 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput236), .C1(
        P2_REG0_REG_8__SCAN_IN), .C2(keyinput136), .A(n15236), .ZN(n15239) );
  AOI22_X1 U16809 ( .A1(P1_D_REG_18__SCAN_IN), .A2(keyinput157), .B1(
        P3_REG0_REG_3__SCAN_IN), .B2(keyinput217), .ZN(n15237) );
  OAI221_X1 U16810 ( .B1(P1_D_REG_18__SCAN_IN), .B2(keyinput157), .C1(
        P3_REG0_REG_3__SCAN_IN), .C2(keyinput217), .A(n15237), .ZN(n15238) );
  NOR4_X1 U16811 ( .A1(n15241), .A2(n15240), .A3(n15239), .A4(n15238), .ZN(
        n15269) );
  AOI22_X1 U16812 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(keyinput139), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput187), .ZN(n15242) );
  OAI221_X1 U16813 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(keyinput139), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput187), .A(n15242), .ZN(n15249)
         );
  AOI22_X1 U16814 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(keyinput208), .B1(
        P2_REG2_REG_15__SCAN_IN), .B2(keyinput148), .ZN(n15243) );
  OAI221_X1 U16815 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(keyinput208), .C1(
        P2_REG2_REG_15__SCAN_IN), .C2(keyinput148), .A(n15243), .ZN(n15248) );
  AOI22_X1 U16816 ( .A1(SI_8_), .A2(keyinput210), .B1(P3_IR_REG_15__SCAN_IN), 
        .B2(keyinput201), .ZN(n15244) );
  OAI221_X1 U16817 ( .B1(SI_8_), .B2(keyinput210), .C1(P3_IR_REG_15__SCAN_IN), 
        .C2(keyinput201), .A(n15244), .ZN(n15247) );
  AOI22_X1 U16818 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(keyinput172), .B1(
        P2_REG1_REG_20__SCAN_IN), .B2(keyinput214), .ZN(n15245) );
  OAI221_X1 U16819 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(keyinput172), .C1(
        P2_REG1_REG_20__SCAN_IN), .C2(keyinput214), .A(n15245), .ZN(n15246) );
  NOR4_X1 U16820 ( .A1(n15249), .A2(n15248), .A3(n15247), .A4(n15246), .ZN(
        n15268) );
  AOI22_X1 U16821 ( .A1(P1_D_REG_28__SCAN_IN), .A2(keyinput128), .B1(
        P2_REG1_REG_5__SCAN_IN), .B2(keyinput150), .ZN(n15250) );
  OAI221_X1 U16822 ( .B1(P1_D_REG_28__SCAN_IN), .B2(keyinput128), .C1(
        P2_REG1_REG_5__SCAN_IN), .C2(keyinput150), .A(n15250), .ZN(n15257) );
  AOI22_X1 U16823 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput245), .B1(
        P3_D_REG_3__SCAN_IN), .B2(keyinput255), .ZN(n15251) );
  OAI221_X1 U16824 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput245), .C1(
        P3_D_REG_3__SCAN_IN), .C2(keyinput255), .A(n15251), .ZN(n15256) );
  AOI22_X1 U16825 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput212), .B1(
        P3_REG2_REG_15__SCAN_IN), .B2(keyinput159), .ZN(n15252) );
  OAI221_X1 U16826 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput212), .C1(
        P3_REG2_REG_15__SCAN_IN), .C2(keyinput159), .A(n15252), .ZN(n15255) );
  AOI22_X1 U16827 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput132), .B1(
        P2_D_REG_18__SCAN_IN), .B2(keyinput129), .ZN(n15253) );
  OAI221_X1 U16828 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput132), .C1(
        P2_D_REG_18__SCAN_IN), .C2(keyinput129), .A(n15253), .ZN(n15254) );
  NOR4_X1 U16829 ( .A1(n15257), .A2(n15256), .A3(n15255), .A4(n15254), .ZN(
        n15267) );
  AOI22_X1 U16830 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput181), .B1(
        P3_IR_REG_29__SCAN_IN), .B2(keyinput134), .ZN(n15258) );
  OAI221_X1 U16831 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput181), .C1(
        P3_IR_REG_29__SCAN_IN), .C2(keyinput134), .A(n15258), .ZN(n15265) );
  AOI22_X1 U16832 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput250), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput216), .ZN(n15259) );
  OAI221_X1 U16833 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput250), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput216), .A(n15259), .ZN(n15264) );
  AOI22_X1 U16834 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(keyinput135), .B1(
        P3_IR_REG_28__SCAN_IN), .B2(keyinput229), .ZN(n15260) );
  OAI221_X1 U16835 ( .B1(P1_DATAO_REG_3__SCAN_IN), .B2(keyinput135), .C1(
        P3_IR_REG_28__SCAN_IN), .C2(keyinput229), .A(n15260), .ZN(n15263) );
  AOI22_X1 U16836 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(keyinput202), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput232), .ZN(n15261) );
  OAI221_X1 U16837 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(keyinput202), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput232), .A(n15261), .ZN(n15262) );
  NOR4_X1 U16838 ( .A1(n15265), .A2(n15264), .A3(n15263), .A4(n15262), .ZN(
        n15266) );
  NAND4_X1 U16839 ( .A1(n15269), .A2(n15268), .A3(n15267), .A4(n15266), .ZN(
        n15418) );
  AOI22_X1 U16840 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(keyinput184), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(keyinput176), .ZN(n15270) );
  OAI221_X1 U16841 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(keyinput184), .C1(
        P2_DATAO_REG_5__SCAN_IN), .C2(keyinput176), .A(n15270), .ZN(n15277) );
  AOI22_X1 U16842 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput243), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput246), .ZN(n15271) );
  OAI221_X1 U16843 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput243), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput246), .A(n15271), .ZN(n15276) );
  AOI22_X1 U16844 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(keyinput189), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput156), .ZN(n15272) );
  OAI221_X1 U16845 ( .B1(P1_REG3_REG_15__SCAN_IN), .B2(keyinput189), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput156), .A(n15272), .ZN(n15275) );
  AOI22_X1 U16846 ( .A1(P3_D_REG_31__SCAN_IN), .A2(keyinput175), .B1(
        P3_D_REG_22__SCAN_IN), .B2(keyinput215), .ZN(n15273) );
  OAI221_X1 U16847 ( .B1(P3_D_REG_31__SCAN_IN), .B2(keyinput175), .C1(
        P3_D_REG_22__SCAN_IN), .C2(keyinput215), .A(n15273), .ZN(n15274) );
  NOR4_X1 U16848 ( .A1(n15277), .A2(n15276), .A3(n15275), .A4(n15274), .ZN(
        n15307) );
  AOI22_X1 U16849 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(keyinput213), .B1(
        P1_REG1_REG_21__SCAN_IN), .B2(keyinput130), .ZN(n15278) );
  OAI221_X1 U16850 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(keyinput213), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput130), .A(n15278), .ZN(n15285) );
  AOI22_X1 U16851 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(keyinput155), .B1(
        P1_REG1_REG_5__SCAN_IN), .B2(keyinput144), .ZN(n15279) );
  OAI221_X1 U16852 ( .B1(P1_REG1_REG_31__SCAN_IN), .B2(keyinput155), .C1(
        P1_REG1_REG_5__SCAN_IN), .C2(keyinput144), .A(n15279), .ZN(n15284) );
  AOI22_X1 U16853 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(keyinput240), .B1(
        P2_REG0_REG_2__SCAN_IN), .B2(keyinput251), .ZN(n15280) );
  OAI221_X1 U16854 ( .B1(P1_REG1_REG_29__SCAN_IN), .B2(keyinput240), .C1(
        P2_REG0_REG_2__SCAN_IN), .C2(keyinput251), .A(n15280), .ZN(n15283) );
  AOI22_X1 U16855 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(keyinput234), .B1(
        P2_REG0_REG_30__SCAN_IN), .B2(keyinput220), .ZN(n15281) );
  OAI221_X1 U16856 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(keyinput234), .C1(
        P2_REG0_REG_30__SCAN_IN), .C2(keyinput220), .A(n15281), .ZN(n15282) );
  NOR4_X1 U16857 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15306) );
  AOI22_X1 U16858 ( .A1(P1_D_REG_9__SCAN_IN), .A2(keyinput164), .B1(
        P3_REG1_REG_0__SCAN_IN), .B2(keyinput226), .ZN(n15286) );
  OAI221_X1 U16859 ( .B1(P1_D_REG_9__SCAN_IN), .B2(keyinput164), .C1(
        P3_REG1_REG_0__SCAN_IN), .C2(keyinput226), .A(n15286), .ZN(n15293) );
  AOI22_X1 U16860 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(keyinput138), .B1(
        P3_IR_REG_5__SCAN_IN), .B2(keyinput154), .ZN(n15287) );
  OAI221_X1 U16861 ( .B1(P3_DATAO_REG_20__SCAN_IN), .B2(keyinput138), .C1(
        P3_IR_REG_5__SCAN_IN), .C2(keyinput154), .A(n15287), .ZN(n15292) );
  AOI22_X1 U16862 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(keyinput168), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(keyinput171), .ZN(n15288) );
  OAI221_X1 U16863 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(keyinput168), .C1(
        P1_DATAO_REG_15__SCAN_IN), .C2(keyinput171), .A(n15288), .ZN(n15291)
         );
  AOI22_X1 U16864 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(keyinput223), .B1(
        P3_ADDR_REG_19__SCAN_IN), .B2(keyinput142), .ZN(n15289) );
  OAI221_X1 U16865 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(keyinput223), .C1(
        P3_ADDR_REG_19__SCAN_IN), .C2(keyinput142), .A(n15289), .ZN(n15290) );
  NOR4_X1 U16866 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15305) );
  AOI22_X1 U16867 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput221), .B1(
        P3_REG2_REG_29__SCAN_IN), .B2(keyinput174), .ZN(n15294) );
  OAI221_X1 U16868 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput221), .C1(
        P3_REG2_REG_29__SCAN_IN), .C2(keyinput174), .A(n15294), .ZN(n15303) );
  AOI22_X1 U16869 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput222), .B1(
        P3_REG1_REG_10__SCAN_IN), .B2(keyinput194), .ZN(n15295) );
  OAI221_X1 U16870 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput222), .C1(
        P3_REG1_REG_10__SCAN_IN), .C2(keyinput194), .A(n15295), .ZN(n15302) );
  AOI22_X1 U16871 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput196), .B1(
        P2_D_REG_11__SCAN_IN), .B2(keyinput147), .ZN(n15296) );
  OAI221_X1 U16872 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput196), .C1(
        P2_D_REG_11__SCAN_IN), .C2(keyinput147), .A(n15296), .ZN(n15301) );
  INV_X1 U16873 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U16874 ( .A1(n15299), .A2(keyinput182), .B1(n15298), .B2(
        keyinput239), .ZN(n15297) );
  OAI221_X1 U16875 ( .B1(n15299), .B2(keyinput182), .C1(n15298), .C2(
        keyinput239), .A(n15297), .ZN(n15300) );
  NOR4_X1 U16876 ( .A1(n15303), .A2(n15302), .A3(n15301), .A4(n15300), .ZN(
        n15304) );
  NAND4_X1 U16877 ( .A1(n15307), .A2(n15306), .A3(n15305), .A4(n15304), .ZN(
        n15417) );
  AOI22_X1 U16878 ( .A1(n15516), .A2(keyinput242), .B1(keyinput237), .B2(
        n15309), .ZN(n15308) );
  OAI221_X1 U16879 ( .B1(n15516), .B2(keyinput242), .C1(n15309), .C2(
        keyinput237), .A(n15308), .ZN(n15318) );
  INV_X1 U16880 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U16881 ( .A1(n15311), .A2(keyinput188), .B1(n15459), .B2(
        keyinput233), .ZN(n15310) );
  OAI221_X1 U16882 ( .B1(n15311), .B2(keyinput188), .C1(n15459), .C2(
        keyinput233), .A(n15310), .ZN(n15317) );
  XOR2_X1 U16883 ( .A(n8907), .B(keyinput141), .Z(n15315) );
  XOR2_X1 U16884 ( .A(n7705), .B(keyinput206), .Z(n15314) );
  XNOR2_X1 U16885 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput218), .ZN(n15313)
         );
  XNOR2_X1 U16886 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput170), .ZN(n15312)
         );
  NAND4_X1 U16887 ( .A1(n15315), .A2(n15314), .A3(n15313), .A4(n15312), .ZN(
        n15316) );
  NOR3_X1 U16888 ( .A1(n15318), .A2(n15317), .A3(n15316), .ZN(n15361) );
  AOI22_X1 U16889 ( .A1(n15321), .A2(keyinput228), .B1(keyinput227), .B2(
        n15320), .ZN(n15319) );
  OAI221_X1 U16890 ( .B1(n15321), .B2(keyinput228), .C1(n15320), .C2(
        keyinput227), .A(n15319), .ZN(n15331) );
  AOI22_X1 U16891 ( .A1(n15323), .A2(keyinput209), .B1(n10100), .B2(
        keyinput173), .ZN(n15322) );
  OAI221_X1 U16892 ( .B1(n15323), .B2(keyinput209), .C1(n10100), .C2(
        keyinput173), .A(n15322), .ZN(n15330) );
  AOI22_X1 U16893 ( .A1(n15326), .A2(keyinput252), .B1(n15325), .B2(
        keyinput177), .ZN(n15324) );
  OAI221_X1 U16894 ( .B1(n15326), .B2(keyinput252), .C1(n15325), .C2(
        keyinput177), .A(n15324), .ZN(n15329) );
  AOI22_X1 U16895 ( .A1(n15443), .A2(keyinput180), .B1(keyinput152), .B2(
        n15483), .ZN(n15327) );
  OAI221_X1 U16896 ( .B1(n15443), .B2(keyinput180), .C1(n15483), .C2(
        keyinput152), .A(n15327), .ZN(n15328) );
  NOR4_X1 U16897 ( .A1(n15331), .A2(n15330), .A3(n15329), .A4(n15328), .ZN(
        n15360) );
  AOI22_X1 U16898 ( .A1(n9652), .A2(keyinput199), .B1(n15333), .B2(keyinput248), .ZN(n15332) );
  OAI221_X1 U16899 ( .B1(n9652), .B2(keyinput199), .C1(n15333), .C2(
        keyinput248), .A(n15332), .ZN(n15338) );
  XNOR2_X1 U16900 ( .A(n15334), .B(keyinput137), .ZN(n15337) );
  XNOR2_X1 U16901 ( .A(n15335), .B(keyinput146), .ZN(n15336) );
  OR3_X1 U16902 ( .A1(n15338), .A2(n15337), .A3(n15336), .ZN(n15346) );
  AOI22_X1 U16903 ( .A1(n15341), .A2(keyinput241), .B1(n15340), .B2(
        keyinput225), .ZN(n15339) );
  OAI221_X1 U16904 ( .B1(n15341), .B2(keyinput241), .C1(n15340), .C2(
        keyinput225), .A(n15339), .ZN(n15345) );
  AOI22_X1 U16905 ( .A1(n14596), .A2(keyinput230), .B1(keyinput178), .B2(
        n15343), .ZN(n15342) );
  OAI221_X1 U16906 ( .B1(n14596), .B2(keyinput230), .C1(n15343), .C2(
        keyinput178), .A(n15342), .ZN(n15344) );
  NOR3_X1 U16907 ( .A1(n15346), .A2(n15345), .A3(n15344), .ZN(n15359) );
  AOI22_X1 U16908 ( .A1(n10048), .A2(keyinput238), .B1(keyinput235), .B2(
        n15491), .ZN(n15347) );
  OAI221_X1 U16909 ( .B1(n10048), .B2(keyinput238), .C1(n15491), .C2(
        keyinput235), .A(n15347), .ZN(n15357) );
  AOI22_X1 U16910 ( .A1(n15350), .A2(keyinput193), .B1(n15349), .B2(
        keyinput169), .ZN(n15348) );
  OAI221_X1 U16911 ( .B1(n15350), .B2(keyinput193), .C1(n15349), .C2(
        keyinput169), .A(n15348), .ZN(n15356) );
  XOR2_X1 U16912 ( .A(n15431), .B(keyinput254), .Z(n15354) );
  XNOR2_X1 U16913 ( .A(keyinput204), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n15353)
         );
  XNOR2_X1 U16914 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput186), .ZN(n15352) );
  XNOR2_X1 U16915 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput253), .ZN(n15351)
         );
  NAND4_X1 U16916 ( .A1(n15354), .A2(n15353), .A3(n15352), .A4(n15351), .ZN(
        n15355) );
  NOR3_X1 U16917 ( .A1(n15357), .A2(n15356), .A3(n15355), .ZN(n15358) );
  NAND4_X1 U16918 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15416) );
  XNOR2_X1 U16919 ( .A(n15362), .B(keyinput153), .ZN(n15366) );
  XNOR2_X1 U16920 ( .A(n15363), .B(keyinput200), .ZN(n15365) );
  XNOR2_X1 U16921 ( .A(keyinput145), .B(n11158), .ZN(n15364) );
  NOR3_X1 U16922 ( .A1(n15366), .A2(n15365), .A3(n15364), .ZN(n15369) );
  INV_X1 U16923 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n15446) );
  XOR2_X1 U16924 ( .A(n15446), .B(keyinput140), .Z(n15368) );
  XNOR2_X1 U16925 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput224), .ZN(n15367)
         );
  NAND3_X1 U16926 ( .A1(n15369), .A2(n15368), .A3(n15367), .ZN(n15375) );
  INV_X1 U16927 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U16928 ( .A1(n15429), .A2(keyinput158), .B1(n15371), .B2(
        keyinput165), .ZN(n15370) );
  OAI221_X1 U16929 ( .B1(n15429), .B2(keyinput158), .C1(n15371), .C2(
        keyinput165), .A(n15370), .ZN(n15374) );
  XNOR2_X1 U16930 ( .A(n15372), .B(keyinput211), .ZN(n15373) );
  NOR3_X1 U16931 ( .A1(n15375), .A2(n15374), .A3(n15373), .ZN(n15414) );
  AOI22_X1 U16932 ( .A1(n15478), .A2(keyinput160), .B1(n15377), .B2(
        keyinput167), .ZN(n15376) );
  OAI221_X1 U16933 ( .B1(n15478), .B2(keyinput160), .C1(n15377), .C2(
        keyinput167), .A(n15376), .ZN(n15386) );
  AOI22_X1 U16934 ( .A1(n15496), .A2(keyinput191), .B1(n9527), .B2(keyinput166), .ZN(n15378) );
  OAI221_X1 U16935 ( .B1(n15496), .B2(keyinput191), .C1(n9527), .C2(
        keyinput166), .A(n15378), .ZN(n15385) );
  INV_X1 U16936 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15380) );
  AOI22_X1 U16937 ( .A1(n15380), .A2(keyinput143), .B1(n14055), .B2(
        keyinput219), .ZN(n15379) );
  OAI221_X1 U16938 ( .B1(n15380), .B2(keyinput143), .C1(n14055), .C2(
        keyinput219), .A(n15379), .ZN(n15384) );
  XOR2_X1 U16939 ( .A(n15507), .B(keyinput205), .Z(n15382) );
  XNOR2_X1 U16940 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput183), .ZN(n15381) );
  NAND2_X1 U16941 ( .A1(n15382), .A2(n15381), .ZN(n15383) );
  NOR4_X1 U16942 ( .A1(n15386), .A2(n15385), .A3(n15384), .A4(n15383), .ZN(
        n15413) );
  INV_X1 U16943 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U16944 ( .A1(n15486), .A2(keyinput207), .B1(n15506), .B2(
        keyinput133), .ZN(n15387) );
  OAI221_X1 U16945 ( .B1(n15486), .B2(keyinput207), .C1(n15506), .C2(
        keyinput133), .A(n15387), .ZN(n15398) );
  INV_X1 U16946 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U16947 ( .A1(n15389), .A2(keyinput185), .B1(n15444), .B2(
        keyinput198), .ZN(n15388) );
  OAI221_X1 U16948 ( .B1(n15389), .B2(keyinput185), .C1(n15444), .C2(
        keyinput198), .A(n15388), .ZN(n15397) );
  AOI22_X1 U16949 ( .A1(n15392), .A2(keyinput231), .B1(keyinput192), .B2(
        n15391), .ZN(n15390) );
  OAI221_X1 U16950 ( .B1(n15392), .B2(keyinput231), .C1(n15391), .C2(
        keyinput192), .A(n15390), .ZN(n15396) );
  INV_X1 U16951 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15524) );
  XOR2_X1 U16952 ( .A(n15524), .B(keyinput149), .Z(n15394) );
  XNOR2_X1 U16953 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput249), .ZN(n15393)
         );
  NAND2_X1 U16954 ( .A1(n15394), .A2(n15393), .ZN(n15395) );
  NOR4_X1 U16955 ( .A1(n15398), .A2(n15397), .A3(n15396), .A4(n15395), .ZN(
        n15412) );
  AOI22_X1 U16956 ( .A1(n15504), .A2(keyinput162), .B1(n15400), .B2(
        keyinput203), .ZN(n15399) );
  OAI221_X1 U16957 ( .B1(n15504), .B2(keyinput162), .C1(n15400), .C2(
        keyinput203), .A(n15399), .ZN(n15410) );
  AOI22_X1 U16958 ( .A1(n15402), .A2(keyinput190), .B1(P3_U3151), .B2(
        keyinput161), .ZN(n15401) );
  OAI221_X1 U16959 ( .B1(n15402), .B2(keyinput190), .C1(P3_U3151), .C2(
        keyinput161), .A(n15401), .ZN(n15409) );
  XOR2_X1 U16960 ( .A(n15449), .B(keyinput247), .Z(n15405) );
  XNOR2_X1 U16961 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput163), .ZN(n15404)
         );
  XNOR2_X1 U16962 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput197), .ZN(n15403) );
  NAND3_X1 U16963 ( .A1(n15405), .A2(n15404), .A3(n15403), .ZN(n15408) );
  XNOR2_X1 U16964 ( .A(n15406), .B(keyinput131), .ZN(n15407) );
  NOR4_X1 U16965 ( .A1(n15410), .A2(n15409), .A3(n15408), .A4(n15407), .ZN(
        n15411) );
  NAND4_X1 U16966 ( .A1(n15414), .A2(n15413), .A3(n15412), .A4(n15411), .ZN(
        n15415) );
  NOR4_X1 U16967 ( .A1(n15418), .A2(n15417), .A3(n15416), .A4(n15415), .ZN(
        n15612) );
  AOI22_X1 U16968 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput84), .B1(
        P3_IR_REG_15__SCAN_IN), .B2(keyinput73), .ZN(n15419) );
  OAI221_X1 U16969 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput84), .C1(
        P3_IR_REG_15__SCAN_IN), .C2(keyinput73), .A(n15419), .ZN(n15427) );
  AOI22_X1 U16970 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput99), .B1(
        P3_IR_REG_14__SCAN_IN), .B2(keyinput69), .ZN(n15420) );
  OAI221_X1 U16971 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput99), .C1(
        P3_IR_REG_14__SCAN_IN), .C2(keyinput69), .A(n15420), .ZN(n15426) );
  AOI22_X1 U16972 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(keyinput6), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput104), .ZN(n15421) );
  OAI221_X1 U16973 ( .B1(P3_IR_REG_29__SCAN_IN), .B2(keyinput6), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput104), .A(n15421), .ZN(n15425) );
  AOI22_X1 U16974 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(keyinput46), .B1(n15423), 
        .B2(keyinput92), .ZN(n15422) );
  OAI221_X1 U16975 ( .B1(P3_REG2_REG_29__SCAN_IN), .B2(keyinput46), .C1(n15423), .C2(keyinput92), .A(n15422), .ZN(n15424) );
  NOR4_X1 U16976 ( .A1(n15427), .A2(n15426), .A3(n15425), .A4(n15424), .ZN(
        n15473) );
  AOI22_X1 U16977 ( .A1(n10596), .A2(keyinput74), .B1(n15429), .B2(keyinput30), 
        .ZN(n15428) );
  OAI221_X1 U16978 ( .B1(n10596), .B2(keyinput74), .C1(n15429), .C2(keyinput30), .A(n15428), .ZN(n15441) );
  AOI22_X1 U16979 ( .A1(n15432), .A2(keyinput23), .B1(n15431), .B2(keyinput126), .ZN(n15430) );
  OAI221_X1 U16980 ( .B1(n15432), .B2(keyinput23), .C1(n15431), .C2(
        keyinput126), .A(n15430), .ZN(n15440) );
  AOI22_X1 U16981 ( .A1(n15435), .A2(keyinput106), .B1(n15434), .B2(keyinput0), 
        .ZN(n15433) );
  OAI221_X1 U16982 ( .B1(n15435), .B2(keyinput106), .C1(n15434), .C2(keyinput0), .A(n15433), .ZN(n15439) );
  XNOR2_X1 U16983 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput116), .ZN(n15437)
         );
  XNOR2_X1 U16984 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput9), .ZN(n15436) );
  NAND2_X1 U16985 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  NOR4_X1 U16986 ( .A1(n15441), .A2(n15440), .A3(n15439), .A4(n15438), .ZN(
        n15472) );
  AOI22_X1 U16987 ( .A1(n15444), .A2(keyinput70), .B1(n15443), .B2(keyinput52), 
        .ZN(n15442) );
  OAI221_X1 U16988 ( .B1(n15444), .B2(keyinput70), .C1(n15443), .C2(keyinput52), .A(n15442), .ZN(n15457) );
  AOI22_X1 U16989 ( .A1(n15447), .A2(keyinput14), .B1(keyinput12), .B2(n15446), 
        .ZN(n15445) );
  OAI221_X1 U16990 ( .B1(n15447), .B2(keyinput14), .C1(n15446), .C2(keyinput12), .A(n15445), .ZN(n15456) );
  AOI22_X1 U16991 ( .A1(n15450), .A2(keyinput27), .B1(n15449), .B2(keyinput119), .ZN(n15448) );
  OAI221_X1 U16992 ( .B1(n15450), .B2(keyinput27), .C1(n15449), .C2(
        keyinput119), .A(n15448), .ZN(n15455) );
  XOR2_X1 U16993 ( .A(n15451), .B(keyinput66), .Z(n15453) );
  XNOR2_X1 U16994 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput122), .ZN(n15452) );
  NAND2_X1 U16995 ( .A1(n15453), .A2(n15452), .ZN(n15454) );
  NOR4_X1 U16996 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15471) );
  AOI22_X1 U16997 ( .A1(n15460), .A2(keyinput88), .B1(keyinput105), .B2(n15459), .ZN(n15458) );
  OAI221_X1 U16998 ( .B1(n15460), .B2(keyinput88), .C1(n15459), .C2(
        keyinput105), .A(n15458), .ZN(n15469) );
  AOI22_X1 U16999 ( .A1(n8938), .A2(keyinput16), .B1(n9254), .B2(keyinput11), 
        .ZN(n15461) );
  OAI221_X1 U17000 ( .B1(n8938), .B2(keyinput16), .C1(n9254), .C2(keyinput11), 
        .A(n15461), .ZN(n15468) );
  XNOR2_X1 U17001 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput48), .ZN(n15464)
         );
  XNOR2_X1 U17002 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput90), .ZN(n15463) );
  XNOR2_X1 U17003 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput72), .ZN(n15462) );
  NAND3_X1 U17004 ( .A1(n15464), .A2(n15463), .A3(n15462), .ZN(n15467) );
  XNOR2_X1 U17005 ( .A(n15465), .B(keyinput117), .ZN(n15466) );
  NOR4_X1 U17006 ( .A1(n15469), .A2(n15468), .A3(n15467), .A4(n15466), .ZN(
        n15470) );
  NAND4_X1 U17007 ( .A1(n15473), .A2(n15472), .A3(n15471), .A4(n15470), .ZN(
        n15611) );
  AOI22_X1 U17008 ( .A1(n15476), .A2(keyinput4), .B1(n15475), .B2(keyinput86), 
        .ZN(n15474) );
  OAI221_X1 U17009 ( .B1(n15476), .B2(keyinput4), .C1(n15475), .C2(keyinput86), 
        .A(n15474), .ZN(n15481) );
  XNOR2_X1 U17010 ( .A(n15477), .B(keyinput40), .ZN(n15480) );
  XNOR2_X1 U17011 ( .A(n15478), .B(keyinput32), .ZN(n15479) );
  OR3_X1 U17012 ( .A1(n15481), .A2(n15480), .A3(n15479), .ZN(n15489) );
  AOI22_X1 U17013 ( .A1(n15483), .A2(keyinput24), .B1(n10100), .B2(keyinput45), 
        .ZN(n15482) );
  OAI221_X1 U17014 ( .B1(n15483), .B2(keyinput24), .C1(n10100), .C2(keyinput45), .A(n15482), .ZN(n15488) );
  AOI22_X1 U17015 ( .A1(n15486), .A2(keyinput79), .B1(n15485), .B2(keyinput95), 
        .ZN(n15484) );
  OAI221_X1 U17016 ( .B1(n15486), .B2(keyinput79), .C1(n15485), .C2(keyinput95), .A(n15484), .ZN(n15487) );
  NOR3_X1 U17017 ( .A1(n15489), .A2(n15488), .A3(n15487), .ZN(n15534) );
  AOI22_X1 U17018 ( .A1(n9137), .A2(keyinput8), .B1(keyinput107), .B2(n15491), 
        .ZN(n15490) );
  OAI221_X1 U17019 ( .B1(n9137), .B2(keyinput8), .C1(n15491), .C2(keyinput107), 
        .A(n15490), .ZN(n15502) );
  AOI22_X1 U17020 ( .A1(n15493), .A2(keyinput1), .B1(keyinput71), .B2(n9652), 
        .ZN(n15492) );
  OAI221_X1 U17021 ( .B1(n15493), .B2(keyinput1), .C1(n9652), .C2(keyinput71), 
        .A(n15492), .ZN(n15501) );
  AOI22_X1 U17022 ( .A1(n15495), .A2(keyinput112), .B1(n8907), .B2(keyinput13), 
        .ZN(n15494) );
  OAI221_X1 U17023 ( .B1(n15495), .B2(keyinput112), .C1(n8907), .C2(keyinput13), .A(n15494), .ZN(n15500) );
  XOR2_X1 U17024 ( .A(n15496), .B(keyinput63), .Z(n15498) );
  XNOR2_X1 U17025 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput7), .ZN(n15497) );
  NAND2_X1 U17026 ( .A1(n15498), .A2(n15497), .ZN(n15499) );
  NOR4_X1 U17027 ( .A1(n15502), .A2(n15501), .A3(n15500), .A4(n15499), .ZN(
        n15533) );
  AOI22_X1 U17028 ( .A1(n9201), .A2(keyinput56), .B1(keyinput34), .B2(n15504), 
        .ZN(n15503) );
  OAI221_X1 U17029 ( .B1(n9201), .B2(keyinput56), .C1(n15504), .C2(keyinput34), 
        .A(n15503), .ZN(n15514) );
  AOI22_X1 U17030 ( .A1(n15507), .A2(keyinput77), .B1(n15506), .B2(keyinput5), 
        .ZN(n15505) );
  OAI221_X1 U17031 ( .B1(n15507), .B2(keyinput77), .C1(n15506), .C2(keyinput5), 
        .A(n15505), .ZN(n15513) );
  XOR2_X1 U17032 ( .A(n8361), .B(keyinput123), .Z(n15511) );
  XNOR2_X1 U17033 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput55), .ZN(n15510) );
  XNOR2_X1 U17034 ( .A(P3_REG2_REG_15__SCAN_IN), .B(keyinput31), .ZN(n15509)
         );
  XNOR2_X1 U17035 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput121), .ZN(n15508)
         );
  NAND4_X1 U17036 ( .A1(n15511), .A2(n15510), .A3(n15509), .A4(n15508), .ZN(
        n15512) );
  NOR3_X1 U17037 ( .A1(n15514), .A2(n15513), .A3(n15512), .ZN(n15532) );
  AOI22_X1 U17038 ( .A1(n15517), .A2(keyinput2), .B1(n15516), .B2(keyinput114), 
        .ZN(n15515) );
  OAI221_X1 U17039 ( .B1(n15517), .B2(keyinput2), .C1(n15516), .C2(keyinput114), .A(n15515), .ZN(n15522) );
  XNOR2_X1 U17040 ( .A(n15518), .B(keyinput42), .ZN(n15521) );
  XNOR2_X1 U17041 ( .A(keyinput22), .B(n15519), .ZN(n15520) );
  OR3_X1 U17042 ( .A1(n15522), .A2(n15521), .A3(n15520), .ZN(n15530) );
  XNOR2_X1 U17043 ( .A(n15523), .B(keyinput36), .ZN(n15529) );
  XNOR2_X1 U17044 ( .A(keyinput21), .B(n15524), .ZN(n15528) );
  XNOR2_X1 U17045 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput115), .ZN(n15526)
         );
  XNOR2_X1 U17046 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput96), .ZN(n15525)
         );
  NAND2_X1 U17047 ( .A1(n15526), .A2(n15525), .ZN(n15527) );
  NOR4_X1 U17048 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n15531) );
  NAND4_X1 U17049 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15610) );
  OAI22_X1 U17050 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(keyinput98), .B1(
        keyinput76), .B2(P1_REG1_REG_7__SCAN_IN), .ZN(n15535) );
  AOI221_X1 U17051 ( .B1(P3_REG1_REG_0__SCAN_IN), .B2(keyinput98), .C1(
        P1_REG1_REG_7__SCAN_IN), .C2(keyinput76), .A(n15535), .ZN(n15542) );
  OAI22_X1 U17052 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput43), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput94), .ZN(n15536) );
  AOI221_X1 U17053 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput43), .C1(
        keyinput94), .C2(P1_IR_REG_27__SCAN_IN), .A(n15536), .ZN(n15541) );
  OAI22_X1 U17054 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput33), .B1(SI_5_), 
        .B2(keyinput51), .ZN(n15537) );
  AOI221_X1 U17055 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput33), .C1(
        keyinput51), .C2(SI_5_), .A(n15537), .ZN(n15540) );
  OAI22_X1 U17056 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(keyinput26), .B1(keyinput83), .B2(P1_D_REG_12__SCAN_IN), .ZN(n15538) );
  AOI221_X1 U17057 ( .B1(P3_IR_REG_5__SCAN_IN), .B2(keyinput26), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput83), .A(n15538), .ZN(n15539) );
  NAND4_X1 U17058 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        n15570) );
  OAI22_X1 U17059 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput64), .B1(
        keyinput35), .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n15543) );
  AOI221_X1 U17060 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput64), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput35), .A(n15543), .ZN(n15550) );
  OAI22_X1 U17061 ( .A1(P3_D_REG_5__SCAN_IN), .A2(keyinput3), .B1(keyinput61), 
        .B2(P1_REG3_REG_15__SCAN_IN), .ZN(n15544) );
  AOI221_X1 U17062 ( .B1(P3_D_REG_5__SCAN_IN), .B2(keyinput3), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput61), .A(n15544), .ZN(n15549) );
  OAI22_X1 U17063 ( .A1(P3_D_REG_31__SCAN_IN), .A2(keyinput47), .B1(
        P1_D_REG_30__SCAN_IN), .B2(keyinput18), .ZN(n15545) );
  AOI221_X1 U17064 ( .B1(P3_D_REG_31__SCAN_IN), .B2(keyinput47), .C1(
        keyinput18), .C2(P1_D_REG_30__SCAN_IN), .A(n15545), .ZN(n15548) );
  OAI22_X1 U17065 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(keyinput81), .B1(
        keyinput110), .B2(P1_REG2_REG_8__SCAN_IN), .ZN(n15546) );
  AOI221_X1 U17066 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(keyinput81), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(keyinput110), .A(n15546), .ZN(n15547) );
  NAND4_X1 U17067 ( .A1(n15550), .A2(n15549), .A3(n15548), .A4(n15547), .ZN(
        n15569) );
  OAI22_X1 U17068 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput50), .B1(
        keyinput85), .B2(P2_ADDR_REG_13__SCAN_IN), .ZN(n15551) );
  AOI221_X1 U17069 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput50), .C1(
        P2_ADDR_REG_13__SCAN_IN), .C2(keyinput85), .A(n15551), .ZN(n15558) );
  OAI22_X1 U17070 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput118), .B1(
        keyinput82), .B2(SI_8_), .ZN(n15552) );
  AOI221_X1 U17071 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput118), .C1(SI_8_), .C2(keyinput82), .A(n15552), .ZN(n15557) );
  OAI22_X1 U17072 ( .A1(P3_D_REG_17__SCAN_IN), .A2(keyinput100), .B1(
        P2_REG2_REG_15__SCAN_IN), .B2(keyinput20), .ZN(n15553) );
  AOI221_X1 U17073 ( .B1(P3_D_REG_17__SCAN_IN), .B2(keyinput100), .C1(
        keyinput20), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15553), .ZN(n15556) );
  OAI22_X1 U17074 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(keyinput91), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput102), .ZN(n15554) );
  AOI221_X1 U17075 ( .B1(P1_REG2_REG_23__SCAN_IN), .B2(keyinput91), .C1(
        keyinput102), .C2(P1_REG2_REG_14__SCAN_IN), .A(n15554), .ZN(n15555) );
  NAND4_X1 U17076 ( .A1(n15558), .A2(n15557), .A3(n15556), .A4(n15555), .ZN(
        n15568) );
  OAI22_X1 U17077 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(keyinput80), .B1(
        P3_DATAO_REG_15__SCAN_IN), .B2(keyinput113), .ZN(n15559) );
  AOI221_X1 U17078 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(keyinput80), .C1(
        keyinput113), .C2(P3_DATAO_REG_15__SCAN_IN), .A(n15559), .ZN(n15566)
         );
  OAI22_X1 U17079 ( .A1(P3_D_REG_11__SCAN_IN), .A2(keyinput120), .B1(
        P1_REG3_REG_8__SCAN_IN), .B2(keyinput38), .ZN(n15560) );
  AOI221_X1 U17080 ( .B1(P3_D_REG_11__SCAN_IN), .B2(keyinput120), .C1(
        keyinput38), .C2(P1_REG3_REG_8__SCAN_IN), .A(n15560), .ZN(n15565) );
  OAI22_X1 U17081 ( .A1(P3_D_REG_27__SCAN_IN), .A2(keyinput41), .B1(
        P1_REG2_REG_5__SCAN_IN), .B2(keyinput97), .ZN(n15561) );
  AOI221_X1 U17082 ( .B1(P3_D_REG_27__SCAN_IN), .B2(keyinput41), .C1(
        keyinput97), .C2(P1_REG2_REG_5__SCAN_IN), .A(n15561), .ZN(n15564) );
  OAI22_X1 U17083 ( .A1(P3_REG0_REG_3__SCAN_IN), .A2(keyinput89), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput28), .ZN(n15562) );
  AOI221_X1 U17084 ( .B1(P3_REG0_REG_3__SCAN_IN), .B2(keyinput89), .C1(
        keyinput28), .C2(P1_D_REG_29__SCAN_IN), .A(n15562), .ZN(n15563) );
  NAND4_X1 U17085 ( .A1(n15566), .A2(n15565), .A3(n15564), .A4(n15563), .ZN(
        n15567) );
  NOR4_X1 U17086 ( .A1(n15570), .A2(n15569), .A3(n15568), .A4(n15567), .ZN(
        n15608) );
  OAI22_X1 U17087 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput57), .B1(keyinput49), .B2(P1_D_REG_3__SCAN_IN), .ZN(n15571) );
  AOI221_X1 U17088 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput57), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput49), .A(n15571), .ZN(n15578) );
  OAI22_X1 U17089 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(keyinput25), .B1(keyinput15), .B2(P3_ADDR_REG_7__SCAN_IN), .ZN(n15572) );
  AOI221_X1 U17090 ( .B1(P3_IR_REG_8__SCAN_IN), .B2(keyinput25), .C1(
        P3_ADDR_REG_7__SCAN_IN), .C2(keyinput15), .A(n15572), .ZN(n15577) );
  OAI22_X1 U17091 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput78), .B1(
        keyinput124), .B2(P1_REG0_REG_28__SCAN_IN), .ZN(n15573) );
  AOI221_X1 U17092 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput78), .C1(
        P1_REG0_REG_28__SCAN_IN), .C2(keyinput124), .A(n15573), .ZN(n15576) );
  OAI22_X1 U17093 ( .A1(P2_D_REG_11__SCAN_IN), .A2(keyinput19), .B1(
        P1_REG1_REG_27__SCAN_IN), .B2(keyinput65), .ZN(n15574) );
  AOI221_X1 U17094 ( .B1(P2_D_REG_11__SCAN_IN), .B2(keyinput19), .C1(
        keyinput65), .C2(P1_REG1_REG_27__SCAN_IN), .A(n15574), .ZN(n15575) );
  NAND4_X1 U17095 ( .A1(n15578), .A2(n15577), .A3(n15576), .A4(n15575), .ZN(
        n15606) );
  OAI22_X1 U17096 ( .A1(P3_D_REG_2__SCAN_IN), .A2(keyinput39), .B1(keyinput17), 
        .B2(P2_REG3_REG_17__SCAN_IN), .ZN(n15579) );
  AOI221_X1 U17097 ( .B1(P3_D_REG_2__SCAN_IN), .B2(keyinput39), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput17), .A(n15579), .ZN(n15586) );
  OAI22_X1 U17098 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput68), .B1(
        keyinput125), .B2(P1_REG3_REG_4__SCAN_IN), .ZN(n15580) );
  AOI221_X1 U17099 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput68), .C1(
        P1_REG3_REG_4__SCAN_IN), .C2(keyinput125), .A(n15580), .ZN(n15585) );
  OAI22_X1 U17100 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(keyinput101), .B1(
        keyinput60), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n15581) );
  AOI221_X1 U17101 ( .B1(P3_IR_REG_28__SCAN_IN), .B2(keyinput101), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput60), .A(n15581), .ZN(n15584) );
  OAI22_X1 U17102 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput75), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(keyinput109), .ZN(n15582) );
  AOI221_X1 U17103 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput75), .C1(
        keyinput109), .C2(P3_DATAO_REG_14__SCAN_IN), .A(n15582), .ZN(n15583)
         );
  NAND4_X1 U17104 ( .A1(n15586), .A2(n15585), .A3(n15584), .A4(n15583), .ZN(
        n15605) );
  OAI22_X1 U17105 ( .A1(P3_REG0_REG_29__SCAN_IN), .A2(keyinput103), .B1(
        keyinput53), .B2(P1_REG1_REG_12__SCAN_IN), .ZN(n15587) );
  AOI221_X1 U17106 ( .B1(P3_REG0_REG_29__SCAN_IN), .B2(keyinput103), .C1(
        P1_REG1_REG_12__SCAN_IN), .C2(keyinput53), .A(n15587), .ZN(n15594) );
  OAI22_X1 U17107 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput93), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput54), .ZN(n15588) );
  AOI221_X1 U17108 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput93), .C1(
        keyinput54), .C2(P1_REG1_REG_18__SCAN_IN), .A(n15588), .ZN(n15593) );
  OAI22_X1 U17109 ( .A1(P1_D_REG_25__SCAN_IN), .A2(keyinput37), .B1(
        P3_WR_REG_SCAN_IN), .B2(keyinput67), .ZN(n15589) );
  AOI221_X1 U17110 ( .B1(P1_D_REG_25__SCAN_IN), .B2(keyinput37), .C1(
        keyinput67), .C2(P3_WR_REG_SCAN_IN), .A(n15589), .ZN(n15592) );
  OAI22_X1 U17111 ( .A1(P3_D_REG_3__SCAN_IN), .A2(keyinput127), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput59), .ZN(n15590) );
  AOI221_X1 U17112 ( .B1(P3_D_REG_3__SCAN_IN), .B2(keyinput127), .C1(
        keyinput59), .C2(P1_DATAO_REG_21__SCAN_IN), .A(n15590), .ZN(n15591) );
  NAND4_X1 U17113 ( .A1(n15594), .A2(n15593), .A3(n15592), .A4(n15591), .ZN(
        n15604) );
  OAI22_X1 U17114 ( .A1(P3_D_REG_22__SCAN_IN), .A2(keyinput87), .B1(
        keyinput108), .B2(P1_REG0_REG_30__SCAN_IN), .ZN(n15595) );
  AOI221_X1 U17115 ( .B1(P3_D_REG_22__SCAN_IN), .B2(keyinput87), .C1(
        P1_REG0_REG_30__SCAN_IN), .C2(keyinput108), .A(n15595), .ZN(n15602) );
  OAI22_X1 U17116 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput62), .B1(
        P3_DATAO_REG_20__SCAN_IN), .B2(keyinput10), .ZN(n15596) );
  AOI221_X1 U17117 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput62), .C1(
        keyinput10), .C2(P3_DATAO_REG_20__SCAN_IN), .A(n15596), .ZN(n15601) );
  OAI22_X1 U17118 ( .A1(P1_D_REG_18__SCAN_IN), .A2(keyinput29), .B1(
        P1_REG3_REG_20__SCAN_IN), .B2(keyinput44), .ZN(n15597) );
  AOI221_X1 U17119 ( .B1(P1_D_REG_18__SCAN_IN), .B2(keyinput29), .C1(
        keyinput44), .C2(P1_REG3_REG_20__SCAN_IN), .A(n15597), .ZN(n15600) );
  OAI22_X1 U17120 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(keyinput58), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput111), .ZN(n15598) );
  AOI221_X1 U17121 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(keyinput58), .C1(
        keyinput111), .C2(P2_REG3_REG_26__SCAN_IN), .A(n15598), .ZN(n15599) );
  NAND4_X1 U17122 ( .A1(n15602), .A2(n15601), .A3(n15600), .A4(n15599), .ZN(
        n15603) );
  NOR4_X1 U17123 ( .A1(n15606), .A2(n15605), .A3(n15604), .A4(n15603), .ZN(
        n15607) );
  NAND2_X1 U17124 ( .A1(n15608), .A2(n15607), .ZN(n15609) );
  NOR4_X1 U17125 ( .A1(n15612), .A2(n15611), .A3(n15610), .A4(n15609), .ZN(
        n15613) );
  XNOR2_X1 U17126 ( .A(n15614), .B(n15613), .ZN(P3_U3240) );
  XOR2_X1 U17127 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15615), .Z(SUB_1596_U53) );
  AOI21_X1 U17128 ( .B1(n15618), .B2(n15617), .A(n15616), .ZN(SUB_1596_U59) );
  OAI21_X1 U17129 ( .B1(n15621), .B2(n15620), .A(n15619), .ZN(SUB_1596_U58) );
  AOI21_X1 U17130 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(SUB_1596_U56) );
  AOI21_X1 U17131 ( .B1(n15627), .B2(n15626), .A(n15625), .ZN(n15628) );
  XOR2_X1 U17132 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15628), .Z(SUB_1596_U60) );
  AOI21_X1 U17133 ( .B1(n15631), .B2(n15630), .A(n15629), .ZN(SUB_1596_U5) );
  NAND2_X1 U10514 ( .A1(n12429), .A2(n12275), .ZN(n12397) );
  INV_X2 U7388 ( .A(n13488), .ZN(n13066) );
  INV_X2 U7547 ( .A(n13030), .ZN(n13488) );
  CLKBUF_X1 U7416 ( .A(n8605), .Z(n11699) );
  CLKBUF_X1 U7423 ( .A(n8786), .Z(n11317) );
  CLKBUF_X3 U7715 ( .A(n9095), .Z(n9096) );
  CLKBUF_X1 U9092 ( .A(n11704), .Z(n11671) );
endmodule

