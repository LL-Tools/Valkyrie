

module b14_C_AntiSAT_k_256_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991;

  INV_X1 U2461 ( .A(n2896), .ZN(n3028) );
  INV_X1 U2462 ( .A(n3030), .ZN(n2872) );
  AOI21_X1 U2463 ( .B1(n3111), .B2(n3115), .A(n2232), .ZN(n3117) );
  INV_X1 U2464 ( .A(IR_REG_31__SCAN_IN), .ZN(n2784) );
  NOR2_X1 U2465 ( .A1(n3123), .A2(n3124), .ZN(n3122) );
  AOI21_X2 U2466 ( .B1(n3631), .B2(n3633), .A(n3632), .ZN(n3697) );
  OAI21_X2 U2467 ( .B1(n4173), .B2(n4153), .A(n2705), .ZN(n4121) );
  OAI21_X2 U2468 ( .B1(n3132), .B2(n3131), .A(n2902), .ZN(n3183) );
  NOR2_X2 U2469 ( .A1(n3122), .A2(n2483), .ZN(n3132) );
  INV_X1 U2470 ( .A(n2719), .ZN(n2218) );
  AOI21_X2 U2471 ( .B1(n3494), .B2(n2452), .A(n2449), .ZN(n3547) );
  OAI21_X2 U2472 ( .B1(n3386), .B2(n2933), .A(n2932), .ZN(n3494) );
  NOR2_X1 U2473 ( .A1(n4202), .A2(n4560), .ZN(n4504) );
  NAND4_X1 U2474 ( .A1(n2548), .A2(n2547), .A3(n2546), .A4(n2545), .ZN(n3898)
         );
  INV_X2 U2475 ( .A(n2867), .ZN(n3104) );
  BUF_X2 U2477 ( .A(n2220), .Z(n3086) );
  AND2_X1 U2478 ( .A1(n2864), .A2(n2863), .ZN(n2895) );
  INV_X1 U2479 ( .A(n2719), .ZN(n2513) );
  NOR2_X1 U2480 ( .A1(n2504), .A2(n4319), .ZN(n2526) );
  BUF_X1 U2481 ( .A(n2862), .Z(n3146) );
  NAND2_X1 U2482 ( .A1(n4472), .A2(n2268), .ZN(n3959) );
  NAND2_X1 U2483 ( .A1(n4473), .A2(n4474), .ZN(n4472) );
  NAND2_X1 U2484 ( .A1(n3424), .A2(n2929), .ZN(n3385) );
  NAND2_X1 U2485 ( .A1(n2465), .A2(n2464), .ZN(n3424) );
  NAND2_X1 U2486 ( .A1(n3448), .A2(n4444), .ZN(n3952) );
  NAND2_X1 U2487 ( .A1(n3315), .A2(n2468), .ZN(n2465) );
  NAND2_X1 U2488 ( .A1(n4385), .A2(n3440), .ZN(n4397) );
  NAND2_X1 U2489 ( .A1(n2896), .A2(n4560), .ZN(n2887) );
  NAND2_X1 U2490 ( .A1(n4368), .A2(n2240), .ZN(n3439) );
  CLKBUF_X3 U2492 ( .A(n2895), .Z(n3015) );
  NAND2_X1 U2493 ( .A1(n4369), .A2(n4370), .ZN(n4368) );
  INV_X1 U2494 ( .A(n2895), .ZN(n2219) );
  NAND3_X1 U2495 ( .A1(n4324), .A2(n3072), .A3(n4323), .ZN(n2864) );
  NAND2_X1 U2496 ( .A1(n2273), .A2(n2272), .ZN(n4369) );
  INV_X1 U2497 ( .A(n2879), .ZN(n4500) );
  OR2_X1 U2498 ( .A1(n3934), .A2(n3437), .ZN(n2273) );
  INV_X2 U2499 ( .A(n3082), .ZN(n3806) );
  AND2_X1 U2500 ( .A1(n2817), .A2(n2870), .ZN(n2482) );
  NAND2_X1 U2501 ( .A1(n4335), .A2(n2311), .ZN(n3436) );
  NAND2_X1 U2502 ( .A1(n2770), .A2(IR_REG_31__SCAN_IN), .ZN(n2771) );
  XNOR2_X1 U2503 ( .A(n2780), .B(n2820), .ZN(n2870) );
  MUX2_X1 U2504 ( .A(IR_REG_31__SCAN_IN), .B(n2502), .S(IR_REG_29__SCAN_IN), 
        .Z(n2503) );
  NAND2_X1 U2505 ( .A1(n2501), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  OR2_X1 U2506 ( .A1(n2779), .A2(n2784), .ZN(n2773) );
  AND2_X1 U2507 ( .A1(n2779), .A2(n2778), .ZN(n2821) );
  AND2_X1 U2508 ( .A1(n2702), .A2(n4727), .ZN(n2779) );
  NOR2_X1 U2509 ( .A1(n2825), .A2(n2358), .ZN(n2267) );
  INV_X1 U2510 ( .A(n2540), .ZN(n2490) );
  AND3_X1 U2511 ( .A1(n2479), .A2(n2601), .A3(n2426), .ZN(n2425) );
  AND2_X1 U2512 ( .A1(n2493), .A2(n2235), .ZN(n2360) );
  AND2_X1 U2513 ( .A1(n2549), .A2(n2489), .ZN(n2479) );
  AND3_X1 U2514 ( .A1(n2295), .A2(n2294), .A3(n2293), .ZN(n2493) );
  INV_X1 U2515 ( .A(IR_REG_22__SCAN_IN), .ZN(n2820) );
  INV_X1 U2516 ( .A(IR_REG_19__SCAN_IN), .ZN(n2776) );
  INV_X1 U2517 ( .A(IR_REG_23__SCAN_IN), .ZN(n2840) );
  INV_X1 U2518 ( .A(IR_REG_3__SCAN_IN), .ZN(n2549) );
  NOR2_X1 U2519 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2601)
         );
  INV_X1 U2520 ( .A(IR_REG_16__SCAN_IN), .ZN(n2692) );
  INV_X1 U2521 ( .A(IR_REG_15__SCAN_IN), .ZN(n4726) );
  BUF_X4 U2522 ( .A(n2526), .Z(n2220) );
  AOI21_X2 U2523 ( .B1(n3697), .B2(n3698), .A(n3699), .ZN(n3592) );
  AOI21_X2 U2524 ( .B1(n3294), .B2(n3295), .A(n2477), .ZN(n3315) );
  AND2_X4 U2525 ( .A1(n3074), .A2(n4319), .ZN(n2527) );
  OR2_X4 U2526 ( .A1(n4319), .A2(n3074), .ZN(n2535) );
  NOR2_X1 U2527 ( .A1(n3508), .A2(n3377), .ZN(n2632) );
  AOI21_X1 U2528 ( .B1(n2348), .B2(n2347), .A(n2613), .ZN(n2346) );
  INV_X1 U2529 ( .A(n2352), .ZN(n2347) );
  AOI21_X1 U2530 ( .B1(n2328), .B2(n3816), .A(n2227), .ZN(n2327) );
  NOR2_X1 U2531 ( .A1(n4428), .A2(n2263), .ZN(n3473) );
  OR2_X1 U2532 ( .A1(n3307), .A2(n3303), .ZN(n2794) );
  INV_X1 U2533 ( .A(IR_REG_13__SCAN_IN), .ZN(n2426) );
  NOR2_X1 U2534 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2496)
         );
  AND4_X1 U2535 ( .A1(n2840), .A2(n2692), .A3(n2494), .A4(n2820), .ZN(n2497)
         );
  NOR2_X1 U2536 ( .A1(n3351), .A2(n2469), .ZN(n2468) );
  INV_X1 U2537 ( .A(n3317), .ZN(n2469) );
  NOR2_X1 U2538 ( .A1(n2446), .A2(n2443), .ZN(n2442) );
  INV_X1 U2539 ( .A(n2978), .ZN(n2443) );
  INV_X1 U2540 ( .A(n2447), .ZN(n2446) );
  XNOR2_X1 U2541 ( .A(n3473), .B(n2310), .ZN(n4439) );
  OR2_X1 U2542 ( .A1(n4439), .A2(n4440), .ZN(n2290) );
  NOR2_X1 U2543 ( .A1(n3959), .A2(n3960), .ZN(n3966) );
  AND2_X1 U2544 ( .A1(n3817), .A2(n2259), .ZN(n2328) );
  OR2_X1 U2545 ( .A1(n4170), .A2(n4196), .ZN(n2696) );
  NOR2_X1 U2546 ( .A1(n3888), .A2(n3534), .ZN(n2660) );
  NAND2_X1 U2547 ( .A1(n3890), .A2(n3407), .ZN(n2644) );
  AOI21_X1 U2548 ( .B1(n2346), .B2(n2349), .A(n2243), .ZN(n2345) );
  NAND2_X1 U2549 ( .A1(n2336), .A2(n2306), .ZN(n2541) );
  NAND2_X1 U2550 ( .A1(n3449), .A2(IR_REG_28__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2551 ( .A1(n3450), .A2(n2498), .ZN(n2336) );
  NAND2_X1 U2552 ( .A1(n4476), .A2(n4477), .ZN(n4475) );
  AND2_X1 U2553 ( .A1(n4088), .A2(n4085), .ZN(n3854) );
  AND2_X1 U2554 ( .A1(n2373), .A2(n3854), .ZN(n2372) );
  NAND2_X1 U2555 ( .A1(n2376), .A2(n2374), .ZN(n2373) );
  AOI21_X1 U2556 ( .B1(n2460), .B2(n2456), .A(n2455), .ZN(n2454) );
  INV_X1 U2557 ( .A(n3503), .ZN(n2455) );
  INV_X1 U2558 ( .A(n3491), .ZN(n2456) );
  NAND2_X1 U2559 ( .A1(n2454), .A2(n2461), .ZN(n2451) );
  NAND2_X1 U2560 ( .A1(n2457), .A2(n3490), .ZN(n2450) );
  CLKBUF_X1 U2561 ( .A(n2887), .Z(n3029) );
  NAND2_X1 U2562 ( .A1(n2313), .A2(n4337), .ZN(n2311) );
  NOR2_X1 U2563 ( .A1(n4981), .A2(n2314), .ZN(n3956) );
  AND2_X1 U2564 ( .A1(n4516), .A2(REG2_REG_15__SCAN_IN), .ZN(n2314) );
  INV_X1 U2565 ( .A(n2541), .ZN(n3082) );
  INV_X1 U2566 ( .A(n3856), .ZN(n2402) );
  INV_X1 U2567 ( .A(n4013), .ZN(n2403) );
  OR2_X1 U2568 ( .A1(n4031), .A2(n3725), .ZN(n2809) );
  NOR2_X1 U2569 ( .A1(n2368), .A2(n2363), .ZN(n2362) );
  INV_X1 U2570 ( .A(n3747), .ZN(n2363) );
  INV_X1 U2571 ( .A(n3765), .ZN(n2367) );
  INV_X1 U2572 ( .A(n3766), .ZN(n2366) );
  NOR2_X1 U2573 ( .A1(n2592), .A2(n2353), .ZN(n2352) );
  INV_X1 U2574 ( .A(n2581), .ZN(n2353) );
  NAND2_X1 U2575 ( .A1(n2790), .A2(n3740), .ZN(n2384) );
  INV_X1 U2576 ( .A(n2385), .ZN(n2381) );
  NOR2_X1 U2577 ( .A1(n3140), .A2(n2386), .ZN(n2385) );
  INV_X1 U2578 ( .A(n3740), .ZN(n2386) );
  NAND2_X1 U2579 ( .A1(n3733), .A2(n3731), .ZN(n3792) );
  INV_X1 U2580 ( .A(n3792), .ZN(n3196) );
  NAND2_X1 U2581 ( .A1(n2509), .A2(n2359), .ZN(n2358) );
  INV_X1 U2582 ( .A(IR_REG_4__SCAN_IN), .ZN(n2489) );
  INV_X1 U2583 ( .A(IR_REG_5__SCAN_IN), .ZN(n2492) );
  INV_X1 U2584 ( .A(IR_REG_9__SCAN_IN), .ZN(n2491) );
  INV_X1 U2585 ( .A(IR_REG_12__SCAN_IN), .ZN(n2293) );
  INV_X1 U2586 ( .A(IR_REG_2__SCAN_IN), .ZN(n2488) );
  OR2_X1 U2587 ( .A1(n3252), .A2(n3251), .ZN(n2472) );
  NAND2_X1 U2588 ( .A1(n3026), .A2(n3027), .ZN(n2440) );
  NOR2_X1 U2589 ( .A1(n2572), .A2(n2571), .ZN(n2583) );
  INV_X1 U2590 ( .A(n4132), .ZN(n3626) );
  NAND2_X1 U2591 ( .A1(n2717), .A2(REG3_REG_23__SCAN_IN), .ZN(n2727) );
  OR2_X1 U2592 ( .A1(n2594), .A2(n2593), .ZN(n2605) );
  NAND2_X1 U2593 ( .A1(n2979), .A2(n2978), .ZN(n3666) );
  NOR2_X1 U2594 ( .A1(n2990), .A2(n2448), .ZN(n2447) );
  INV_X1 U2595 ( .A(n3679), .ZN(n2992) );
  NOR2_X1 U2596 ( .A1(n2466), .A2(n3427), .ZN(n2464) );
  AOI22_X1 U2597 ( .A1(n2894), .A2(n2889), .B1(n3043), .B2(n2888), .ZN(n2892)
         );
  XNOR2_X1 U2598 ( .A(n2886), .B(n3030), .ZN(n2891) );
  NAND2_X1 U2599 ( .A1(n2418), .A2(n2422), .ZN(n3685) );
  INV_X1 U2600 ( .A(n2423), .ZN(n2422) );
  OAI21_X1 U2601 ( .B1(n3646), .B2(n2424), .A(n3687), .ZN(n2423) );
  AND2_X1 U2602 ( .A1(n3015), .A2(n3042), .ZN(n3878) );
  OAI211_X1 U2603 ( .C1(n2414), .C2(n4584), .A(n2411), .B(n2410), .ZN(n3925)
         );
  OR2_X1 U2604 ( .A1(n2412), .A2(n4584), .ZN(n2411) );
  XNOR2_X1 U2605 ( .A(n3456), .B(n4330), .ZN(n3933) );
  NAND2_X1 U2606 ( .A1(n4374), .A2(n2236), .ZN(n3460) );
  NAND2_X1 U2607 ( .A1(n4396), .A2(n3441), .ZN(n3442) );
  OAI22_X1 U2608 ( .A1(n4392), .A2(n4390), .B1(REG1_REG_7__SCAN_IN), .B2(n4524), .ZN(n3462) );
  NOR2_X1 U2609 ( .A1(n4411), .A2(n3467), .ZN(n3470) );
  AND2_X1 U2610 ( .A1(n3466), .A2(REG1_REG_9__SCAN_IN), .ZN(n3467) );
  OR2_X1 U2611 ( .A1(n4421), .A2(n4836), .ZN(n2279) );
  NAND2_X1 U2612 ( .A1(n2290), .A2(n2239), .ZN(n2406) );
  NAND2_X1 U2613 ( .A1(n2406), .A2(n2405), .ZN(n3943) );
  INV_X1 U2614 ( .A(n3476), .ZN(n2405) );
  NAND2_X1 U2615 ( .A1(n2409), .A2(REG1_REG_14__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U2616 ( .A1(n3945), .A2(n2409), .ZN(n2407) );
  INV_X1 U2617 ( .A(n4977), .ZN(n2409) );
  XNOR2_X1 U2618 ( .A(n3956), .B(n2670), .ZN(n4463) );
  NAND2_X1 U2619 ( .A1(n4463), .A2(n4462), .ZN(n4461) );
  NOR2_X1 U2620 ( .A1(n4976), .A2(n2291), .ZN(n3946) );
  AND2_X1 U2621 ( .A1(n4516), .A2(REG1_REG_15__SCAN_IN), .ZN(n2291) );
  OAI21_X1 U2622 ( .B1(n2327), .B2(n2326), .A(n2254), .ZN(n2325) );
  OR2_X1 U2623 ( .A1(n2762), .A2(n3051), .ZN(n3982) );
  OR2_X1 U2624 ( .A1(n3816), .A2(n2322), .ZN(n2321) );
  NAND2_X1 U2625 ( .A1(n2747), .A2(n2746), .ZN(n2322) );
  OR2_X1 U2626 ( .A1(n2737), .A2(n3638), .ZN(n2748) );
  AND2_X1 U2627 ( .A1(n4148), .A2(n4131), .ZN(n2712) );
  AND2_X1 U2628 ( .A1(n2249), .A2(n4104), .ZN(n2356) );
  AND2_X1 U2629 ( .A1(n4151), .A2(n4175), .ZN(n2703) );
  AND2_X1 U2630 ( .A1(n2662), .A2(REG3_REG_16__SCAN_IN), .ZN(n2683) );
  AND2_X1 U2631 ( .A1(n4347), .A2(n3563), .ZN(n2681) );
  INV_X1 U2632 ( .A(n3889), .ZN(n3537) );
  NAND2_X1 U2633 ( .A1(n2222), .A2(n2341), .ZN(n2340) );
  NOR2_X1 U2634 ( .A1(n3824), .A2(n2343), .ZN(n2342) );
  INV_X1 U2635 ( .A(n2644), .ZN(n2343) );
  OAI21_X1 U2636 ( .B1(n3371), .B2(n2390), .A(n2388), .ZN(n3531) );
  AOI21_X1 U2637 ( .B1(n2391), .B2(n2389), .A(n2341), .ZN(n2388) );
  INV_X1 U2638 ( .A(n2391), .ZN(n2390) );
  INV_X1 U2639 ( .A(n2393), .ZN(n2389) );
  NAND2_X1 U2640 ( .A1(n2387), .A2(n2391), .ZN(n3840) );
  NAND2_X1 U2641 ( .A1(n3371), .A2(n2393), .ZN(n2387) );
  INV_X1 U2642 ( .A(n3890), .ZN(n3550) );
  OAI21_X1 U2643 ( .B1(n3371), .B2(n3768), .A(n3763), .ZN(n3406) );
  OR2_X1 U2644 ( .A1(n2605), .A2(n3420), .ZN(n2614) );
  INV_X1 U2645 ( .A(n3892), .ZN(n3365) );
  INV_X1 U2646 ( .A(n3893), .ZN(n3332) );
  AOI21_X1 U2647 ( .B1(n2399), .B2(n2397), .A(n2396), .ZN(n2395) );
  INV_X1 U2648 ( .A(n2399), .ZN(n2398) );
  INV_X1 U2649 ( .A(n3753), .ZN(n2396) );
  NOR2_X1 U2650 ( .A1(n2237), .A2(n2331), .ZN(n2330) );
  NAND2_X1 U2651 ( .A1(n3728), .A2(n3730), .ZN(n4492) );
  AND2_X1 U2652 ( .A1(n2867), .A2(n4533), .ZN(n4483) );
  NAND2_X1 U2653 ( .A1(n4483), .A2(n4492), .ZN(n4485) );
  OR2_X1 U2654 ( .A1(n4022), .A2(n2857), .ZN(n3999) );
  INV_X1 U2655 ( .A(n4169), .ZN(n4175) );
  NAND2_X1 U2656 ( .A1(n4197), .A2(n2301), .ZN(n4174) );
  NOR2_X1 U2657 ( .A1(n4268), .A2(n3563), .ZN(n4197) );
  AND2_X1 U2658 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2510)
         );
  CLKBUF_X1 U2659 ( .A(n2864), .Z(n2869) );
  AND2_X1 U2660 ( .A1(n2439), .A2(n2430), .ZN(n2429) );
  AND2_X1 U2661 ( .A1(n3591), .A2(n4353), .ZN(n2430) );
  OR2_X1 U2662 ( .A1(n2434), .A2(n3722), .ZN(n2432) );
  OAI21_X1 U2663 ( .B1(n2439), .B2(n2436), .A(n2435), .ZN(n2434) );
  NOR2_X1 U2664 ( .A1(n3591), .A2(n2437), .ZN(n2436) );
  NAND2_X1 U2665 ( .A1(n2439), .A2(n2440), .ZN(n2435) );
  NAND2_X1 U2666 ( .A1(n3034), .A2(n2440), .ZN(n2438) );
  INV_X1 U2667 ( .A(n3887), .ZN(n4173) );
  INV_X1 U2668 ( .A(n4343), .ZN(n3714) );
  INV_X1 U2669 ( .A(n4071), .ZN(n4106) );
  INV_X1 U2670 ( .A(n3160), .ZN(n4533) );
  INV_X1 U2671 ( .A(n4196), .ZN(n3693) );
  INV_X1 U2672 ( .A(n3276), .ZN(n3895) );
  NAND2_X1 U2673 ( .A1(n4375), .A2(n4376), .ZN(n4374) );
  NAND2_X1 U2674 ( .A1(n4397), .A2(n4398), .ZN(n4396) );
  NAND2_X1 U2675 ( .A1(n4408), .A2(REG2_REG_8__SCAN_IN), .ZN(n4407) );
  NOR2_X1 U2676 ( .A1(n2234), .A2(n4412), .ZN(n4411) );
  XNOR2_X1 U2677 ( .A(n3470), .B(n3469), .ZN(n4421) );
  XNOR2_X1 U2678 ( .A(n3946), .B(n2670), .ZN(n4466) );
  NAND2_X1 U2679 ( .A1(n4466), .A2(n4465), .ZN(n4464) );
  NAND2_X1 U2680 ( .A1(n4479), .A2(n2285), .ZN(n2284) );
  NOR2_X1 U2681 ( .A1(n2287), .A2(n3948), .ZN(n2285) );
  INV_X1 U2682 ( .A(n3965), .ZN(n2287) );
  NAND2_X1 U2683 ( .A1(n4475), .A2(n2269), .ZN(n3949) );
  XNOR2_X1 U2684 ( .A(n2309), .B(n3969), .ZN(n3974) );
  NAND2_X1 U2685 ( .A1(n2324), .A2(n2327), .ZN(n3996) );
  NAND2_X1 U2686 ( .A1(n4029), .A2(n2328), .ZN(n2324) );
  NAND2_X1 U2687 ( .A1(n2296), .A2(n4345), .ZN(n4268) );
  INV_X1 U2688 ( .A(n3645), .ZN(n2424) );
  NOR2_X1 U2689 ( .A1(n2424), .A2(n2420), .ZN(n2419) );
  INV_X1 U2690 ( .A(n2961), .ZN(n2420) );
  INV_X1 U2691 ( .A(n3925), .ZN(n2417) );
  NOR2_X1 U2692 ( .A1(n3923), .A2(n2241), .ZN(n3455) );
  AND2_X1 U2693 ( .A1(n3794), .A2(n4048), .ZN(n3863) );
  NAND2_X1 U2694 ( .A1(n2370), .A2(n2369), .ZN(n4066) );
  AOI21_X1 U2695 ( .B1(n2372), .B2(n2375), .A(n3855), .ZN(n2369) );
  INV_X1 U2696 ( .A(n2376), .ZN(n2375) );
  AOI21_X1 U2697 ( .B1(n3726), .B2(n4143), .A(n2377), .ZN(n2376) );
  INV_X1 U2698 ( .A(n3849), .ZN(n4143) );
  OR2_X1 U2699 ( .A1(n3558), .A2(n3780), .ZN(n4139) );
  NOR2_X1 U2700 ( .A1(n3404), .A2(n2394), .ZN(n2393) );
  AOI21_X1 U2701 ( .B1(n2393), .B2(n3768), .A(n2392), .ZN(n2391) );
  INV_X1 U2702 ( .A(n3333), .ZN(n2350) );
  AND2_X1 U2703 ( .A1(n3746), .A2(n2400), .ZN(n2399) );
  INV_X1 U2704 ( .A(n3754), .ZN(n2397) );
  INV_X1 U2705 ( .A(n2333), .ZN(n2331) );
  OR2_X1 U2706 ( .A1(n3897), .A2(n3153), .ZN(n2333) );
  NAND2_X1 U2707 ( .A1(n2554), .A2(n2334), .ZN(n2332) );
  NOR2_X1 U2708 ( .A1(n2562), .A2(n2335), .ZN(n2334) );
  NAND2_X1 U2709 ( .A1(n4490), .A2(n2888), .ZN(n3731) );
  NAND2_X1 U2710 ( .A1(n2879), .A2(n2875), .ZN(n3728) );
  AND2_X1 U2711 ( .A1(n4325), .A2(n2816), .ZN(n3083) );
  NOR2_X1 U2712 ( .A1(n4070), .A2(n4092), .ZN(n2303) );
  AND2_X1 U2713 ( .A1(n3693), .A2(n4175), .ZN(n2301) );
  OR2_X1 U2714 ( .A1(n3376), .A2(n3377), .ZN(n3375) );
  NOR2_X1 U2715 ( .A1(n2300), .A2(n3224), .ZN(n2298) );
  NAND2_X1 U2716 ( .A1(n3298), .A2(n3267), .ZN(n2300) );
  INV_X1 U2717 ( .A(n3165), .ZN(n2299) );
  INV_X1 U2718 ( .A(IR_REG_20__SCAN_IN), .ZN(n2777) );
  INV_X1 U2719 ( .A(IR_REG_8__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U2720 ( .A1(n2453), .A2(n2458), .ZN(n2452) );
  NAND2_X1 U2721 ( .A1(n2451), .A2(n2450), .ZN(n2449) );
  INV_X1 U2722 ( .A(n2454), .ZN(n2453) );
  OAI21_X1 U2723 ( .B1(n3351), .B2(n2467), .A(n2925), .ZN(n2466) );
  INV_X1 U2724 ( .A(n2440), .ZN(n2437) );
  OAI22_X1 U2725 ( .A1(n3152), .A2(n3019), .B1(n3028), .B2(n3180), .ZN(n2903)
         );
  OAI22_X1 U2726 ( .A1(n3550), .A2(n3029), .B1(n3019), .B2(n3511), .ZN(n3503)
         );
  NAND2_X1 U2727 ( .A1(n2220), .A2(REG2_REG_1__SCAN_IN), .ZN(n2515) );
  OR2_X1 U2728 ( .A1(n2535), .A2(n2512), .ZN(n2518) );
  INV_X1 U2729 ( .A(n2957), .ZN(n2958) );
  OR2_X1 U2730 ( .A1(n2634), .A2(n4718), .ZN(n2651) );
  NAND2_X1 U2731 ( .A1(n2220), .A2(REG2_REG_0__SCAN_IN), .ZN(n2521) );
  AOI21_X1 U2732 ( .B1(n2338), .B2(n2416), .A(n2288), .ZN(n3923) );
  NAND2_X1 U2733 ( .A1(n3454), .A2(REG1_REG_1__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U2734 ( .A1(n2417), .A2(n2289), .ZN(n2288) );
  NAND2_X1 U2735 ( .A1(n3902), .A2(n2415), .ZN(n2289) );
  NAND2_X1 U2736 ( .A1(n2315), .A2(REG1_REG_1__SCAN_IN), .ZN(n3924) );
  OAI211_X1 U2737 ( .C1(REG1_REG_1__SCAN_IN), .C2(n2315), .A(n3924), .B(n3454), 
        .ZN(n3926) );
  OR2_X1 U2738 ( .A1(n3917), .A2(n2247), .ZN(n2313) );
  XNOR2_X1 U2739 ( .A(n3455), .B(n4337), .ZN(n4334) );
  INV_X1 U2740 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3420) );
  NAND2_X1 U2741 ( .A1(n4415), .A2(n3444), .ZN(n3445) );
  INV_X1 U2742 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U2743 ( .A1(n4433), .A2(n2264), .ZN(n3447) );
  OAI22_X1 U2744 ( .A1(n3952), .A2(n3951), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4328), .ZN(n3953) );
  AND2_X1 U2745 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  NAND2_X1 U2746 ( .A1(n4461), .A2(n3957), .ZN(n4473) );
  NOR2_X1 U2747 ( .A1(n3966), .A2(n2271), .ZN(n2309) );
  AOI21_X1 U2748 ( .B1(n2809), .B2(n2253), .A(n2401), .ZN(n3987) );
  OR2_X1 U2749 ( .A1(n2258), .A2(n3984), .ZN(n2401) );
  NOR2_X1 U2750 ( .A1(n3999), .A2(n4000), .ZN(n4210) );
  NAND2_X1 U2751 ( .A1(n4016), .A2(n3856), .ZN(n3986) );
  NAND2_X1 U2752 ( .A1(n2809), .A2(n3836), .ZN(n4014) );
  AND2_X1 U2753 ( .A1(n2769), .A2(n2768), .ZN(n4019) );
  AND2_X1 U2754 ( .A1(n3806), .A2(DATAI_24_), .ZN(n4070) );
  AOI21_X1 U2755 ( .B1(n2356), .B2(n2712), .A(n2256), .ZN(n2355) );
  AND2_X1 U2756 ( .A1(n2733), .A2(n2732), .ZN(n4095) );
  NOR2_X1 U2757 ( .A1(n2708), .A2(n2707), .ZN(n2713) );
  NAND2_X1 U2758 ( .A1(n2371), .A2(n2376), .ZN(n4129) );
  NAND2_X1 U2759 ( .A1(n4139), .A2(n3726), .ZN(n2371) );
  AND2_X1 U2760 ( .A1(n4197), .A2(n2265), .ZN(n4123) );
  AND2_X1 U2761 ( .A1(n2701), .A2(n2700), .ZN(n4151) );
  NAND2_X1 U2762 ( .A1(n2683), .A2(n2487), .ZN(n2698) );
  NOR2_X1 U2763 ( .A1(n4272), .A2(n3534), .ZN(n2296) );
  NAND2_X1 U2764 ( .A1(n3843), .A2(n3848), .ZN(n3826) );
  NAND2_X1 U2765 ( .A1(n2339), .A2(n2223), .ZN(n2661) );
  NOR2_X1 U2766 ( .A1(n3375), .A2(n3407), .ZN(n3414) );
  AOI21_X1 U2767 ( .B1(n3759), .B2(n2367), .A(n2366), .ZN(n2365) );
  AND2_X1 U2768 ( .A1(n3497), .A2(n3391), .ZN(n2621) );
  NOR2_X1 U2769 ( .A1(n2614), .A2(n4918), .ZN(n2622) );
  NAND2_X1 U2770 ( .A1(n2364), .A2(n3759), .ZN(n3360) );
  NAND2_X1 U2771 ( .A1(n3327), .A2(n3765), .ZN(n2364) );
  NAND2_X1 U2772 ( .A1(n2794), .A2(n3747), .ZN(n3327) );
  NAND2_X1 U2773 ( .A1(n2351), .A2(n2591), .ZN(n3334) );
  NAND2_X1 U2774 ( .A1(n2582), .A2(n2352), .ZN(n2351) );
  AND2_X1 U2775 ( .A1(n2575), .A2(n2574), .ZN(n3276) );
  INV_X1 U2776 ( .A(n4493), .ZN(n4167) );
  AOI21_X1 U2777 ( .B1(n2382), .B2(n2381), .A(n2380), .ZN(n2378) );
  INV_X1 U2778 ( .A(n3752), .ZN(n2380) );
  AND3_X1 U2779 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2780 ( .A1(n2563), .A2(REG3_REG_6__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U2781 ( .A1(n2379), .A2(n2382), .ZN(n3223) );
  NAND2_X1 U2782 ( .A1(n3168), .A2(n2385), .ZN(n2379) );
  INV_X1 U2783 ( .A(n3898), .ZN(n3152) );
  OAI21_X1 U2784 ( .B1(n3168), .B2(n2790), .A(n3740), .ZN(n3148) );
  NOR2_X1 U2785 ( .A1(n3165), .A2(n3153), .ZN(n3231) );
  OR2_X1 U2786 ( .A1(n3218), .A2(n3169), .ZN(n3165) );
  NAND2_X1 U2787 ( .A1(n3083), .A2(n4321), .ZN(n4188) );
  INV_X1 U2788 ( .A(n4489), .ZN(n4185) );
  NAND2_X1 U2789 ( .A1(n4038), .A2(n4023), .ZN(n4022) );
  AND2_X1 U2790 ( .A1(n4113), .A2(n2302), .ZN(n4038) );
  AND2_X1 U2791 ( .A1(n2230), .A2(n4040), .ZN(n2302) );
  INV_X1 U2792 ( .A(n4070), .ZN(n4076) );
  NAND2_X1 U2793 ( .A1(n4113), .A2(n2303), .ZN(n4075) );
  AND2_X1 U2794 ( .A1(n4123), .A2(n4114), .ZN(n4113) );
  NAND2_X1 U2795 ( .A1(n4113), .A2(n4097), .ZN(n4096) );
  NAND2_X1 U2796 ( .A1(n4197), .A2(n2229), .ZN(n4152) );
  INV_X1 U2797 ( .A(n2296), .ZN(n3576) );
  NAND2_X1 U2798 ( .A1(n3367), .A2(n3391), .ZN(n3376) );
  NOR2_X1 U2799 ( .A1(n3304), .A2(n3309), .ZN(n3336) );
  AND2_X1 U2800 ( .A1(n3336), .A2(n3423), .ZN(n3367) );
  NAND2_X1 U2801 ( .A1(n2299), .A2(n2297), .ZN(n3304) );
  AND2_X1 U2802 ( .A1(n2298), .A2(n3322), .ZN(n2297) );
  NAND2_X1 U2803 ( .A1(n2299), .A2(n2298), .ZN(n3279) );
  NOR3_X1 U2804 ( .A1(n3165), .A2(n3224), .A3(n3153), .ZN(n4561) );
  NAND2_X1 U2805 ( .A1(n4485), .A2(n2524), .ZN(n3197) );
  AND3_X1 U2806 ( .A1(n2856), .A2(n2855), .A3(n2854), .ZN(n3063) );
  NAND2_X1 U2807 ( .A1(n2509), .A2(n2242), .ZN(n2474) );
  INV_X1 U2808 ( .A(IR_REG_29__SCAN_IN), .ZN(n4871) );
  NOR2_X1 U2809 ( .A1(n2267), .A2(n2244), .ZN(n3450) );
  AND3_X1 U2810 ( .A1(n2425), .A2(n2359), .A3(n2490), .ZN(n2304) );
  OR2_X1 U2811 ( .A1(n2821), .A2(n2784), .ZN(n2780) );
  INV_X1 U2812 ( .A(IR_REG_21__SCAN_IN), .ZN(n2775) );
  INV_X1 U2813 ( .A(IR_REG_17__SCAN_IN), .ZN(n2691) );
  AND3_X1 U2814 ( .A1(n2235), .A2(n2479), .A3(n2601), .ZN(n2427) );
  INV_X1 U2815 ( .A(IR_REG_7__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U2816 ( .A1(n2278), .A2(n2413), .ZN(n2412) );
  NOR2_X1 U2817 ( .A1(n2784), .A2(IR_REG_2__SCAN_IN), .ZN(n2278) );
  OAI21_X1 U2818 ( .B1(n2533), .B2(n2784), .A(IR_REG_2__SCAN_IN), .ZN(n2414)
         );
  INV_X1 U2819 ( .A(n3245), .ZN(n3298) );
  AOI22_X1 U2820 ( .A1(n2473), .A2(n3252), .B1(n3251), .B2(n2221), .ZN(n2470)
         );
  OR2_X1 U2821 ( .A1(n2221), .A2(n3251), .ZN(n2473) );
  AND2_X1 U2822 ( .A1(n2755), .A2(n2762), .ZN(n4024) );
  NAND2_X1 U2823 ( .A1(n2465), .A2(n2463), .ZN(n3426) );
  INV_X1 U2824 ( .A(n2466), .ZN(n2463) );
  INV_X1 U2825 ( .A(n3735), .ZN(n3216) );
  INV_X1 U2826 ( .A(n2889), .ZN(n4490) );
  NAND2_X1 U2827 ( .A1(n3665), .A2(n3668), .ZN(n3622) );
  INV_X1 U2828 ( .A(n3891), .ZN(n3497) );
  INV_X1 U2829 ( .A(n3896), .ZN(n3266) );
  AOI21_X1 U2830 ( .B1(n3315), .B2(n3317), .A(n3316), .ZN(n3350) );
  NAND2_X1 U2831 ( .A1(n2459), .A2(n3491), .ZN(n3506) );
  OR2_X1 U2832 ( .A1(n3494), .A2(n3490), .ZN(n2459) );
  AOI21_X1 U2833 ( .B1(n2447), .B2(n2445), .A(n2252), .ZN(n2444) );
  INV_X1 U2834 ( .A(n3667), .ZN(n2445) );
  INV_X1 U2835 ( .A(n3362), .ZN(n3391) );
  NAND2_X1 U2836 ( .A1(n2927), .A2(n2928), .ZN(n2929) );
  NAND2_X1 U2837 ( .A1(n2881), .A2(n2880), .ZN(n2883) );
  XNOR2_X1 U2838 ( .A(n2891), .B(n2890), .ZN(n3124) );
  OR2_X1 U2839 ( .A1(n3058), .A2(n3049), .ZN(n3704) );
  NAND2_X1 U2840 ( .A1(n2421), .A2(n3645), .ZN(n3686) );
  NAND2_X1 U2841 ( .A1(n3644), .A2(n3646), .ZN(n2421) );
  AND2_X1 U2842 ( .A1(n3059), .A2(n3102), .ZN(n4358) );
  INV_X1 U2843 ( .A(n4034), .ZN(n4074) );
  OR2_X1 U2844 ( .A1(n3058), .A2(n3044), .ZN(n4343) );
  INV_X1 U2845 ( .A(n3534), .ZN(n3717) );
  INV_X1 U2846 ( .A(n4358), .ZN(n3720) );
  NAND2_X1 U2847 ( .A1(n2724), .A2(n2723), .ZN(n4071) );
  NAND4_X1 U2848 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3887)
         );
  INV_X1 U2849 ( .A(n4151), .ZN(n4186) );
  NAND4_X1 U2850 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .ZN(n4170)
         );
  NAND4_X1 U2851 ( .A1(n2676), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(n4347)
         );
  NAND4_X1 U2852 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n3508)
         );
  NAND4_X1 U2853 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n3892)
         );
  NAND4_X1 U2854 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n3893)
         );
  NAND4_X1 U2855 ( .A1(n2588), .A2(n2587), .A3(n2586), .A4(n2585), .ZN(n3894)
         );
  CLKBUF_X2 U2856 ( .A(U4043), .Z(n3901) );
  OAI21_X1 U2857 ( .B1(n2315), .B2(n3435), .A(n2292), .ZN(n3904) );
  NAND2_X1 U2858 ( .A1(n2315), .A2(n3435), .ZN(n2292) );
  XNOR2_X1 U2859 ( .A(n2313), .B(n2312), .ZN(n4336) );
  NAND2_X1 U2860 ( .A1(n4336), .A2(REG2_REG_3__SCAN_IN), .ZN(n4335) );
  OAI22_X1 U2861 ( .A1(n3933), .A2(n3459), .B1(n3458), .B2(n3457), .ZN(n4375)
         );
  NAND2_X1 U2862 ( .A1(n4386), .A2(REG2_REG_6__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U2863 ( .A1(n4383), .A2(n3461), .ZN(n4392) );
  NAND2_X1 U2864 ( .A1(n4407), .A2(n3443), .ZN(n4416) );
  NAND2_X1 U2865 ( .A1(n4416), .A2(n4417), .ZN(n4415) );
  INV_X1 U2866 ( .A(n2279), .ZN(n4420) );
  AND2_X1 U2867 ( .A1(n2279), .A2(n2246), .ZN(n4430) );
  XNOR2_X1 U2868 ( .A(n3447), .B(n2310), .ZN(n4445) );
  NAND2_X1 U2869 ( .A1(n4445), .A2(REG2_REG_12__SCAN_IN), .ZN(n4444) );
  INV_X1 U2870 ( .A(n2290), .ZN(n4438) );
  INV_X1 U2871 ( .A(n2406), .ZN(n3477) );
  XNOR2_X1 U2872 ( .A(n3944), .B(n4518), .ZN(n4449) );
  NOR2_X1 U2873 ( .A1(n4449), .A2(n4762), .ZN(n4448) );
  NAND2_X1 U2874 ( .A1(n4464), .A2(n3947), .ZN(n4476) );
  INV_X1 U2875 ( .A(n4450), .ZN(n4985) );
  OR2_X1 U2876 ( .A1(n2275), .A2(n3966), .ZN(n2274) );
  NAND2_X1 U2877 ( .A1(n2276), .A2(n4985), .ZN(n2275) );
  NAND2_X1 U2878 ( .A1(n3959), .A2(n3960), .ZN(n2276) );
  NAND2_X1 U2879 ( .A1(n2233), .A2(n3961), .ZN(n2277) );
  AOI21_X1 U2880 ( .B1(n3949), .B2(n3948), .A(n4975), .ZN(n3961) );
  AND2_X1 U2881 ( .A1(n3433), .A2(n3085), .ZN(n4980) );
  INV_X1 U2882 ( .A(n2286), .ZN(n2283) );
  AOI22_X1 U2883 ( .A1(n2231), .A2(n3948), .B1(n3965), .B2(n2266), .ZN(n2286)
         );
  AOI21_X1 U2884 ( .B1(n2318), .B2(n2226), .A(n2245), .ZN(n3998) );
  NAND2_X1 U2885 ( .A1(n2323), .A2(n2320), .ZN(n4012) );
  AND2_X1 U2886 ( .A1(n2321), .A2(n3817), .ZN(n2320) );
  AND2_X1 U2887 ( .A1(n2748), .A2(n2738), .ZN(n4059) );
  NAND2_X1 U2888 ( .A1(n2357), .A2(n2356), .ZN(n4103) );
  OR2_X1 U2889 ( .A1(n4121), .A2(n2712), .ZN(n2357) );
  NAND2_X1 U2890 ( .A1(n3414), .A2(n3551), .ZN(n4272) );
  AOI21_X1 U2891 ( .B1(n2645), .B2(n2644), .A(n2222), .ZN(n3518) );
  NAND2_X1 U2892 ( .A1(n2339), .A2(n2340), .ZN(n3517) );
  NAND2_X1 U2893 ( .A1(n2582), .A2(n2581), .ZN(n3277) );
  INV_X1 U2894 ( .A(n4182), .ZN(n4204) );
  OR2_X1 U2895 ( .A1(n3081), .A2(n3046), .ZN(n4124) );
  INV_X1 U2896 ( .A(n4504), .ZN(n4179) );
  INV_X1 U2897 ( .A(DATAI_0_), .ZN(n2307) );
  INV_X1 U2898 ( .A(n4124), .ZN(n4499) );
  AND2_X2 U2899 ( .A1(n3063), .A2(n3062), .ZN(n4595) );
  AND2_X1 U2900 ( .A1(n4197), .A2(n3693), .ZN(n4176) );
  AND2_X1 U2901 ( .A1(n2836), .A2(n2837), .ZN(n3078) );
  NAND2_X1 U2902 ( .A1(n3077), .A2(n3142), .ZN(n4509) );
  INV_X1 U2903 ( .A(n3048), .ZN(n4321) );
  AND2_X1 U2904 ( .A1(n3084), .A2(STATE_REG_SCAN_IN), .ZN(n4510) );
  INV_X1 U2905 ( .A(n3453), .ZN(n4526) );
  NAND2_X1 U2906 ( .A1(n2414), .A2(n2412), .ZN(n4331) );
  OR2_X1 U2907 ( .A1(n2438), .A2(n3722), .ZN(n2433) );
  AND2_X1 U2908 ( .A1(n2432), .A2(n3061), .ZN(n2431) );
  NAND2_X1 U2909 ( .A1(n4479), .A2(n2283), .ZN(n2282) );
  OR2_X1 U2910 ( .A1(n3949), .A2(n2284), .ZN(n2281) );
  OR2_X1 U2911 ( .A1(n4007), .A2(n4257), .ZN(n3066) );
  AND2_X1 U2912 ( .A1(n2860), .A2(n2859), .ZN(n2861) );
  OR2_X1 U2913 ( .A1(n4007), .A2(n4312), .ZN(n2860) );
  NAND2_X1 U2914 ( .A1(n2317), .A2(n2316), .ZN(U3351) );
  NAND2_X1 U2915 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2316) );
  AND2_X1 U2916 ( .A1(n2911), .A2(n2910), .ZN(n2221) );
  INV_X1 U2917 ( .A(n4337), .ZN(n2312) );
  NAND2_X1 U2918 ( .A1(n2490), .A2(n2479), .ZN(n2560) );
  XNOR2_X1 U2919 ( .A(n2878), .B(n3030), .ZN(n2881) );
  AND2_X1 U2920 ( .A1(n3550), .A2(n3511), .ZN(n2222) );
  INV_X1 U2921 ( .A(n2349), .ZN(n2348) );
  NAND2_X1 U2922 ( .A1(n2591), .A2(n2350), .ZN(n2349) );
  AND2_X1 U2923 ( .A1(n2340), .A2(n2255), .ZN(n2223) );
  AND2_X1 U2924 ( .A1(n2357), .A2(n2249), .ZN(n2224) );
  AND2_X1 U2925 ( .A1(n2328), .A2(n3995), .ZN(n2225) );
  INV_X1 U2926 ( .A(n3995), .ZN(n2326) );
  NAND2_X1 U2927 ( .A1(n2257), .A2(n2427), .ZN(n2640) );
  AND2_X1 U2928 ( .A1(n2225), .A2(n2329), .ZN(n2226) );
  AND2_X1 U2929 ( .A1(n2761), .A2(n2760), .ZN(n4037) );
  AND2_X1 U2930 ( .A1(n3886), .A2(n4017), .ZN(n2227) );
  AND2_X1 U2931 ( .A1(n2225), .A2(n2319), .ZN(n2228) );
  AND2_X1 U2932 ( .A1(n3040), .A2(n3039), .ZN(n4353) );
  INV_X1 U2933 ( .A(n4353), .ZN(n3722) );
  INV_X1 U2934 ( .A(n4147), .ZN(n4153) );
  AND2_X1 U2935 ( .A1(n2301), .A2(n4153), .ZN(n2229) );
  AND2_X1 U2936 ( .A1(n2303), .A2(n4053), .ZN(n2230) );
  NOR2_X1 U2937 ( .A1(n2266), .A2(n3965), .ZN(n2231) );
  NOR2_X1 U2938 ( .A1(n2869), .A2(n3902), .ZN(n2232) );
  OR2_X1 U2939 ( .A1(n3948), .A2(n3949), .ZN(n2233) );
  NAND3_X1 U2940 ( .A1(n2532), .A2(n2531), .A3(n2530), .ZN(n2889) );
  NOR2_X1 U2941 ( .A1(n4402), .A2(n3464), .ZN(n2234) );
  NAND4_X1 U2942 ( .A1(n2539), .A2(n2538), .A3(n2537), .A4(n2536), .ZN(n3899)
         );
  NAND2_X1 U2943 ( .A1(n2962), .A2(n2961), .ZN(n3644) );
  NAND4_X1 U2944 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n2867)
         );
  INV_X1 U2945 ( .A(n2535), .ZN(n2739) );
  NAND2_X1 U2946 ( .A1(n3666), .A2(n3667), .ZN(n3665) );
  AND3_X1 U2947 ( .A1(n2600), .A2(n2492), .A3(n2491), .ZN(n2235) );
  OR2_X1 U2948 ( .A1(n4526), .A2(n4890), .ZN(n2236) );
  NOR2_X1 U2949 ( .A1(n3896), .A2(n3224), .ZN(n2237) );
  NOR2_X1 U2950 ( .A1(n4448), .A2(n3945), .ZN(n2238) );
  OAI22_X1 U2951 ( .A1(n2887), .A2(n3125), .B1(n2219), .B2(n2879), .ZN(n2880)
         );
  OR2_X1 U2952 ( .A1(n3473), .A2(n2310), .ZN(n2239) );
  OR2_X1 U2953 ( .A1(n4526), .A2(n3438), .ZN(n2240) );
  AND2_X1 U2954 ( .A1(n4331), .A2(REG1_REG_2__SCAN_IN), .ZN(n2241) );
  INV_X1 U2955 ( .A(n2461), .ZN(n2460) );
  AND2_X1 U2956 ( .A1(n2498), .A2(n2359), .ZN(n2242) );
  AND2_X1 U2957 ( .A1(n3365), .A2(n3423), .ZN(n2243) );
  AND2_X1 U2958 ( .A1(n2784), .A2(n2509), .ZN(n2244) );
  OR2_X1 U2959 ( .A1(n2228), .A2(n2325), .ZN(n2245) );
  OAI21_X1 U2960 ( .B1(n3332), .B2(n3354), .A(n2485), .ZN(n2613) );
  INV_X1 U2961 ( .A(IR_REG_27__SCAN_IN), .ZN(n2509) );
  OR2_X1 U2962 ( .A1(n3470), .A2(n3469), .ZN(n2246) );
  AND2_X1 U2963 ( .A1(n4331), .A2(REG2_REG_2__SCAN_IN), .ZN(n2247) );
  INV_X1 U2964 ( .A(n2383), .ZN(n2382) );
  OAI21_X1 U2965 ( .B1(n3140), .B2(n2384), .A(n3751), .ZN(n2383) );
  AND2_X1 U2966 ( .A1(n2277), .A2(n2274), .ZN(n2248) );
  INV_X1 U2967 ( .A(IR_REG_26__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U2968 ( .A1(n4108), .A2(n3624), .ZN(n2249) );
  AND2_X1 U2969 ( .A1(n4113), .A2(n2230), .ZN(n2250) );
  INV_X1 U2970 ( .A(n3463), .ZN(n2404) );
  INV_X1 U2971 ( .A(n3224), .ZN(n3257) );
  AND2_X1 U2972 ( .A1(n2427), .A2(n2490), .ZN(n2611) );
  AOI21_X1 U2973 ( .B1(n4161), .B2(n2704), .A(n2703), .ZN(n4137) );
  AND2_X1 U2974 ( .A1(n2403), .A2(n3836), .ZN(n2251) );
  INV_X1 U2975 ( .A(IR_REG_24__SCAN_IN), .ZN(n2822) );
  INV_X1 U2976 ( .A(n3763), .ZN(n2394) );
  AND2_X1 U2977 ( .A1(n3619), .A2(n3620), .ZN(n2252) );
  INV_X1 U2978 ( .A(n3772), .ZN(n2392) );
  AND2_X1 U2979 ( .A1(n2251), .A2(n3985), .ZN(n2253) );
  INV_X1 U2980 ( .A(n2746), .ZN(n2319) );
  AND2_X1 U2981 ( .A1(n2804), .A2(n2803), .ZN(n3726) );
  INV_X1 U2982 ( .A(n3726), .ZN(n2374) );
  INV_X1 U2983 ( .A(IR_REG_10__SCAN_IN), .ZN(n2295) );
  OR2_X1 U2984 ( .A1(n4019), .A2(n3994), .ZN(n2254) );
  NAND2_X1 U2985 ( .A1(n3537), .A2(n3551), .ZN(n2255) );
  INV_X1 U2986 ( .A(IR_REG_28__SCAN_IN), .ZN(n2498) );
  INV_X1 U2987 ( .A(n2458), .ZN(n2457) );
  NAND2_X1 U2988 ( .A1(n3504), .A2(n3491), .ZN(n2458) );
  NOR2_X1 U2989 ( .A1(n3626), .A2(n4114), .ZN(n2256) );
  INV_X1 U2990 ( .A(n2747), .ZN(n2329) );
  AND2_X1 U2991 ( .A1(n2490), .A2(n2493), .ZN(n2257) );
  AND2_X1 U2992 ( .A1(n3985), .A2(n2402), .ZN(n2258) );
  OR2_X1 U2993 ( .A1(n3886), .A2(n4017), .ZN(n2259) );
  NOR2_X1 U2994 ( .A1(n3601), .A2(n3600), .ZN(n2260) );
  AND2_X1 U2995 ( .A1(n2642), .A2(n2478), .ZN(n2702) );
  NOR2_X1 U2996 ( .A1(n3816), .A2(n2319), .ZN(n2261) );
  INV_X1 U2997 ( .A(n3474), .ZN(n2310) );
  NAND2_X1 U2998 ( .A1(n2332), .A2(n2333), .ZN(n3222) );
  INV_X1 U2999 ( .A(n3759), .ZN(n2368) );
  NAND2_X1 U3000 ( .A1(n2471), .A2(n2470), .ZN(n3294) );
  NAND2_X1 U3001 ( .A1(n2827), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  NOR2_X1 U3002 ( .A1(n3262), .A2(n2221), .ZN(n2262) );
  INV_X1 U3003 ( .A(n3668), .ZN(n2448) );
  INV_X1 U3004 ( .A(n3850), .ZN(n2377) );
  AND2_X1 U3005 ( .A1(n3472), .A2(REG1_REG_11__SCAN_IN), .ZN(n2263) );
  INV_X1 U3006 ( .A(n4053), .ZN(n4058) );
  AND2_X1 U3007 ( .A1(n3530), .A2(n3749), .ZN(n3824) );
  INV_X1 U3008 ( .A(n3824), .ZN(n2341) );
  OR2_X1 U3009 ( .A1(n4520), .A2(n4917), .ZN(n2264) );
  INV_X1 U3010 ( .A(IR_REG_11__SCAN_IN), .ZN(n2294) );
  AND2_X1 U3011 ( .A1(n2229), .A2(n3624), .ZN(n2265) );
  AND2_X1 U3012 ( .A1(n3967), .A2(REG1_REG_18__SCAN_IN), .ZN(n2266) );
  OR2_X1 U3013 ( .A1(n4367), .A2(n4322), .ZN(n4975) );
  INV_X1 U3014 ( .A(n4017), .ZN(n4023) );
  OR2_X1 U3015 ( .A1(n3958), .A2(REG2_REG_17__SCAN_IN), .ZN(n2268) );
  OR2_X1 U3016 ( .A1(n3958), .A2(REG1_REG_17__SCAN_IN), .ZN(n2269) );
  INV_X1 U3017 ( .A(n3316), .ZN(n2467) );
  INV_X1 U3018 ( .A(n4040), .ZN(n4033) );
  AND2_X1 U3019 ( .A1(n4479), .A2(n2231), .ZN(n2270) );
  INV_X1 U3020 ( .A(IR_REG_0__SCAN_IN), .ZN(n2308) );
  INV_X1 U3021 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2415) );
  INV_X1 U3022 ( .A(DATAI_1_), .ZN(n2337) );
  AND2_X1 U3023 ( .A1(n3967), .A2(REG2_REG_18__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U3024 ( .A1(n3436), .A2(n4330), .ZN(n2272) );
  XNOR2_X1 U3025 ( .A(n3436), .B(n4330), .ZN(n3934) );
  MUX2_X1 U3026 ( .A(n4773), .B(REG2_REG_2__SCAN_IN), .S(n4331), .Z(n3920) );
  NOR2_X2 U3027 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2533)
         );
  NAND4_X1 U3028 ( .A1(n2281), .A2(n2280), .A3(n3975), .A4(n2282), .ZN(U3259)
         );
  NAND2_X1 U3029 ( .A1(n3949), .A2(n2270), .ZN(n2280) );
  NOR2_X1 U3030 ( .A1(n4403), .A2(n4404), .ZN(n4402) );
  XNOR2_X1 U3031 ( .A(n3462), .B(n2404), .ZN(n4403) );
  XNOR2_X2 U3032 ( .A(n2514), .B(IR_REG_1__SCAN_IN), .ZN(n2315) );
  AND2_X1 U3033 ( .A1(n2425), .A2(n2490), .ZN(n2305) );
  NAND3_X1 U3034 ( .A1(n2480), .A2(n2360), .A3(n2304), .ZN(n2511) );
  NAND2_X1 U3035 ( .A1(n2642), .A2(n2480), .ZN(n2825) );
  AND2_X2 U3036 ( .A1(n2305), .A2(n2360), .ZN(n2642) );
  INV_X1 U3037 ( .A(n2511), .ZN(n2833) );
  MUX2_X1 U3038 ( .A(n2308), .B(n2307), .S(n2541), .Z(n3160) );
  INV_X1 U3039 ( .A(n2315), .ZN(n2338) );
  NAND2_X1 U3040 ( .A1(n2315), .A2(REG2_REG_1__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U3041 ( .A1(n2315), .A2(STATE_REG_SCAN_IN), .ZN(n2317) );
  MUX2_X1 U3042 ( .A(REG1_REG_1__SCAN_IN), .B(n2415), .S(n2315), .Z(n3903) );
  NAND2_X1 U3043 ( .A1(n4456), .A2(n2315), .ZN(n3905) );
  INV_X1 U3044 ( .A(n4047), .ZN(n2318) );
  OAI21_X1 U3045 ( .B1(n4047), .B2(n2747), .A(n2746), .ZN(n4029) );
  NAND2_X1 U3046 ( .A1(n4047), .A2(n2261), .ZN(n2323) );
  NAND2_X1 U3047 ( .A1(n2332), .A2(n2330), .ZN(n2570) );
  NAND2_X1 U3048 ( .A1(n2554), .A2(n2553), .ZN(n3139) );
  INV_X1 U3049 ( .A(n2553), .ZN(n2335) );
  MUX2_X1 U3050 ( .A(n2338), .B(n2337), .S(n2541), .Z(n2879) );
  NAND2_X1 U3051 ( .A1(n2645), .A2(n2342), .ZN(n2339) );
  INV_X1 U3052 ( .A(n2661), .ZN(n3538) );
  NAND2_X1 U3053 ( .A1(n2582), .A2(n2346), .ZN(n2344) );
  NAND2_X1 U3054 ( .A1(n2344), .A2(n2345), .ZN(n3359) );
  NAND2_X1 U3055 ( .A1(n4121), .A2(n2356), .ZN(n2354) );
  NAND2_X1 U3056 ( .A1(n2354), .A2(n2355), .ZN(n4084) );
  NAND3_X1 U3057 ( .A1(n3792), .A2(n4485), .A3(n2524), .ZN(n3195) );
  NAND2_X1 U3058 ( .A1(n3573), .A2(n3826), .ZN(n3572) );
  NAND2_X1 U3059 ( .A1(n4193), .A2(n2696), .ZN(n4161) );
  NAND2_X1 U3060 ( .A1(n2361), .A2(n2365), .ZN(n2795) );
  NAND2_X1 U3061 ( .A1(n2794), .A2(n2362), .ZN(n2361) );
  NAND2_X1 U3062 ( .A1(n4139), .A2(n2372), .ZN(n2370) );
  NAND2_X1 U3063 ( .A1(n3125), .A2(n4500), .ZN(n3730) );
  AND4_X2 U3064 ( .A1(n2518), .A2(n2515), .A3(n2517), .A4(n2516), .ZN(n3125)
         );
  OAI21_X1 U3065 ( .B1(n3168), .B2(n2383), .A(n2378), .ZN(n2791) );
  OAI21_X1 U3066 ( .B1(n3238), .B2(n2398), .A(n2395), .ZN(n3307) );
  OAI21_X1 U3067 ( .B1(n3238), .B2(n2793), .A(n3754), .ZN(n3272) );
  NAND2_X1 U3068 ( .A1(n2793), .A2(n3754), .ZN(n2400) );
  NAND2_X1 U3069 ( .A1(n2809), .A2(n2251), .ZN(n4016) );
  OAI21_X1 U3070 ( .B1(n2408), .B2(n4449), .A(n2407), .ZN(n4976) );
  INV_X1 U3071 ( .A(n2533), .ZN(n2413) );
  NAND3_X1 U3072 ( .A1(n2412), .A2(n2414), .A3(n4584), .ZN(n2410) );
  NAND2_X1 U3073 ( .A1(n2962), .A2(n2419), .ZN(n2418) );
  OAI211_X1 U3074 ( .C1(n3592), .C2(n2433), .A(n2428), .B(n2431), .ZN(U3217)
         );
  NAND2_X1 U3075 ( .A1(n3592), .A2(n2429), .ZN(n2428) );
  INV_X1 U3076 ( .A(n3034), .ZN(n2439) );
  NAND2_X1 U3077 ( .A1(n2979), .A2(n2442), .ZN(n2441) );
  NAND2_X1 U3078 ( .A1(n2441), .A2(n2444), .ZN(n3677) );
  NAND2_X1 U3079 ( .A1(n2462), .A2(n2940), .ZN(n2461) );
  NAND2_X1 U3080 ( .A1(n3490), .A2(n3491), .ZN(n2462) );
  NAND2_X1 U3081 ( .A1(n3262), .A2(n2472), .ZN(n2471) );
  INV_X1 U3082 ( .A(n2499), .ZN(n2786) );
  NOR2_X2 U3083 ( .A1(n2825), .A2(n2474), .ZN(n2499) );
  XNOR2_X1 U3084 ( .A(n3996), .B(n2326), .ZN(n4004) );
  OR2_X1 U3085 ( .A1(n2535), .A2(n2525), .ZN(n2532) );
  NAND2_X1 U3086 ( .A1(n2839), .A2(n2828), .ZN(n2829) );
  OAI21_X1 U3087 ( .B1(n3385), .B2(n2931), .A(n3387), .ZN(n2932) );
  NAND2_X1 U3088 ( .A1(n2873), .A2(n2872), .ZN(n2874) );
  OR2_X1 U3089 ( .A1(n3053), .A2(n3052), .ZN(n2475) );
  NOR2_X1 U3090 ( .A1(n3060), .A2(n4358), .ZN(n2476) );
  INV_X1 U3091 ( .A(n3979), .ZN(n4200) );
  AND2_X2 U3092 ( .A1(n3144), .A2(n3063), .ZN(n4580) );
  AND2_X1 U3093 ( .A1(n2915), .A2(n2914), .ZN(n2477) );
  NOR2_X1 U3094 ( .A1(IR_REG_14__SCAN_IN), .A2(n2693), .ZN(n2478) );
  INV_X1 U3095 ( .A(n3713), .ZN(n3560) );
  NAND4_X1 U3096 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n3713)
         );
  AND4_X1 U3097 ( .A1(n2497), .A2(n2481), .A3(n2496), .A4(n2495), .ZN(n2480)
         );
  AND4_X1 U3098 ( .A1(n4822), .A2(n4726), .A3(n2776), .A4(n2822), .ZN(n2481)
         );
  AND2_X1 U3099 ( .A1(n2893), .A2(n2892), .ZN(n2483) );
  OR2_X1 U3100 ( .A1(n3455), .A2(n2312), .ZN(n2484) );
  NAND2_X1 U3101 ( .A1(n3892), .A2(n3328), .ZN(n2485) );
  INV_X1 U3102 ( .A(n3575), .ZN(n4345) );
  INV_X1 U3103 ( .A(IR_REG_25__SCAN_IN), .ZN(n2494) );
  NOR2_X1 U3104 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2495)
         );
  NOR2_X1 U3105 ( .A1(n3004), .A2(n3006), .ZN(n3002) );
  AND2_X1 U3106 ( .A1(n3805), .A2(n4065), .ZN(n3852) );
  AND2_X1 U3107 ( .A1(n4162), .A2(n2800), .ZN(n3849) );
  INV_X1 U3108 ( .A(IR_REG_14__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U3109 ( .A1(n2526), .A2(REG2_REG_2__SCAN_IN), .ZN(n2529) );
  OR2_X1 U3110 ( .A1(n4074), .A2(n4053), .ZN(n2746) );
  OR2_X1 U3111 ( .A1(n3409), .A2(n3496), .ZN(n2631) );
  INV_X1 U3112 ( .A(IR_REG_18__SCAN_IN), .ZN(n4727) );
  INV_X1 U3113 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2571) );
  INV_X1 U3114 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2593) );
  INV_X1 U3115 ( .A(n3468), .ZN(n3469) );
  AND2_X1 U3116 ( .A1(n3982), .A2(n2763), .ZN(n4005) );
  NAND2_X1 U3117 ( .A1(n2782), .A2(n2816), .ZN(n2862) );
  INV_X1 U3118 ( .A(n3650), .ZN(n3563) );
  INV_X1 U3119 ( .A(n3523), .ZN(n3551) );
  INV_X1 U3120 ( .A(n3328), .ZN(n3423) );
  INV_X1 U3121 ( .A(n3309), .ZN(n3354) );
  OR2_X1 U3122 ( .A1(n2698), .A2(n2697), .ZN(n2708) );
  NOR2_X1 U3123 ( .A1(n2651), .A2(n2486), .ZN(n2662) );
  AND2_X1 U3124 ( .A1(n2713), .A2(REG3_REG_22__SCAN_IN), .ZN(n2717) );
  OR2_X1 U3125 ( .A1(n2535), .A2(n2519), .ZN(n2523) );
  INV_X1 U3126 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4918) );
  INV_X1 U3127 ( .A(n3624), .ZN(n4131) );
  NAND2_X1 U3128 ( .A1(n3713), .A2(n3575), .ZN(n2671) );
  INV_X1 U3129 ( .A(n3888), .ZN(n4344) );
  INV_X1 U3130 ( .A(n4191), .ZN(n4493) );
  INV_X1 U3131 ( .A(n4486), .ZN(n4107) );
  AND2_X1 U3132 ( .A1(n3806), .A2(DATAI_20_), .ZN(n4147) );
  INV_X1 U3133 ( .A(n3894), .ZN(n3312) );
  NAND2_X1 U3134 ( .A1(n2659), .A2(IR_REG_31__SCAN_IN), .ZN(n2679) );
  INV_X1 U3135 ( .A(n3704), .ZN(n4348) );
  OR2_X1 U3136 ( .A1(n2727), .A2(n3660), .ZN(n2737) );
  INV_X1 U3137 ( .A(n3599), .ZN(n3678) );
  NOR2_X1 U3138 ( .A1(n2748), .A2(n3703), .ZN(n2754) );
  INV_X1 U3139 ( .A(n4095), .ZN(n3096) );
  INV_X1 U3140 ( .A(n4975), .ZN(n4479) );
  NAND2_X1 U3141 ( .A1(n3572), .A2(n2671), .ZN(n3557) );
  NAND2_X1 U3142 ( .A1(n3867), .A2(n2810), .ZN(n4191) );
  AOI21_X1 U3143 ( .B1(n2853), .B2(n4899), .A(n3078), .ZN(n3062) );
  INV_X1 U3144 ( .A(n4569), .ZN(n4572) );
  INV_X1 U3145 ( .A(n3407), .ZN(n3511) );
  INV_X1 U3146 ( .A(n4560), .ZN(n4577) );
  INV_X1 U3147 ( .A(IR_REG_30__SCAN_IN), .ZN(n3588) );
  AND2_X1 U31480 ( .A1(n2589), .A2(n2580), .ZN(n4524) );
  NOR2_X1 U31490 ( .A1(n2475), .A2(n2476), .ZN(n3061) );
  OR2_X1 U3150 ( .A1(n2749), .A2(n2754), .ZN(n4041) );
  INV_X1 U3151 ( .A(n4037), .ZN(n3886) );
  NAND2_X1 U3152 ( .A1(n2745), .A2(n2744), .ZN(n4034) );
  NAND4_X1 U3153 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .ZN(n3889)
         );
  INV_X1 U3154 ( .A(n4524), .ZN(n4401) );
  OR2_X1 U3155 ( .A1(n4367), .A2(n4321), .ZN(n4989) );
  OR2_X1 U3156 ( .A1(n4507), .A2(n3147), .ZN(n4182) );
  AND2_X1 U3157 ( .A1(n3145), .A2(n4124), .ZN(n4507) );
  INV_X1 U3158 ( .A(n4595), .ZN(n4593) );
  INV_X1 U3159 ( .A(n4359), .ZN(n4287) );
  INV_X1 U3160 ( .A(n4580), .ZN(n4578) );
  INV_X1 U3161 ( .A(n4509), .ZN(n4508) );
  INV_X1 U3162 ( .A(n4319), .ZN(n4320) );
  NAND2_X1 U3163 ( .A1(n2583), .A2(REG3_REG_8__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U3164 ( .A1(n2622), .A2(REG3_REG_12__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3165 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2486) );
  AND2_X1 U3166 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2487) );
  INV_X1 U3167 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2697) );
  XNOR2_X1 U3168 ( .A(n2708), .B(REG3_REG_20__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U3169 ( .A1(n2533), .A2(n2488), .ZN(n2540) );
  NAND2_X1 U3170 ( .A1(n2499), .A2(n4871), .ZN(n2501) );
  XNOR2_X2 U3171 ( .A(n2500), .B(n3588), .ZN(n4319) );
  NAND2_X1 U3172 ( .A1(n2786), .A2(IR_REG_31__SCAN_IN), .ZN(n2502) );
  NAND2_X2 U3173 ( .A1(n2501), .A2(n2503), .ZN(n3074) );
  NAND2_X1 U3174 ( .A1(n4155), .A2(n2739), .ZN(n2508) );
  INV_X1 U3175 ( .A(n3074), .ZN(n2504) );
  NAND2_X2 U3176 ( .A1(n4319), .A2(n2504), .ZN(n2719) );
  NAND2_X1 U3177 ( .A1(n2218), .A2(REG1_REG_20__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3178 ( .A1(n3086), .A2(REG2_REG_20__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3179 ( .A1(n2740), .A2(REG0_REG_20__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3180 ( .A1(n2511), .A2(n2510), .ZN(n3449) );
  INV_X1 U3181 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U3182 ( .A1(n2513), .A2(REG1_REG_1__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U3183 ( .A1(n2527), .A2(REG0_REG_1__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3184 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2514)
         );
  NAND4_X1 U3185 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n2875)
         );
  INV_X1 U3186 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3187 ( .A1(n2513), .A2(REG1_REG_0__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3188 ( .A1(n2527), .A2(REG0_REG_0__SCAN_IN), .ZN(n2520) );
  INV_X1 U3189 ( .A(n3125), .ZN(n3900) );
  NAND2_X1 U3190 ( .A1(n3900), .A2(n4500), .ZN(n2524) );
  INV_X1 U3191 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U3192 ( .A1(n2513), .A2(REG1_REG_2__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U3193 ( .A1(n2527), .A2(REG0_REG_2__SCAN_IN), .ZN(n2528) );
  AND2_X1 U3194 ( .A1(n2529), .A2(n2528), .ZN(n2530) );
  MUX2_X1 U3195 ( .A(n4331), .B(DATAI_2_), .S(n2541), .Z(n2888) );
  INV_X1 U3196 ( .A(n2888), .ZN(n3192) );
  NAND2_X1 U3197 ( .A1(n2889), .A2(n3192), .ZN(n3733) );
  NAND2_X1 U3198 ( .A1(n4490), .A2(n3192), .ZN(n2534) );
  NAND2_X1 U3199 ( .A1(n3195), .A2(n2534), .ZN(n3205) );
  NAND2_X1 U3200 ( .A1(n2220), .A2(REG2_REG_3__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U3201 ( .A1(n2527), .A2(REG0_REG_3__SCAN_IN), .ZN(n2538) );
  INV_X2 U3202 ( .A(n2535), .ZN(n2764) );
  INV_X1 U3203 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3204 ( .A1(n2764), .A2(n3136), .ZN(n2537) );
  NAND2_X1 U3205 ( .A1(n2513), .A2(REG1_REG_3__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U3206 ( .A1(n2540), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  XNOR2_X1 U3207 ( .A(n2550), .B(IR_REG_3__SCAN_IN), .ZN(n4337) );
  MUX2_X1 U3208 ( .A(n4337), .B(DATAI_3_), .S(n2541), .Z(n3735) );
  NOR2_X1 U3209 ( .A1(n3899), .A2(n3735), .ZN(n2543) );
  NAND2_X1 U32100 ( .A1(n3899), .A2(n3735), .ZN(n2542) );
  OAI21_X2 U32110 ( .B1(n3205), .B2(n2543), .A(n2542), .ZN(n3167) );
  NAND2_X1 U32120 ( .A1(n2218), .A2(REG1_REG_4__SCAN_IN), .ZN(n2548) );
  INV_X1 U32130 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2544) );
  XNOR2_X1 U32140 ( .A(n2544), .B(REG3_REG_3__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U32150 ( .A1(n2764), .A2(n3186), .ZN(n2547) );
  NAND2_X1 U32160 ( .A1(n2527), .A2(REG0_REG_4__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32170 ( .A1(n2220), .A2(REG2_REG_4__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32180 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  NAND2_X1 U32190 ( .A1(n2551), .A2(IR_REG_31__SCAN_IN), .ZN(n2552) );
  XNOR2_X1 U32200 ( .A(n2552), .B(IR_REG_4__SCAN_IN), .ZN(n4330) );
  MUX2_X1 U32210 ( .A(n4330), .B(DATAI_4_), .S(n3806), .Z(n3169) );
  NAND2_X1 U32220 ( .A1(n3152), .A2(n3169), .ZN(n3737) );
  INV_X1 U32230 ( .A(n3169), .ZN(n3180) );
  NAND2_X1 U32240 ( .A1(n3898), .A2(n3180), .ZN(n3740) );
  NAND2_X1 U32250 ( .A1(n3737), .A2(n3740), .ZN(n3823) );
  NAND2_X1 U32260 ( .A1(n3167), .A2(n3823), .ZN(n2554) );
  NAND2_X1 U32270 ( .A1(n3898), .A2(n3169), .ZN(n2553) );
  NAND2_X1 U32280 ( .A1(n2218), .A2(REG1_REG_5__SCAN_IN), .ZN(n2559) );
  AOI21_X1 U32290 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2555) );
  NOR2_X1 U32300 ( .A1(n2555), .A2(n2563), .ZN(n3154) );
  NAND2_X1 U32310 ( .A1(n2764), .A2(n3154), .ZN(n2558) );
  NAND2_X1 U32320 ( .A1(n2740), .A2(REG0_REG_5__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U32330 ( .A1(n3086), .A2(REG2_REG_5__SCAN_IN), .ZN(n2556) );
  NAND4_X1 U32340 ( .A1(n2559), .A2(n2558), .A3(n2557), .A4(n2556), .ZN(n3897)
         );
  NAND2_X1 U32350 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2561) );
  XNOR2_X1 U32360 ( .A(n2561), .B(IR_REG_5__SCAN_IN), .ZN(n3453) );
  MUX2_X1 U32370 ( .A(n3453), .B(DATAI_5_), .S(n3806), .Z(n3153) );
  AND2_X1 U32380 ( .A1(n3897), .A2(n3153), .ZN(n2562) );
  NAND2_X1 U32390 ( .A1(n2218), .A2(REG1_REG_6__SCAN_IN), .ZN(n2567) );
  OAI21_X1 U32400 ( .B1(n2563), .B2(REG3_REG_6__SCAN_IN), .A(n2572), .ZN(n3232) );
  INV_X1 U32410 ( .A(n3232), .ZN(n3259) );
  NAND2_X1 U32420 ( .A1(n2764), .A2(n3259), .ZN(n2566) );
  NAND2_X1 U32430 ( .A1(n2527), .A2(REG0_REG_6__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U32440 ( .A1(n3086), .A2(REG2_REG_6__SCAN_IN), .ZN(n2564) );
  NAND4_X1 U32450 ( .A1(n2567), .A2(n2566), .A3(n2565), .A4(n2564), .ZN(n3896)
         );
  NOR2_X1 U32460 ( .A1(n2560), .A2(IR_REG_5__SCAN_IN), .ZN(n2602) );
  OR2_X1 U32470 ( .A1(n2602), .A2(n2784), .ZN(n2568) );
  XNOR2_X1 U32480 ( .A(n2568), .B(IR_REG_6__SCAN_IN), .ZN(n4329) );
  MUX2_X1 U32490 ( .A(n4329), .B(DATAI_6_), .S(n3806), .Z(n3224) );
  NAND2_X1 U32500 ( .A1(n3896), .A2(n3224), .ZN(n2569) );
  NAND2_X1 U32510 ( .A1(n2570), .A2(n2569), .ZN(n3242) );
  AOI22_X1 U32520 ( .A1(n2218), .A2(REG1_REG_7__SCAN_IN), .B1(n2740), .B2(
        REG0_REG_7__SCAN_IN), .ZN(n2575) );
  AND2_X1 U32530 ( .A1(n2572), .A2(n2571), .ZN(n2573) );
  NOR2_X1 U32540 ( .A1(n2583), .A2(n2573), .ZN(n3300) );
  AOI22_X1 U32550 ( .A1(n2739), .A2(n3300), .B1(n2220), .B2(
        REG2_REG_7__SCAN_IN), .ZN(n2574) );
  INV_X1 U32560 ( .A(IR_REG_6__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U32570 ( .A1(n2602), .A2(n2576), .ZN(n2577) );
  NAND2_X1 U32580 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32590 ( .A1(n2579), .A2(n2578), .ZN(n2589) );
  OR2_X1 U32600 ( .A1(n2579), .A2(n2578), .ZN(n2580) );
  MUX2_X1 U32610 ( .A(n4524), .B(DATAI_7_), .S(n3806), .Z(n3245) );
  NAND2_X1 U32620 ( .A1(n3276), .A2(n3245), .ZN(n2792) );
  NAND2_X1 U32630 ( .A1(n3895), .A2(n3298), .ZN(n3754) );
  NAND2_X1 U32640 ( .A1(n2792), .A2(n3754), .ZN(n3790) );
  NAND2_X1 U32650 ( .A1(n3242), .A2(n3790), .ZN(n2582) );
  NAND2_X1 U32660 ( .A1(n3895), .A2(n3245), .ZN(n2581) );
  NAND2_X1 U32670 ( .A1(n2218), .A2(REG1_REG_8__SCAN_IN), .ZN(n2588) );
  OR2_X1 U32680 ( .A1(n2583), .A2(REG3_REG_8__SCAN_IN), .ZN(n2584) );
  AND2_X1 U32690 ( .A1(n2594), .A2(n2584), .ZN(n3324) );
  NAND2_X1 U32700 ( .A1(n2739), .A2(n3324), .ZN(n2587) );
  NAND2_X1 U32710 ( .A1(n2527), .A2(REG0_REG_8__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32720 ( .A1(n2220), .A2(REG2_REG_8__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U32730 ( .A1(n2589), .A2(IR_REG_31__SCAN_IN), .ZN(n2590) );
  XNOR2_X1 U32740 ( .A(n2590), .B(IR_REG_8__SCAN_IN), .ZN(n3463) );
  MUX2_X1 U32750 ( .A(n3463), .B(DATAI_8_), .S(n3806), .Z(n3280) );
  AND2_X1 U32760 ( .A1(n3894), .A2(n3280), .ZN(n2592) );
  INV_X1 U32770 ( .A(n3280), .ZN(n3322) );
  NAND2_X1 U32780 ( .A1(n3312), .A2(n3322), .ZN(n2591) );
  NAND2_X1 U32790 ( .A1(n2218), .A2(REG1_REG_9__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U32800 ( .A1(n2594), .A2(n2593), .ZN(n2595) );
  AND2_X1 U32810 ( .A1(n2605), .A2(n2595), .ZN(n3356) );
  NAND2_X1 U32820 ( .A1(n2764), .A2(n3356), .ZN(n2598) );
  NAND2_X1 U32830 ( .A1(n2527), .A2(REG0_REG_9__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U32840 ( .A1(n3086), .A2(REG2_REG_9__SCAN_IN), .ZN(n2596) );
  NAND3_X1 U32850 ( .A1(n2602), .A2(n2601), .A3(n2600), .ZN(n2603) );
  NAND2_X1 U32860 ( .A1(n2603), .A2(IR_REG_31__SCAN_IN), .ZN(n2604) );
  XNOR2_X1 U32870 ( .A(n2604), .B(IR_REG_9__SCAN_IN), .ZN(n3466) );
  MUX2_X1 U32880 ( .A(n3466), .B(DATAI_9_), .S(n3806), .Z(n3309) );
  NOR2_X1 U32890 ( .A1(n3893), .A2(n3309), .ZN(n3333) );
  NAND2_X1 U32900 ( .A1(n2218), .A2(REG1_REG_10__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U32910 ( .A1(n2605), .A2(n3420), .ZN(n2606) );
  AND2_X1 U32920 ( .A1(n2614), .A2(n2606), .ZN(n3430) );
  NAND2_X1 U32930 ( .A1(n2764), .A2(n3430), .ZN(n2609) );
  NAND2_X1 U32940 ( .A1(n2740), .A2(REG0_REG_10__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U32950 ( .A1(n3086), .A2(REG2_REG_10__SCAN_IN), .ZN(n2607) );
  OR2_X1 U32960 ( .A1(n2611), .A2(n2784), .ZN(n2612) );
  XNOR2_X1 U32970 ( .A(n2612), .B(IR_REG_10__SCAN_IN), .ZN(n3468) );
  MUX2_X1 U32980 ( .A(n3468), .B(DATAI_10_), .S(n3806), .Z(n3328) );
  NAND2_X1 U32990 ( .A1(n2218), .A2(REG1_REG_11__SCAN_IN), .ZN(n2619) );
  AND2_X1 U33000 ( .A1(n2614), .A2(n4918), .ZN(n2615) );
  NOR2_X1 U33010 ( .A1(n2622), .A2(n2615), .ZN(n3393) );
  NAND2_X1 U33020 ( .A1(n2739), .A2(n3393), .ZN(n2618) );
  NAND2_X1 U33030 ( .A1(n2740), .A2(REG0_REG_11__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33040 ( .A1(n3086), .A2(REG2_REG_11__SCAN_IN), .ZN(n2616) );
  NAND4_X1 U33050 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n3891)
         );
  NAND2_X1 U33060 ( .A1(n2611), .A2(n2295), .ZN(n2620) );
  NAND2_X1 U33070 ( .A1(n2620), .A2(IR_REG_31__SCAN_IN), .ZN(n2628) );
  XNOR2_X1 U33080 ( .A(n2628), .B(IR_REG_11__SCAN_IN), .ZN(n3472) );
  MUX2_X1 U33090 ( .A(n3472), .B(DATAI_11_), .S(n3806), .Z(n3362) );
  NAND2_X1 U33100 ( .A1(n3497), .A2(n3362), .ZN(n3771) );
  NAND2_X1 U33110 ( .A1(n3891), .A2(n3391), .ZN(n3766) );
  NAND2_X1 U33120 ( .A1(n3771), .A2(n3766), .ZN(n3799) );
  AOI21_X2 U33130 ( .B1(n3359), .B2(n3799), .A(n2621), .ZN(n3381) );
  INV_X1 U33140 ( .A(n3381), .ZN(n2633) );
  NAND2_X1 U33150 ( .A1(n2218), .A2(REG1_REG_12__SCAN_IN), .ZN(n2627) );
  OR2_X1 U33160 ( .A1(n2622), .A2(REG3_REG_12__SCAN_IN), .ZN(n2623) );
  AND2_X1 U33170 ( .A1(n2623), .A2(n2634), .ZN(n3378) );
  NAND2_X1 U33180 ( .A1(n2739), .A2(n3378), .ZN(n2626) );
  NAND2_X1 U33190 ( .A1(n2527), .A2(REG0_REG_12__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33200 ( .A1(n3086), .A2(REG2_REG_12__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U33210 ( .A1(n2628), .A2(n2294), .ZN(n2629) );
  NAND2_X1 U33220 ( .A1(n2629), .A2(IR_REG_31__SCAN_IN), .ZN(n2630) );
  XNOR2_X1 U33230 ( .A(n2630), .B(IR_REG_12__SCAN_IN), .ZN(n3474) );
  MUX2_X1 U33240 ( .A(n3474), .B(DATAI_12_), .S(n3806), .Z(n3377) );
  INV_X1 U33250 ( .A(n3508), .ZN(n3409) );
  INV_X1 U33260 ( .A(n3377), .ZN(n3496) );
  OAI21_X2 U33270 ( .B1(n2633), .B2(n2632), .A(n2631), .ZN(n3405) );
  INV_X1 U33280 ( .A(n3405), .ZN(n2645) );
  NAND2_X1 U33290 ( .A1(n2218), .A2(REG1_REG_13__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U33300 ( .A1(n2634), .A2(n4718), .ZN(n2635) );
  AND2_X1 U33310 ( .A1(n2651), .A2(n2635), .ZN(n3513) );
  NAND2_X1 U33320 ( .A1(n2764), .A2(n3513), .ZN(n2638) );
  NAND2_X1 U33330 ( .A1(n2527), .A2(REG0_REG_13__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U33340 ( .A1(n3086), .A2(REG2_REG_13__SCAN_IN), .ZN(n2636) );
  NAND4_X1 U33350 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n3890)
         );
  NAND2_X1 U33360 ( .A1(n2640), .A2(IR_REG_31__SCAN_IN), .ZN(n2641) );
  MUX2_X1 U33370 ( .A(IR_REG_31__SCAN_IN), .B(n2641), .S(IR_REG_13__SCAN_IN), 
        .Z(n2643) );
  INV_X1 U33380 ( .A(n2642), .ZN(n2658) );
  AND2_X1 U33390 ( .A1(n2643), .A2(n2658), .ZN(n4328) );
  MUX2_X1 U33400 ( .A(n4328), .B(DATAI_13_), .S(n3806), .Z(n3407) );
  NAND2_X1 U33410 ( .A1(n2218), .A2(REG1_REG_14__SCAN_IN), .ZN(n2649) );
  XNOR2_X1 U33420 ( .A(n2651), .B(REG3_REG_14__SCAN_IN), .ZN(n3544) );
  NAND2_X1 U33430 ( .A1(n2764), .A2(n3544), .ZN(n2648) );
  NAND2_X1 U33440 ( .A1(n2527), .A2(REG0_REG_14__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U33450 ( .A1(n2220), .A2(REG2_REG_14__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U33460 ( .A1(n2658), .A2(IR_REG_31__SCAN_IN), .ZN(n2650) );
  XNOR2_X1 U33470 ( .A(n2650), .B(IR_REG_14__SCAN_IN), .ZN(n4455) );
  MUX2_X1 U33480 ( .A(n4455), .B(DATAI_14_), .S(n3806), .Z(n3523) );
  NAND2_X1 U33490 ( .A1(n3537), .A2(n3523), .ZN(n3530) );
  NAND2_X1 U33500 ( .A1(n3889), .A2(n3551), .ZN(n3749) );
  NAND2_X1 U33510 ( .A1(n2218), .A2(REG1_REG_15__SCAN_IN), .ZN(n2657) );
  INV_X1 U33520 ( .A(n2651), .ZN(n2652) );
  AOI21_X1 U3353 ( .B1(n2652), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2653) );
  NOR2_X1 U33540 ( .A1(n2653), .A2(n2662), .ZN(n3719) );
  NAND2_X1 U3355 ( .A1(n2739), .A2(n3719), .ZN(n2656) );
  NAND2_X1 U3356 ( .A1(n2527), .A2(REG0_REG_15__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3357 ( .A1(n3086), .A2(REG2_REG_15__SCAN_IN), .ZN(n2654) );
  NAND4_X1 U3358 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n3888)
         );
  OR2_X1 U3359 ( .A1(n2658), .A2(IR_REG_14__SCAN_IN), .ZN(n2659) );
  XNOR2_X1 U3360 ( .A(n2679), .B(IR_REG_15__SCAN_IN), .ZN(n4516) );
  MUX2_X1 U3361 ( .A(n4516), .B(DATAI_15_), .S(n3806), .Z(n3534) );
  OAI22_X2 U3362 ( .A1(n2661), .A2(n2660), .B1(n4344), .B2(n3717), .ZN(n3573)
         );
  NOR2_X1 U3363 ( .A1(n2662), .A2(REG3_REG_16__SCAN_IN), .ZN(n2663) );
  OR2_X1 U3364 ( .A1(n2683), .A2(n2663), .ZN(n4357) );
  INV_X1 U3365 ( .A(n4357), .ZN(n3574) );
  NAND2_X1 U3366 ( .A1(n2739), .A2(n3574), .ZN(n2667) );
  NAND2_X1 U3367 ( .A1(n2218), .A2(REG1_REG_16__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3368 ( .A1(n2220), .A2(REG2_REG_16__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3369 ( .A1(n2740), .A2(REG0_REG_16__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3370 ( .A1(n2679), .A2(n4726), .ZN(n2668) );
  NAND2_X1 U3371 ( .A1(n2668), .A2(IR_REG_31__SCAN_IN), .ZN(n2669) );
  XNOR2_X1 U3372 ( .A(n2669), .B(n2692), .ZN(n4515) );
  INV_X1 U3373 ( .A(n4515), .ZN(n2670) );
  MUX2_X1 U3374 ( .A(n2670), .B(DATAI_16_), .S(n3806), .Z(n3575) );
  NAND2_X1 U3375 ( .A1(n3560), .A2(n3575), .ZN(n3843) );
  NAND2_X1 U3376 ( .A1(n3713), .A2(n4345), .ZN(n3848) );
  INV_X1 U3377 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2672) );
  XNOR2_X1 U3378 ( .A(n2683), .B(n2672), .ZN(n3652) );
  NAND2_X1 U3379 ( .A1(n2764), .A2(n3652), .ZN(n2676) );
  NAND2_X1 U3380 ( .A1(n2218), .A2(REG1_REG_17__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3381 ( .A1(n3086), .A2(REG2_REG_17__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3382 ( .A1(n2740), .A2(REG0_REG_17__SCAN_IN), .ZN(n2673) );
  INV_X1 U3383 ( .A(n4347), .ZN(n4189) );
  OR2_X1 U3384 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2677)
         );
  NAND2_X1 U3385 ( .A1(IR_REG_31__SCAN_IN), .A2(n2677), .ZN(n2678) );
  NAND2_X1 U3386 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  XNOR2_X1 U3387 ( .A(n2680), .B(IR_REG_17__SCAN_IN), .ZN(n4513) );
  INV_X1 U3388 ( .A(DATAI_17_), .ZN(n4512) );
  MUX2_X1 U3389 ( .A(n4513), .B(n4512), .S(n3806), .Z(n3650) );
  NAND2_X1 U3390 ( .A1(n4189), .A2(n3650), .ZN(n2682) );
  AOI21_X1 U3391 ( .B1(n3557), .B2(n2682), .A(n2681), .ZN(n4195) );
  NAND2_X1 U3392 ( .A1(n2218), .A2(REG1_REG_18__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3393 ( .A1(n2683), .A2(REG3_REG_17__SCAN_IN), .ZN(n2685) );
  INV_X1 U3394 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3395 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  AND2_X1 U3396 ( .A1(n2686), .A2(n2698), .ZN(n4199) );
  NAND2_X1 U3397 ( .A1(n2739), .A2(n4199), .ZN(n2689) );
  NAND2_X1 U3398 ( .A1(n2740), .A2(REG0_REG_18__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U3399 ( .A1(n2220), .A2(REG2_REG_18__SCAN_IN), .ZN(n2687) );
  INV_X1 U3400 ( .A(n4170), .ZN(n3613) );
  NAND3_X1 U3401 ( .A1(n2692), .A2(n4726), .A3(n2691), .ZN(n2693) );
  INV_X1 U3402 ( .A(n2702), .ZN(n2694) );
  NAND2_X1 U3403 ( .A1(n2694), .A2(IR_REG_31__SCAN_IN), .ZN(n2695) );
  XNOR2_X1 U3404 ( .A(n2695), .B(IR_REG_18__SCAN_IN), .ZN(n3967) );
  MUX2_X1 U3405 ( .A(n3967), .B(DATAI_18_), .S(n3806), .Z(n4196) );
  NAND2_X1 U3406 ( .A1(n3613), .A2(n4196), .ZN(n4140) );
  NAND2_X1 U3407 ( .A1(n4170), .A2(n3693), .ZN(n4162) );
  NAND2_X1 U3408 ( .A1(n4140), .A2(n4162), .ZN(n4194) );
  NAND2_X1 U3409 ( .A1(n4195), .A2(n4194), .ZN(n4193) );
  AOI22_X1 U3410 ( .A1(n2218), .A2(REG1_REG_19__SCAN_IN), .B1(n2740), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3411 ( .A1(n2698), .A2(n2697), .ZN(n2699) );
  AND2_X1 U3412 ( .A1(n2708), .A2(n2699), .ZN(n4177) );
  AOI22_X1 U3413 ( .A1(n2764), .A2(n4177), .B1(n3086), .B2(
        REG2_REG_19__SCAN_IN), .ZN(n2700) );
  XNOR2_X2 U3414 ( .A(n2773), .B(IR_REG_19__SCAN_IN), .ZN(n4327) );
  MUX2_X1 U3415 ( .A(n4327), .B(DATAI_19_), .S(n3806), .Z(n4169) );
  NAND2_X1 U3416 ( .A1(n4186), .A2(n4169), .ZN(n2704) );
  OAI21_X1 U3417 ( .B1(n4147), .B2(n3887), .A(n4137), .ZN(n2705) );
  INV_X1 U3418 ( .A(n2708), .ZN(n2706) );
  AOI21_X1 U3419 ( .B1(n2706), .B2(REG3_REG_20__SCAN_IN), .A(
        REG3_REG_21__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U3420 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2707) );
  OR2_X1 U3421 ( .A1(n2709), .A2(n2713), .ZN(n4125) );
  AOI22_X1 U3422 ( .A1(n2218), .A2(REG1_REG_21__SCAN_IN), .B1(n2740), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3423 ( .A1(n2220), .A2(REG2_REG_21__SCAN_IN), .ZN(n2710) );
  OAI211_X1 U3424 ( .C1(n4125), .C2(n2535), .A(n2711), .B(n2710), .ZN(n4148)
         );
  NAND2_X1 U3425 ( .A1(n3806), .A2(DATAI_21_), .ZN(n3624) );
  INV_X1 U3426 ( .A(n4148), .ZN(n4108) );
  NOR2_X1 U3427 ( .A1(n2713), .A2(REG3_REG_22__SCAN_IN), .ZN(n2714) );
  OR2_X1 U3428 ( .A1(n2717), .A2(n2714), .ZN(n3680) );
  AOI22_X1 U3429 ( .A1(n2218), .A2(REG1_REG_22__SCAN_IN), .B1(n2740), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3430 ( .A1(n3086), .A2(REG2_REG_22__SCAN_IN), .ZN(n2715) );
  OAI211_X1 U3431 ( .C1(n3680), .C2(n2535), .A(n2716), .B(n2715), .ZN(n4132)
         );
  NAND2_X1 U3432 ( .A1(n3806), .A2(DATAI_22_), .ZN(n4114) );
  OR2_X1 U3433 ( .A1(n4132), .A2(n4114), .ZN(n4088) );
  NAND2_X1 U3434 ( .A1(n4132), .A2(n4114), .ZN(n2805) );
  NAND2_X1 U3435 ( .A1(n4088), .A2(n2805), .ZN(n4104) );
  OR2_X1 U3436 ( .A1(n2717), .A2(REG3_REG_23__SCAN_IN), .ZN(n2718) );
  AND2_X1 U3437 ( .A1(n2727), .A2(n2718), .ZN(n4098) );
  NAND2_X1 U3438 ( .A1(n4098), .A2(n2739), .ZN(n2724) );
  INV_X1 U3439 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4239) );
  NAND2_X1 U3440 ( .A1(n2740), .A2(REG0_REG_23__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3441 ( .A1(n3086), .A2(REG2_REG_23__SCAN_IN), .ZN(n2720) );
  OAI211_X1 U3442 ( .C1(n2719), .C2(n4239), .A(n2721), .B(n2720), .ZN(n2722)
         );
  INV_X1 U3443 ( .A(n2722), .ZN(n2723) );
  NAND2_X1 U3444 ( .A1(n3806), .A2(DATAI_23_), .ZN(n4097) );
  NAND2_X1 U3445 ( .A1(n4106), .A2(n4097), .ZN(n2726) );
  NOR2_X1 U3446 ( .A1(n4106), .A2(n4097), .ZN(n2725) );
  AOI21_X1 U3447 ( .B1(n4084), .B2(n2726), .A(n2725), .ZN(n4064) );
  INV_X1 U3448 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3660) );
  NAND2_X1 U3449 ( .A1(n2727), .A2(n3660), .ZN(n2728) );
  NAND2_X1 U3450 ( .A1(n2737), .A2(n2728), .ZN(n4078) );
  OR2_X1 U3451 ( .A1(n4078), .A2(n2535), .ZN(n2733) );
  INV_X1 U3452 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U3453 ( .A1(n2740), .A2(REG0_REG_24__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U3454 ( .A1(n2220), .A2(REG2_REG_24__SCAN_IN), .ZN(n2729) );
  OAI211_X1 U3455 ( .C1(n2719), .C2(n4235), .A(n2730), .B(n2729), .ZN(n2731)
         );
  INV_X1 U3456 ( .A(n2731), .ZN(n2732) );
  NAND2_X1 U3457 ( .A1(n3096), .A2(n4070), .ZN(n2734) );
  NAND2_X1 U34580 ( .A1(n4064), .A2(n2734), .ZN(n2736) );
  NAND2_X1 U34590 ( .A1(n4095), .A2(n4076), .ZN(n2735) );
  NAND2_X1 U3460 ( .A1(n2736), .A2(n2735), .ZN(n4047) );
  INV_X1 U3461 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U3462 ( .A1(n2737), .A2(n3638), .ZN(n2738) );
  NAND2_X1 U3463 ( .A1(n4059), .A2(n2739), .ZN(n2745) );
  INV_X1 U3464 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U3465 ( .A1(n3086), .A2(REG2_REG_25__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U3466 ( .A1(n2740), .A2(REG0_REG_25__SCAN_IN), .ZN(n2741) );
  OAI211_X1 U34670 ( .C1(n2719), .C2(n4834), .A(n2742), .B(n2741), .ZN(n2743)
         );
  INV_X1 U3468 ( .A(n2743), .ZN(n2744) );
  NAND2_X1 U34690 ( .A1(n3806), .A2(DATAI_25_), .ZN(n4053) );
  NOR2_X1 U3470 ( .A1(n4034), .A2(n4058), .ZN(n2747) );
  INV_X1 U34710 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3703) );
  AND2_X1 U3472 ( .A1(n2748), .A2(n3703), .ZN(n2749) );
  INV_X1 U34730 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U3474 ( .A1(n3086), .A2(REG2_REG_26__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U34750 ( .A1(n2527), .A2(REG0_REG_26__SCAN_IN), .ZN(n2750) );
  OAI211_X1 U3476 ( .C1(n2719), .C2(n4771), .A(n2751), .B(n2750), .ZN(n2752)
         );
  INV_X1 U34770 ( .A(n2752), .ZN(n2753) );
  OAI21_X1 U3478 ( .B1(n4041), .B2(n2535), .A(n2753), .ZN(n4055) );
  NAND2_X1 U34790 ( .A1(n3806), .A2(DATAI_26_), .ZN(n4040) );
  AND2_X1 U3480 ( .A1(n4055), .A2(n4033), .ZN(n3816) );
  INV_X1 U34810 ( .A(n4055), .ZN(n3593) );
  NAND2_X1 U3482 ( .A1(n3593), .A2(n4040), .ZN(n3817) );
  OR2_X1 U34830 ( .A1(n2754), .A2(REG3_REG_27__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U3484 ( .A1(n2754), .A2(REG3_REG_27__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U34850 ( .A1(n4024), .A2(n2764), .ZN(n2761) );
  INV_X1 U3486 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U34870 ( .A1(n3086), .A2(REG2_REG_27__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U3488 ( .A1(n2740), .A2(REG0_REG_27__SCAN_IN), .ZN(n2756) );
  OAI211_X1 U34890 ( .C1(n2719), .C2(n2758), .A(n2757), .B(n2756), .ZN(n2759)
         );
  INV_X1 U3490 ( .A(n2759), .ZN(n2760) );
  AND2_X1 U34910 ( .A1(n3806), .A2(DATAI_27_), .ZN(n4017) );
  INV_X1 U3492 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U34930 ( .A1(n2762), .A2(n3051), .ZN(n2763) );
  NAND2_X1 U3494 ( .A1(n4005), .A2(n2764), .ZN(n2769) );
  INV_X1 U34950 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U3496 ( .A1(n3086), .A2(REG2_REG_28__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U34970 ( .A1(n2527), .A2(REG0_REG_28__SCAN_IN), .ZN(n2765) );
  OAI211_X1 U3498 ( .C1(n2719), .C2(n3065), .A(n2766), .B(n2765), .ZN(n2767)
         );
  INV_X1 U34990 ( .A(n2767), .ZN(n2768) );
  INV_X1 U3500 ( .A(n4019), .ZN(n3885) );
  AND2_X1 U35010 ( .A1(n3806), .A2(DATAI_28_), .ZN(n2857) );
  INV_X1 U3502 ( .A(n2857), .ZN(n3994) );
  NAND2_X1 U35030 ( .A1(n3885), .A2(n3994), .ZN(n3985) );
  NAND2_X1 U3504 ( .A1(n4019), .A2(n2857), .ZN(n3983) );
  NAND2_X1 U35050 ( .A1(n3985), .A2(n3983), .ZN(n3995) );
  NAND2_X1 U35060 ( .A1(n2773), .A2(n2776), .ZN(n2770) );
  XNOR2_X2 U35070 ( .A(n2771), .B(n2777), .ZN(n2782) );
  OAI21_X1 U35080 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U35090 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  XNOR2_X2 U35100 ( .A(n2774), .B(n2775), .ZN(n2816) );
  AND3_X1 U35110 ( .A1(n2777), .A2(n2776), .A3(n2775), .ZN(n2778) );
  INV_X1 U35120 ( .A(n2870), .ZN(n4325) );
  XNOR2_X1 U35130 ( .A(n3146), .B(n4325), .ZN(n2781) );
  INV_X1 U35140 ( .A(n4327), .ZN(n3972) );
  NAND2_X1 U35150 ( .A1(n2781), .A2(n3972), .ZN(n3519) );
  NAND3_X1 U35160 ( .A1(n2782), .A2(n4327), .A3(n2870), .ZN(n4528) );
  NAND2_X1 U35170 ( .A1(n3519), .A2(n4528), .ZN(n4569) );
  NOR2_X1 U35180 ( .A1(n2267), .A2(n2784), .ZN(n2783) );
  MUX2_X1 U35190 ( .A(n2784), .B(n2783), .S(IR_REG_28__SCAN_IN), .Z(n2785) );
  INV_X1 U35200 ( .A(n2785), .ZN(n2787) );
  NAND2_X1 U35210 ( .A1(n2787), .A2(n2786), .ZN(n3048) );
  NAND2_X1 U35220 ( .A1(n3104), .A2(n4533), .ZN(n4491) );
  OR2_X1 U35230 ( .A1(n4492), .A2(n4491), .ZN(n4495) );
  NAND2_X1 U35240 ( .A1(n4495), .A2(n3730), .ZN(n2788) );
  NAND2_X1 U35250 ( .A1(n2788), .A2(n3196), .ZN(n3207) );
  NAND2_X1 U35260 ( .A1(n3207), .A2(n3731), .ZN(n2789) );
  XNOR2_X1 U35270 ( .A(n3899), .B(n3735), .ZN(n3811) );
  NAND2_X1 U35280 ( .A1(n2789), .A2(n3811), .ZN(n3209) );
  NAND2_X1 U35290 ( .A1(n2897), .A2(n3735), .ZN(n3736) );
  NAND2_X1 U35300 ( .A1(n3209), .A2(n3736), .ZN(n3168) );
  INV_X1 U35310 ( .A(n3737), .ZN(n2790) );
  INV_X1 U35320 ( .A(n3153), .ZN(n3267) );
  AND2_X1 U35330 ( .A1(n3897), .A2(n3267), .ZN(n3140) );
  INV_X1 U35340 ( .A(n3897), .ZN(n3226) );
  NAND2_X1 U35350 ( .A1(n3226), .A2(n3153), .ZN(n3751) );
  NAND2_X1 U35360 ( .A1(n3896), .A2(n3257), .ZN(n3752) );
  NAND2_X1 U35370 ( .A1(n3266), .A2(n3224), .ZN(n3742) );
  NAND2_X1 U35380 ( .A1(n2791), .A2(n3742), .ZN(n3238) );
  INV_X1 U35390 ( .A(n2792), .ZN(n2793) );
  NAND2_X1 U35400 ( .A1(n3312), .A2(n3280), .ZN(n3746) );
  NAND2_X1 U35410 ( .A1(n3894), .A2(n3322), .ZN(n3753) );
  AND2_X1 U35420 ( .A1(n3893), .A2(n3354), .ZN(n3303) );
  NAND2_X1 U35430 ( .A1(n3332), .A2(n3309), .ZN(n3747) );
  NAND2_X1 U35440 ( .A1(n3892), .A2(n3423), .ZN(n3765) );
  NAND2_X1 U35450 ( .A1(n3365), .A2(n3328), .ZN(n3759) );
  NAND2_X1 U35460 ( .A1(n2795), .A2(n3771), .ZN(n3371) );
  NOR2_X1 U35470 ( .A1(n3508), .A2(n3496), .ZN(n3768) );
  NAND2_X1 U35480 ( .A1(n3508), .A2(n3496), .ZN(n3763) );
  AND2_X1 U35490 ( .A1(n3890), .A2(n3511), .ZN(n3404) );
  NAND2_X1 U35500 ( .A1(n3550), .A2(n3407), .ZN(n3772) );
  NAND2_X1 U35510 ( .A1(n4344), .A2(n3534), .ZN(n3773) );
  NAND2_X1 U35520 ( .A1(n3888), .A2(n3717), .ZN(n3750) );
  NAND2_X1 U35530 ( .A1(n3773), .A2(n3750), .ZN(n3791) );
  INV_X1 U35540 ( .A(n3530), .ZN(n3842) );
  NOR2_X1 U35550 ( .A1(n3791), .A2(n3842), .ZN(n2796) );
  NAND2_X1 U35560 ( .A1(n3531), .A2(n2796), .ZN(n2797) );
  NAND2_X1 U35570 ( .A1(n2797), .A2(n3750), .ZN(n3568) );
  INV_X1 U35580 ( .A(n3826), .ZN(n2798) );
  NAND2_X1 U35590 ( .A1(n3568), .A2(n2798), .ZN(n2799) );
  NAND2_X1 U35600 ( .A1(n2799), .A2(n3848), .ZN(n3558) );
  AND2_X1 U35610 ( .A1(n4347), .A2(n3650), .ZN(n3780) );
  NAND2_X1 U35620 ( .A1(n4186), .A2(n4175), .ZN(n2800) );
  NAND2_X1 U35630 ( .A1(n4189), .A2(n3563), .ZN(n4138) );
  NAND2_X1 U35640 ( .A1(n4140), .A2(n4138), .ZN(n2801) );
  NAND2_X1 U35650 ( .A1(n2801), .A2(n3849), .ZN(n2804) );
  NAND2_X1 U35660 ( .A1(n4151), .A2(n4169), .ZN(n4142) );
  NAND2_X1 U35670 ( .A1(n4173), .A2(n4147), .ZN(n2802) );
  AND2_X1 U35680 ( .A1(n4142), .A2(n2802), .ZN(n2803) );
  NAND2_X1 U35690 ( .A1(n3887), .A2(n4153), .ZN(n3850) );
  OR2_X1 U35700 ( .A1(n4148), .A2(n3624), .ZN(n4085) );
  NAND2_X1 U35710 ( .A1(n4071), .A2(n4097), .ZN(n2806) );
  AND2_X1 U35720 ( .A1(n2806), .A2(n2805), .ZN(n3785) );
  AND2_X1 U35730 ( .A1(n4148), .A2(n3624), .ZN(n3819) );
  NAND2_X1 U35740 ( .A1(n4088), .A2(n3819), .ZN(n2807) );
  NAND2_X1 U35750 ( .A1(n3785), .A2(n2807), .ZN(n3855) );
  NAND2_X1 U35760 ( .A1(n4095), .A2(n4070), .ZN(n3805) );
  OR2_X1 U35770 ( .A1(n4071), .A2(n4097), .ZN(n4065) );
  NAND2_X1 U35780 ( .A1(n4066), .A2(n3852), .ZN(n4049) );
  NAND2_X1 U35790 ( .A1(n4034), .A2(n4053), .ZN(n3794) );
  NAND2_X1 U35800 ( .A1(n3096), .A2(n4076), .ZN(n4048) );
  NAND2_X1 U35810 ( .A1(n4049), .A2(n3863), .ZN(n2808) );
  NAND2_X1 U3582 ( .A1(n4074), .A2(n4058), .ZN(n3795) );
  NAND2_X1 U3583 ( .A1(n2808), .A2(n3795), .ZN(n4031) );
  NOR2_X1 U3584 ( .A1(n4055), .A2(n4040), .ZN(n3725) );
  NAND2_X1 U3585 ( .A1(n4055), .A2(n4040), .ZN(n3836) );
  NAND2_X1 U3586 ( .A1(n3886), .A2(n4023), .ZN(n3787) );
  NAND2_X1 U3587 ( .A1(n4037), .A2(n4017), .ZN(n3856) );
  NAND2_X1 U3588 ( .A1(n3787), .A2(n3856), .ZN(n4013) );
  XOR2_X1 U3589 ( .A(n3995), .B(n3986), .Z(n2811) );
  INV_X1 U3590 ( .A(n2782), .ZN(n4326) );
  NAND2_X1 U3591 ( .A1(n4326), .A2(n2816), .ZN(n3867) );
  NAND2_X1 U3592 ( .A1(n4325), .A2(n4327), .ZN(n2810) );
  NAND2_X1 U3593 ( .A1(n2811), .A2(n4167), .ZN(n2819) );
  INV_X1 U3594 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4770) );
  NAND2_X1 U3595 ( .A1(n2527), .A2(REG0_REG_29__SCAN_IN), .ZN(n2813) );
  NAND2_X1 U3596 ( .A1(n3086), .A2(REG2_REG_29__SCAN_IN), .ZN(n2812) );
  OAI211_X1 U3597 ( .C1(n2719), .C2(n4770), .A(n2813), .B(n2812), .ZN(n2814)
         );
  INV_X1 U3598 ( .A(n2814), .ZN(n2815) );
  OAI21_X1 U3599 ( .B1(n3982), .B2(n2535), .A(n2815), .ZN(n3884) );
  NAND2_X1 U3600 ( .A1(n3083), .A2(n3048), .ZN(n4489) );
  INV_X1 U3601 ( .A(n2816), .ZN(n2817) );
  AND2_X2 U3602 ( .A1(n2482), .A2(n4326), .ZN(n4486) );
  AOI22_X1 U3603 ( .A1(n3884), .A2(n4185), .B1(n2857), .B2(n4486), .ZN(n2818)
         );
  OAI211_X1 U3604 ( .C1(n4037), .C2(n4188), .A(n2819), .B(n2818), .ZN(n4009)
         );
  AOI21_X1 U3605 ( .B1(n4004), .B2(n4569), .A(n4009), .ZN(n3064) );
  NAND2_X1 U3606 ( .A1(n2821), .A2(n2820), .ZN(n2827) );
  NAND2_X1 U3607 ( .A1(n2840), .A2(n2822), .ZN(n2823) );
  OAI21_X1 U3608 ( .B1(n2827), .B2(n2823), .A(IR_REG_31__SCAN_IN), .ZN(n2824)
         );
  MUX2_X1 U3609 ( .A(IR_REG_31__SCAN_IN), .B(n2824), .S(IR_REG_25__SCAN_IN), 
        .Z(n2826) );
  NAND2_X1 U3610 ( .A1(n2826), .A2(n2825), .ZN(n2838) );
  NAND2_X1 U3611 ( .A1(n2838), .A2(B_REG_SCAN_IN), .ZN(n2830) );
  OR2_X1 U3612 ( .A1(n2784), .A2(n2840), .ZN(n2828) );
  XNOR2_X2 U3613 ( .A(n2829), .B(n2822), .ZN(n3072) );
  MUX2_X1 U3614 ( .A(n2830), .B(B_REG_SCAN_IN), .S(n3072), .Z(n2835) );
  NAND2_X1 U3615 ( .A1(n2825), .A2(IR_REG_31__SCAN_IN), .ZN(n2831) );
  MUX2_X1 U3616 ( .A(IR_REG_31__SCAN_IN), .B(n2831), .S(IR_REG_26__SCAN_IN), 
        .Z(n2832) );
  INV_X1 U3617 ( .A(n2832), .ZN(n2834) );
  NOR2_X1 U3618 ( .A1(n2834), .A2(n2833), .ZN(n4323) );
  NAND2_X1 U3619 ( .A1(n2835), .A2(n4323), .ZN(n3077) );
  INV_X1 U3620 ( .A(n3077), .ZN(n2853) );
  INV_X1 U3621 ( .A(D_REG_0__SCAN_IN), .ZN(n4899) );
  INV_X1 U3622 ( .A(n3072), .ZN(n2836) );
  INV_X1 U3623 ( .A(n4323), .ZN(n2837) );
  INV_X1 U3624 ( .A(n3062), .ZN(n3144) );
  NAND2_X1 U3625 ( .A1(n2838), .A2(n2837), .ZN(n3079) );
  OAI21_X1 U3626 ( .B1(n3077), .B2(D_REG_1__SCAN_IN), .A(n3079), .ZN(n2856) );
  INV_X1 U3627 ( .A(n2838), .ZN(n4324) );
  XNOR2_X1 U3628 ( .A(n2839), .B(n2840), .ZN(n3084) );
  NAND2_X1 U3629 ( .A1(n2869), .A2(n4510), .ZN(n3081) );
  OR2_X1 U3630 ( .A1(n4528), .A2(n2816), .ZN(n3046) );
  NAND2_X1 U3631 ( .A1(n2782), .A2(n3972), .ZN(n2841) );
  NAND2_X1 U3632 ( .A1(n3083), .A2(n2841), .ZN(n3141) );
  NAND2_X1 U3633 ( .A1(n3046), .A2(n3141), .ZN(n2842) );
  NOR2_X1 U3634 ( .A1(n3081), .A2(n2842), .ZN(n2855) );
  NOR2_X1 U3635 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_8__SCAN_IN), .ZN(n2846) );
  NOR4_X1 U3636 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2845) );
  NOR4_X1 U3637 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2844) );
  NOR4_X1 U3638 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2843) );
  AND4_X1 U3639 ( .A1(n2846), .A2(n2845), .A3(n2844), .A4(n2843), .ZN(n2852)
         );
  NOR4_X1 U3640 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2850) );
  NOR4_X1 U3641 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2849) );
  NOR4_X1 U3642 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2848) );
  NOR4_X1 U3643 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2847) );
  AND4_X1 U3644 ( .A1(n2850), .A2(n2849), .A3(n2848), .A4(n2847), .ZN(n2851)
         );
  NAND2_X1 U3645 ( .A1(n2852), .A2(n2851), .ZN(n3035) );
  NAND2_X1 U3646 ( .A1(n2853), .A2(n3035), .ZN(n2854) );
  NAND2_X1 U3647 ( .A1(n2879), .A2(n3160), .ZN(n4502) );
  NOR2_X1 U3648 ( .A1(n4502), .A2(n2888), .ZN(n4540) );
  NAND2_X1 U3649 ( .A1(n4540), .A2(n3216), .ZN(n3218) );
  INV_X1 U3650 ( .A(n4022), .ZN(n2858) );
  OAI21_X1 U3651 ( .B1(n2858), .B2(n3994), .A(n3999), .ZN(n4007) );
  NAND2_X2 U3652 ( .A1(n2782), .A2(n2482), .ZN(n4560) );
  NAND2_X1 U3653 ( .A1(n4580), .A2(n4577), .ZN(n4312) );
  INV_X1 U3654 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U3655 ( .A1(n4578), .A2(REG0_REG_28__SCAN_IN), .ZN(n2859) );
  OAI21_X1 U3656 ( .B1(n3064), .B2(n4578), .A(n2861), .ZN(U3514) );
  AND2_X4 U3657 ( .A1(n2862), .A2(n2864), .ZN(n2896) );
  INV_X1 U3658 ( .A(n2862), .ZN(n2863) );
  OAI22_X1 U3659 ( .A1(n3497), .A2(n3029), .B1(n2219), .B2(n3391), .ZN(n2931)
         );
  INV_X1 U3660 ( .A(n2931), .ZN(n3386) );
  NAND2_X1 U3661 ( .A1(n2867), .A2(n3043), .ZN(n2866) );
  NAND2_X1 U3662 ( .A1(n2896), .A2(n4533), .ZN(n2865) );
  NAND2_X1 U3663 ( .A1(n2866), .A2(n2865), .ZN(n3111) );
  NAND2_X1 U3664 ( .A1(n3043), .A2(n4533), .ZN(n2868) );
  OAI21_X1 U3665 ( .B1(n3104), .B2(n2887), .A(n2868), .ZN(n3115) );
  NAND2_X1 U3666 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3902) );
  INV_X1 U3667 ( .A(n3111), .ZN(n2873) );
  NOR2_X1 U3668 ( .A1(n2870), .A2(n4327), .ZN(n3041) );
  INV_X1 U3669 ( .A(n3041), .ZN(n2871) );
  NAND2_X4 U3670 ( .A1(n2871), .A2(n3146), .ZN(n3030) );
  NAND2_X1 U3671 ( .A1(n3117), .A2(n2874), .ZN(n3108) );
  NAND2_X1 U3672 ( .A1(n2875), .A2(n2895), .ZN(n2877) );
  NAND2_X1 U3673 ( .A1(n2896), .A2(n4500), .ZN(n2876) );
  NAND2_X1 U3674 ( .A1(n2877), .A2(n2876), .ZN(n2878) );
  INV_X1 U3675 ( .A(n2880), .ZN(n2882) );
  XNOR2_X1 U3676 ( .A(n2881), .B(n2882), .ZN(n3106) );
  NAND2_X1 U3677 ( .A1(n3108), .A2(n3106), .ZN(n3107) );
  NAND2_X1 U3678 ( .A1(n3107), .A2(n2883), .ZN(n3123) );
  NAND2_X1 U3679 ( .A1(n2889), .A2(n3043), .ZN(n2885) );
  NAND2_X1 U3680 ( .A1(n2896), .A2(n2888), .ZN(n2884) );
  NAND2_X1 U3681 ( .A1(n2885), .A2(n2884), .ZN(n2886) );
  INV_X2 U3682 ( .A(n2887), .ZN(n2894) );
  INV_X1 U3683 ( .A(n2892), .ZN(n2890) );
  INV_X1 U3684 ( .A(n2891), .ZN(n2893) );
  AOI22_X1 U3685 ( .A1(n2894), .A2(n3899), .B1(n3043), .B2(n3735), .ZN(n2900)
         );
  INV_X1 U3686 ( .A(n3899), .ZN(n2897) );
  OAI22_X1 U3687 ( .A1(n2897), .A2(n2219), .B1(n3028), .B2(n3216), .ZN(n2898)
         );
  XNOR2_X1 U3688 ( .A(n2898), .B(n3030), .ZN(n2899) );
  XOR2_X1 U3689 ( .A(n2900), .B(n2899), .Z(n3131) );
  INV_X1 U3690 ( .A(n2899), .ZN(n2901) );
  NAND2_X1 U3691 ( .A1(n2901), .A2(n2900), .ZN(n2902) );
  XNOR2_X1 U3692 ( .A(n2903), .B(n3030), .ZN(n2905) );
  OAI22_X1 U3693 ( .A1(n3152), .A2(n3029), .B1(n3019), .B2(n3180), .ZN(n2904)
         );
  XNOR2_X1 U3694 ( .A(n2905), .B(n2904), .ZN(n3181) );
  NOR2_X1 U3695 ( .A1(n3183), .A2(n3181), .ZN(n3182) );
  AND2_X1 U3696 ( .A1(n2905), .A2(n2904), .ZN(n2906) );
  NOR2_X1 U3697 ( .A1(n3182), .A2(n2906), .ZN(n3264) );
  NAND2_X1 U3698 ( .A1(n3897), .A2(n3015), .ZN(n2908) );
  NAND2_X1 U3699 ( .A1(n2896), .A2(n3153), .ZN(n2907) );
  NAND2_X1 U3700 ( .A1(n2908), .A2(n2907), .ZN(n2909) );
  XNOR2_X1 U3701 ( .A(n2909), .B(n3030), .ZN(n2911) );
  OAI22_X1 U3702 ( .A1(n3226), .A2(n3029), .B1(n3019), .B2(n3267), .ZN(n2910)
         );
  XNOR2_X1 U3703 ( .A(n2911), .B(n2910), .ZN(n3263) );
  NOR2_X1 U3704 ( .A1(n3264), .A2(n3263), .ZN(n3262) );
  OAI22_X1 U3705 ( .A1(n3266), .A2(n3029), .B1(n3019), .B2(n3257), .ZN(n3251)
         );
  OAI22_X1 U3706 ( .A1(n3266), .A2(n3019), .B1(n3028), .B2(n3257), .ZN(n2912)
         );
  XNOR2_X1 U3707 ( .A(n2912), .B(n3030), .ZN(n3252) );
  OAI22_X1 U3708 ( .A1(n3276), .A2(n3029), .B1(n3019), .B2(n3298), .ZN(n2914)
         );
  OAI22_X1 U3709 ( .A1(n3276), .A2(n3019), .B1(n3028), .B2(n3298), .ZN(n2913)
         );
  XNOR2_X1 U3710 ( .A(n2913), .B(n3030), .ZN(n2915) );
  XOR2_X1 U3711 ( .A(n2914), .B(n2915), .Z(n3295) );
  NAND2_X1 U3712 ( .A1(n3894), .A2(n3015), .ZN(n2917) );
  NAND2_X1 U3713 ( .A1(n2896), .A2(n3280), .ZN(n2916) );
  NAND2_X1 U3714 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  XNOR2_X1 U3715 ( .A(n2918), .B(n2872), .ZN(n2919) );
  AOI22_X1 U3716 ( .A1(n2894), .A2(n3894), .B1(n3015), .B2(n3280), .ZN(n2920)
         );
  OR2_X1 U3717 ( .A1(n2919), .A2(n2920), .ZN(n3317) );
  AND2_X1 U3718 ( .A1(n2920), .A2(n2919), .ZN(n3316) );
  AOI22_X1 U3719 ( .A1(n2894), .A2(n3893), .B1(n3015), .B2(n3309), .ZN(n2923)
         );
  OAI22_X1 U3720 ( .A1(n3332), .A2(n3019), .B1(n3028), .B2(n3354), .ZN(n2921)
         );
  XNOR2_X1 U3721 ( .A(n2921), .B(n3030), .ZN(n2922) );
  XOR2_X1 U3722 ( .A(n2923), .B(n2922), .Z(n3351) );
  INV_X1 U3723 ( .A(n2922), .ZN(n2924) );
  NAND2_X1 U3724 ( .A1(n2924), .A2(n2923), .ZN(n2925) );
  OAI22_X1 U3725 ( .A1(n3365), .A2(n3019), .B1(n3028), .B2(n3423), .ZN(n2926)
         );
  XNOR2_X1 U3726 ( .A(n2926), .B(n3030), .ZN(n2927) );
  OAI22_X1 U3727 ( .A1(n3365), .A2(n3029), .B1(n3019), .B2(n3423), .ZN(n2928)
         );
  XNOR2_X1 U3728 ( .A(n2927), .B(n2928), .ZN(n3427) );
  INV_X1 U3729 ( .A(n3385), .ZN(n2933) );
  OAI22_X1 U3730 ( .A1(n3497), .A2(n3019), .B1(n3028), .B2(n3391), .ZN(n2930)
         );
  XNOR2_X1 U3731 ( .A(n2930), .B(n3030), .ZN(n3387) );
  AOI22_X1 U3732 ( .A1(n2894), .A2(n3508), .B1(n3015), .B2(n3377), .ZN(n2938)
         );
  NAND2_X1 U3733 ( .A1(n3508), .A2(n3015), .ZN(n2935) );
  NAND2_X1 U3734 ( .A1(n2896), .A2(n3377), .ZN(n2934) );
  NAND2_X1 U3735 ( .A1(n2935), .A2(n2934), .ZN(n2936) );
  XNOR2_X1 U3736 ( .A(n2936), .B(n2872), .ZN(n2937) );
  NOR2_X1 U3737 ( .A1(n2938), .A2(n2937), .ZN(n3490) );
  NAND2_X1 U3738 ( .A1(n2938), .A2(n2937), .ZN(n3491) );
  OAI22_X1 U3739 ( .A1(n3550), .A2(n3019), .B1(n3028), .B2(n3511), .ZN(n2939)
         );
  XOR2_X1 U3740 ( .A(n3030), .B(n2939), .Z(n2940) );
  INV_X1 U3741 ( .A(n2940), .ZN(n3504) );
  AOI22_X1 U3742 ( .A1(n2894), .A2(n3889), .B1(n3015), .B2(n3523), .ZN(n2945)
         );
  NAND2_X1 U3743 ( .A1(n3889), .A2(n3015), .ZN(n2942) );
  NAND2_X1 U3744 ( .A1(n2896), .A2(n3523), .ZN(n2941) );
  NAND2_X1 U3745 ( .A1(n2942), .A2(n2941), .ZN(n2943) );
  XNOR2_X1 U3746 ( .A(n2943), .B(n2872), .ZN(n2944) );
  OR2_X1 U3747 ( .A1(n2945), .A2(n2944), .ZN(n3546) );
  NAND2_X1 U3748 ( .A1(n3547), .A2(n3546), .ZN(n2946) );
  NAND2_X1 U3749 ( .A1(n2945), .A2(n2944), .ZN(n3545) );
  NAND2_X1 U3750 ( .A1(n2946), .A2(n3545), .ZN(n2956) );
  OAI22_X1 U3751 ( .A1(n4344), .A2(n3019), .B1(n3028), .B2(n3717), .ZN(n2947)
         );
  XOR2_X1 U3752 ( .A(n3030), .B(n2947), .Z(n2957) );
  NAND2_X1 U3753 ( .A1(n2956), .A2(n2957), .ZN(n3711) );
  NAND2_X1 U3754 ( .A1(n2894), .A2(n3888), .ZN(n2949) );
  NAND2_X1 U3755 ( .A1(n3015), .A2(n3534), .ZN(n2948) );
  NAND2_X1 U3756 ( .A1(n2949), .A2(n2948), .ZN(n4349) );
  NAND2_X1 U3757 ( .A1(n3711), .A2(n4349), .ZN(n2960) );
  AOI22_X1 U3758 ( .A1(n2894), .A2(n3713), .B1(n3015), .B2(n3575), .ZN(n2954)
         );
  NAND2_X1 U3759 ( .A1(n3713), .A2(n3015), .ZN(n2951) );
  NAND2_X1 U3760 ( .A1(n2896), .A2(n3575), .ZN(n2950) );
  NAND2_X1 U3761 ( .A1(n2951), .A2(n2950), .ZN(n2952) );
  XNOR2_X1 U3762 ( .A(n2952), .B(n2872), .ZN(n2953) );
  NAND2_X1 U3763 ( .A1(n2954), .A2(n2953), .ZN(n2961) );
  OAI21_X1 U3764 ( .B1(n2954), .B2(n2953), .A(n2961), .ZN(n2955) );
  INV_X1 U3765 ( .A(n2955), .ZN(n4351) );
  INV_X1 U3766 ( .A(n2956), .ZN(n2959) );
  NAND2_X1 U3767 ( .A1(n2959), .A2(n2958), .ZN(n3710) );
  NAND3_X1 U3768 ( .A1(n2960), .A2(n4351), .A3(n3710), .ZN(n2962) );
  AOI22_X1 U3769 ( .A1(n2894), .A2(n4347), .B1(n3015), .B2(n3563), .ZN(n2967)
         );
  NAND2_X1 U3770 ( .A1(n4347), .A2(n3015), .ZN(n2964) );
  NAND2_X1 U3771 ( .A1(n2896), .A2(n3563), .ZN(n2963) );
  NAND2_X1 U3772 ( .A1(n2964), .A2(n2963), .ZN(n2965) );
  XNOR2_X1 U3773 ( .A(n2965), .B(n2872), .ZN(n2966) );
  OR2_X1 U3774 ( .A1(n2967), .A2(n2966), .ZN(n3646) );
  NAND2_X1 U3775 ( .A1(n2967), .A2(n2966), .ZN(n3645) );
  NAND2_X1 U3776 ( .A1(n4170), .A2(n3015), .ZN(n2969) );
  NAND2_X1 U3777 ( .A1(n2896), .A2(n4196), .ZN(n2968) );
  NAND2_X1 U3778 ( .A1(n2969), .A2(n2968), .ZN(n2970) );
  XNOR2_X1 U3779 ( .A(n2970), .B(n2872), .ZN(n2972) );
  AOI22_X1 U3780 ( .A1(n2894), .A2(n4170), .B1(n3015), .B2(n4196), .ZN(n2971)
         );
  OR2_X1 U3781 ( .A1(n2972), .A2(n2971), .ZN(n3687) );
  NAND2_X1 U3782 ( .A1(n2972), .A2(n2971), .ZN(n3689) );
  NAND2_X1 U3783 ( .A1(n3685), .A2(n3689), .ZN(n3610) );
  OAI22_X1 U3784 ( .A1(n4151), .A2(n3019), .B1(n3028), .B2(n4175), .ZN(n2973)
         );
  XNOR2_X1 U3785 ( .A(n2973), .B(n3030), .ZN(n2975) );
  NOR2_X1 U3786 ( .A1(n3019), .A2(n4175), .ZN(n2974) );
  AOI21_X1 U3787 ( .B1(n4186), .B2(n2894), .A(n2974), .ZN(n2976) );
  XNOR2_X1 U3788 ( .A(n2975), .B(n2976), .ZN(n3611) );
  NAND2_X1 U3789 ( .A1(n3610), .A2(n3611), .ZN(n2979) );
  INV_X1 U3790 ( .A(n2975), .ZN(n2977) );
  NAND2_X1 U3791 ( .A1(n2977), .A2(n2976), .ZN(n2978) );
  NAND2_X1 U3792 ( .A1(n3887), .A2(n3015), .ZN(n2981) );
  NAND2_X1 U3793 ( .A1(n2896), .A2(n4147), .ZN(n2980) );
  NAND2_X1 U3794 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  XNOR2_X1 U3795 ( .A(n2982), .B(n2872), .ZN(n2984) );
  AOI22_X1 U3796 ( .A1(n2894), .A2(n3887), .B1(n3015), .B2(n4147), .ZN(n2983)
         );
  OR2_X1 U3797 ( .A1(n2984), .A2(n2983), .ZN(n3667) );
  NAND2_X1 U3798 ( .A1(n2984), .A2(n2983), .ZN(n3668) );
  NAND2_X1 U3799 ( .A1(n4148), .A2(n3015), .ZN(n2986) );
  NAND2_X1 U3800 ( .A1(n2896), .A2(n4131), .ZN(n2985) );
  NAND2_X1 U3801 ( .A1(n2986), .A2(n2985), .ZN(n2987) );
  XNOR2_X1 U3802 ( .A(n2987), .B(n3030), .ZN(n3619) );
  NAND2_X1 U3803 ( .A1(n2894), .A2(n4148), .ZN(n2989) );
  NAND2_X1 U3804 ( .A1(n3015), .A2(n4131), .ZN(n2988) );
  NAND2_X1 U3805 ( .A1(n2989), .A2(n2988), .ZN(n3620) );
  NOR2_X1 U3806 ( .A1(n3619), .A2(n3620), .ZN(n2990) );
  INV_X1 U3807 ( .A(n3677), .ZN(n2993) );
  OAI22_X1 U3808 ( .A1(n3626), .A2(n2219), .B1(n3028), .B2(n4114), .ZN(n2991)
         );
  XNOR2_X1 U3809 ( .A(n2991), .B(n3030), .ZN(n2995) );
  OAI22_X1 U3810 ( .A1(n3626), .A2(n3029), .B1(n3019), .B2(n4114), .ZN(n2994)
         );
  XNOR2_X1 U3811 ( .A(n2995), .B(n2994), .ZN(n3679) );
  NAND2_X1 U3812 ( .A1(n2993), .A2(n2992), .ZN(n3599) );
  NOR2_X1 U3813 ( .A1(n2995), .A2(n2994), .ZN(n3601) );
  NAND2_X1 U3814 ( .A1(n4071), .A2(n3015), .ZN(n2997) );
  INV_X1 U3815 ( .A(n4097), .ZN(n4092) );
  NAND2_X1 U3816 ( .A1(n2896), .A2(n4092), .ZN(n2996) );
  NAND2_X1 U3817 ( .A1(n2997), .A2(n2996), .ZN(n2998) );
  XNOR2_X1 U3818 ( .A(n2998), .B(n2872), .ZN(n3001) );
  NOR2_X1 U3819 ( .A1(n3019), .A2(n4097), .ZN(n2999) );
  AOI21_X1 U3820 ( .B1(n4071), .B2(n2894), .A(n2999), .ZN(n3000) );
  XNOR2_X1 U3821 ( .A(n3001), .B(n3000), .ZN(n3600) );
  NAND2_X1 U3822 ( .A1(n3599), .A2(n2260), .ZN(n3602) );
  NOR2_X1 U3823 ( .A1(n3001), .A2(n3000), .ZN(n3004) );
  OAI22_X1 U3824 ( .A1(n4095), .A2(n3029), .B1(n2219), .B2(n4076), .ZN(n3006)
         );
  NAND2_X1 U3825 ( .A1(n3602), .A2(n3002), .ZN(n3656) );
  OAI22_X1 U3826 ( .A1(n4095), .A2(n3019), .B1(n3028), .B2(n4076), .ZN(n3003)
         );
  XNOR2_X1 U3827 ( .A(n3003), .B(n3030), .ZN(n3657) );
  NAND2_X1 U3828 ( .A1(n3656), .A2(n3657), .ZN(n3008) );
  INV_X1 U3829 ( .A(n3004), .ZN(n3005) );
  NAND2_X1 U3830 ( .A1(n3602), .A2(n3005), .ZN(n3007) );
  NAND2_X1 U3831 ( .A1(n3007), .A2(n3006), .ZN(n3655) );
  NAND2_X1 U3832 ( .A1(n3008), .A2(n3655), .ZN(n3631) );
  NAND2_X1 U3833 ( .A1(n4034), .A2(n3015), .ZN(n3010) );
  NAND2_X1 U3834 ( .A1(n2896), .A2(n4058), .ZN(n3009) );
  NAND2_X1 U3835 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  XNOR2_X1 U3836 ( .A(n3011), .B(n2872), .ZN(n3014) );
  NOR2_X1 U3837 ( .A1(n3019), .A2(n4053), .ZN(n3012) );
  AOI21_X1 U3838 ( .B1(n4034), .B2(n2894), .A(n3012), .ZN(n3013) );
  NAND2_X1 U3839 ( .A1(n3014), .A2(n3013), .ZN(n3633) );
  NOR2_X1 U3840 ( .A1(n3014), .A2(n3013), .ZN(n3632) );
  NAND2_X1 U3841 ( .A1(n4055), .A2(n3015), .ZN(n3017) );
  NAND2_X1 U3842 ( .A1(n2896), .A2(n4033), .ZN(n3016) );
  NAND2_X1 U3843 ( .A1(n3017), .A2(n3016), .ZN(n3018) );
  XNOR2_X1 U3844 ( .A(n3018), .B(n2872), .ZN(n3024) );
  INV_X1 U3845 ( .A(n3024), .ZN(n3022) );
  NOR2_X1 U3846 ( .A1(n3019), .A2(n4040), .ZN(n3020) );
  AOI21_X1 U3847 ( .B1(n4055), .B2(n2894), .A(n3020), .ZN(n3023) );
  INV_X1 U3848 ( .A(n3023), .ZN(n3021) );
  NAND2_X1 U3849 ( .A1(n3022), .A2(n3021), .ZN(n3698) );
  AND2_X1 U3850 ( .A1(n3024), .A2(n3023), .ZN(n3699) );
  OAI22_X1 U3851 ( .A1(n4037), .A2(n3029), .B1(n3019), .B2(n4023), .ZN(n3027)
         );
  OAI22_X1 U3852 ( .A1(n4037), .A2(n3019), .B1(n4023), .B2(n3028), .ZN(n3025)
         );
  XNOR2_X1 U3853 ( .A(n3025), .B(n3030), .ZN(n3026) );
  XOR2_X1 U3854 ( .A(n3027), .B(n3026), .Z(n3591) );
  OAI22_X1 U3855 ( .A1(n4019), .A2(n3019), .B1(n3028), .B2(n3994), .ZN(n3033)
         );
  OAI22_X1 U3856 ( .A1(n4019), .A2(n3029), .B1(n3019), .B2(n3994), .ZN(n3031)
         );
  XNOR2_X1 U3857 ( .A(n3031), .B(n3030), .ZN(n3032) );
  XOR2_X1 U3858 ( .A(n3033), .B(n3032), .Z(n3034) );
  INV_X1 U3859 ( .A(D_REG_1__SCAN_IN), .ZN(n4902) );
  NOR2_X1 U3860 ( .A1(n3035), .A2(n4902), .ZN(n3036) );
  OAI21_X1 U3861 ( .B1(n3077), .B2(n3036), .A(n3079), .ZN(n3037) );
  INV_X1 U3862 ( .A(n3037), .ZN(n3143) );
  NAND2_X1 U3863 ( .A1(n3143), .A2(n3062), .ZN(n3058) );
  INV_X1 U3864 ( .A(n3058), .ZN(n3040) );
  AOI21_X1 U3865 ( .B1(n4327), .B2(n2482), .A(n3083), .ZN(n3038) );
  NAND2_X1 U3866 ( .A1(n4107), .A2(n3038), .ZN(n3054) );
  NOR2_X1 U3867 ( .A1(n3081), .A2(n3054), .ZN(n3039) );
  AND2_X1 U3868 ( .A1(n4510), .A2(n3041), .ZN(n3042) );
  NAND2_X1 U3869 ( .A1(n3878), .A2(n4321), .ZN(n3044) );
  INV_X1 U3870 ( .A(n3081), .ZN(n3142) );
  NAND2_X1 U3871 ( .A1(n3142), .A2(n4486), .ZN(n3045) );
  OR2_X1 U3872 ( .A1(n3058), .A2(n3045), .ZN(n3047) );
  AND2_X2 U3873 ( .A1(n3047), .A2(n4124), .ZN(n3705) );
  OAI22_X1 U3874 ( .A1(n4037), .A2(n4343), .B1(n3705), .B2(n3994), .ZN(n3053)
         );
  NAND2_X1 U3875 ( .A1(n3878), .A2(n3048), .ZN(n3049) );
  NAND2_X1 U3876 ( .A1(n3884), .A2(n4348), .ZN(n3050) );
  OAI21_X1 U3877 ( .B1(STATE_REG_SCAN_IN), .B2(n3051), .A(n3050), .ZN(n3052)
         );
  INV_X1 U3878 ( .A(n4005), .ZN(n3060) );
  NAND2_X1 U3879 ( .A1(n3054), .A2(n4107), .ZN(n3055) );
  NAND2_X1 U3880 ( .A1(n3058), .A2(n3055), .ZN(n3056) );
  NAND2_X1 U3881 ( .A1(n3056), .A2(n3141), .ZN(n3101) );
  NAND2_X1 U3882 ( .A1(n2869), .A2(n3084), .ZN(n3057) );
  OAI21_X1 U3883 ( .B1(n3101), .B2(n3057), .A(STATE_REG_SCAN_IN), .ZN(n3059)
         );
  NAND2_X1 U3884 ( .A1(n3058), .A2(n3878), .ZN(n3102) );
  MUX2_X2 U3885 ( .A(n3065), .B(n3064), .S(n4595), .Z(n3067) );
  NAND2_X1 U3886 ( .A1(n4595), .A2(n4577), .ZN(n4257) );
  NAND2_X1 U3887 ( .A1(n3067), .A2(n3066), .ZN(U3546) );
  INV_X1 U3888 ( .A(n4510), .ZN(n3068) );
  NOR2_X2 U3889 ( .A1(n2869), .A2(n3068), .ZN(U4043) );
  INV_X2 U3890 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3891 ( .A(DATAI_18_), .ZN(n3070) );
  NAND2_X1 U3892 ( .A1(n3967), .A2(STATE_REG_SCAN_IN), .ZN(n3069) );
  OAI21_X1 U3893 ( .B1(STATE_REG_SCAN_IN), .B2(n3070), .A(n3069), .ZN(U3334)
         );
  INV_X1 U3894 ( .A(DATAI_21_), .ZN(n4706) );
  NAND2_X1 U3895 ( .A1(n2816), .A2(STATE_REG_SCAN_IN), .ZN(n3071) );
  OAI21_X1 U3896 ( .B1(STATE_REG_SCAN_IN), .B2(n4706), .A(n3071), .ZN(U3331)
         );
  INV_X1 U3897 ( .A(DATAI_24_), .ZN(n4885) );
  NAND2_X1 U3898 ( .A1(n3072), .A2(STATE_REG_SCAN_IN), .ZN(n3073) );
  OAI21_X1 U3899 ( .B1(STATE_REG_SCAN_IN), .B2(n4885), .A(n3073), .ZN(U3328)
         );
  INV_X1 U3900 ( .A(DATAI_29_), .ZN(n3076) );
  NAND2_X1 U3901 ( .A1(n2504), .A2(STATE_REG_SCAN_IN), .ZN(n3075) );
  OAI21_X1 U3902 ( .B1(STATE_REG_SCAN_IN), .B2(n3076), .A(n3075), .ZN(U3323)
         );
  AOI22_X1 U3903 ( .A1(n4509), .A2(n4899), .B1(n3078), .B2(n4510), .ZN(U3458)
         );
  INV_X1 U3904 ( .A(n3079), .ZN(n3080) );
  AOI22_X1 U3905 ( .A1(n4509), .A2(n4902), .B1(n3080), .B2(n4510), .ZN(U3459)
         );
  OR2_X1 U3906 ( .A1(n3084), .A2(U3149), .ZN(n3882) );
  NAND2_X1 U3907 ( .A1(n3081), .A2(n3882), .ZN(n3433) );
  AOI21_X1 U3908 ( .B1(n3084), .B2(n3083), .A(n3082), .ZN(n3432) );
  INV_X1 U3909 ( .A(n3432), .ZN(n3085) );
  NOR2_X1 U3910 ( .A1(n4980), .A2(n3901), .ZN(U3148) );
  INV_X1 U3911 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3091) );
  INV_X1 U3912 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3913 ( .A1(n3086), .A2(REG2_REG_30__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3914 ( .A1(n2527), .A2(REG0_REG_30__SCAN_IN), .ZN(n3087) );
  OAI211_X1 U3915 ( .C1(n2719), .C2(n3089), .A(n3088), .B(n3087), .ZN(n3990)
         );
  NAND2_X1 U3916 ( .A1(U4043), .A2(n3990), .ZN(n3090) );
  OAI21_X1 U3917 ( .B1(n3901), .B2(n3091), .A(n3090), .ZN(U3580) );
  INV_X1 U3918 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4876) );
  NAND2_X1 U3919 ( .A1(U4043), .A2(n3508), .ZN(n3092) );
  OAI21_X1 U3920 ( .B1(n3901), .B2(n4876), .A(n3092), .ZN(U3562) );
  INV_X1 U3921 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U3922 ( .A1(U4043), .A2(n2889), .ZN(n3093) );
  OAI21_X1 U3923 ( .B1(n3901), .B2(n4793), .A(n3093), .ZN(U3552) );
  INV_X1 U3924 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U3925 ( .A1(n4071), .A2(U4043), .ZN(n3094) );
  OAI21_X1 U3926 ( .B1(n3901), .B2(n4920), .A(n3094), .ZN(U3573) );
  INV_X1 U3927 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U3928 ( .A1(n4186), .A2(U4043), .ZN(n3095) );
  OAI21_X1 U3929 ( .B1(n3901), .B2(n4850), .A(n3095), .ZN(U3569) );
  INV_X1 U3930 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U3931 ( .A1(n3096), .A2(U4043), .ZN(n3097) );
  OAI21_X1 U3932 ( .B1(n3901), .B2(n4796), .A(n3097), .ZN(U3574) );
  INV_X1 U3933 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U3934 ( .A1(n3901), .A2(n4347), .ZN(n3098) );
  OAI21_X1 U3935 ( .B1(n3901), .B2(n4792), .A(n3098), .ZN(U3567) );
  INV_X1 U3936 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U3937 ( .A1(n3901), .A2(n3713), .ZN(n3099) );
  OAI21_X1 U3938 ( .B1(n3901), .B2(n4840), .A(n3099), .ZN(U3566) );
  INV_X1 U3939 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U3940 ( .A1(n4148), .A2(U4043), .ZN(n3100) );
  OAI21_X1 U3941 ( .B1(n3901), .B2(n4849), .A(n3100), .ZN(U3571) );
  INV_X1 U3942 ( .A(n3101), .ZN(n3103) );
  NAND3_X1 U3943 ( .A1(n3103), .A2(n3142), .A3(n3102), .ZN(n3128) );
  INV_X1 U3944 ( .A(n3128), .ZN(n3121) );
  INV_X1 U3945 ( .A(n3705), .ZN(n3119) );
  OAI22_X1 U3946 ( .A1(n3104), .A2(n4343), .B1(n3704), .B2(n4490), .ZN(n3105)
         );
  AOI21_X1 U3947 ( .B1(n4500), .B2(n3119), .A(n3105), .ZN(n3110) );
  OAI211_X1 U3948 ( .C1(n3106), .C2(n3108), .A(n3107), .B(n4353), .ZN(n3109)
         );
  OAI211_X1 U3949 ( .C1(n3121), .C2(n2512), .A(n3110), .B(n3109), .ZN(U3219)
         );
  INV_X1 U3950 ( .A(n2869), .ZN(n3112) );
  OAI21_X1 U3951 ( .B1(IR_REG_0__SCAN_IN), .B2(REG1_REG_0__SCAN_IN), .A(n3112), 
        .ZN(n3113) );
  NAND2_X1 U3952 ( .A1(n2873), .A2(n3113), .ZN(n3114) );
  OR2_X1 U3953 ( .A1(n3115), .A2(n3114), .ZN(n3116) );
  NAND2_X1 U3954 ( .A1(n3117), .A2(n3116), .ZN(n3909) );
  OAI22_X1 U3955 ( .A1(n3722), .A2(n3909), .B1(n3125), .B2(n3704), .ZN(n3118)
         );
  AOI21_X1 U3956 ( .B1(n4533), .B2(n3119), .A(n3118), .ZN(n3120) );
  OAI21_X1 U3957 ( .B1(n3121), .B2(n2519), .A(n3120), .ZN(U3229) );
  AOI21_X1 U3958 ( .B1(n3124), .B2(n3123), .A(n3122), .ZN(n3130) );
  OAI22_X1 U3959 ( .A1(n2897), .A2(n3704), .B1(n4343), .B2(n3125), .ZN(n3127)
         );
  NOR2_X1 U3960 ( .A1(n3705), .A2(n3192), .ZN(n3126) );
  AOI211_X1 U3961 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3128), .A(n3127), .B(n3126), 
        .ZN(n3129) );
  OAI21_X1 U3962 ( .B1(n3130), .B2(n3722), .A(n3129), .ZN(U3234) );
  XOR2_X1 U3963 ( .A(n3132), .B(n3131), .Z(n3138) );
  NOR2_X1 U3964 ( .A1(STATE_REG_SCAN_IN), .A2(n3136), .ZN(n4332) );
  AOI21_X1 U3965 ( .B1(n4348), .B2(n3898), .A(n4332), .ZN(n3134) );
  NAND2_X1 U3966 ( .A1(n3714), .A2(n2889), .ZN(n3133) );
  OAI211_X1 U3967 ( .C1(n3705), .C2(n3216), .A(n3134), .B(n3133), .ZN(n3135)
         );
  AOI21_X1 U3968 ( .B1(n3720), .B2(n3136), .A(n3135), .ZN(n3137) );
  OAI21_X1 U3969 ( .B1(n3138), .B2(n3722), .A(n3137), .ZN(U3215) );
  INV_X1 U3970 ( .A(n3140), .ZN(n3739) );
  NAND2_X1 U3971 ( .A1(n3739), .A2(n3751), .ZN(n3798) );
  XNOR2_X1 U3972 ( .A(n3139), .B(n3798), .ZN(n4556) );
  NAND4_X1 U3973 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3145)
         );
  OR2_X1 U3974 ( .A1(n3146), .A2(n3972), .ZN(n3158) );
  AND2_X1 U3975 ( .A1(n3519), .A2(n3158), .ZN(n3147) );
  XNOR2_X1 U3976 ( .A(n3148), .B(n3798), .ZN(n3149) );
  NAND2_X1 U3977 ( .A1(n3149), .A2(n4191), .ZN(n3151) );
  AOI22_X1 U3978 ( .A1(n3896), .A2(n4185), .B1(n4486), .B2(n3153), .ZN(n3150)
         );
  OAI211_X1 U3979 ( .C1(n3152), .C2(n4188), .A(n3151), .B(n3150), .ZN(n4558)
         );
  NAND2_X1 U3980 ( .A1(n4558), .A2(n3979), .ZN(n3157) );
  OR2_X1 U3981 ( .A1(n4507), .A2(n4327), .ZN(n4202) );
  AOI21_X1 U3982 ( .B1(n3153), .B2(n3165), .A(n3231), .ZN(n4559) );
  INV_X1 U3983 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3438) );
  INV_X1 U3984 ( .A(n3154), .ZN(n3271) );
  OAI22_X1 U3985 ( .A1(n3979), .A2(n3438), .B1(n3271), .B2(n4124), .ZN(n3155)
         );
  AOI21_X1 U3986 ( .B1(n4504), .B2(n4559), .A(n3155), .ZN(n3156) );
  OAI211_X1 U3987 ( .C1(n4556), .C2(n4182), .A(n3157), .B(n3156), .ZN(U3285)
         );
  NAND2_X1 U3988 ( .A1(n2867), .A2(n3160), .ZN(n3727) );
  AND2_X1 U3989 ( .A1(n4491), .A2(n3727), .ZN(n4529) );
  OR2_X1 U3990 ( .A1(n4507), .A2(n3158), .ZN(n3527) );
  AOI21_X1 U3991 ( .B1(n2482), .B2(n3972), .A(n4486), .ZN(n3161) );
  AOI21_X1 U3992 ( .B1(n4493), .B2(n3519), .A(n4529), .ZN(n3159) );
  AOI21_X1 U3993 ( .B1(n4185), .B2(n3900), .A(n3159), .ZN(n4530) );
  OAI21_X1 U3994 ( .B1(n3161), .B2(n3160), .A(n4530), .ZN(n3162) );
  AOI22_X1 U3995 ( .A1(n3162), .A2(n3979), .B1(REG3_REG_0__SCAN_IN), .B2(n4499), .ZN(n3164) );
  NAND2_X1 U3996 ( .A1(n4200), .A2(REG2_REG_0__SCAN_IN), .ZN(n3163) );
  OAI211_X1 U3997 ( .C1(n4529), .C2(n3527), .A(n3164), .B(n3163), .ZN(U3290)
         );
  INV_X1 U3998 ( .A(n3218), .ZN(n3166) );
  OAI211_X1 U3999 ( .C1(n3166), .C2(n3180), .A(n4577), .B(n3165), .ZN(n4551)
         );
  NOR2_X1 U4000 ( .A1(n4551), .A2(n4327), .ZN(n3174) );
  XNOR2_X1 U4001 ( .A(n3167), .B(n3823), .ZN(n3175) );
  XOR2_X1 U4002 ( .A(n3823), .B(n3168), .Z(n3172) );
  AOI22_X1 U4003 ( .A1(n3897), .A2(n4185), .B1(n3169), .B2(n4486), .ZN(n3170)
         );
  OAI21_X1 U4004 ( .B1(n2897), .B2(n4188), .A(n3170), .ZN(n3171) );
  AOI21_X1 U4005 ( .B1(n3172), .B2(n4191), .A(n3171), .ZN(n3173) );
  OAI21_X1 U4006 ( .B1(n3519), .B2(n3175), .A(n3173), .ZN(n4552) );
  AOI211_X1 U4007 ( .C1(n4499), .C2(n3186), .A(n3174), .B(n4552), .ZN(n3177)
         );
  INV_X1 U4008 ( .A(n3175), .ZN(n4554) );
  INV_X1 U4009 ( .A(n3527), .ZN(n4503) );
  AOI22_X1 U4010 ( .A1(n4554), .A2(n4503), .B1(REG2_REG_4__SCAN_IN), .B2(n4200), .ZN(n3176) );
  OAI21_X1 U4011 ( .B1(n3177), .B2(n4200), .A(n3176), .ZN(U3286) );
  AND2_X1 U4012 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3932) );
  AOI21_X1 U4013 ( .B1(n4348), .B2(n3897), .A(n3932), .ZN(n3179) );
  NAND2_X1 U4014 ( .A1(n3714), .A2(n3899), .ZN(n3178) );
  OAI211_X1 U4015 ( .C1(n3705), .C2(n3180), .A(n3179), .B(n3178), .ZN(n3185)
         );
  AOI211_X1 U4016 ( .C1(n3181), .C2(n3183), .A(n3722), .B(n3182), .ZN(n3184)
         );
  AOI211_X1 U4017 ( .C1(n3186), .C2(n3720), .A(n3185), .B(n3184), .ZN(n3187)
         );
  INV_X1 U4018 ( .A(n3187), .ZN(U3227) );
  INV_X1 U4019 ( .A(n4502), .ZN(n3188) );
  NOR2_X1 U4020 ( .A1(n3188), .A2(n3192), .ZN(n4541) );
  NOR3_X1 U4021 ( .A1(n4179), .A2(n4540), .A3(n4541), .ZN(n3204) );
  NAND3_X1 U4022 ( .A1(n3792), .A2(n3730), .A3(n4495), .ZN(n3189) );
  NAND2_X1 U4023 ( .A1(n3207), .A2(n3189), .ZN(n3194) );
  INV_X1 U4024 ( .A(n4188), .ZN(n4487) );
  NAND2_X1 U4025 ( .A1(n3900), .A2(n4487), .ZN(n3191) );
  NAND2_X1 U4026 ( .A1(n3899), .A2(n4185), .ZN(n3190) );
  OAI211_X1 U4027 ( .C1(n4107), .C2(n3192), .A(n3191), .B(n3190), .ZN(n3193)
         );
  AOI21_X1 U4028 ( .B1(n3194), .B2(n4191), .A(n3193), .ZN(n3200) );
  NAND2_X1 U4029 ( .A1(n3197), .A2(n3196), .ZN(n3198) );
  NAND2_X1 U4030 ( .A1(n3195), .A2(n3198), .ZN(n4544) );
  INV_X1 U4031 ( .A(n3519), .ZN(n4498) );
  NAND2_X1 U4032 ( .A1(n4544), .A2(n4498), .ZN(n3199) );
  NAND2_X1 U4033 ( .A1(n3200), .A2(n3199), .ZN(n4542) );
  MUX2_X1 U4034 ( .A(REG2_REG_2__SCAN_IN), .B(n4542), .S(n3979), .Z(n3203) );
  INV_X1 U4035 ( .A(n4544), .ZN(n3201) );
  OAI22_X1 U4036 ( .A1(n3527), .A2(n3201), .B1(n2525), .B2(n4124), .ZN(n3202)
         );
  OR3_X1 U4037 ( .A1(n3204), .A2(n3203), .A3(n3202), .ZN(U3288) );
  INV_X1 U4038 ( .A(n3811), .ZN(n3206) );
  XNOR2_X1 U4039 ( .A(n3205), .B(n3206), .ZN(n4548) );
  NAND2_X1 U4040 ( .A1(n4548), .A2(n4498), .ZN(n3215) );
  NAND3_X1 U4041 ( .A1(n3207), .A2(n3731), .A3(n3206), .ZN(n3208) );
  NAND2_X1 U4042 ( .A1(n3209), .A2(n3208), .ZN(n3213) );
  NAND2_X1 U40430 ( .A1(n2889), .A2(n4487), .ZN(n3211) );
  NAND2_X1 U4044 ( .A1(n3898), .A2(n4185), .ZN(n3210) );
  OAI211_X1 U4045 ( .C1(n4107), .C2(n3216), .A(n3211), .B(n3210), .ZN(n3212)
         );
  AOI21_X1 U4046 ( .B1(n3213), .B2(n4191), .A(n3212), .ZN(n3214) );
  AND2_X1 U4047 ( .A1(n3215), .A2(n3214), .ZN(n4550) );
  OR2_X1 U4048 ( .A1(n4540), .A2(n3216), .ZN(n3217) );
  NAND2_X1 U4049 ( .A1(n3218), .A2(n3217), .ZN(n4546) );
  AOI22_X1 U4050 ( .A1(n4507), .A2(REG2_REG_3__SCAN_IN), .B1(n4499), .B2(n3136), .ZN(n3219) );
  OAI21_X1 U4051 ( .B1(n4179), .B2(n4546), .A(n3219), .ZN(n3220) );
  AOI21_X1 U4052 ( .B1(n4503), .B2(n4548), .A(n3220), .ZN(n3221) );
  OAI21_X1 U4053 ( .B1(n4507), .B2(n4550), .A(n3221), .ZN(U3287) );
  NAND2_X1 U4054 ( .A1(n3742), .A2(n3752), .ZN(n3825) );
  XOR2_X1 U4055 ( .A(n3825), .B(n3222), .Z(n3230) );
  XOR2_X1 U4056 ( .A(n3825), .B(n3223), .Z(n3228) );
  AOI22_X1 U4057 ( .A1(n3895), .A2(n4185), .B1(n3224), .B2(n4486), .ZN(n3225)
         );
  OAI21_X1 U4058 ( .B1(n3226), .B2(n4188), .A(n3225), .ZN(n3227) );
  AOI21_X1 U4059 ( .B1(n3228), .B2(n4191), .A(n3227), .ZN(n3229) );
  OAI21_X1 U4060 ( .B1(n3230), .B2(n3519), .A(n3229), .ZN(n4563) );
  INV_X1 U4061 ( .A(n4563), .ZN(n3237) );
  INV_X1 U4062 ( .A(n3230), .ZN(n4565) );
  NOR2_X1 U4063 ( .A1(n3231), .A2(n3257), .ZN(n4562) );
  NOR3_X1 U4064 ( .A1(n4179), .A2(n4561), .A3(n4562), .ZN(n3235) );
  INV_X1 U4065 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3233) );
  OAI22_X1 U4066 ( .A1(n3979), .A2(n3233), .B1(n3232), .B2(n4124), .ZN(n3234)
         );
  AOI211_X1 U4067 ( .C1(n4565), .C2(n4503), .A(n3235), .B(n3234), .ZN(n3236)
         );
  OAI21_X1 U4068 ( .B1(n3237), .B2(n4200), .A(n3236), .ZN(U3284) );
  XOR2_X1 U4069 ( .A(n3790), .B(n3238), .Z(n3239) );
  NAND2_X1 U4070 ( .A1(n3239), .A2(n4191), .ZN(n3241) );
  AOI22_X1 U4071 ( .A1(n3894), .A2(n4185), .B1(n4486), .B2(n3245), .ZN(n3240)
         );
  OAI211_X1 U4072 ( .C1(n3266), .C2(n4188), .A(n3241), .B(n3240), .ZN(n4567)
         );
  INV_X1 U4073 ( .A(n4567), .ZN(n3250) );
  XOR2_X1 U4074 ( .A(n3242), .B(n3790), .Z(n4570) );
  INV_X1 U4075 ( .A(n4561), .ZN(n3244) );
  INV_X1 U4076 ( .A(n3279), .ZN(n3243) );
  AOI211_X1 U4077 ( .C1(n3245), .C2(n3244), .A(n4560), .B(n3243), .ZN(n4568)
         );
  INV_X1 U4078 ( .A(n4568), .ZN(n3247) );
  AOI22_X1 U4079 ( .A1(n4200), .A2(REG2_REG_7__SCAN_IN), .B1(n3300), .B2(n4499), .ZN(n3246) );
  OAI21_X1 U4080 ( .B1(n3247), .B2(n4202), .A(n3246), .ZN(n3248) );
  AOI21_X1 U4081 ( .B1(n4570), .B2(n4204), .A(n3248), .ZN(n3249) );
  OAI21_X1 U4082 ( .B1(n3250), .B2(n4200), .A(n3249), .ZN(U3283) );
  XNOR2_X1 U4083 ( .A(n3252), .B(n3251), .ZN(n3253) );
  XNOR2_X1 U4084 ( .A(n2262), .B(n3253), .ZN(n3261) );
  INV_X1 U4085 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3254) );
  NOR2_X1 U4086 ( .A1(STATE_REG_SCAN_IN), .A2(n3254), .ZN(n4379) );
  AOI21_X1 U4087 ( .B1(n3714), .B2(n3897), .A(n4379), .ZN(n3256) );
  NAND2_X1 U4088 ( .A1(n4348), .A2(n3895), .ZN(n3255) );
  OAI211_X1 U4089 ( .C1(n3705), .C2(n3257), .A(n3256), .B(n3255), .ZN(n3258)
         );
  AOI21_X1 U4090 ( .B1(n3720), .B2(n3259), .A(n3258), .ZN(n3260) );
  OAI21_X1 U4091 ( .B1(n3261), .B2(n3722), .A(n3260), .ZN(U3236) );
  AOI211_X1 U4092 ( .C1(n3264), .C2(n3263), .A(n3722), .B(n3262), .ZN(n3265)
         );
  INV_X1 U4093 ( .A(n3265), .ZN(n3270) );
  AND2_X1 U4094 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4373) );
  OAI22_X1 U4095 ( .A1(n3705), .A2(n3267), .B1(n3266), .B2(n3704), .ZN(n3268)
         );
  AOI211_X1 U4096 ( .C1(n3714), .C2(n3898), .A(n4373), .B(n3268), .ZN(n3269)
         );
  OAI211_X1 U4097 ( .C1(n4358), .C2(n3271), .A(n3270), .B(n3269), .ZN(U3224)
         );
  NAND2_X1 U4098 ( .A1(n3746), .A2(n3753), .ZN(n3821) );
  XNOR2_X1 U4099 ( .A(n3272), .B(n3821), .ZN(n3273) );
  NAND2_X1 U4100 ( .A1(n3273), .A2(n4167), .ZN(n3275) );
  AOI22_X1 U4101 ( .A1(n3893), .A2(n4185), .B1(n3280), .B2(n4486), .ZN(n3274)
         );
  OAI211_X1 U4102 ( .C1(n3276), .C2(n4188), .A(n3275), .B(n3274), .ZN(n3286)
         );
  INV_X1 U4103 ( .A(n3286), .ZN(n3285) );
  XOR2_X1 U4104 ( .A(n3277), .B(n3821), .Z(n3287) );
  INV_X1 U4105 ( .A(n3304), .ZN(n3278) );
  AOI21_X1 U4106 ( .B1(n3280), .B2(n3279), .A(n3278), .ZN(n3291) );
  INV_X1 U4107 ( .A(n3291), .ZN(n3282) );
  AOI22_X1 U4108 ( .A1(n4200), .A2(REG2_REG_8__SCAN_IN), .B1(n3324), .B2(n4499), .ZN(n3281) );
  OAI21_X1 U4109 ( .B1(n3282), .B2(n4179), .A(n3281), .ZN(n3283) );
  AOI21_X1 U4110 ( .B1(n3287), .B2(n4204), .A(n3283), .ZN(n3284) );
  OAI21_X1 U4111 ( .B1(n4507), .B2(n3285), .A(n3284), .ZN(U3282) );
  AOI21_X1 U4112 ( .B1(n3287), .B2(n4569), .A(n3286), .ZN(n3293) );
  INV_X1 U4113 ( .A(n4312), .ZN(n3398) );
  INV_X1 U4114 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3288) );
  NOR2_X1 U4115 ( .A1(n4580), .A2(n3288), .ZN(n3289) );
  AOI21_X1 U4116 ( .B1(n3291), .B2(n3398), .A(n3289), .ZN(n3290) );
  OAI21_X1 U4117 ( .B1(n3293), .B2(n4578), .A(n3290), .ZN(U3483) );
  INV_X1 U4118 ( .A(n4257), .ZN(n3400) );
  AOI22_X1 U4119 ( .A1(n3291), .A2(n3400), .B1(n4593), .B2(REG1_REG_8__SCAN_IN), .ZN(n3292) );
  OAI21_X1 U4120 ( .B1(n3293), .B2(n4593), .A(n3292), .ZN(U3526) );
  XNOR2_X1 U4121 ( .A(n3294), .B(n3295), .ZN(n3302) );
  AND2_X1 U4122 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4394) );
  AOI21_X1 U4123 ( .B1(n4348), .B2(n3894), .A(n4394), .ZN(n3297) );
  NAND2_X1 U4124 ( .A1(n3714), .A2(n3896), .ZN(n3296) );
  OAI211_X1 U4125 ( .C1(n3705), .C2(n3298), .A(n3297), .B(n3296), .ZN(n3299)
         );
  AOI21_X1 U4126 ( .B1(n3720), .B2(n3300), .A(n3299), .ZN(n3301) );
  OAI21_X1 U4127 ( .B1(n3302), .B2(n3722), .A(n3301), .ZN(U3210) );
  INV_X1 U4128 ( .A(n3303), .ZN(n3761) );
  NAND2_X1 U4129 ( .A1(n3761), .A2(n3747), .ZN(n3800) );
  XOR2_X1 U4130 ( .A(n3334), .B(n3800), .Z(n4573) );
  AOI21_X1 U4131 ( .B1(n3309), .B2(n3304), .A(n3336), .ZN(n4576) );
  INV_X1 U4132 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3434) );
  INV_X1 U4133 ( .A(n3356), .ZN(n3305) );
  OAI22_X1 U4134 ( .A1(n3979), .A2(n3434), .B1(n3305), .B2(n4124), .ZN(n3306)
         );
  AOI21_X1 U4135 ( .B1(n4576), .B2(n4504), .A(n3306), .ZN(n3314) );
  XNOR2_X1 U4136 ( .A(n3307), .B(n3800), .ZN(n3308) );
  NAND2_X1 U4137 ( .A1(n3308), .A2(n4191), .ZN(n3311) );
  AOI22_X1 U4138 ( .A1(n3892), .A2(n4185), .B1(n4486), .B2(n3309), .ZN(n3310)
         );
  OAI211_X1 U4139 ( .C1(n3312), .C2(n4188), .A(n3311), .B(n3310), .ZN(n4575)
         );
  NAND2_X1 U4140 ( .A1(n4575), .A2(n3979), .ZN(n3313) );
  OAI211_X1 U4141 ( .C1(n4573), .C2(n4182), .A(n3314), .B(n3313), .ZN(U3281)
         );
  NAND2_X1 U4142 ( .A1(n2467), .A2(n3317), .ZN(n3318) );
  XNOR2_X1 U4143 ( .A(n3315), .B(n3318), .ZN(n3326) );
  INV_X1 U4144 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3319) );
  NOR2_X1 U4145 ( .A1(STATE_REG_SCAN_IN), .A2(n3319), .ZN(n4406) );
  AOI21_X1 U4146 ( .B1(n4348), .B2(n3893), .A(n4406), .ZN(n3321) );
  NAND2_X1 U4147 ( .A1(n3714), .A2(n3895), .ZN(n3320) );
  OAI211_X1 U4148 ( .C1(n3705), .C2(n3322), .A(n3321), .B(n3320), .ZN(n3323)
         );
  AOI21_X1 U4149 ( .B1(n3720), .B2(n3324), .A(n3323), .ZN(n3325) );
  OAI21_X1 U4150 ( .B1(n3326), .B2(n3722), .A(n3325), .ZN(U3218) );
  NAND2_X1 U4151 ( .A1(n3759), .A2(n3765), .ZN(n3796) );
  XOR2_X1 U4152 ( .A(n3796), .B(n3327), .Z(n3331) );
  AOI22_X1 U4153 ( .A1(n3891), .A2(n4185), .B1(n4486), .B2(n3328), .ZN(n3329)
         );
  OAI21_X1 U4154 ( .B1(n3332), .B2(n4188), .A(n3329), .ZN(n3330) );
  AOI21_X1 U4155 ( .B1(n3331), .B2(n4191), .A(n3330), .ZN(n3342) );
  OAI22_X1 U4156 ( .A1(n3334), .A2(n3333), .B1(n3332), .B2(n3354), .ZN(n3335)
         );
  XNOR2_X1 U4157 ( .A(n3335), .B(n3796), .ZN(n3343) );
  INV_X1 U4158 ( .A(n3343), .ZN(n3340) );
  NOR2_X1 U4159 ( .A1(n3336), .A2(n3423), .ZN(n3337) );
  OR2_X1 U4160 ( .A1(n3367), .A2(n3337), .ZN(n3346) );
  AOI22_X1 U4161 ( .A1(n4507), .A2(REG2_REG_10__SCAN_IN), .B1(n3430), .B2(
        n4499), .ZN(n3338) );
  OAI21_X1 U4162 ( .B1(n3346), .B2(n4179), .A(n3338), .ZN(n3339) );
  AOI21_X1 U4163 ( .B1(n3340), .B2(n4204), .A(n3339), .ZN(n3341) );
  OAI21_X1 U4164 ( .B1(n3342), .B2(n4200), .A(n3341), .ZN(U3280) );
  OAI21_X1 U4165 ( .B1(n4572), .B2(n3343), .A(n3342), .ZN(n3348) );
  INV_X1 U4166 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4836) );
  OAI22_X1 U4167 ( .A1(n3346), .A2(n4257), .B1(n4595), .B2(n4836), .ZN(n3344)
         );
  AOI21_X1 U4168 ( .B1(n3348), .B2(n4595), .A(n3344), .ZN(n3345) );
  INV_X1 U4169 ( .A(n3345), .ZN(U3528) );
  INV_X1 U4170 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4853) );
  OAI22_X1 U4171 ( .A1(n3346), .A2(n4312), .B1(n4580), .B2(n4853), .ZN(n3347)
         );
  AOI21_X1 U4172 ( .B1(n3348), .B2(n4580), .A(n3347), .ZN(n3349) );
  INV_X1 U4173 ( .A(n3349), .ZN(U3487) );
  XOR2_X1 U4174 ( .A(n3351), .B(n3350), .Z(n3358) );
  AND2_X1 U4175 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4414) );
  AOI21_X1 U4176 ( .B1(n4348), .B2(n3892), .A(n4414), .ZN(n3353) );
  NAND2_X1 U4177 ( .A1(n3714), .A2(n3894), .ZN(n3352) );
  OAI211_X1 U4178 ( .C1(n3705), .C2(n3354), .A(n3353), .B(n3352), .ZN(n3355)
         );
  AOI21_X1 U4179 ( .B1(n3720), .B2(n3356), .A(n3355), .ZN(n3357) );
  OAI21_X1 U4180 ( .B1(n3358), .B2(n3722), .A(n3357), .ZN(U3228) );
  XNOR2_X1 U4181 ( .A(n3359), .B(n3799), .ZN(n4277) );
  XOR2_X1 U4182 ( .A(n3360), .B(n3799), .Z(n3361) );
  NAND2_X1 U4183 ( .A1(n3361), .A2(n4167), .ZN(n3364) );
  AOI22_X1 U4184 ( .A1(n3508), .A2(n4185), .B1(n4486), .B2(n3362), .ZN(n3363)
         );
  OAI211_X1 U4185 ( .C1(n3365), .C2(n4188), .A(n3364), .B(n3363), .ZN(n3366)
         );
  AOI21_X1 U4186 ( .B1(n4498), .B2(n4277), .A(n3366), .ZN(n4279) );
  OAI21_X1 U4187 ( .B1(n3367), .B2(n3391), .A(n3376), .ZN(n4280) );
  AOI22_X1 U4188 ( .A1(n4200), .A2(REG2_REG_11__SCAN_IN), .B1(n3393), .B2(
        n4499), .ZN(n3368) );
  OAI21_X1 U4189 ( .B1(n4280), .B2(n4179), .A(n3368), .ZN(n3369) );
  AOI21_X1 U4190 ( .B1(n4277), .B2(n4503), .A(n3369), .ZN(n3370) );
  OAI21_X1 U4191 ( .B1(n4279), .B2(n4200), .A(n3370), .ZN(U3279) );
  OR2_X1 U4192 ( .A1(n2394), .A2(n3768), .ZN(n3797) );
  XOR2_X1 U4193 ( .A(n3797), .B(n3371), .Z(n3372) );
  NAND2_X1 U4194 ( .A1(n3372), .A2(n4167), .ZN(n3374) );
  AOI22_X1 U4195 ( .A1(n3890), .A2(n4185), .B1(n4486), .B2(n3377), .ZN(n3373)
         );
  OAI211_X1 U4196 ( .C1(n3497), .C2(n4188), .A(n3374), .B(n3373), .ZN(n3396)
         );
  INV_X1 U4197 ( .A(n3396), .ZN(n3384) );
  INV_X1 U4198 ( .A(n3375), .ZN(n3415) );
  AOI21_X1 U4199 ( .B1(n3377), .B2(n3376), .A(n3415), .ZN(n3401) );
  INV_X1 U4200 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3379) );
  INV_X1 U4201 ( .A(n3378), .ZN(n3502) );
  OAI22_X1 U4202 ( .A1(n3979), .A2(n3379), .B1(n3502), .B2(n4124), .ZN(n3380)
         );
  AOI21_X1 U4203 ( .B1(n3401), .B2(n4504), .A(n3380), .ZN(n3383) );
  XOR2_X1 U4204 ( .A(n3381), .B(n3797), .Z(n3397) );
  NAND2_X1 U4205 ( .A1(n3397), .A2(n4204), .ZN(n3382) );
  OAI211_X1 U4206 ( .C1(n3384), .C2(n4507), .A(n3383), .B(n3382), .ZN(U3278)
         );
  XNOR2_X1 U4207 ( .A(n3387), .B(n3386), .ZN(n3388) );
  XNOR2_X1 U4208 ( .A(n3385), .B(n3388), .ZN(n3395) );
  NOR2_X1 U4209 ( .A1(STATE_REG_SCAN_IN), .A2(n4918), .ZN(n4432) );
  AOI21_X1 U4210 ( .B1(n3714), .B2(n3892), .A(n4432), .ZN(n3390) );
  NAND2_X1 U4211 ( .A1(n4348), .A2(n3508), .ZN(n3389) );
  OAI211_X1 U4212 ( .C1(n3705), .C2(n3391), .A(n3390), .B(n3389), .ZN(n3392)
         );
  AOI21_X1 U4213 ( .B1(n3720), .B2(n3393), .A(n3392), .ZN(n3394) );
  OAI21_X1 U4214 ( .B1(n3395), .B2(n3722), .A(n3394), .ZN(U3233) );
  AOI21_X1 U4215 ( .B1(n3397), .B2(n4569), .A(n3396), .ZN(n3403) );
  AOI22_X1 U4216 ( .A1(n3401), .A2(n3398), .B1(REG0_REG_12__SCAN_IN), .B2(
        n4578), .ZN(n3399) );
  OAI21_X1 U4217 ( .B1(n3403), .B2(n4578), .A(n3399), .ZN(U3491) );
  AOI22_X1 U4218 ( .A1(n3401), .A2(n3400), .B1(REG1_REG_12__SCAN_IN), .B2(
        n4593), .ZN(n3402) );
  OAI21_X1 U4219 ( .B1(n3403), .B2(n4593), .A(n3402), .ZN(U3530) );
  INV_X1 U4220 ( .A(n3404), .ZN(n3764) );
  NAND2_X1 U4221 ( .A1(n3764), .A2(n3772), .ZN(n3801) );
  XNOR2_X1 U4222 ( .A(n3405), .B(n3801), .ZN(n3413) );
  XNOR2_X1 U4223 ( .A(n3406), .B(n3801), .ZN(n3411) );
  AOI22_X1 U4224 ( .A1(n3889), .A2(n4185), .B1(n4486), .B2(n3407), .ZN(n3408)
         );
  OAI21_X1 U4225 ( .B1(n3409), .B2(n4188), .A(n3408), .ZN(n3410) );
  AOI21_X1 U4226 ( .B1(n3411), .B2(n4167), .A(n3410), .ZN(n3412) );
  OAI21_X1 U4227 ( .B1(n3413), .B2(n3519), .A(n3412), .ZN(n3482) );
  INV_X1 U4228 ( .A(n3482), .ZN(n3419) );
  INV_X1 U4229 ( .A(n3413), .ZN(n3483) );
  INV_X1 U4230 ( .A(n3414), .ZN(n3524) );
  OAI21_X1 U4231 ( .B1(n3415), .B2(n3511), .A(n3524), .ZN(n3489) );
  AOI22_X1 U4232 ( .A1(n4200), .A2(REG2_REG_13__SCAN_IN), .B1(n3513), .B2(
        n4499), .ZN(n3416) );
  OAI21_X1 U4233 ( .B1(n3489), .B2(n4179), .A(n3416), .ZN(n3417) );
  AOI21_X1 U4234 ( .B1(n3483), .B2(n4503), .A(n3417), .ZN(n3418) );
  OAI21_X1 U4235 ( .B1(n3419), .B2(n4507), .A(n3418), .ZN(U3277) );
  NOR2_X1 U4236 ( .A1(STATE_REG_SCAN_IN), .A2(n3420), .ZN(n4422) );
  AOI21_X1 U4237 ( .B1(n3714), .B2(n3893), .A(n4422), .ZN(n3422) );
  NAND2_X1 U4238 ( .A1(n4348), .A2(n3891), .ZN(n3421) );
  OAI211_X1 U4239 ( .C1(n3705), .C2(n3423), .A(n3422), .B(n3421), .ZN(n3429)
         );
  INV_X1 U4240 ( .A(n3424), .ZN(n3425) );
  AOI211_X1 U4241 ( .C1(n3427), .C2(n3426), .A(n3722), .B(n3425), .ZN(n3428)
         );
  AOI211_X1 U4242 ( .C1(n3430), .C2(n3720), .A(n3429), .B(n3428), .ZN(n3431)
         );
  INV_X1 U4243 ( .A(n3431), .ZN(U3214) );
  NAND2_X1 U4244 ( .A1(n3433), .A2(n3432), .ZN(n4367) );
  INV_X1 U4245 ( .A(n4328), .ZN(n3481) );
  INV_X1 U4246 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4917) );
  INV_X1 U4247 ( .A(n3472), .ZN(n4520) );
  AOI22_X1 U4248 ( .A1(n3472), .A2(REG2_REG_11__SCAN_IN), .B1(n4917), .B2(
        n4520), .ZN(n4435) );
  NAND2_X1 U4249 ( .A1(n3466), .A2(REG2_REG_9__SCAN_IN), .ZN(n3444) );
  INV_X1 U4250 ( .A(n3466), .ZN(n4522) );
  AOI22_X1 U4251 ( .A1(n3466), .A2(REG2_REG_9__SCAN_IN), .B1(n3434), .B2(n4522), .ZN(n4417) );
  NAND2_X1 U4252 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4524), .ZN(n3441) );
  INV_X1 U4253 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4880) );
  AOI22_X1 U4254 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4524), .B1(n4401), .B2(n4880), .ZN(n4398) );
  AOI22_X1 U4255 ( .A1(n3453), .A2(REG2_REG_5__SCAN_IN), .B1(n3438), .B2(n4526), .ZN(n4370) );
  INV_X1 U4256 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4773) );
  INV_X1 U4257 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3435) );
  NAND3_X1 U4258 ( .A1(n3904), .A2(REG2_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n3919) );
  AOI21_X1 U4259 ( .B1(n3919), .B2(n3918), .A(n3920), .ZN(n3917) );
  INV_X1 U4260 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3437) );
  INV_X1 U4261 ( .A(n4330), .ZN(n3457) );
  NAND2_X1 U4262 ( .A1(n3439), .A2(n4329), .ZN(n3440) );
  INV_X1 U4263 ( .A(n4329), .ZN(n4381) );
  XNOR2_X1 U4264 ( .A(n3439), .B(n4381), .ZN(n4386) );
  NAND2_X1 U4265 ( .A1(n3463), .A2(n3442), .ZN(n3443) );
  XNOR2_X1 U4266 ( .A(n3442), .B(n2404), .ZN(n4408) );
  NAND2_X1 U4267 ( .A1(n3468), .A2(n3445), .ZN(n3446) );
  XNOR2_X1 U4268 ( .A(n3445), .B(n3469), .ZN(n4425) );
  NAND2_X1 U4269 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4425), .ZN(n4424) );
  NAND2_X1 U4270 ( .A1(n3446), .A2(n4424), .ZN(n4434) );
  NAND2_X1 U4271 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  NAND2_X1 U4272 ( .A1(n3474), .A2(n3447), .ZN(n3448) );
  INV_X1 U4273 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4842) );
  AND2_X1 U4274 ( .A1(n4328), .A2(REG2_REG_13__SCAN_IN), .ZN(n3951) );
  AOI21_X1 U4275 ( .B1(n4842), .B2(n3481), .A(n3951), .ZN(n3452) );
  AND2_X1 U4276 ( .A1(n3450), .A2(n3449), .ZN(n4322) );
  NAND2_X1 U4277 ( .A1(n4321), .A2(n4322), .ZN(n3910) );
  OR2_X1 U4278 ( .A1(n4367), .A2(n3910), .ZN(n4450) );
  AOI21_X1 U4279 ( .B1(n3452), .B2(n3952), .A(n4450), .ZN(n3451) );
  OAI21_X1 U4280 ( .B1(n3952), .B2(n3452), .A(n3451), .ZN(n3480) );
  NOR2_X1 U4281 ( .A1(STATE_REG_SCAN_IN), .A2(n4718), .ZN(n3507) );
  INV_X1 U4282 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4837) );
  NOR2_X1 U4283 ( .A1(n4837), .A2(n4401), .ZN(n4390) );
  INV_X1 U4284 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4890) );
  AOI22_X1 U4285 ( .A1(n3453), .A2(REG1_REG_5__SCAN_IN), .B1(n4890), .B2(n4526), .ZN(n4376) );
  INV_X1 U4286 ( .A(n3902), .ZN(n3454) );
  INV_X1 U4287 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U4288 ( .A1(REG1_REG_3__SCAN_IN), .A2(n4334), .ZN(n4333) );
  NAND2_X1 U4289 ( .A1(n4333), .A2(n2484), .ZN(n3456) );
  INV_X1 U4290 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3459) );
  INV_X1 U4291 ( .A(n3456), .ZN(n3458) );
  NAND2_X1 U4292 ( .A1(n3460), .A2(n4329), .ZN(n3461) );
  XNOR2_X1 U4293 ( .A(n3460), .B(n4381), .ZN(n4384) );
  NAND2_X1 U4294 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4384), .ZN(n4383) );
  NOR2_X1 U4295 ( .A1(n2404), .A2(n3462), .ZN(n3464) );
  INV_X1 U4296 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U4297 ( .A1(n3466), .A2(REG1_REG_9__SCAN_IN), .ZN(n3465) );
  OAI21_X1 U4298 ( .B1(n3466), .B2(REG1_REG_9__SCAN_IN), .A(n3465), .ZN(n4412)
         );
  INV_X1 U4299 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4300 ( .A1(n3472), .A2(n3471), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4520), .ZN(n4429) );
  NOR2_X1 U4301 ( .A1(n4430), .A2(n4429), .ZN(n4428) );
  INV_X1 U4302 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4440) );
  NAND2_X1 U4303 ( .A1(n4328), .A2(REG1_REG_13__SCAN_IN), .ZN(n3942) );
  OAI21_X1 U4304 ( .B1(n4328), .B2(REG1_REG_13__SCAN_IN), .A(n3942), .ZN(n3476) );
  INV_X1 U4305 ( .A(n3943), .ZN(n3475) );
  AOI211_X1 U4306 ( .C1(n3477), .C2(n3476), .A(n3475), .B(n4975), .ZN(n3478)
         );
  AOI211_X1 U4307 ( .C1(n4980), .C2(ADDR_REG_13__SCAN_IN), .A(n3507), .B(n3478), .ZN(n3479) );
  OAI211_X1 U4308 ( .C1(n4989), .C2(n3481), .A(n3480), .B(n3479), .ZN(U3253)
         );
  INV_X1 U4309 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3484) );
  INV_X1 U4310 ( .A(n4528), .ZN(n4566) );
  AOI21_X1 U4311 ( .B1(n4566), .B2(n3483), .A(n3482), .ZN(n3486) );
  MUX2_X1 U4312 ( .A(n3484), .B(n3486), .S(n4595), .Z(n3485) );
  OAI21_X1 U4313 ( .B1(n4257), .B2(n3489), .A(n3485), .ZN(U3531) );
  INV_X1 U4314 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3487) );
  MUX2_X1 U4315 ( .A(n3487), .B(n3486), .S(n4580), .Z(n3488) );
  OAI21_X1 U4316 ( .B1(n3489), .B2(n4312), .A(n3488), .ZN(U3493) );
  INV_X1 U4317 ( .A(n3490), .ZN(n3492) );
  NAND2_X1 U4318 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  XNOR2_X1 U4319 ( .A(n3494), .B(n3493), .ZN(n3495) );
  NAND2_X1 U4320 ( .A1(n3495), .A2(n4353), .ZN(n3501) );
  OAI22_X1 U4321 ( .A1(n3705), .A2(n3496), .B1(n3550), .B2(n3704), .ZN(n3499)
         );
  NAND2_X1 U4322 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4441) );
  OAI21_X1 U4323 ( .B1(n4343), .B2(n3497), .A(n4441), .ZN(n3498) );
  NOR2_X1 U4324 ( .A1(n3499), .A2(n3498), .ZN(n3500) );
  OAI211_X1 U4325 ( .C1(n4358), .C2(n3502), .A(n3501), .B(n3500), .ZN(U3221)
         );
  XNOR2_X1 U4326 ( .A(n3504), .B(n3503), .ZN(n3505) );
  XNOR2_X1 U4327 ( .A(n3506), .B(n3505), .ZN(n3515) );
  AOI21_X1 U4328 ( .B1(n3714), .B2(n3508), .A(n3507), .ZN(n3510) );
  NAND2_X1 U4329 ( .A1(n4348), .A2(n3889), .ZN(n3509) );
  OAI211_X1 U4330 ( .C1(n3705), .C2(n3511), .A(n3510), .B(n3509), .ZN(n3512)
         );
  AOI21_X1 U4331 ( .B1(n3720), .B2(n3513), .A(n3512), .ZN(n3514) );
  OAI21_X1 U4332 ( .B1(n3515), .B2(n3722), .A(n3514), .ZN(U3231) );
  OAI21_X1 U4333 ( .B1(n3824), .B2(n3840), .A(n3531), .ZN(n3522) );
  AOI22_X1 U4334 ( .A1(n3888), .A2(n4185), .B1(n4486), .B2(n3523), .ZN(n3516)
         );
  OAI21_X1 U4335 ( .B1(n3550), .B2(n4188), .A(n3516), .ZN(n3521) );
  AOI21_X1 U4336 ( .B1(n3518), .B2(n3824), .A(n3517), .ZN(n4276) );
  NOR2_X1 U4337 ( .A1(n4276), .A2(n3519), .ZN(n3520) );
  AOI211_X1 U4338 ( .C1(n4191), .C2(n3522), .A(n3521), .B(n3520), .ZN(n4275)
         );
  AOI22_X1 U4339 ( .A1(n4200), .A2(REG2_REG_14__SCAN_IN), .B1(n3544), .B2(
        n4499), .ZN(n3526) );
  NAND2_X1 U4340 ( .A1(n3524), .A2(n3523), .ZN(n4273) );
  NAND3_X1 U4341 ( .A1(n4273), .A2(n4504), .A3(n4272), .ZN(n3525) );
  OAI211_X1 U4342 ( .C1(n4276), .C2(n3527), .A(n3526), .B(n3525), .ZN(n3528)
         );
  INV_X1 U4343 ( .A(n3528), .ZN(n3529) );
  OAI21_X1 U4344 ( .B1(n4275), .B2(n4507), .A(n3529), .ZN(U3276) );
  NAND2_X1 U4345 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  XOR2_X1 U4346 ( .A(n3791), .B(n3532), .Z(n3533) );
  NAND2_X1 U4347 ( .A1(n3533), .A2(n4167), .ZN(n3536) );
  AOI22_X1 U4348 ( .A1(n3713), .A2(n4185), .B1(n4486), .B2(n3534), .ZN(n3535)
         );
  OAI211_X1 U4349 ( .C1(n3537), .C2(n4188), .A(n3536), .B(n3535), .ZN(n3581)
         );
  INV_X1 U4350 ( .A(n3581), .ZN(n3543) );
  XOR2_X1 U4351 ( .A(n3538), .B(n3791), .Z(n3582) );
  INV_X1 U4352 ( .A(n4272), .ZN(n3539) );
  OAI21_X1 U4353 ( .B1(n3539), .B2(n3717), .A(n3576), .ZN(n3587) );
  AOI22_X1 U4354 ( .A1(n4200), .A2(REG2_REG_15__SCAN_IN), .B1(n3719), .B2(
        n4499), .ZN(n3540) );
  OAI21_X1 U4355 ( .B1(n3587), .B2(n4179), .A(n3540), .ZN(n3541) );
  AOI21_X1 U4356 ( .B1(n3582), .B2(n4204), .A(n3541), .ZN(n3542) );
  OAI21_X1 U4357 ( .B1(n4200), .B2(n3543), .A(n3542), .ZN(U3275) );
  INV_X1 U4358 ( .A(n3544), .ZN(n3556) );
  NAND2_X1 U4359 ( .A1(n3546), .A2(n3545), .ZN(n3548) );
  XOR2_X1 U4360 ( .A(n3548), .B(n3547), .Z(n3549) );
  NAND2_X1 U4361 ( .A1(n3549), .A2(n4353), .ZN(n3555) );
  OAI22_X1 U4362 ( .A1(n3705), .A2(n3551), .B1(n3550), .B2(n4343), .ZN(n3553)
         );
  NAND2_X1 U4363 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4457) );
  OAI21_X1 U4364 ( .B1(n3704), .B2(n4344), .A(n4457), .ZN(n3552) );
  NOR2_X1 U4365 ( .A1(n3553), .A2(n3552), .ZN(n3554) );
  OAI211_X1 U4366 ( .C1(n4358), .C2(n3556), .A(n3555), .B(n3554), .ZN(U3212)
         );
  INV_X1 U4367 ( .A(n3780), .ZN(n3847) );
  NAND2_X1 U4368 ( .A1(n3847), .A2(n4138), .ZN(n3822) );
  XNOR2_X1 U4369 ( .A(n3557), .B(n3822), .ZN(n4266) );
  XNOR2_X1 U4370 ( .A(n3558), .B(n3822), .ZN(n3562) );
  AOI22_X1 U4371 ( .A1(n4170), .A2(n4185), .B1(n4486), .B2(n3563), .ZN(n3559)
         );
  OAI21_X1 U4372 ( .B1(n3560), .B2(n4188), .A(n3559), .ZN(n3561) );
  AOI21_X1 U4373 ( .B1(n3562), .B2(n4191), .A(n3561), .ZN(n4265) );
  AOI22_X1 U4374 ( .A1(n4200), .A2(REG2_REG_17__SCAN_IN), .B1(n3652), .B2(
        n4499), .ZN(n3565) );
  INV_X1 U4375 ( .A(n4197), .ZN(n4263) );
  NAND2_X1 U4376 ( .A1(n4268), .A2(n3563), .ZN(n4262) );
  NAND3_X1 U4377 ( .A1(n4263), .A2(n4504), .A3(n4262), .ZN(n3564) );
  OAI211_X1 U4378 ( .C1(n4265), .C2(n4507), .A(n3565), .B(n3564), .ZN(n3566)
         );
  INV_X1 U4379 ( .A(n3566), .ZN(n3567) );
  OAI21_X1 U4380 ( .B1(n4266), .B2(n4182), .A(n3567), .ZN(U3273) );
  XNOR2_X1 U4381 ( .A(n3568), .B(n3826), .ZN(n3571) );
  AOI22_X1 U4382 ( .A1(n4347), .A2(n4185), .B1(n4486), .B2(n3575), .ZN(n3569)
         );
  OAI21_X1 U4383 ( .B1(n4344), .B2(n4188), .A(n3569), .ZN(n3570) );
  AOI21_X1 U4384 ( .B1(n3571), .B2(n4191), .A(n3570), .ZN(n4270) );
  OAI21_X1 U4385 ( .B1(n3573), .B2(n3826), .A(n3572), .ZN(n4271) );
  AOI22_X1 U4386 ( .A1(n4200), .A2(REG2_REG_16__SCAN_IN), .B1(n3574), .B2(
        n4499), .ZN(n3578) );
  NAND2_X1 U4387 ( .A1(n3576), .A2(n3575), .ZN(n4267) );
  NAND3_X1 U4388 ( .A1(n4268), .A2(n4504), .A3(n4267), .ZN(n3577) );
  OAI211_X1 U4389 ( .C1(n4271), .C2(n4182), .A(n3578), .B(n3577), .ZN(n3579)
         );
  INV_X1 U4390 ( .A(n3579), .ZN(n3580) );
  OAI21_X1 U4391 ( .B1(n4200), .B2(n4270), .A(n3580), .ZN(U3274) );
  INV_X1 U4392 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4855) );
  AOI21_X1 U4393 ( .B1(n3582), .B2(n4569), .A(n3581), .ZN(n3584) );
  MUX2_X1 U4394 ( .A(n4855), .B(n3584), .S(n4595), .Z(n3583) );
  OAI21_X1 U4395 ( .B1(n4257), .B2(n3587), .A(n3583), .ZN(U3533) );
  INV_X1 U4396 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3585) );
  MUX2_X1 U4397 ( .A(n3585), .B(n3584), .S(n4580), .Z(n3586) );
  OAI21_X1 U4398 ( .B1(n3587), .B2(n4312), .A(n3586), .ZN(U3497) );
  NAND3_X1 U4399 ( .A1(n3588), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3590) );
  INV_X1 U4400 ( .A(DATAI_31_), .ZN(n3589) );
  OAI22_X1 U4401 ( .A1(n2501), .A2(n3590), .B1(STATE_REG_SCAN_IN), .B2(n3589), 
        .ZN(U3321) );
  XNOR2_X1 U4402 ( .A(n3592), .B(n3591), .ZN(n3598) );
  OAI22_X1 U4403 ( .A1(n3593), .A2(n4343), .B1(n3705), .B2(n4023), .ZN(n3596)
         );
  INV_X1 U4404 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3594) );
  OAI22_X1 U4405 ( .A1(n4019), .A2(n3704), .B1(STATE_REG_SCAN_IN), .B2(n3594), 
        .ZN(n3595) );
  AOI211_X1 U4406 ( .C1(n4024), .C2(n3720), .A(n3596), .B(n3595), .ZN(n3597)
         );
  OAI21_X1 U4407 ( .B1(n3598), .B2(n3722), .A(n3597), .ZN(U3211) );
  INV_X1 U4408 ( .A(n4098), .ZN(n3609) );
  OAI21_X1 U4409 ( .B1(n3678), .B2(n3601), .A(n3600), .ZN(n3603) );
  NAND3_X1 U4410 ( .A1(n3603), .A2(n3602), .A3(n4353), .ZN(n3608) );
  OAI22_X1 U4411 ( .A1(n3705), .A2(n4097), .B1(n4095), .B2(n3704), .ZN(n3606)
         );
  INV_X1 U4412 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3604) );
  OAI22_X1 U4413 ( .A1(n4343), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n3604), 
        .ZN(n3605) );
  NOR2_X1 U4414 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  OAI211_X1 U4415 ( .C1(n4358), .C2(n3609), .A(n3608), .B(n3607), .ZN(U3213)
         );
  INV_X1 U4416 ( .A(n4177), .ZN(n3618) );
  XNOR2_X1 U4417 ( .A(n3610), .B(n3611), .ZN(n3612) );
  NAND2_X1 U4418 ( .A1(n3612), .A2(n4353), .ZN(n3617) );
  OAI22_X1 U4419 ( .A1(n3705), .A2(n4175), .B1(n3613), .B2(n4343), .ZN(n3615)
         );
  NAND2_X1 U4420 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3971) );
  OAI21_X1 U4421 ( .B1(n3704), .B2(n4173), .A(n3971), .ZN(n3614) );
  NOR2_X1 U4422 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  OAI211_X1 U4423 ( .C1(n4358), .C2(n3618), .A(n3617), .B(n3616), .ZN(U3216)
         );
  XOR2_X1 U4424 ( .A(n3620), .B(n3619), .Z(n3621) );
  XNOR2_X1 U4425 ( .A(n3622), .B(n3621), .ZN(n3623) );
  NAND2_X1 U4426 ( .A1(n3623), .A2(n4353), .ZN(n3630) );
  OAI22_X1 U4427 ( .A1(n3705), .A2(n3624), .B1(n4173), .B2(n4343), .ZN(n3628)
         );
  INV_X1 U4428 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3625) );
  OAI22_X1 U4429 ( .A1(n3704), .A2(n3626), .B1(STATE_REG_SCAN_IN), .B2(n3625), 
        .ZN(n3627) );
  NOR2_X1 U4430 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  OAI211_X1 U4431 ( .C1(n4358), .C2(n4125), .A(n3630), .B(n3629), .ZN(U3220)
         );
  INV_X1 U4432 ( .A(n4059), .ZN(n3643) );
  INV_X1 U4433 ( .A(n3632), .ZN(n3634) );
  NAND2_X1 U4434 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  XNOR2_X1 U4435 ( .A(n3631), .B(n3635), .ZN(n3636) );
  NAND2_X1 U4436 ( .A1(n3636), .A2(n4353), .ZN(n3642) );
  NAND2_X1 U4437 ( .A1(n4055), .A2(n4348), .ZN(n3637) );
  OAI21_X1 U4438 ( .B1(STATE_REG_SCAN_IN), .B2(n3638), .A(n3637), .ZN(n3640)
         );
  OAI22_X1 U4439 ( .A1(n3705), .A2(n4053), .B1(n4095), .B2(n4343), .ZN(n3639)
         );
  NOR2_X1 U4440 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  OAI211_X1 U4441 ( .C1(n4358), .C2(n3643), .A(n3642), .B(n3641), .ZN(U3222)
         );
  NAND2_X1 U4442 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  XNOR2_X1 U4443 ( .A(n3644), .B(n3647), .ZN(n3654) );
  AND2_X1 U4444 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4471) );
  AOI21_X1 U4445 ( .B1(n3714), .B2(n3713), .A(n4471), .ZN(n3649) );
  NAND2_X1 U4446 ( .A1(n4348), .A2(n4170), .ZN(n3648) );
  OAI211_X1 U4447 ( .C1(n3650), .C2(n3705), .A(n3649), .B(n3648), .ZN(n3651)
         );
  AOI21_X1 U4448 ( .B1(n3720), .B2(n3652), .A(n3651), .ZN(n3653) );
  OAI21_X1 U4449 ( .B1(n3654), .B2(n3722), .A(n3653), .ZN(U3225) );
  NAND2_X1 U4450 ( .A1(n3655), .A2(n3656), .ZN(n3658) );
  XNOR2_X1 U4451 ( .A(n3658), .B(n3657), .ZN(n3659) );
  NAND2_X1 U4452 ( .A1(n3659), .A2(n4353), .ZN(n3664) );
  OAI22_X1 U4453 ( .A1(n3705), .A2(n4076), .B1(n4074), .B2(n3704), .ZN(n3662)
         );
  OAI22_X1 U4454 ( .A1(n4343), .A2(n4106), .B1(STATE_REG_SCAN_IN), .B2(n3660), 
        .ZN(n3661) );
  NOR2_X1 U4455 ( .A1(n3662), .A2(n3661), .ZN(n3663) );
  OAI211_X1 U4456 ( .C1(n4358), .C2(n4078), .A(n3664), .B(n3663), .ZN(U3226)
         );
  INV_X1 U4457 ( .A(n4155), .ZN(n3676) );
  NOR2_X1 U4458 ( .A1(n3665), .A2(n2448), .ZN(n3670) );
  AOI21_X1 U4459 ( .B1(n3668), .B2(n3667), .A(n3666), .ZN(n3669) );
  OAI21_X1 U4460 ( .B1(n3670), .B2(n3669), .A(n4353), .ZN(n3675) );
  OAI22_X1 U4461 ( .A1(n3705), .A2(n4153), .B1(n4151), .B2(n4343), .ZN(n3673)
         );
  INV_X1 U4462 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3671) );
  OAI22_X1 U4463 ( .A1(n3704), .A2(n4108), .B1(STATE_REG_SCAN_IN), .B2(n3671), 
        .ZN(n3672) );
  NOR2_X1 U4464 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  OAI211_X1 U4465 ( .C1(n4358), .C2(n3676), .A(n3675), .B(n3674), .ZN(U3230)
         );
  AOI21_X1 U4466 ( .B1(n3679), .B2(n3677), .A(n3678), .ZN(n3684) );
  INV_X1 U4467 ( .A(n3680), .ZN(n4112) );
  INV_X1 U4468 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4877) );
  OAI22_X1 U4469 ( .A1(n4343), .A2(n4108), .B1(STATE_REG_SCAN_IN), .B2(n4877), 
        .ZN(n3682) );
  OAI22_X1 U4470 ( .A1(n3705), .A2(n4114), .B1(n4106), .B2(n3704), .ZN(n3681)
         );
  AOI211_X1 U4471 ( .C1(n3720), .C2(n4112), .A(n3682), .B(n3681), .ZN(n3683)
         );
  OAI21_X1 U4472 ( .B1(n3684), .B2(n3722), .A(n3683), .ZN(U3232) );
  INV_X1 U4473 ( .A(n3685), .ZN(n3690) );
  AOI21_X1 U4474 ( .B1(n3689), .B2(n3687), .A(n3686), .ZN(n3688) );
  AOI21_X1 U4475 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n3696) );
  AND2_X1 U4476 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3962) );
  AOI21_X1 U4477 ( .B1(n4348), .B2(n4186), .A(n3962), .ZN(n3692) );
  NAND2_X1 U4478 ( .A1(n3714), .A2(n4347), .ZN(n3691) );
  OAI211_X1 U4479 ( .C1(n3705), .C2(n3693), .A(n3692), .B(n3691), .ZN(n3694)
         );
  AOI21_X1 U4480 ( .B1(n3720), .B2(n4199), .A(n3694), .ZN(n3695) );
  OAI21_X1 U4481 ( .B1(n3696), .B2(n3722), .A(n3695), .ZN(U3235) );
  INV_X1 U4482 ( .A(n3698), .ZN(n3700) );
  NOR2_X1 U4483 ( .A1(n3700), .A2(n3699), .ZN(n3701) );
  XNOR2_X1 U4484 ( .A(n3697), .B(n3701), .ZN(n3702) );
  NAND2_X1 U4485 ( .A1(n3702), .A2(n4353), .ZN(n3709) );
  OAI22_X1 U4486 ( .A1(n4037), .A2(n3704), .B1(STATE_REG_SCAN_IN), .B2(n3703), 
        .ZN(n3707) );
  OAI22_X1 U4487 ( .A1(n3705), .A2(n4040), .B1(n4074), .B2(n4343), .ZN(n3706)
         );
  NOR2_X1 U4488 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  OAI211_X1 U4489 ( .C1(n4358), .C2(n4041), .A(n3709), .B(n3708), .ZN(U3237)
         );
  NAND2_X1 U4490 ( .A1(n3710), .A2(n3711), .ZN(n3712) );
  XOR2_X1 U4491 ( .A(n4349), .B(n3712), .Z(n3723) );
  AND2_X1 U4492 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4979) );
  AOI21_X1 U4493 ( .B1(n4348), .B2(n3713), .A(n4979), .ZN(n3716) );
  NAND2_X1 U4494 ( .A1(n3714), .A2(n3889), .ZN(n3715) );
  OAI211_X1 U4495 ( .C1(n3705), .C2(n3717), .A(n3716), .B(n3715), .ZN(n3718)
         );
  AOI21_X1 U4496 ( .B1(n3720), .B2(n3719), .A(n3718), .ZN(n3721) );
  OAI21_X1 U4497 ( .B1(n3723), .B2(n3722), .A(n3721), .ZN(U3238) );
  INV_X1 U4498 ( .A(n3795), .ZN(n3724) );
  NOR2_X1 U4499 ( .A1(n3725), .A2(n3724), .ZN(n3858) );
  INV_X1 U4500 ( .A(n3852), .ZN(n3786) );
  INV_X1 U4501 ( .A(n4491), .ZN(n3729) );
  OAI211_X1 U4502 ( .C1(n3729), .C2(n2816), .A(n3728), .B(n3727), .ZN(n3732)
         );
  NAND3_X1 U4503 ( .A1(n3732), .A2(n3731), .A3(n3730), .ZN(n3734) );
  OAI211_X1 U4504 ( .C1(n2897), .C2(n3735), .A(n3734), .B(n3733), .ZN(n3738)
         );
  NAND3_X1 U4505 ( .A1(n3738), .A2(n3737), .A3(n3736), .ZN(n3741) );
  NAND4_X1 U4506 ( .A1(n3741), .A2(n3740), .A3(n3752), .A4(n3739), .ZN(n3744)
         );
  INV_X1 U4507 ( .A(n3790), .ZN(n3743) );
  NAND3_X1 U4508 ( .A1(n3744), .A2(n3743), .A3(n3742), .ZN(n3745) );
  NAND3_X1 U4509 ( .A1(n3745), .A2(n3754), .A3(n3753), .ZN(n3748) );
  AND3_X1 U4510 ( .A1(n3748), .A2(n3747), .A3(n3746), .ZN(n3758) );
  NAND2_X1 U4511 ( .A1(n3750), .A2(n3749), .ZN(n3757) );
  AND2_X1 U4512 ( .A1(n3757), .A2(n3773), .ZN(n3845) );
  INV_X1 U4513 ( .A(n3751), .ZN(n3755) );
  NAND4_X1 U4514 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3756)
         );
  OAI22_X1 U4515 ( .A1(n3758), .A2(n3757), .B1(n3845), .B2(n3756), .ZN(n3762)
         );
  INV_X1 U4516 ( .A(n3845), .ZN(n3760) );
  AOI22_X1 U4517 ( .A1(n3762), .A2(n3761), .B1(n2368), .B2(n3760), .ZN(n3777)
         );
  NAND2_X1 U4518 ( .A1(n3764), .A2(n3763), .ZN(n3769) );
  INV_X1 U4519 ( .A(n3769), .ZN(n3767) );
  NAND3_X1 U4520 ( .A1(n3767), .A2(n3766), .A3(n3765), .ZN(n3776) );
  INV_X1 U4521 ( .A(n3768), .ZN(n3770) );
  AOI21_X1 U4522 ( .B1(n3771), .B2(n3770), .A(n3769), .ZN(n3774) );
  INV_X1 U4523 ( .A(n3773), .ZN(n3841) );
  NOR4_X1 U4524 ( .A1(n3774), .A2(n3842), .A3(n2392), .A4(n3841), .ZN(n3775)
         );
  OAI22_X1 U4525 ( .A1(n3777), .A2(n3776), .B1(n3845), .B2(n3775), .ZN(n3779)
         );
  INV_X1 U4526 ( .A(n3843), .ZN(n3778) );
  AOI21_X1 U4527 ( .B1(n3779), .B2(n3848), .A(n3778), .ZN(n3781) );
  NOR4_X1 U4528 ( .A1(n3781), .A2(n2377), .A3(n3780), .A4(n4143), .ZN(n3782)
         );
  AOI21_X1 U4529 ( .B1(n3850), .B2(n2374), .A(n3782), .ZN(n3783) );
  OAI21_X1 U4530 ( .B1(n3783), .B2(n3819), .A(n3854), .ZN(n3784) );
  OAI221_X1 U4531 ( .B1(n3786), .B2(n3785), .C1(n3786), .C2(n3784), .A(n3863), 
        .ZN(n3789) );
  NAND2_X1 U4532 ( .A1(n3806), .A2(DATAI_29_), .ZN(n3976) );
  NAND2_X1 U4533 ( .A1(n3884), .A2(n3976), .ZN(n3834) );
  NAND4_X1 U4534 ( .A1(n3834), .A2(n3985), .A3(n3787), .A4(n3836), .ZN(n3788)
         );
  AOI21_X1 U4535 ( .B1(n3858), .B2(n3789), .A(n3788), .ZN(n3832) );
  NOR4_X1 U4536 ( .A1(n3792), .A2(n4492), .A3(n3791), .A4(n3790), .ZN(n3793)
         );
  XNOR2_X1 U4537 ( .A(n3887), .B(n4147), .ZN(n4144) );
  XNOR2_X1 U4538 ( .A(n4151), .B(n4169), .ZN(n4160) );
  INV_X1 U4539 ( .A(n4160), .ZN(n4165) );
  NAND3_X1 U4540 ( .A1(n3793), .A2(n4144), .A3(n4165), .ZN(n3815) );
  NAND2_X1 U4541 ( .A1(n3795), .A2(n3794), .ZN(n4050) );
  INV_X1 U4542 ( .A(n4050), .ZN(n3804) );
  NOR4_X1 U4543 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n2816), .ZN(n3803)
         );
  NOR4_X1 U4544 ( .A1(n3801), .A2(n3800), .A3(n4194), .A4(n3799), .ZN(n3802)
         );
  NAND3_X1 U4545 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3814) );
  NAND2_X1 U4546 ( .A1(n4048), .A2(n3805), .ZN(n4068) );
  INV_X1 U4547 ( .A(n4068), .ZN(n3812) );
  INV_X1 U4548 ( .A(n3990), .ZN(n3807) );
  NAND2_X1 U4549 ( .A1(n3806), .A2(DATAI_30_), .ZN(n4209) );
  INV_X1 U4550 ( .A(n4209), .ZN(n4215) );
  NAND2_X1 U4551 ( .A1(n3807), .A2(n4215), .ZN(n3810) );
  INV_X1 U4552 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U4553 ( .A1(n2220), .A2(REG2_REG_31__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U4554 ( .A1(n2740), .A2(REG0_REG_31__SCAN_IN), .ZN(n3808) );
  OAI211_X1 U4555 ( .C1(n2719), .C2(n4206), .A(n3809), .B(n3808), .ZN(n3977)
         );
  NAND2_X1 U4556 ( .A1(n3806), .A2(DATAI_31_), .ZN(n3978) );
  NAND2_X1 U4557 ( .A1(n3977), .A2(n3978), .ZN(n3869) );
  AND2_X1 U4558 ( .A1(n3810), .A2(n3869), .ZN(n3859) );
  NAND4_X1 U4559 ( .A1(n3812), .A2(n3811), .A3(n4529), .A4(n3859), .ZN(n3813)
         );
  OR4_X1 U4560 ( .A1(n4013), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3830) );
  INV_X1 U4561 ( .A(n3816), .ZN(n3818) );
  NAND2_X1 U4562 ( .A1(n3818), .A2(n3817), .ZN(n4030) );
  XNOR2_X1 U4563 ( .A(n4071), .B(n4092), .ZN(n4089) );
  INV_X1 U4564 ( .A(n3819), .ZN(n3820) );
  AND2_X1 U4565 ( .A1(n3820), .A2(n4085), .ZN(n4122) );
  INV_X1 U4566 ( .A(n4122), .ZN(n4128) );
  NOR4_X1 U4567 ( .A1(n4128), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3828)
         );
  NOR4_X1 U4568 ( .A1(n4104), .A2(n2341), .A3(n3826), .A4(n3825), .ZN(n3827)
         );
  NAND4_X1 U4569 ( .A1(n4030), .A2(n4089), .A3(n3828), .A4(n3827), .ZN(n3829)
         );
  OR2_X1 U4570 ( .A1(n3884), .A2(n3976), .ZN(n3857) );
  NAND2_X1 U4571 ( .A1(n3857), .A2(n3834), .ZN(n3997) );
  NOR4_X1 U4572 ( .A1(n3995), .A2(n3830), .A3(n3829), .A4(n3997), .ZN(n3831)
         );
  MUX2_X1 U4573 ( .A(n3832), .B(n3831), .S(n4326), .Z(n3833) );
  INV_X1 U4574 ( .A(n3833), .ZN(n3876) );
  NAND2_X1 U4575 ( .A1(n3990), .A2(n4209), .ZN(n3866) );
  OAI21_X1 U4576 ( .B1(n3977), .B2(n3978), .A(n3866), .ZN(n3875) );
  AND2_X1 U4577 ( .A1(n3983), .A2(n3856), .ZN(n3835) );
  NAND2_X1 U4578 ( .A1(n3834), .A2(n3985), .ZN(n3837) );
  OAI211_X1 U4579 ( .C1(n3835), .C2(n3837), .A(n3859), .B(n3857), .ZN(n3871)
         );
  INV_X1 U4580 ( .A(n3836), .ZN(n3838) );
  NOR3_X1 U4581 ( .A1(n4013), .A2(n3838), .A3(n3837), .ZN(n3839) );
  NOR2_X1 U4582 ( .A1(n3871), .A2(n3839), .ZN(n3865) );
  NOR3_X1 U4583 ( .A1(n3842), .A2(n3841), .A3(n3840), .ZN(n3844) );
  OAI21_X1 U4584 ( .B1(n3845), .B2(n3844), .A(n3843), .ZN(n3846) );
  AND4_X1 U4585 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3851)
         );
  OAI21_X1 U4586 ( .B1(n3851), .B2(n2374), .A(n3850), .ZN(n3853) );
  OAI221_X1 U4587 ( .B1(n3855), .B2(n3854), .C1(n3855), .C2(n3853), .A(n3852), 
        .ZN(n3862) );
  NAND4_X1 U4588 ( .A1(n3858), .A2(n3857), .A3(n3983), .A4(n3856), .ZN(n3861)
         );
  INV_X1 U4589 ( .A(n3859), .ZN(n3860) );
  AOI211_X1 U4590 ( .C1(n3863), .C2(n3862), .A(n3861), .B(n3860), .ZN(n3864)
         );
  OAI22_X1 U4591 ( .A1(n3865), .A2(n3864), .B1(n3977), .B2(n4209), .ZN(n3873)
         );
  AOI21_X1 U4592 ( .B1(n3866), .B2(n3977), .A(n3978), .ZN(n3868) );
  NOR2_X1 U4593 ( .A1(n3868), .A2(n3867), .ZN(n3872) );
  AOI21_X1 U4594 ( .B1(n3875), .B2(n3869), .A(n4326), .ZN(n3870) );
  AOI22_X1 U4595 ( .A1(n3873), .A2(n3872), .B1(n3871), .B2(n3870), .ZN(n3874)
         );
  OAI21_X1 U4596 ( .B1(n3876), .B2(n3875), .A(n3874), .ZN(n3877) );
  XNOR2_X1 U4597 ( .A(n3877), .B(n4327), .ZN(n3883) );
  INV_X1 U4598 ( .A(n3878), .ZN(n3879) );
  NOR2_X1 U4599 ( .A1(n3879), .A2(n3910), .ZN(n3881) );
  OAI21_X1 U4600 ( .B1(n3882), .B2(n4325), .A(B_REG_SCAN_IN), .ZN(n3880) );
  OAI22_X1 U4601 ( .A1(n3883), .A2(n3882), .B1(n3881), .B2(n3880), .ZN(U3239)
         );
  MUX2_X1 U4602 ( .A(DATAO_REG_31__SCAN_IN), .B(n3977), .S(n3901), .Z(U3581)
         );
  MUX2_X1 U4603 ( .A(DATAO_REG_29__SCAN_IN), .B(n3884), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4604 ( .A(DATAO_REG_28__SCAN_IN), .B(n3885), .S(n3901), .Z(U3578)
         );
  MUX2_X1 U4605 ( .A(DATAO_REG_27__SCAN_IN), .B(n3886), .S(n3901), .Z(U3577)
         );
  MUX2_X1 U4606 ( .A(DATAO_REG_26__SCAN_IN), .B(n4055), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4607 ( .A(DATAO_REG_25__SCAN_IN), .B(n4034), .S(n3901), .Z(U3575)
         );
  MUX2_X1 U4608 ( .A(DATAO_REG_22__SCAN_IN), .B(n4132), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4609 ( .A(DATAO_REG_20__SCAN_IN), .B(n3887), .S(n3901), .Z(U3570)
         );
  MUX2_X1 U4610 ( .A(DATAO_REG_18__SCAN_IN), .B(n4170), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4611 ( .A(DATAO_REG_15__SCAN_IN), .B(n3888), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4612 ( .A(DATAO_REG_14__SCAN_IN), .B(n3889), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4613 ( .A(DATAO_REG_13__SCAN_IN), .B(n3890), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4614 ( .A(DATAO_REG_11__SCAN_IN), .B(n3891), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4615 ( .A(DATAO_REG_10__SCAN_IN), .B(n3892), .S(n3901), .Z(U3560)
         );
  MUX2_X1 U4616 ( .A(DATAO_REG_9__SCAN_IN), .B(n3893), .S(n3901), .Z(U3559) );
  MUX2_X1 U4617 ( .A(DATAO_REG_8__SCAN_IN), .B(n3894), .S(n3901), .Z(U3558) );
  MUX2_X1 U4618 ( .A(DATAO_REG_7__SCAN_IN), .B(n3895), .S(U4043), .Z(U3557) );
  MUX2_X1 U4619 ( .A(DATAO_REG_6__SCAN_IN), .B(n3896), .S(n3901), .Z(U3556) );
  MUX2_X1 U4620 ( .A(DATAO_REG_5__SCAN_IN), .B(n3897), .S(U4043), .Z(U3555) );
  MUX2_X1 U4621 ( .A(DATAO_REG_4__SCAN_IN), .B(n3898), .S(n3901), .Z(U3554) );
  MUX2_X1 U4622 ( .A(DATAO_REG_3__SCAN_IN), .B(n3899), .S(n3901), .Z(U3553) );
  MUX2_X1 U4623 ( .A(DATAO_REG_1__SCAN_IN), .B(n3900), .S(n3901), .Z(U3551) );
  MUX2_X1 U4624 ( .A(DATAO_REG_0__SCAN_IN), .B(n2867), .S(n3901), .Z(U3550) );
  OAI211_X1 U4625 ( .C1(n3454), .C2(n3903), .A(n4479), .B(n3926), .ZN(n3908)
         );
  AND2_X1 U4626 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3911)
         );
  OAI211_X1 U4627 ( .C1(n3911), .C2(n3904), .A(n4985), .B(n3919), .ZN(n3907)
         );
  AOI22_X1 U4628 ( .A1(n4980), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3906) );
  INV_X1 U4629 ( .A(n4989), .ZN(n4456) );
  NAND4_X1 U4630 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(U3241)
         );
  INV_X1 U4631 ( .A(n4322), .ZN(n4363) );
  NAND3_X1 U4632 ( .A1(n3909), .A2(n4321), .A3(n4363), .ZN(n3914) );
  INV_X1 U4633 ( .A(n3910), .ZN(n3912) );
  OAI21_X1 U4634 ( .B1(REG2_REG_0__SCAN_IN), .B2(n4363), .A(n4321), .ZN(n4362)
         );
  AOI22_X1 U4635 ( .A1(n3912), .A2(n3911), .B1(n4362), .B2(n2308), .ZN(n3913)
         );
  NAND3_X1 U4636 ( .A1(n3914), .A2(U4043), .A3(n3913), .ZN(n3940) );
  INV_X1 U4637 ( .A(n4980), .ZN(n4459) );
  INV_X1 U4638 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n3915) );
  OAI22_X1 U4639 ( .A1(n4459), .A2(n3915), .B1(STATE_REG_SCAN_IN), .B2(n2525), 
        .ZN(n3916) );
  AOI21_X1 U4640 ( .B1(n4331), .B2(n4456), .A(n3916), .ZN(n3931) );
  INV_X1 U4641 ( .A(n3917), .ZN(n3922) );
  NAND3_X1 U4642 ( .A1(n3920), .A2(n3919), .A3(n3918), .ZN(n3921) );
  NAND3_X1 U4643 ( .A1(n4985), .A2(n3922), .A3(n3921), .ZN(n3930) );
  INV_X1 U4644 ( .A(n3923), .ZN(n3928) );
  NAND3_X1 U4645 ( .A1(n3926), .A2(n3925), .A3(n3924), .ZN(n3927) );
  NAND3_X1 U4646 ( .A1(n4479), .A2(n3928), .A3(n3927), .ZN(n3929) );
  NAND4_X1 U4647 ( .A1(n3940), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(U3242)
         );
  AOI21_X1 U4648 ( .B1(n4980), .B2(ADDR_REG_4__SCAN_IN), .A(n3932), .ZN(n3939)
         );
  XNOR2_X1 U4649 ( .A(n3933), .B(REG1_REG_4__SCAN_IN), .ZN(n3936) );
  XNOR2_X1 U4650 ( .A(n3934), .B(REG2_REG_4__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4651 ( .A1(n4479), .A2(n3936), .B1(n4985), .B2(n3935), .ZN(n3938)
         );
  NAND2_X1 U4652 ( .A1(n4456), .A2(n4330), .ZN(n3937) );
  NAND4_X1 U4653 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(U3244)
         );
  INV_X1 U4654 ( .A(n3967), .ZN(n3964) );
  INV_X1 U4655 ( .A(n4513), .ZN(n3958) );
  INV_X1 U4656 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4657 ( .A1(n4513), .A2(n3941), .B1(REG1_REG_17__SCAN_IN), .B2(
        n3958), .ZN(n4477) );
  INV_X1 U4658 ( .A(n4455), .ZN(n4518) );
  NOR2_X1 U4659 ( .A1(n3944), .A2(n4518), .ZN(n3945) );
  INV_X1 U4660 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4762) );
  INV_X1 U4661 ( .A(n4516), .ZN(n4988) );
  AOI22_X1 U4662 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4988), .B1(n4516), .B2(
        n4855), .ZN(n4977) );
  NAND2_X1 U4663 ( .A1(n3946), .A2(n4515), .ZN(n3947) );
  INV_X1 U4664 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4465) );
  XNOR2_X1 U4665 ( .A(n3967), .B(REG1_REG_18__SCAN_IN), .ZN(n3948) );
  XNOR2_X1 U4666 ( .A(n3967), .B(REG2_REG_18__SCAN_IN), .ZN(n3960) );
  NOR2_X1 U4667 ( .A1(REG2_REG_17__SCAN_IN), .A2(n3958), .ZN(n3950) );
  AOI21_X1 U4668 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3958), .A(n3950), .ZN(n4474) );
  NOR2_X1 U4669 ( .A1(n4518), .A2(n3953), .ZN(n3954) );
  INV_X1 U4670 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4776) );
  XOR2_X1 U4671 ( .A(n4455), .B(n3953), .Z(n4452) );
  NOR2_X1 U4672 ( .A1(n4776), .A2(n4452), .ZN(n4451) );
  NOR2_X1 U4673 ( .A1(n3954), .A2(n4451), .ZN(n4982) );
  NAND2_X1 U4674 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4516), .ZN(n3955) );
  OAI21_X1 U4675 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4516), .A(n3955), .ZN(n4983) );
  NOR2_X1 U4676 ( .A1(n4982), .A2(n4983), .ZN(n4981) );
  NAND2_X1 U4677 ( .A1(n3956), .A2(n4515), .ZN(n3957) );
  INV_X1 U4678 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4462) );
  AOI21_X1 U4679 ( .B1(n4980), .B2(ADDR_REG_18__SCAN_IN), .A(n3962), .ZN(n3963) );
  OAI211_X1 U4680 ( .C1(n3964), .C2(n4989), .A(n2248), .B(n3963), .ZN(U3258)
         );
  XNOR2_X1 U4681 ( .A(n4327), .B(REG1_REG_19__SCAN_IN), .ZN(n3965) );
  INV_X1 U4682 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3968) );
  MUX2_X1 U4683 ( .A(REG2_REG_19__SCAN_IN), .B(n3968), .S(n4327), .Z(n3969) );
  NAND2_X1 U4684 ( .A1(n4980), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3970) );
  OAI211_X1 U4685 ( .C1(n4989), .C2(n3972), .A(n3971), .B(n3970), .ZN(n3973)
         );
  AOI21_X1 U4686 ( .B1(n3974), .B2(n4985), .A(n3973), .ZN(n3975) );
  INV_X1 U4687 ( .A(n3976), .ZN(n4000) );
  NAND2_X1 U4688 ( .A1(n4210), .A2(n4209), .ZN(n4212) );
  XOR2_X1 U4689 ( .A(n3978), .B(n4212), .Z(n4284) );
  INV_X1 U4690 ( .A(n4507), .ZN(n3979) );
  AOI21_X1 U4691 ( .B1(B_REG_SCAN_IN), .B2(n4322), .A(n4489), .ZN(n3989) );
  NAND2_X1 U4692 ( .A1(n3977), .A2(n3989), .ZN(n4213) );
  OAI21_X1 U4693 ( .B1(n3978), .B2(n4107), .A(n4213), .ZN(n4281) );
  NAND2_X1 U4694 ( .A1(n3979), .A2(n4281), .ZN(n3981) );
  NAND2_X1 U4695 ( .A1(n4200), .A2(REG2_REG_31__SCAN_IN), .ZN(n3980) );
  OAI211_X1 U4696 ( .C1(n4284), .C2(n4179), .A(n3981), .B(n3980), .ZN(U3260)
         );
  INV_X1 U4697 ( .A(n3982), .ZN(n3993) );
  INV_X1 U4698 ( .A(n3983), .ZN(n3984) );
  XNOR2_X1 U4699 ( .A(n3987), .B(n3997), .ZN(n3988) );
  NAND2_X1 U4700 ( .A1(n3988), .A2(n4167), .ZN(n3992) );
  AOI22_X1 U4701 ( .A1(n3990), .A2(n3989), .B1(n4486), .B2(n4000), .ZN(n3991)
         );
  OAI211_X1 U4702 ( .C1(n4019), .C2(n4188), .A(n3992), .B(n3991), .ZN(n4218)
         );
  AOI21_X1 U4703 ( .B1(n3993), .B2(n4499), .A(n4218), .ZN(n4003) );
  XNOR2_X1 U4704 ( .A(n3998), .B(n3997), .ZN(n4217) );
  NAND2_X1 U4705 ( .A1(n4217), .A2(n4204), .ZN(n4002) );
  AOI21_X1 U4706 ( .B1(n4000), .B2(n3999), .A(n4210), .ZN(n4219) );
  AOI22_X1 U4707 ( .A1(n4219), .A2(n4504), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4200), .ZN(n4001) );
  OAI211_X1 U4708 ( .C1(n4507), .C2(n4003), .A(n4002), .B(n4001), .ZN(U3354)
         );
  INV_X1 U4709 ( .A(n4004), .ZN(n4011) );
  AOI22_X1 U4710 ( .A1(n4005), .A2(n4499), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4200), .ZN(n4006) );
  OAI21_X1 U4711 ( .B1(n4007), .B2(n4179), .A(n4006), .ZN(n4008) );
  AOI21_X1 U4712 ( .B1(n4009), .B2(n3979), .A(n4008), .ZN(n4010) );
  OAI21_X1 U4713 ( .B1(n4011), .B2(n4182), .A(n4010), .ZN(U3262) );
  XNOR2_X1 U4714 ( .A(n4012), .B(n4013), .ZN(n4222) );
  NAND2_X1 U4715 ( .A1(n4014), .A2(n4013), .ZN(n4015) );
  NAND2_X1 U4716 ( .A1(n4016), .A2(n4015), .ZN(n4021) );
  AOI22_X1 U4717 ( .A1(n4055), .A2(n4487), .B1(n4017), .B2(n4486), .ZN(n4018)
         );
  OAI21_X1 U4718 ( .B1(n4019), .B2(n4489), .A(n4018), .ZN(n4020) );
  AOI21_X1 U4719 ( .B1(n4021), .B2(n4191), .A(n4020), .ZN(n4223) );
  NOR2_X1 U4720 ( .A1(n4223), .A2(n4507), .ZN(n4027) );
  OAI21_X1 U4721 ( .B1(n4038), .B2(n4023), .A(n4022), .ZN(n4225) );
  AOI22_X1 U4722 ( .A1(REG2_REG_27__SCAN_IN), .A2(n4507), .B1(n4024), .B2(
        n4499), .ZN(n4025) );
  OAI21_X1 U4723 ( .B1(n4225), .B2(n4179), .A(n4025), .ZN(n4026) );
  AOI211_X1 U4724 ( .C1(n4222), .C2(n4204), .A(n4027), .B(n4026), .ZN(n4028)
         );
  INV_X1 U4725 ( .A(n4028), .ZN(U3263) );
  XNOR2_X1 U4726 ( .A(n4029), .B(n4030), .ZN(n4227) );
  INV_X1 U4727 ( .A(n4227), .ZN(n4046) );
  XNOR2_X1 U4728 ( .A(n4031), .B(n4030), .ZN(n4032) );
  NAND2_X1 U4729 ( .A1(n4032), .A2(n4167), .ZN(n4036) );
  AOI22_X1 U4730 ( .A1(n4034), .A2(n4487), .B1(n4033), .B2(n4486), .ZN(n4035)
         );
  OAI211_X1 U4731 ( .C1(n4037), .C2(n4489), .A(n4036), .B(n4035), .ZN(n4226)
         );
  INV_X1 U4732 ( .A(n4038), .ZN(n4039) );
  OAI21_X1 U4733 ( .B1(n2250), .B2(n4040), .A(n4039), .ZN(n4293) );
  NOR2_X1 U4734 ( .A1(n4293), .A2(n4179), .ZN(n4044) );
  INV_X1 U4735 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4042) );
  OAI22_X1 U4736 ( .A1(n3979), .A2(n4042), .B1(n4041), .B2(n4124), .ZN(n4043)
         );
  AOI211_X1 U4737 ( .C1(n4226), .C2(n3979), .A(n4044), .B(n4043), .ZN(n4045)
         );
  OAI21_X1 U4738 ( .B1(n4046), .B2(n4182), .A(n4045), .ZN(U3264) );
  XOR2_X1 U4739 ( .A(n4050), .B(n4047), .Z(n4232) );
  NAND2_X1 U4740 ( .A1(n4049), .A2(n4048), .ZN(n4051) );
  XNOR2_X1 U4741 ( .A(n4051), .B(n4050), .ZN(n4052) );
  NAND2_X1 U4742 ( .A1(n4052), .A2(n4167), .ZN(n4057) );
  OAI22_X1 U4743 ( .A1(n4095), .A2(n4188), .B1(n4053), .B2(n4107), .ZN(n4054)
         );
  AOI21_X1 U4744 ( .B1(n4055), .B2(n4185), .A(n4054), .ZN(n4056) );
  NAND2_X1 U4745 ( .A1(n4057), .A2(n4056), .ZN(n4229) );
  AOI21_X1 U4746 ( .B1(n4058), .B2(n4075), .A(n2250), .ZN(n4230) );
  INV_X1 U4747 ( .A(n4230), .ZN(n4061) );
  AOI22_X1 U4748 ( .A1(n4507), .A2(REG2_REG_25__SCAN_IN), .B1(n4059), .B2(
        n4499), .ZN(n4060) );
  OAI21_X1 U4749 ( .B1(n4061), .B2(n4179), .A(n4060), .ZN(n4062) );
  AOI21_X1 U4750 ( .B1(n4229), .B2(n3979), .A(n4062), .ZN(n4063) );
  OAI21_X1 U4751 ( .B1(n4232), .B2(n4182), .A(n4063), .ZN(U3265) );
  XNOR2_X1 U4752 ( .A(n4064), .B(n4068), .ZN(n4234) );
  INV_X1 U4753 ( .A(n4234), .ZN(n4083) );
  NAND2_X1 U4754 ( .A1(n4066), .A2(n4065), .ZN(n4067) );
  XOR2_X1 U4755 ( .A(n4068), .B(n4067), .Z(n4069) );
  NAND2_X1 U4756 ( .A1(n4069), .A2(n4167), .ZN(n4073) );
  AOI22_X1 U4757 ( .A1(n4071), .A2(n4487), .B1(n4486), .B2(n4070), .ZN(n4072)
         );
  OAI211_X1 U4758 ( .C1(n4074), .C2(n4489), .A(n4073), .B(n4072), .ZN(n4233)
         );
  INV_X1 U4759 ( .A(n4096), .ZN(n4077) );
  OAI21_X1 U4760 ( .B1(n4077), .B2(n4076), .A(n4075), .ZN(n4298) );
  INV_X1 U4761 ( .A(n4078), .ZN(n4079) );
  AOI22_X1 U4762 ( .A1(n4507), .A2(REG2_REG_24__SCAN_IN), .B1(n4079), .B2(
        n4499), .ZN(n4080) );
  OAI21_X1 U4763 ( .B1(n4298), .B2(n4179), .A(n4080), .ZN(n4081) );
  AOI21_X1 U4764 ( .B1(n4233), .B2(n3979), .A(n4081), .ZN(n4082) );
  OAI21_X1 U4765 ( .B1(n4083), .B2(n4182), .A(n4082), .ZN(U3266) );
  XNOR2_X1 U4766 ( .A(n4084), .B(n4089), .ZN(n4238) );
  INV_X1 U4767 ( .A(n4238), .ZN(n4102) );
  INV_X1 U4768 ( .A(n4129), .ZN(n4087) );
  INV_X1 U4769 ( .A(n4085), .ZN(n4086) );
  AOI21_X1 U4770 ( .B1(n4087), .B2(n4122), .A(n4086), .ZN(n4105) );
  OAI21_X1 U4771 ( .B1(n4105), .B2(n4104), .A(n4088), .ZN(n4090) );
  XNOR2_X1 U4772 ( .A(n4090), .B(n4089), .ZN(n4091) );
  NAND2_X1 U4773 ( .A1(n4091), .A2(n4167), .ZN(n4094) );
  AOI22_X1 U4774 ( .A1(n4132), .A2(n4487), .B1(n4486), .B2(n4092), .ZN(n4093)
         );
  OAI211_X1 U4775 ( .C1(n4095), .C2(n4489), .A(n4094), .B(n4093), .ZN(n4237)
         );
  OAI21_X1 U4776 ( .B1(n4113), .B2(n4097), .A(n4096), .ZN(n4302) );
  AOI22_X1 U4777 ( .A1(n4507), .A2(REG2_REG_23__SCAN_IN), .B1(n4098), .B2(
        n4499), .ZN(n4099) );
  OAI21_X1 U4778 ( .B1(n4302), .B2(n4179), .A(n4099), .ZN(n4100) );
  AOI21_X1 U4779 ( .B1(n4237), .B2(n3979), .A(n4100), .ZN(n4101) );
  OAI21_X1 U4780 ( .B1(n4102), .B2(n4182), .A(n4101), .ZN(U3267) );
  OAI21_X1 U4781 ( .B1(n2224), .B2(n4104), .A(n4103), .ZN(n4245) );
  XNOR2_X1 U4782 ( .A(n4105), .B(n4104), .ZN(n4111) );
  NOR2_X1 U4783 ( .A1(n4106), .A2(n4489), .ZN(n4110) );
  OAI22_X1 U4784 ( .A1(n4108), .A2(n4188), .B1(n4114), .B2(n4107), .ZN(n4109)
         );
  AOI211_X1 U4785 ( .C1(n4111), .C2(n4191), .A(n4110), .B(n4109), .ZN(n4244)
         );
  AOI22_X1 U4786 ( .A1(n4507), .A2(REG2_REG_22__SCAN_IN), .B1(n4112), .B2(
        n4499), .ZN(n4118) );
  INV_X1 U4787 ( .A(n4113), .ZN(n4242) );
  INV_X1 U4788 ( .A(n4123), .ZN(n4116) );
  INV_X1 U4789 ( .A(n4114), .ZN(n4115) );
  NAND2_X1 U4790 ( .A1(n4116), .A2(n4115), .ZN(n4241) );
  NAND3_X1 U4791 ( .A1(n4242), .A2(n4504), .A3(n4241), .ZN(n4117) );
  OAI211_X1 U4792 ( .C1(n4244), .C2(n4507), .A(n4118), .B(n4117), .ZN(n4119)
         );
  INV_X1 U4793 ( .A(n4119), .ZN(n4120) );
  OAI21_X1 U4794 ( .B1(n4245), .B2(n4182), .A(n4120), .ZN(U3268) );
  XOR2_X1 U4795 ( .A(n4122), .B(n4121), .Z(n4249) );
  AOI21_X1 U4796 ( .B1(n4131), .B2(n4152), .A(n4123), .ZN(n4247) );
  INV_X1 U4797 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4126) );
  OAI22_X1 U4798 ( .A1(n3979), .A2(n4126), .B1(n4125), .B2(n4124), .ZN(n4127)
         );
  AOI21_X1 U4799 ( .B1(n4247), .B2(n4504), .A(n4127), .ZN(n4136) );
  XNOR2_X1 U4800 ( .A(n4129), .B(n4128), .ZN(n4130) );
  NAND2_X1 U4801 ( .A1(n4130), .A2(n4167), .ZN(n4134) );
  AOI22_X1 U4802 ( .A1(n4132), .A2(n4185), .B1(n4486), .B2(n4131), .ZN(n4133)
         );
  OAI211_X1 U4803 ( .C1(n4173), .C2(n4188), .A(n4134), .B(n4133), .ZN(n4246)
         );
  NAND2_X1 U4804 ( .A1(n4246), .A2(n3979), .ZN(n4135) );
  OAI211_X1 U4805 ( .C1(n4249), .C2(n4182), .A(n4136), .B(n4135), .ZN(U3269)
         );
  XNOR2_X1 U4806 ( .A(n4137), .B(n4144), .ZN(n4251) );
  INV_X1 U4807 ( .A(n4251), .ZN(n4159) );
  NAND2_X1 U4808 ( .A1(n4139), .A2(n4138), .ZN(n4184) );
  INV_X1 U4809 ( .A(n4140), .ZN(n4141) );
  NOR2_X1 U4810 ( .A1(n4184), .A2(n4141), .ZN(n4164) );
  OAI21_X1 U4811 ( .B1(n4164), .B2(n4143), .A(n4142), .ZN(n4145) );
  XNOR2_X1 U4812 ( .A(n4145), .B(n4144), .ZN(n4146) );
  NAND2_X1 U4813 ( .A1(n4146), .A2(n4167), .ZN(n4150) );
  AOI22_X1 U4814 ( .A1(n4148), .A2(n4185), .B1(n4486), .B2(n4147), .ZN(n4149)
         );
  OAI211_X1 U4815 ( .C1(n4151), .C2(n4188), .A(n4150), .B(n4149), .ZN(n4250)
         );
  INV_X1 U4816 ( .A(n4174), .ZN(n4154) );
  OAI21_X1 U4817 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4308) );
  AOI22_X1 U4818 ( .A1(n4507), .A2(REG2_REG_20__SCAN_IN), .B1(n4155), .B2(
        n4499), .ZN(n4156) );
  OAI21_X1 U4819 ( .B1(n4308), .B2(n4179), .A(n4156), .ZN(n4157) );
  AOI21_X1 U4820 ( .B1(n4250), .B2(n3979), .A(n4157), .ZN(n4158) );
  OAI21_X1 U4821 ( .B1(n4159), .B2(n4182), .A(n4158), .ZN(U3270) );
  XNOR2_X1 U4822 ( .A(n4161), .B(n4160), .ZN(n4254) );
  INV_X1 U4823 ( .A(n4254), .ZN(n4183) );
  INV_X1 U4824 ( .A(n4162), .ZN(n4163) );
  NOR2_X1 U4825 ( .A1(n4164), .A2(n4163), .ZN(n4166) );
  XNOR2_X1 U4826 ( .A(n4166), .B(n4165), .ZN(n4168) );
  NAND2_X1 U4827 ( .A1(n4168), .A2(n4167), .ZN(n4172) );
  AOI22_X1 U4828 ( .A1(n4170), .A2(n4487), .B1(n4486), .B2(n4169), .ZN(n4171)
         );
  OAI211_X1 U4829 ( .C1(n4173), .C2(n4489), .A(n4172), .B(n4171), .ZN(n4253)
         );
  OAI21_X1 U4830 ( .B1(n4176), .B2(n4175), .A(n4174), .ZN(n4313) );
  AOI22_X1 U4831 ( .A1(n4200), .A2(REG2_REG_19__SCAN_IN), .B1(n4177), .B2(
        n4499), .ZN(n4178) );
  OAI21_X1 U4832 ( .B1(n4313), .B2(n4179), .A(n4178), .ZN(n4180) );
  AOI21_X1 U4833 ( .B1(n4253), .B2(n3979), .A(n4180), .ZN(n4181) );
  OAI21_X1 U4834 ( .B1(n4183), .B2(n4182), .A(n4181), .ZN(U3271) );
  XOR2_X1 U4835 ( .A(n4194), .B(n4184), .Z(n4192) );
  AOI22_X1 U4836 ( .A1(n4186), .A2(n4185), .B1(n4196), .B2(n4486), .ZN(n4187)
         );
  OAI21_X1 U4837 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4190) );
  AOI21_X1 U4838 ( .B1(n4192), .B2(n4191), .A(n4190), .ZN(n4260) );
  OAI21_X1 U4839 ( .B1(n4195), .B2(n4194), .A(n4193), .ZN(n4258) );
  XNOR2_X1 U4840 ( .A(n4197), .B(n4196), .ZN(n4198) );
  NAND2_X1 U4841 ( .A1(n4198), .A2(n4577), .ZN(n4259) );
  AOI22_X1 U4842 ( .A1(n4200), .A2(REG2_REG_18__SCAN_IN), .B1(n4199), .B2(
        n4499), .ZN(n4201) );
  OAI21_X1 U4843 ( .B1(n4259), .B2(n4202), .A(n4201), .ZN(n4203) );
  AOI21_X1 U4844 ( .B1(n4258), .B2(n4204), .A(n4203), .ZN(n4205) );
  OAI21_X1 U4845 ( .B1(n4200), .B2(n4260), .A(n4205), .ZN(U3272) );
  NOR2_X1 U4846 ( .A1(n4595), .A2(n4206), .ZN(n4207) );
  AOI21_X1 U4847 ( .B1(n4595), .B2(n4281), .A(n4207), .ZN(n4208) );
  OAI21_X1 U4848 ( .B1(n4284), .B2(n4257), .A(n4208), .ZN(U3549) );
  OR2_X1 U4849 ( .A1(n4210), .A2(n4209), .ZN(n4211) );
  AND2_X1 U4850 ( .A1(n4212), .A2(n4211), .ZN(n4359) );
  INV_X1 U4851 ( .A(n4213), .ZN(n4214) );
  AOI21_X1 U4852 ( .B1(n4215), .B2(n4486), .A(n4214), .ZN(n4361) );
  MUX2_X1 U4853 ( .A(n3089), .B(n4361), .S(n4595), .Z(n4216) );
  OAI21_X1 U4854 ( .B1(n4287), .B2(n4257), .A(n4216), .ZN(U3548) );
  NAND2_X1 U4855 ( .A1(n4217), .A2(n4569), .ZN(n4221) );
  AOI21_X1 U4856 ( .B1(n4577), .B2(n4219), .A(n4218), .ZN(n4220) );
  NAND2_X1 U4857 ( .A1(n4221), .A2(n4220), .ZN(n4288) );
  MUX2_X1 U4858 ( .A(REG1_REG_29__SCAN_IN), .B(n4288), .S(n4595), .Z(U3547) );
  NAND2_X1 U4859 ( .A1(n4222), .A2(n4569), .ZN(n4224) );
  OAI211_X1 U4860 ( .C1(n4560), .C2(n4225), .A(n4224), .B(n4223), .ZN(n4289)
         );
  MUX2_X1 U4861 ( .A(REG1_REG_27__SCAN_IN), .B(n4289), .S(n4595), .Z(U3545) );
  AOI21_X1 U4862 ( .B1(n4227), .B2(n4569), .A(n4226), .ZN(n4290) );
  MUX2_X1 U4863 ( .A(n4771), .B(n4290), .S(n4595), .Z(n4228) );
  OAI21_X1 U4864 ( .B1(n4257), .B2(n4293), .A(n4228), .ZN(U3544) );
  AOI21_X1 U4865 ( .B1(n4577), .B2(n4230), .A(n4229), .ZN(n4231) );
  OAI21_X1 U4866 ( .B1(n4232), .B2(n4572), .A(n4231), .ZN(n4294) );
  MUX2_X1 U4867 ( .A(REG1_REG_25__SCAN_IN), .B(n4294), .S(n4595), .Z(U3543) );
  AOI21_X1 U4868 ( .B1(n4234), .B2(n4569), .A(n4233), .ZN(n4295) );
  MUX2_X1 U4869 ( .A(n4235), .B(n4295), .S(n4595), .Z(n4236) );
  OAI21_X1 U4870 ( .B1(n4257), .B2(n4298), .A(n4236), .ZN(U3542) );
  AOI21_X1 U4871 ( .B1(n4238), .B2(n4569), .A(n4237), .ZN(n4299) );
  MUX2_X1 U4872 ( .A(n4239), .B(n4299), .S(n4595), .Z(n4240) );
  OAI21_X1 U4873 ( .B1(n4257), .B2(n4302), .A(n4240), .ZN(U3541) );
  NAND3_X1 U4874 ( .A1(n4242), .A2(n4577), .A3(n4241), .ZN(n4243) );
  OAI211_X1 U4875 ( .C1(n4245), .C2(n4572), .A(n4244), .B(n4243), .ZN(n4303)
         );
  MUX2_X1 U4876 ( .A(REG1_REG_22__SCAN_IN), .B(n4303), .S(n4595), .Z(U3540) );
  AOI21_X1 U4877 ( .B1(n4577), .B2(n4247), .A(n4246), .ZN(n4248) );
  OAI21_X1 U4878 ( .B1(n4249), .B2(n4572), .A(n4248), .ZN(n4304) );
  MUX2_X1 U4879 ( .A(REG1_REG_21__SCAN_IN), .B(n4304), .S(n4595), .Z(U3539) );
  INV_X1 U4880 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4852) );
  AOI21_X1 U4881 ( .B1(n4251), .B2(n4569), .A(n4250), .ZN(n4305) );
  MUX2_X1 U4882 ( .A(n4852), .B(n4305), .S(n4595), .Z(n4252) );
  OAI21_X1 U4883 ( .B1(n4257), .B2(n4308), .A(n4252), .ZN(U3538) );
  INV_X1 U4884 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4255) );
  AOI21_X1 U4885 ( .B1(n4254), .B2(n4569), .A(n4253), .ZN(n4309) );
  MUX2_X1 U4886 ( .A(n4255), .B(n4309), .S(n4595), .Z(n4256) );
  OAI21_X1 U4887 ( .B1(n4257), .B2(n4313), .A(n4256), .ZN(U3537) );
  INV_X1 U4888 ( .A(n4258), .ZN(n4261) );
  OAI211_X1 U4889 ( .C1(n4261), .C2(n4572), .A(n4260), .B(n4259), .ZN(n4314)
         );
  MUX2_X1 U4890 ( .A(REG1_REG_18__SCAN_IN), .B(n4314), .S(n4595), .Z(U3536) );
  NAND3_X1 U4891 ( .A1(n4263), .A2(n4577), .A3(n4262), .ZN(n4264) );
  OAI211_X1 U4892 ( .C1(n4266), .C2(n4572), .A(n4265), .B(n4264), .ZN(n4315)
         );
  MUX2_X1 U4893 ( .A(REG1_REG_17__SCAN_IN), .B(n4315), .S(n4595), .Z(U3535) );
  NAND3_X1 U4894 ( .A1(n4268), .A2(n4577), .A3(n4267), .ZN(n4269) );
  OAI211_X1 U4895 ( .C1(n4271), .C2(n4572), .A(n4270), .B(n4269), .ZN(n4316)
         );
  MUX2_X1 U4896 ( .A(REG1_REG_16__SCAN_IN), .B(n4316), .S(n4595), .Z(U3534) );
  NAND3_X1 U4897 ( .A1(n4273), .A2(n4577), .A3(n4272), .ZN(n4274) );
  OAI211_X1 U4898 ( .C1(n4276), .C2(n4528), .A(n4275), .B(n4274), .ZN(n4317)
         );
  MUX2_X1 U4899 ( .A(REG1_REG_14__SCAN_IN), .B(n4317), .S(n4595), .Z(U3532) );
  NAND2_X1 U4900 ( .A1(n4277), .A2(n4566), .ZN(n4278) );
  OAI211_X1 U4901 ( .C1(n4560), .C2(n4280), .A(n4279), .B(n4278), .ZN(n4318)
         );
  MUX2_X1 U4902 ( .A(REG1_REG_11__SCAN_IN), .B(n4318), .S(n4595), .Z(U3529) );
  NAND2_X1 U4903 ( .A1(n4580), .A2(n4281), .ZN(n4283) );
  NAND2_X1 U4904 ( .A1(n4578), .A2(REG0_REG_31__SCAN_IN), .ZN(n4282) );
  OAI211_X1 U4905 ( .C1(n4284), .C2(n4312), .A(n4283), .B(n4282), .ZN(U3517)
         );
  INV_X1 U4906 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4285) );
  MUX2_X1 U4907 ( .A(n4285), .B(n4361), .S(n4580), .Z(n4286) );
  OAI21_X1 U4908 ( .B1(n4287), .B2(n4312), .A(n4286), .ZN(U3516) );
  MUX2_X1 U4909 ( .A(REG0_REG_29__SCAN_IN), .B(n4288), .S(n4580), .Z(U3515) );
  MUX2_X1 U4910 ( .A(REG0_REG_27__SCAN_IN), .B(n4289), .S(n4580), .Z(U3513) );
  INV_X1 U4911 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4291) );
  MUX2_X1 U4912 ( .A(n4291), .B(n4290), .S(n4580), .Z(n4292) );
  OAI21_X1 U4913 ( .B1(n4293), .B2(n4312), .A(n4292), .ZN(U3512) );
  MUX2_X1 U4914 ( .A(REG0_REG_25__SCAN_IN), .B(n4294), .S(n4580), .Z(U3511) );
  INV_X1 U4915 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4296) );
  MUX2_X1 U4916 ( .A(n4296), .B(n4295), .S(n4580), .Z(n4297) );
  OAI21_X1 U4917 ( .B1(n4298), .B2(n4312), .A(n4297), .ZN(U3510) );
  INV_X1 U4918 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4300) );
  MUX2_X1 U4919 ( .A(n4300), .B(n4299), .S(n4580), .Z(n4301) );
  OAI21_X1 U4920 ( .B1(n4302), .B2(n4312), .A(n4301), .ZN(U3509) );
  MUX2_X1 U4921 ( .A(REG0_REG_22__SCAN_IN), .B(n4303), .S(n4580), .Z(U3508) );
  MUX2_X1 U4922 ( .A(REG0_REG_21__SCAN_IN), .B(n4304), .S(n4580), .Z(U3507) );
  INV_X1 U4923 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4306) );
  MUX2_X1 U4924 ( .A(n4306), .B(n4305), .S(n4580), .Z(n4307) );
  OAI21_X1 U4925 ( .B1(n4308), .B2(n4312), .A(n4307), .ZN(U3506) );
  INV_X1 U4926 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4310) );
  MUX2_X1 U4927 ( .A(n4310), .B(n4309), .S(n4580), .Z(n4311) );
  OAI21_X1 U4928 ( .B1(n4313), .B2(n4312), .A(n4311), .ZN(U3505) );
  MUX2_X1 U4929 ( .A(REG0_REG_18__SCAN_IN), .B(n4314), .S(n4580), .Z(U3503) );
  MUX2_X1 U4930 ( .A(REG0_REG_17__SCAN_IN), .B(n4315), .S(n4580), .Z(U3501) );
  MUX2_X1 U4931 ( .A(REG0_REG_16__SCAN_IN), .B(n4316), .S(n4580), .Z(U3499) );
  MUX2_X1 U4932 ( .A(REG0_REG_14__SCAN_IN), .B(n4317), .S(n4580), .Z(U3495) );
  MUX2_X1 U4933 ( .A(REG0_REG_11__SCAN_IN), .B(n4318), .S(n4580), .Z(U3489) );
  MUX2_X1 U4934 ( .A(n4320), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4935 ( .A(DATAI_28_), .B(n4321), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4936 ( .A(DATAI_27_), .B(n4322), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4937 ( .A(n4323), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4938 ( .A(DATAI_25_), .B(n4324), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4939 ( .A(DATAI_22_), .B(n4325), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4940 ( .A(DATAI_20_), .B(n4326), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4941 ( .A(DATAI_19_), .B(n4327), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4942 ( .A(n4328), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U4943 ( .A(n4329), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4944 ( .A(DATAI_4_), .B(n4330), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4945 ( .A(DATAI_3_), .B(n4337), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4946 ( .A(n4331), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI21_X1 U4947 ( .B1(n4980), .B2(ADDR_REG_3__SCAN_IN), .A(n4332), .ZN(n4341)
         );
  OAI211_X1 U4948 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4334), .A(n4479), .B(n4333), 
        .ZN(n4340) );
  OAI211_X1 U4949 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4336), .A(n4985), .B(n4335), 
        .ZN(n4339) );
  NAND2_X1 U4950 ( .A1(n4456), .A2(n4337), .ZN(n4338) );
  NAND4_X1 U4951 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(U3243)
         );
  INV_X1 U4952 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4342) );
  NOR2_X1 U4953 ( .A1(STATE_REG_SCAN_IN), .A2(n4342), .ZN(n4460) );
  OAI22_X1 U4954 ( .A1(n3705), .A2(n4345), .B1(n4344), .B2(n4343), .ZN(n4346)
         );
  AOI211_X1 U4955 ( .C1(n4348), .C2(n4347), .A(n4460), .B(n4346), .ZN(n4356)
         );
  INV_X1 U4956 ( .A(n3710), .ZN(n4350) );
  OAI21_X1 U4957 ( .B1(n4350), .B2(n4349), .A(n3711), .ZN(n4352) );
  XNOR2_X1 U4958 ( .A(n4352), .B(n4351), .ZN(n4354) );
  NAND2_X1 U4959 ( .A1(n4354), .A2(n4353), .ZN(n4355) );
  OAI211_X1 U4960 ( .C1(n4358), .C2(n4357), .A(n4356), .B(n4355), .ZN(U3223)
         );
  AOI22_X1 U4961 ( .A1(n4359), .A2(n4504), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4200), .ZN(n4360) );
  OAI21_X1 U4962 ( .B1(n4507), .B2(n4361), .A(n4360), .ZN(U3261) );
  INV_X1 U4963 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4581) );
  AOI21_X1 U4964 ( .B1(n4581), .B2(n4363), .A(n4362), .ZN(n4364) );
  XOR2_X1 U4965 ( .A(n4364), .B(n2308), .Z(n4366) );
  AOI22_X1 U4966 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4980), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4365) );
  OAI21_X1 U4967 ( .B1(n4367), .B2(n4366), .A(n4365), .ZN(U3240) );
  INV_X1 U4968 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4820) );
  OAI211_X1 U4969 ( .C1(n4370), .C2(n4369), .A(n4985), .B(n4368), .ZN(n4371)
         );
  OAI21_X1 U4970 ( .B1(n4820), .B2(n4459), .A(n4371), .ZN(n4372) );
  NOR2_X1 U4971 ( .A1(n4373), .A2(n4372), .ZN(n4378) );
  OAI211_X1 U4972 ( .C1(n4376), .C2(n4375), .A(n4479), .B(n4374), .ZN(n4377)
         );
  OAI211_X1 U4973 ( .C1(n4989), .C2(n4526), .A(n4378), .B(n4377), .ZN(U3245)
         );
  AOI21_X1 U4974 ( .B1(n4980), .B2(ADDR_REG_6__SCAN_IN), .A(n4379), .ZN(n4380)
         );
  OAI21_X1 U4975 ( .B1(n4989), .B2(n4381), .A(n4380), .ZN(n4382) );
  INV_X1 U4976 ( .A(n4382), .ZN(n4389) );
  OAI211_X1 U4977 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4384), .A(n4479), .B(n4383), 
        .ZN(n4388) );
  OAI211_X1 U4978 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4386), .A(n4985), .B(n4385), 
        .ZN(n4387) );
  NAND3_X1 U4979 ( .A1(n4389), .A2(n4388), .A3(n4387), .ZN(U3246) );
  AOI21_X1 U4980 ( .B1(n4837), .B2(n4401), .A(n4390), .ZN(n4393) );
  OAI21_X1 U4981 ( .B1(n4393), .B2(n4392), .A(n4479), .ZN(n4391) );
  AOI21_X1 U4982 ( .B1(n4393), .B2(n4392), .A(n4391), .ZN(n4395) );
  AOI211_X1 U4983 ( .C1(n4980), .C2(ADDR_REG_7__SCAN_IN), .A(n4395), .B(n4394), 
        .ZN(n4400) );
  OAI211_X1 U4984 ( .C1(n4398), .C2(n4397), .A(n4985), .B(n4396), .ZN(n4399)
         );
  OAI211_X1 U4985 ( .C1(n4989), .C2(n4401), .A(n4400), .B(n4399), .ZN(U3247)
         );
  AOI211_X1 U4986 ( .C1(n4404), .C2(n4403), .A(n4402), .B(n4975), .ZN(n4405)
         );
  AOI211_X1 U4987 ( .C1(ADDR_REG_8__SCAN_IN), .C2(n4980), .A(n4406), .B(n4405), 
        .ZN(n4410) );
  OAI211_X1 U4988 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4408), .A(n4985), .B(n4407), 
        .ZN(n4409) );
  OAI211_X1 U4989 ( .C1(n4989), .C2(n2404), .A(n4410), .B(n4409), .ZN(U3248)
         );
  AOI211_X1 U4990 ( .C1(n2234), .C2(n4412), .A(n4411), .B(n4975), .ZN(n4413)
         );
  AOI211_X1 U4991 ( .C1(n4980), .C2(ADDR_REG_9__SCAN_IN), .A(n4414), .B(n4413), 
        .ZN(n4419) );
  OAI211_X1 U4992 ( .C1(n4417), .C2(n4416), .A(n4985), .B(n4415), .ZN(n4418)
         );
  OAI211_X1 U4993 ( .C1(n4989), .C2(n4522), .A(n4419), .B(n4418), .ZN(U3249)
         );
  AOI211_X1 U4994 ( .C1(n4836), .C2(n4421), .A(n4420), .B(n4975), .ZN(n4423)
         );
  AOI211_X1 U4995 ( .C1(n4980), .C2(ADDR_REG_10__SCAN_IN), .A(n4423), .B(n4422), .ZN(n4427) );
  OAI211_X1 U4996 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4425), .A(n4985), .B(n4424), .ZN(n4426) );
  OAI211_X1 U4997 ( .C1(n4989), .C2(n3469), .A(n4427), .B(n4426), .ZN(U3250)
         );
  AOI211_X1 U4998 ( .C1(n4430), .C2(n4429), .A(n4428), .B(n4975), .ZN(n4431)
         );
  AOI211_X1 U4999 ( .C1(n4980), .C2(ADDR_REG_11__SCAN_IN), .A(n4432), .B(n4431), .ZN(n4437) );
  OAI211_X1 U5000 ( .C1(n4435), .C2(n4434), .A(n4985), .B(n4433), .ZN(n4436)
         );
  OAI211_X1 U5001 ( .C1(n4989), .C2(n4520), .A(n4437), .B(n4436), .ZN(U3251)
         );
  AOI211_X1 U5002 ( .C1(n4440), .C2(n4439), .A(n4438), .B(n4975), .ZN(n4443)
         );
  INV_X1 U5003 ( .A(n4441), .ZN(n4442) );
  AOI211_X1 U5004 ( .C1(n4980), .C2(ADDR_REG_12__SCAN_IN), .A(n4443), .B(n4442), .ZN(n4447) );
  OAI211_X1 U5005 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4445), .A(n4985), .B(n4444), .ZN(n4446) );
  OAI211_X1 U5006 ( .C1(n4989), .C2(n2310), .A(n4447), .B(n4446), .ZN(U3252)
         );
  INV_X1 U5007 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4923) );
  AOI211_X1 U5008 ( .C1(n4762), .C2(n4449), .A(n4448), .B(n4975), .ZN(n4454)
         );
  AOI211_X1 U5009 ( .C1(n4776), .C2(n4452), .A(n4451), .B(n4450), .ZN(n4453)
         );
  AOI211_X1 U5010 ( .C1(n4456), .C2(n4455), .A(n4454), .B(n4453), .ZN(n4458)
         );
  OAI211_X1 U5011 ( .C1(n4459), .C2(n4923), .A(n4458), .B(n4457), .ZN(U3254)
         );
  AOI21_X1 U5012 ( .B1(n4980), .B2(ADDR_REG_16__SCAN_IN), .A(n4460), .ZN(n4470) );
  OAI21_X1 U5013 ( .B1(n4463), .B2(n4462), .A(n4461), .ZN(n4468) );
  OAI21_X1 U5014 ( .B1(n4466), .B2(n4465), .A(n4464), .ZN(n4467) );
  AOI22_X1 U5015 ( .A1(n4985), .A2(n4468), .B1(n4479), .B2(n4467), .ZN(n4469)
         );
  OAI211_X1 U5016 ( .C1(n4515), .C2(n4989), .A(n4470), .B(n4469), .ZN(U3256)
         );
  AOI21_X1 U5017 ( .B1(n4980), .B2(ADDR_REG_17__SCAN_IN), .A(n4471), .ZN(n4482) );
  OAI21_X1 U5018 ( .B1(n4474), .B2(n4473), .A(n4472), .ZN(n4480) );
  OAI21_X1 U5019 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(n4478) );
  AOI22_X1 U5020 ( .A1(n4985), .A2(n4480), .B1(n4479), .B2(n4478), .ZN(n4481)
         );
  OAI211_X1 U5021 ( .C1(n4513), .C2(n4989), .A(n4482), .B(n4481), .ZN(U3257)
         );
  OR2_X1 U5022 ( .A1(n4492), .A2(n4483), .ZN(n4484) );
  AND2_X1 U5023 ( .A1(n4485), .A2(n4484), .ZN(n4536) );
  AOI22_X1 U5024 ( .A1(n2867), .A2(n4487), .B1(n4500), .B2(n4486), .ZN(n4488)
         );
  OAI21_X1 U5025 ( .B1(n4490), .B2(n4489), .A(n4488), .ZN(n4497) );
  NAND2_X1 U5026 ( .A1(n4492), .A2(n4491), .ZN(n4494) );
  AOI21_X1 U5027 ( .B1(n4495), .B2(n4494), .A(n4493), .ZN(n4496) );
  AOI211_X1 U5028 ( .C1(n4536), .C2(n4498), .A(n4497), .B(n4496), .ZN(n4538)
         );
  AOI22_X1 U5029 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4507), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4499), .ZN(n4506) );
  NAND2_X1 U5030 ( .A1(n4500), .A2(n4533), .ZN(n4501) );
  AND2_X1 U5031 ( .A1(n4502), .A2(n4501), .ZN(n4535) );
  AOI22_X1 U5032 ( .A1(n4504), .A2(n4535), .B1(n4503), .B2(n4536), .ZN(n4505)
         );
  OAI211_X1 U5033 ( .C1(n4507), .C2(n4538), .A(n4506), .B(n4505), .ZN(U3289)
         );
  AND2_X1 U5034 ( .A1(D_REG_31__SCAN_IN), .A2(n4509), .ZN(U3291) );
  INV_X1 U5035 ( .A(D_REG_30__SCAN_IN), .ZN(n4743) );
  NOR2_X1 U5036 ( .A1(n4508), .A2(n4743), .ZN(U3292) );
  AND2_X1 U5037 ( .A1(D_REG_29__SCAN_IN), .A2(n4509), .ZN(U3293) );
  AND2_X1 U5038 ( .A1(D_REG_28__SCAN_IN), .A2(n4509), .ZN(U3294) );
  INV_X1 U5039 ( .A(D_REG_27__SCAN_IN), .ZN(n4843) );
  NOR2_X1 U5040 ( .A1(n4508), .A2(n4843), .ZN(U3295) );
  INV_X1 U5041 ( .A(D_REG_26__SCAN_IN), .ZN(n4870) );
  NOR2_X1 U5042 ( .A1(n4508), .A2(n4870), .ZN(U3296) );
  AND2_X1 U5043 ( .A1(D_REG_25__SCAN_IN), .A2(n4509), .ZN(U3297) );
  INV_X1 U5044 ( .A(D_REG_24__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U5045 ( .A1(n4508), .A2(n4886), .ZN(U3298) );
  AND2_X1 U5046 ( .A1(D_REG_23__SCAN_IN), .A2(n4509), .ZN(U3299) );
  INV_X1 U5047 ( .A(D_REG_22__SCAN_IN), .ZN(n4859) );
  NOR2_X1 U5048 ( .A1(n4508), .A2(n4859), .ZN(U3300) );
  AND2_X1 U5049 ( .A1(D_REG_21__SCAN_IN), .A2(n4509), .ZN(U3301) );
  AND2_X1 U5050 ( .A1(D_REG_20__SCAN_IN), .A2(n4509), .ZN(U3302) );
  AND2_X1 U5051 ( .A1(D_REG_19__SCAN_IN), .A2(n4509), .ZN(U3303) );
  AND2_X1 U5052 ( .A1(D_REG_18__SCAN_IN), .A2(n4509), .ZN(U3304) );
  AND2_X1 U5053 ( .A1(D_REG_17__SCAN_IN), .A2(n4509), .ZN(U3305) );
  INV_X1 U5054 ( .A(D_REG_16__SCAN_IN), .ZN(n4858) );
  NOR2_X1 U5055 ( .A1(n4508), .A2(n4858), .ZN(U3306) );
  INV_X1 U5056 ( .A(D_REG_15__SCAN_IN), .ZN(n4735) );
  NOR2_X1 U5057 ( .A1(n4508), .A2(n4735), .ZN(U3307) );
  AND2_X1 U5058 ( .A1(D_REG_14__SCAN_IN), .A2(n4509), .ZN(U3308) );
  AND2_X1 U5059 ( .A1(D_REG_13__SCAN_IN), .A2(n4509), .ZN(U3309) );
  AND2_X1 U5060 ( .A1(D_REG_12__SCAN_IN), .A2(n4509), .ZN(U3310) );
  AND2_X1 U5061 ( .A1(D_REG_11__SCAN_IN), .A2(n4509), .ZN(U3311) );
  INV_X1 U5062 ( .A(D_REG_10__SCAN_IN), .ZN(n4736) );
  NOR2_X1 U5063 ( .A1(n4508), .A2(n4736), .ZN(U3312) );
  AND2_X1 U5064 ( .A1(D_REG_9__SCAN_IN), .A2(n4509), .ZN(U3313) );
  AND2_X1 U5065 ( .A1(n4509), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  AND2_X1 U5066 ( .A1(D_REG_7__SCAN_IN), .A2(n4509), .ZN(U3315) );
  AND2_X1 U5067 ( .A1(n4509), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  INV_X1 U5068 ( .A(D_REG_5__SCAN_IN), .ZN(n4889) );
  NOR2_X1 U5069 ( .A1(n4508), .A2(n4889), .ZN(U3317) );
  AND2_X1 U5070 ( .A1(D_REG_4__SCAN_IN), .A2(n4509), .ZN(U3318) );
  AND2_X1 U5071 ( .A1(D_REG_3__SCAN_IN), .A2(n4509), .ZN(U3319) );
  AND2_X1 U5072 ( .A1(D_REG_2__SCAN_IN), .A2(n4509), .ZN(U3320) );
  INV_X1 U5073 ( .A(DATAI_23_), .ZN(n4511) );
  AOI21_X1 U5074 ( .B1(U3149), .B2(n4511), .A(n4510), .ZN(U3329) );
  AOI22_X1 U5075 ( .A1(STATE_REG_SCAN_IN), .A2(n4513), .B1(n4512), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5076 ( .A(DATAI_16_), .ZN(n4514) );
  AOI22_X1 U5077 ( .A1(STATE_REG_SCAN_IN), .A2(n4515), .B1(n4514), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5078 ( .A1(U3149), .A2(n4516), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4517) );
  INV_X1 U5079 ( .A(n4517), .ZN(U3337) );
  INV_X1 U5080 ( .A(DATAI_14_), .ZN(n4709) );
  AOI22_X1 U5081 ( .A1(STATE_REG_SCAN_IN), .A2(n4518), .B1(n4709), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5082 ( .A(DATAI_12_), .ZN(n4519) );
  AOI22_X1 U5083 ( .A1(STATE_REG_SCAN_IN), .A2(n2310), .B1(n4519), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5084 ( .A(DATAI_11_), .ZN(n4708) );
  AOI22_X1 U5085 ( .A1(STATE_REG_SCAN_IN), .A2(n4520), .B1(n4708), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5086 ( .A(DATAI_10_), .ZN(n4907) );
  AOI22_X1 U5087 ( .A1(STATE_REG_SCAN_IN), .A2(n3469), .B1(n4907), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5088 ( .A(DATAI_9_), .ZN(n4521) );
  AOI22_X1 U5089 ( .A1(STATE_REG_SCAN_IN), .A2(n4522), .B1(n4521), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5090 ( .A(DATAI_8_), .ZN(n4523) );
  AOI22_X1 U5091 ( .A1(STATE_REG_SCAN_IN), .A2(n2404), .B1(n4523), .B2(U3149), 
        .ZN(U3344) );
  OAI22_X1 U5092 ( .A1(U3149), .A2(n4524), .B1(DATAI_7_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4525) );
  INV_X1 U5093 ( .A(n4525), .ZN(U3345) );
  INV_X1 U5094 ( .A(DATAI_5_), .ZN(n4823) );
  AOI22_X1 U5095 ( .A1(STATE_REG_SCAN_IN), .A2(n4526), .B1(n4823), .B2(U3149), 
        .ZN(U3347) );
  OAI22_X1 U5096 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4527) );
  INV_X1 U5097 ( .A(n4527), .ZN(U3352) );
  NOR2_X1 U5098 ( .A1(n4529), .A2(n4528), .ZN(n4532) );
  INV_X1 U5099 ( .A(n4530), .ZN(n4531) );
  AOI211_X1 U5100 ( .C1(n4533), .C2(n2482), .A(n4532), .B(n4531), .ZN(n4582)
         );
  INV_X1 U5101 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5102 ( .A1(n4580), .A2(n4582), .B1(n4534), .B2(n4578), .ZN(U3467)
         );
  AOI22_X1 U5103 ( .A1(n4536), .A2(n4566), .B1(n4577), .B2(n4535), .ZN(n4537)
         );
  AND2_X1 U5104 ( .A1(n4538), .A2(n4537), .ZN(n4583) );
  INV_X1 U5105 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5106 ( .A1(n4580), .A2(n4583), .B1(n4539), .B2(n4578), .ZN(U3469)
         );
  NOR3_X1 U5107 ( .A1(n4541), .A2(n4540), .A3(n4560), .ZN(n4543) );
  AOI211_X1 U5108 ( .C1(n4566), .C2(n4544), .A(n4543), .B(n4542), .ZN(n4585)
         );
  INV_X1 U5109 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5110 ( .A1(n4580), .A2(n4585), .B1(n4545), .B2(n4578), .ZN(U3471)
         );
  NOR2_X1 U5111 ( .A1(n4546), .A2(n4560), .ZN(n4547) );
  AOI21_X1 U5112 ( .B1(n4548), .B2(n4566), .A(n4547), .ZN(n4549) );
  AND2_X1 U5113 ( .A1(n4550), .A2(n4549), .ZN(n4587) );
  INV_X1 U5114 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4904) );
  AOI22_X1 U5115 ( .A1(n4580), .A2(n4587), .B1(n4904), .B2(n4578), .ZN(U3473)
         );
  INV_X1 U5116 ( .A(n4551), .ZN(n4553) );
  AOI211_X1 U5117 ( .C1(n4554), .C2(n4566), .A(n4553), .B(n4552), .ZN(n4588)
         );
  INV_X1 U5118 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5119 ( .A1(n4580), .A2(n4588), .B1(n4555), .B2(n4578), .ZN(U3475)
         );
  NOR2_X1 U5120 ( .A1(n4556), .A2(n4572), .ZN(n4557) );
  AOI211_X1 U5121 ( .C1(n4577), .C2(n4559), .A(n4558), .B(n4557), .ZN(n4589)
         );
  INV_X1 U5122 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U5123 ( .A1(n4580), .A2(n4589), .B1(n4742), .B2(n4578), .ZN(U3477)
         );
  NOR3_X1 U5124 ( .A1(n4562), .A2(n4561), .A3(n4560), .ZN(n4564) );
  AOI211_X1 U5125 ( .C1(n4566), .C2(n4565), .A(n4564), .B(n4563), .ZN(n4591)
         );
  INV_X1 U5126 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5127 ( .A1(n4580), .A2(n4591), .B1(n4745), .B2(n4578), .ZN(U3479)
         );
  AOI211_X1 U5128 ( .C1(n4570), .C2(n4569), .A(n4568), .B(n4567), .ZN(n4592)
         );
  INV_X1 U5129 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5130 ( .A1(n4580), .A2(n4592), .B1(n4571), .B2(n4578), .ZN(U3481)
         );
  NOR2_X1 U5131 ( .A1(n4573), .A2(n4572), .ZN(n4574) );
  AOI211_X1 U5132 ( .C1(n4577), .C2(n4576), .A(n4575), .B(n4574), .ZN(n4594)
         );
  INV_X1 U5133 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5134 ( .A1(n4580), .A2(n4594), .B1(n4579), .B2(n4578), .ZN(U3485)
         );
  AOI22_X1 U5135 ( .A1(n4595), .A2(n4582), .B1(n4581), .B2(n4593), .ZN(U3518)
         );
  AOI22_X1 U5136 ( .A1(n4595), .A2(n4583), .B1(n2415), .B2(n4593), .ZN(U3519)
         );
  AOI22_X1 U5137 ( .A1(n4595), .A2(n4585), .B1(n4584), .B2(n4593), .ZN(U3520)
         );
  INV_X1 U5138 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5139 ( .A1(n4595), .A2(n4587), .B1(n4586), .B2(n4593), .ZN(U3521)
         );
  AOI22_X1 U5140 ( .A1(n4595), .A2(n4588), .B1(n3459), .B2(n4593), .ZN(U3522)
         );
  AOI22_X1 U5141 ( .A1(n4595), .A2(n4589), .B1(n4890), .B2(n4593), .ZN(U3523)
         );
  INV_X1 U5142 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U5143 ( .A1(n4595), .A2(n4591), .B1(n4590), .B2(n4593), .ZN(U3524)
         );
  AOI22_X1 U5144 ( .A1(n4595), .A2(n4592), .B1(n4837), .B2(n4593), .ZN(U3525)
         );
  INV_X1 U5145 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4914) );
  AOI22_X1 U5146 ( .A1(n4595), .A2(n4594), .B1(n4914), .B2(n4593), .ZN(U3527)
         );
  OAI22_X1 U5147 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput52), .B1(keyinput44), 
        .B2(REG3_REG_17__SCAN_IN), .ZN(n4596) );
  AOI221_X1 U5148 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput52), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput44), .A(n4596), .ZN(n4603) );
  OAI22_X1 U5149 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput20), .B1(keyinput108), .B2(DATAO_REG_24__SCAN_IN), .ZN(n4597) );
  AOI221_X1 U5150 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput20), .C1(
        DATAO_REG_24__SCAN_IN), .C2(keyinput108), .A(n4597), .ZN(n4602) );
  OAI22_X1 U5151 ( .A1(DATAI_21_), .A2(keyinput40), .B1(keyinput36), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4598) );
  AOI221_X1 U5152 ( .B1(DATAI_21_), .B2(keyinput40), .C1(DATAO_REG_30__SCAN_IN), .C2(keyinput36), .A(n4598), .ZN(n4601) );
  OAI22_X1 U5153 ( .A1(REG2_REG_26__SCAN_IN), .A2(keyinput4), .B1(keyinput28), 
        .B2(REG1_REG_22__SCAN_IN), .ZN(n4599) );
  AOI221_X1 U5154 ( .B1(REG2_REG_26__SCAN_IN), .B2(keyinput4), .C1(
        REG1_REG_22__SCAN_IN), .C2(keyinput28), .A(n4599), .ZN(n4600) );
  NAND4_X1 U5155 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(n4631)
         );
  OAI22_X1 U5156 ( .A1(REG2_REG_0__SCAN_IN), .A2(keyinput32), .B1(keyinput80), 
        .B2(ADDR_REG_16__SCAN_IN), .ZN(n4604) );
  AOI221_X1 U5157 ( .B1(REG2_REG_0__SCAN_IN), .B2(keyinput32), .C1(
        ADDR_REG_16__SCAN_IN), .C2(keyinput80), .A(n4604), .ZN(n4611) );
  OAI22_X1 U5158 ( .A1(REG0_REG_15__SCAN_IN), .A2(keyinput116), .B1(
        keyinput111), .B2(REG0_REG_5__SCAN_IN), .ZN(n4605) );
  AOI221_X1 U5159 ( .B1(REG0_REG_15__SCAN_IN), .B2(keyinput116), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput111), .A(n4605), .ZN(n4610) );
  OAI22_X1 U5160 ( .A1(REG1_REG_29__SCAN_IN), .A2(keyinput72), .B1(keyinput25), 
        .B2(D_REG_10__SCAN_IN), .ZN(n4606) );
  AOI221_X1 U5161 ( .B1(REG1_REG_29__SCAN_IN), .B2(keyinput72), .C1(
        D_REG_10__SCAN_IN), .C2(keyinput25), .A(n4606), .ZN(n4609) );
  OAI22_X1 U5162 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput48), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput84), .ZN(n4607) );
  AOI221_X1 U5163 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput48), .C1(keyinput84), 
        .C2(REG0_REG_6__SCAN_IN), .A(n4607), .ZN(n4608) );
  NAND4_X1 U5164 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4630)
         );
  OAI22_X1 U5165 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput125), .B1(keyinput73), .B2(REG0_REG_22__SCAN_IN), .ZN(n4612) );
  AOI221_X1 U5166 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput125), .C1(
        REG0_REG_22__SCAN_IN), .C2(keyinput73), .A(n4612), .ZN(n4619) );
  OAI22_X1 U5167 ( .A1(REG3_REG_18__SCAN_IN), .A2(keyinput77), .B1(keyinput81), 
        .B2(REG3_REG_10__SCAN_IN), .ZN(n4613) );
  AOI221_X1 U5168 ( .B1(REG3_REG_18__SCAN_IN), .B2(keyinput77), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput81), .A(n4613), .ZN(n4618) );
  OAI22_X1 U5169 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput113), .B1(DATAI_18_), 
        .B2(keyinput37), .ZN(n4614) );
  AOI221_X1 U5170 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput113), .C1(keyinput37), 
        .C2(DATAI_18_), .A(n4614), .ZN(n4617) );
  OAI22_X1 U5171 ( .A1(REG2_REG_28__SCAN_IN), .A2(keyinput109), .B1(
        keyinput121), .B2(DATAI_14_), .ZN(n4615) );
  AOI221_X1 U5172 ( .B1(REG2_REG_28__SCAN_IN), .B2(keyinput109), .C1(DATAI_14_), .C2(keyinput121), .A(n4615), .ZN(n4616) );
  NAND4_X1 U5173 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4629)
         );
  OAI22_X1 U5174 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput19), .B1(
        REG1_REG_0__SCAN_IN), .B2(keyinput27), .ZN(n4620) );
  AOI221_X1 U5175 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput19), .C1(keyinput27), 
        .C2(REG1_REG_0__SCAN_IN), .A(n4620), .ZN(n4627) );
  OAI22_X1 U5176 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput23), .B1(keyinput12), 
        .B2(DATAI_2_), .ZN(n4621) );
  AOI221_X1 U5177 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput23), .C1(DATAI_2_), 
        .C2(keyinput12), .A(n4621), .ZN(n4626) );
  OAI22_X1 U5178 ( .A1(D_REG_30__SCAN_IN), .A2(keyinput11), .B1(
        REG1_REG_14__SCAN_IN), .B2(keyinput97), .ZN(n4622) );
  AOI221_X1 U5179 ( .B1(D_REG_30__SCAN_IN), .B2(keyinput11), .C1(keyinput97), 
        .C2(REG1_REG_14__SCAN_IN), .A(n4622), .ZN(n4625) );
  OAI22_X1 U5180 ( .A1(DATAI_20_), .A2(keyinput7), .B1(keyinput31), .B2(
        REG2_REG_2__SCAN_IN), .ZN(n4623) );
  AOI221_X1 U5181 ( .B1(DATAI_20_), .B2(keyinput7), .C1(REG2_REG_2__SCAN_IN), 
        .C2(keyinput31), .A(n4623), .ZN(n4624) );
  NAND4_X1 U5182 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4628)
         );
  NOR4_X1 U5183 ( .A1(n4631), .A2(n4630), .A3(n4629), .A4(n4628), .ZN(n4974)
         );
  AOI22_X1 U5184 ( .A1(DATAI_19_), .A2(keyinput189), .B1(DATAI_20_), .B2(
        keyinput135), .ZN(n4632) );
  OAI221_X1 U5185 ( .B1(DATAI_19_), .B2(keyinput189), .C1(DATAI_20_), .C2(
        keyinput135), .A(n4632), .ZN(n4639) );
  AOI22_X1 U5186 ( .A1(DATAI_18_), .A2(keyinput165), .B1(DATAI_17_), .B2(
        keyinput136), .ZN(n4633) );
  OAI221_X1 U5187 ( .B1(DATAI_18_), .B2(keyinput165), .C1(DATAI_17_), .C2(
        keyinput136), .A(n4633), .ZN(n4638) );
  AOI22_X1 U5188 ( .A1(DATAI_6_), .A2(keyinput251), .B1(DATAI_10_), .B2(
        keyinput157), .ZN(n4634) );
  OAI221_X1 U5189 ( .B1(DATAI_6_), .B2(keyinput251), .C1(DATAI_10_), .C2(
        keyinput157), .A(n4634), .ZN(n4637) );
  AOI22_X1 U5190 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput253), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput177), .ZN(n4635) );
  OAI221_X1 U5191 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput253), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput177), .A(n4635), .ZN(n4636) );
  NOR4_X1 U5192 ( .A1(n4639), .A2(n4638), .A3(n4637), .A4(n4636), .ZN(n4667)
         );
  AOI22_X1 U5193 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput209), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput172), .ZN(n4640) );
  OAI221_X1 U5194 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput209), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput172), .A(n4640), .ZN(n4647) );
  AOI22_X1 U5195 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput231), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput184), .ZN(n4641) );
  OAI221_X1 U5196 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput231), .C1(
        IR_REG_14__SCAN_IN), .C2(keyinput184), .A(n4641), .ZN(n4646) );
  AOI22_X1 U5197 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput241), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput176), .ZN(n4642) );
  OAI221_X1 U5198 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput241), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput176), .A(n4642), .ZN(n4645) );
  AOI22_X1 U5199 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput158), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput183), .ZN(n4643) );
  OAI221_X1 U5200 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput158), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput183), .A(n4643), .ZN(n4644) );
  NOR4_X1 U5201 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4666)
         );
  AOI22_X1 U5202 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput171), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput180), .ZN(n4648) );
  OAI221_X1 U5203 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput171), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput180), .A(n4648), .ZN(n4655) );
  AOI22_X1 U5204 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput222), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput228), .ZN(n4649) );
  OAI221_X1 U5205 ( .B1(D_REG_16__SCAN_IN), .B2(keyinput222), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput228), .A(n4649), .ZN(n4654) );
  AOI22_X1 U5206 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput131), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput199), .ZN(n4650) );
  OAI221_X1 U5207 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput131), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput199), .A(n4650), .ZN(n4653) );
  AOI22_X1 U5208 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput174), .B1(
        REG0_REG_9__SCAN_IN), .B2(keyinput161), .ZN(n4651) );
  OAI221_X1 U5209 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput174), .C1(
        REG0_REG_9__SCAN_IN), .C2(keyinput161), .A(n4651), .ZN(n4652) );
  NOR4_X1 U5210 ( .A1(n4655), .A2(n4654), .A3(n4653), .A4(n4652), .ZN(n4665)
         );
  AOI22_X1 U5211 ( .A1(REG0_REG_12__SCAN_IN), .A2(keyinput238), .B1(
        REG0_REG_15__SCAN_IN), .B2(keyinput244), .ZN(n4656) );
  OAI221_X1 U5212 ( .B1(REG0_REG_12__SCAN_IN), .B2(keyinput238), .C1(
        REG0_REG_15__SCAN_IN), .C2(keyinput244), .A(n4656), .ZN(n4663) );
  AOI22_X1 U5213 ( .A1(REG0_REG_16__SCAN_IN), .A2(keyinput149), .B1(
        REG0_REG_21__SCAN_IN), .B2(keyinput250), .ZN(n4657) );
  OAI221_X1 U5214 ( .B1(REG0_REG_16__SCAN_IN), .B2(keyinput149), .C1(
        REG0_REG_21__SCAN_IN), .C2(keyinput250), .A(n4657), .ZN(n4662) );
  AOI22_X1 U5215 ( .A1(REG0_REG_23__SCAN_IN), .A2(keyinput211), .B1(
        REG0_REG_26__SCAN_IN), .B2(keyinput247), .ZN(n4658) );
  OAI221_X1 U5216 ( .B1(REG0_REG_23__SCAN_IN), .B2(keyinput211), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput247), .A(n4658), .ZN(n4661) );
  AOI22_X1 U5217 ( .A1(REG1_REG_0__SCAN_IN), .A2(keyinput155), .B1(
        REG1_REG_1__SCAN_IN), .B2(keyinput226), .ZN(n4659) );
  OAI221_X1 U5218 ( .B1(REG1_REG_0__SCAN_IN), .B2(keyinput155), .C1(
        REG1_REG_1__SCAN_IN), .C2(keyinput226), .A(n4659), .ZN(n4660) );
  NOR4_X1 U5219 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4664)
         );
  NAND4_X1 U5220 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4809)
         );
  AOI22_X1 U5221 ( .A1(REG1_REG_7__SCAN_IN), .A2(keyinput196), .B1(
        REG1_REG_8__SCAN_IN), .B2(keyinput150), .ZN(n4668) );
  OAI221_X1 U5222 ( .B1(REG1_REG_7__SCAN_IN), .B2(keyinput196), .C1(
        REG1_REG_8__SCAN_IN), .C2(keyinput150), .A(n4668), .ZN(n4675) );
  AOI22_X1 U5223 ( .A1(REG1_REG_16__SCAN_IN), .A2(keyinput194), .B1(
        REG1_REG_9__SCAN_IN), .B2(keyinput145), .ZN(n4669) );
  OAI221_X1 U5224 ( .B1(REG1_REG_16__SCAN_IN), .B2(keyinput194), .C1(
        REG1_REG_9__SCAN_IN), .C2(keyinput145), .A(n4669), .ZN(n4674) );
  AOI22_X1 U5225 ( .A1(REG1_REG_15__SCAN_IN), .A2(keyinput234), .B1(
        REG1_REG_20__SCAN_IN), .B2(keyinput246), .ZN(n4670) );
  OAI221_X1 U5226 ( .B1(REG1_REG_15__SCAN_IN), .B2(keyinput234), .C1(
        REG1_REG_20__SCAN_IN), .C2(keyinput246), .A(n4670), .ZN(n4673) );
  AOI22_X1 U5227 ( .A1(REG1_REG_23__SCAN_IN), .A2(keyinput192), .B1(
        REG1_REG_27__SCAN_IN), .B2(keyinput227), .ZN(n4671) );
  OAI221_X1 U5228 ( .B1(REG1_REG_23__SCAN_IN), .B2(keyinput192), .C1(
        REG1_REG_27__SCAN_IN), .C2(keyinput227), .A(n4671), .ZN(n4672) );
  NOR4_X1 U5229 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4703)
         );
  AOI22_X1 U5230 ( .A1(REG2_REG_4__SCAN_IN), .A2(keyinput206), .B1(
        REG2_REG_0__SCAN_IN), .B2(keyinput160), .ZN(n4676) );
  OAI221_X1 U5231 ( .B1(REG2_REG_4__SCAN_IN), .B2(keyinput206), .C1(
        REG2_REG_0__SCAN_IN), .C2(keyinput160), .A(n4676), .ZN(n4683) );
  AOI22_X1 U5232 ( .A1(REG2_REG_8__SCAN_IN), .A2(keyinput154), .B1(
        REG2_REG_13__SCAN_IN), .B2(keyinput248), .ZN(n4677) );
  OAI221_X1 U5233 ( .B1(REG2_REG_8__SCAN_IN), .B2(keyinput154), .C1(
        REG2_REG_13__SCAN_IN), .C2(keyinput248), .A(n4677), .ZN(n4682) );
  AOI22_X1 U5234 ( .A1(REG2_REG_11__SCAN_IN), .A2(keyinput197), .B1(
        REG2_REG_15__SCAN_IN), .B2(keyinput173), .ZN(n4678) );
  OAI221_X1 U5235 ( .B1(REG2_REG_11__SCAN_IN), .B2(keyinput197), .C1(
        REG2_REG_15__SCAN_IN), .C2(keyinput173), .A(n4678), .ZN(n4681) );
  AOI22_X1 U5236 ( .A1(REG2_REG_18__SCAN_IN), .A2(keyinput204), .B1(
        REG2_REG_22__SCAN_IN), .B2(keyinput133), .ZN(n4679) );
  OAI221_X1 U5237 ( .B1(REG2_REG_18__SCAN_IN), .B2(keyinput204), .C1(
        REG2_REG_22__SCAN_IN), .C2(keyinput133), .A(n4679), .ZN(n4680) );
  NOR4_X1 U5238 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4702)
         );
  AOI22_X1 U5239 ( .A1(ADDR_REG_9__SCAN_IN), .A2(keyinput207), .B1(
        REG2_REG_29__SCAN_IN), .B2(keyinput182), .ZN(n4684) );
  OAI221_X1 U5240 ( .B1(ADDR_REG_9__SCAN_IN), .B2(keyinput207), .C1(
        REG2_REG_29__SCAN_IN), .C2(keyinput182), .A(n4684), .ZN(n4691) );
  AOI22_X1 U5241 ( .A1(ADDR_REG_2__SCAN_IN), .A2(keyinput175), .B1(
        ADDR_REG_4__SCAN_IN), .B2(keyinput198), .ZN(n4685) );
  OAI221_X1 U5242 ( .B1(ADDR_REG_2__SCAN_IN), .B2(keyinput175), .C1(
        ADDR_REG_4__SCAN_IN), .C2(keyinput198), .A(n4685), .ZN(n4690) );
  AOI22_X1 U5243 ( .A1(DATAO_REG_12__SCAN_IN), .A2(keyinput214), .B1(
        DATAO_REG_4__SCAN_IN), .B2(keyinput148), .ZN(n4686) );
  OAI221_X1 U5244 ( .B1(DATAO_REG_12__SCAN_IN), .B2(keyinput214), .C1(
        DATAO_REG_4__SCAN_IN), .C2(keyinput148), .A(n4686), .ZN(n4689) );
  AOI22_X1 U5245 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput164), .B1(
        DATAO_REG_23__SCAN_IN), .B2(keyinput185), .ZN(n4687) );
  OAI221_X1 U5246 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput164), .C1(
        DATAO_REG_23__SCAN_IN), .C2(keyinput185), .A(n4687), .ZN(n4688) );
  NOR4_X1 U5247 ( .A1(n4691), .A2(n4690), .A3(n4689), .A4(n4688), .ZN(n4701)
         );
  AOI22_X1 U5248 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput129), .B1(
        REG3_REG_11__SCAN_IN), .B2(keyinput213), .ZN(n4692) );
  OAI221_X1 U5249 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput129), .C1(
        REG3_REG_11__SCAN_IN), .C2(keyinput213), .A(n4692), .ZN(n4699) );
  AOI22_X1 U5250 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput218), .B1(
        REG3_REG_22__SCAN_IN), .B2(keyinput215), .ZN(n4693) );
  OAI221_X1 U5251 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput218), .C1(
        REG3_REG_22__SCAN_IN), .C2(keyinput215), .A(n4693), .ZN(n4698) );
  AOI22_X1 U5252 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput151), .B1(
        IR_REG_29__SCAN_IN), .B2(keyinput191), .ZN(n4694) );
  OAI221_X1 U5253 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput151), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput191), .A(n4694), .ZN(n4697) );
  AOI22_X1 U5254 ( .A1(ADDR_REG_11__SCAN_IN), .A2(keyinput178), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput130), .ZN(n4695) );
  OAI221_X1 U5255 ( .B1(ADDR_REG_11__SCAN_IN), .B2(keyinput178), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput130), .A(n4695), .ZN(n4696) );
  NOR4_X1 U5256 ( .A1(n4699), .A2(n4698), .A3(n4697), .A4(n4696), .ZN(n4700)
         );
  NAND4_X1 U5257 ( .A1(n4703), .A2(n4702), .A3(n4701), .A4(n4700), .ZN(n4808)
         );
  INV_X1 U5258 ( .A(DATAI_26_), .ZN(n4869) );
  AOI22_X1 U5259 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput138), .B1(n4869), .B2(
        keyinput219), .ZN(n4704) );
  OAI221_X1 U5260 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput138), .C1(n4869), .C2(
        keyinput219), .A(n4704), .ZN(n4715) );
  AOI22_X1 U5261 ( .A1(n4885), .A2(keyinput163), .B1(n4706), .B2(keyinput168), 
        .ZN(n4705) );
  OAI221_X1 U5262 ( .B1(n4885), .B2(keyinput163), .C1(n4706), .C2(keyinput168), 
        .A(n4705), .ZN(n4714) );
  AOI22_X1 U5263 ( .A1(n4709), .A2(keyinput249), .B1(keyinput202), .B2(n4708), 
        .ZN(n4707) );
  OAI221_X1 U5264 ( .B1(n4709), .B2(keyinput249), .C1(n4708), .C2(keyinput202), 
        .A(n4707), .ZN(n4713) );
  INV_X1 U5265 ( .A(DATAI_2_), .ZN(n4711) );
  AOI22_X1 U5266 ( .A1(n4823), .A2(keyinput152), .B1(keyinput140), .B2(n4711), 
        .ZN(n4710) );
  OAI221_X1 U5267 ( .B1(n4823), .B2(keyinput152), .C1(n4711), .C2(keyinput140), 
        .A(n4710), .ZN(n4712) );
  NOR4_X1 U5268 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4755)
         );
  AOI22_X1 U5269 ( .A1(n2337), .A2(keyinput167), .B1(n3136), .B2(keyinput252), 
        .ZN(n4716) );
  OAI221_X1 U5270 ( .B1(n2337), .B2(keyinput167), .C1(n3136), .C2(keyinput252), 
        .A(n4716), .ZN(n4725) );
  AOI22_X1 U5271 ( .A1(n2512), .A2(keyinput170), .B1(n4718), .B2(keyinput181), 
        .ZN(n4717) );
  OAI221_X1 U5272 ( .B1(n2512), .B2(keyinput170), .C1(n4718), .C2(keyinput181), 
        .A(n4717), .ZN(n4724) );
  XOR2_X1 U5273 ( .A(n2308), .B(keyinput235), .Z(n4722) );
  XNOR2_X1 U5274 ( .A(IR_REG_6__SCAN_IN), .B(keyinput233), .ZN(n4721) );
  XNOR2_X1 U5275 ( .A(IR_REG_8__SCAN_IN), .B(keyinput210), .ZN(n4720) );
  XNOR2_X1 U5276 ( .A(IR_REG_13__SCAN_IN), .B(keyinput223), .ZN(n4719) );
  NAND4_X1 U5277 ( .A1(n4722), .A2(n4721), .A3(n4720), .A4(n4719), .ZN(n4723)
         );
  NOR3_X1 U5278 ( .A1(n4725), .A2(n4724), .A3(n4723), .ZN(n4754) );
  XNOR2_X1 U5279 ( .A(n2784), .B(keyinput147), .ZN(n4730) );
  XNOR2_X1 U5280 ( .A(n4726), .B(keyinput128), .ZN(n4729) );
  XNOR2_X1 U5281 ( .A(n4727), .B(keyinput179), .ZN(n4728) );
  NOR3_X1 U5282 ( .A1(n4730), .A2(n4729), .A3(n4728), .ZN(n4733) );
  XNOR2_X1 U5283 ( .A(IR_REG_22__SCAN_IN), .B(keyinput245), .ZN(n4732) );
  XNOR2_X1 U5284 ( .A(IR_REG_20__SCAN_IN), .B(keyinput187), .ZN(n4731) );
  NAND3_X1 U5285 ( .A1(n4733), .A2(n4732), .A3(n4731), .ZN(n4739) );
  AOI22_X1 U5286 ( .A1(n4736), .A2(keyinput153), .B1(n4735), .B2(keyinput254), 
        .ZN(n4734) );
  OAI221_X1 U5287 ( .B1(n4736), .B2(keyinput153), .C1(n4735), .C2(keyinput254), 
        .A(n4734), .ZN(n4738) );
  XNOR2_X1 U5288 ( .A(n4902), .B(keyinput143), .ZN(n4737) );
  NOR3_X1 U5289 ( .A1(n4739), .A2(n4738), .A3(n4737), .ZN(n4753) );
  AOI22_X1 U5290 ( .A1(n4886), .A2(keyinput162), .B1(n4859), .B2(keyinput230), 
        .ZN(n4740) );
  OAI221_X1 U5291 ( .B1(n4886), .B2(keyinput162), .C1(n4859), .C2(keyinput230), 
        .A(n4740), .ZN(n4751) );
  AOI22_X1 U5292 ( .A1(n4743), .A2(keyinput139), .B1(keyinput239), .B2(n4742), 
        .ZN(n4741) );
  OAI221_X1 U5293 ( .B1(n4743), .B2(keyinput139), .C1(n4742), .C2(keyinput239), 
        .A(n4741), .ZN(n4750) );
  AOI22_X1 U5294 ( .A1(n4745), .A2(keyinput212), .B1(n4853), .B2(keyinput255), 
        .ZN(n4744) );
  OAI221_X1 U5295 ( .B1(n4745), .B2(keyinput212), .C1(n4853), .C2(keyinput255), 
        .A(n4744), .ZN(n4749) );
  INV_X1 U5296 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4747) );
  INV_X1 U5297 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4905) );
  AOI22_X1 U5298 ( .A1(n4747), .A2(keyinput169), .B1(n4905), .B2(keyinput134), 
        .ZN(n4746) );
  OAI221_X1 U5299 ( .B1(n4747), .B2(keyinput169), .C1(n4905), .C2(keyinput134), 
        .A(n4746), .ZN(n4748) );
  NOR4_X1 U5300 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n4752)
         );
  NAND4_X1 U5301 ( .A1(n4755), .A2(n4754), .A3(n4753), .A4(n4752), .ZN(n4807)
         );
  INV_X1 U5302 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4758) );
  INV_X1 U5303 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4757) );
  AOI22_X1 U5304 ( .A1(n4758), .A2(keyinput193), .B1(n4757), .B2(keyinput201), 
        .ZN(n4756) );
  OAI221_X1 U5305 ( .B1(n4758), .B2(keyinput193), .C1(n4757), .C2(keyinput201), 
        .A(n4756), .ZN(n4768) );
  AOI22_X1 U5306 ( .A1(n4760), .A2(keyinput146), .B1(keyinput166), .B2(n4890), 
        .ZN(n4759) );
  OAI221_X1 U5307 ( .B1(n4760), .B2(keyinput146), .C1(n4890), .C2(keyinput166), 
        .A(n4759), .ZN(n4767) );
  AOI22_X1 U5308 ( .A1(n4836), .A2(keyinput220), .B1(n4762), .B2(keyinput225), 
        .ZN(n4761) );
  OAI221_X1 U5309 ( .B1(n4836), .B2(keyinput220), .C1(n4762), .C2(keyinput225), 
        .A(n4761), .ZN(n4766) );
  INV_X1 U5310 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5311 ( .A1(n4764), .A2(keyinput156), .B1(n4834), .B2(keyinput188), 
        .ZN(n4763) );
  OAI221_X1 U5312 ( .B1(n4764), .B2(keyinput156), .C1(n4834), .C2(keyinput188), 
        .A(n4763), .ZN(n4765) );
  NOR4_X1 U5313 ( .A1(n4768), .A2(n4767), .A3(n4766), .A4(n4765), .ZN(n4805)
         );
  AOI22_X1 U5314 ( .A1(n4771), .A2(keyinput242), .B1(n4770), .B2(keyinput200), 
        .ZN(n4769) );
  OAI221_X1 U5315 ( .B1(n4771), .B2(keyinput242), .C1(n4770), .C2(keyinput200), 
        .A(n4769), .ZN(n4780) );
  AOI22_X1 U5316 ( .A1(n4773), .A2(keyinput159), .B1(keyinput142), .B2(n3435), 
        .ZN(n4772) );
  OAI221_X1 U5317 ( .B1(n4773), .B2(keyinput159), .C1(n3435), .C2(keyinput142), 
        .A(n4772), .ZN(n4779) );
  AOI22_X1 U5318 ( .A1(n3233), .A2(keyinput217), .B1(keyinput203), .B2(n4880), 
        .ZN(n4774) );
  OAI221_X1 U5319 ( .B1(n3233), .B2(keyinput217), .C1(n4880), .C2(keyinput203), 
        .A(n4774), .ZN(n4778) );
  INV_X1 U5320 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5321 ( .A1(n4776), .A2(keyinput190), .B1(n4915), .B2(keyinput141), 
        .ZN(n4775) );
  OAI221_X1 U5322 ( .B1(n4776), .B2(keyinput190), .C1(n4915), .C2(keyinput141), 
        .A(n4775), .ZN(n4777) );
  NOR4_X1 U5323 ( .A1(n4780), .A2(n4779), .A3(n4778), .A4(n4777), .ZN(n4804)
         );
  INV_X1 U5324 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4824) );
  INV_X1 U5325 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U5326 ( .A1(n4824), .A2(keyinput144), .B1(n4782), .B2(keyinput237), 
        .ZN(n4781) );
  OAI221_X1 U5327 ( .B1(n4824), .B2(keyinput144), .C1(n4782), .C2(keyinput237), 
        .A(n4781), .ZN(n4790) );
  INV_X1 U5328 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4784) );
  INV_X1 U5329 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U5330 ( .A1(n4784), .A2(keyinput208), .B1(n4839), .B2(keyinput232), 
        .ZN(n4783) );
  OAI221_X1 U5331 ( .B1(n4784), .B2(keyinput208), .C1(n4839), .C2(keyinput232), 
        .A(n4783), .ZN(n4789) );
  INV_X1 U5332 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U5333 ( .A1(n4923), .A2(keyinput137), .B1(keyinput229), .B2(n4819), 
        .ZN(n4785) );
  OAI221_X1 U5334 ( .B1(n4923), .B2(keyinput137), .C1(n4819), .C2(keyinput229), 
        .A(n4785), .ZN(n4788) );
  INV_X1 U5335 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5336 ( .A1(n4856), .A2(keyinput243), .B1(keyinput221), .B2(n4820), 
        .ZN(n4786) );
  OAI221_X1 U5337 ( .B1(n4856), .B2(keyinput243), .C1(n4820), .C2(keyinput221), 
        .A(n4786), .ZN(n4787) );
  NOR4_X1 U5338 ( .A1(n4790), .A2(n4789), .A3(n4788), .A4(n4787), .ZN(n4803)
         );
  AOI22_X1 U5339 ( .A1(n4793), .A2(keyinput195), .B1(keyinput186), .B2(n4792), 
        .ZN(n4791) );
  OAI221_X1 U5340 ( .B1(n4793), .B2(keyinput195), .C1(n4792), .C2(keyinput186), 
        .A(n4791), .ZN(n4801) );
  AOI22_X1 U5341 ( .A1(n4840), .A2(keyinput216), .B1(keyinput240), .B2(n4850), 
        .ZN(n4794) );
  OAI221_X1 U5342 ( .B1(n4840), .B2(keyinput216), .C1(n4850), .C2(keyinput240), 
        .A(n4794), .ZN(n4800) );
  AOI22_X1 U5343 ( .A1(n4849), .A2(keyinput224), .B1(keyinput236), .B2(n4796), 
        .ZN(n4795) );
  OAI221_X1 U5344 ( .B1(n4849), .B2(keyinput224), .C1(n4796), .C2(keyinput236), 
        .A(n4795), .ZN(n4799) );
  AOI22_X1 U5345 ( .A1(n2684), .A2(keyinput205), .B1(keyinput132), .B2(n4042), 
        .ZN(n4797) );
  OAI221_X1 U5346 ( .B1(n2684), .B2(keyinput205), .C1(n4042), .C2(keyinput132), 
        .A(n4797), .ZN(n4798) );
  NOR4_X1 U5347 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4802)
         );
  NAND4_X1 U5348 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4806)
         );
  NOR4_X1 U5349 ( .A1(n4809), .A2(n4808), .A3(n4807), .A4(n4806), .ZN(n4935)
         );
  AOI22_X1 U5350 ( .A1(REG0_REG_11__SCAN_IN), .A2(keyinput41), .B1(
        REG0_REG_9__SCAN_IN), .B2(keyinput33), .ZN(n4810) );
  OAI221_X1 U5351 ( .B1(REG0_REG_11__SCAN_IN), .B2(keyinput41), .C1(
        REG0_REG_9__SCAN_IN), .C2(keyinput33), .A(n4810), .ZN(n4817) );
  AOI22_X1 U5352 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput1), .B1(DATAI_19_), 
        .B2(keyinput61), .ZN(n4811) );
  OAI221_X1 U5353 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput1), .C1(DATAI_19_), 
        .C2(keyinput61), .A(n4811), .ZN(n4816) );
  AOI22_X1 U5354 ( .A1(REG0_REG_17__SCAN_IN), .A2(keyinput65), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput49), .ZN(n4812) );
  OAI221_X1 U5355 ( .B1(REG0_REG_17__SCAN_IN), .B2(keyinput65), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput49), .A(n4812), .ZN(n4815) );
  AOI22_X1 U5356 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput53), .B1(n3233), 
        .B2(keyinput89), .ZN(n4813) );
  OAI221_X1 U5357 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput53), .C1(n3233), 
        .C2(keyinput89), .A(n4813), .ZN(n4814) );
  NOR4_X1 U5358 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n4867)
         );
  AOI22_X1 U5359 ( .A1(n4820), .A2(keyinput93), .B1(n4819), .B2(keyinput101), 
        .ZN(n4818) );
  OAI221_X1 U5360 ( .B1(n4820), .B2(keyinput93), .C1(n4819), .C2(keyinput101), 
        .A(n4818), .ZN(n4831) );
  AOI22_X1 U5361 ( .A1(n4823), .A2(keyinput24), .B1(n4822), .B2(keyinput56), 
        .ZN(n4821) );
  OAI221_X1 U5362 ( .B1(n4823), .B2(keyinput24), .C1(n4822), .C2(keyinput56), 
        .A(n4821), .ZN(n4830) );
  XOR2_X1 U5363 ( .A(n4824), .B(keyinput16), .Z(n4828) );
  XNOR2_X1 U5364 ( .A(DATAI_17_), .B(keyinput8), .ZN(n4827) );
  XNOR2_X1 U5365 ( .A(IR_REG_6__SCAN_IN), .B(keyinput105), .ZN(n4826) );
  XNOR2_X1 U5366 ( .A(IR_REG_22__SCAN_IN), .B(keyinput117), .ZN(n4825) );
  NAND4_X1 U5367 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), .ZN(n4829)
         );
  NOR3_X1 U5368 ( .A1(n4831), .A2(n4830), .A3(n4829), .ZN(n4866) );
  INV_X1 U5369 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U5370 ( .A1(n4834), .A2(keyinput60), .B1(keyinput76), .B2(n4833), 
        .ZN(n4832) );
  OAI221_X1 U5371 ( .B1(n4834), .B2(keyinput60), .C1(n4833), .C2(keyinput76), 
        .A(n4832), .ZN(n4847) );
  AOI22_X1 U5372 ( .A1(n4837), .A2(keyinput68), .B1(n4836), .B2(keyinput92), 
        .ZN(n4835) );
  OAI221_X1 U5373 ( .B1(n4837), .B2(keyinput68), .C1(n4836), .C2(keyinput92), 
        .A(n4835), .ZN(n4846) );
  AOI22_X1 U5374 ( .A1(n4840), .A2(keyinput88), .B1(n4839), .B2(keyinput104), 
        .ZN(n4838) );
  OAI221_X1 U5375 ( .B1(n4840), .B2(keyinput88), .C1(n4839), .C2(keyinput104), 
        .A(n4838), .ZN(n4845) );
  AOI22_X1 U5376 ( .A1(n4843), .A2(keyinput100), .B1(keyinput120), .B2(n4842), 
        .ZN(n4841) );
  OAI221_X1 U5377 ( .B1(n4843), .B2(keyinput100), .C1(n4842), .C2(keyinput120), 
        .A(n4841), .ZN(n4844) );
  NOR4_X1 U5378 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4865)
         );
  AOI22_X1 U5379 ( .A1(n4850), .A2(keyinput112), .B1(keyinput96), .B2(n4849), 
        .ZN(n4848) );
  OAI221_X1 U5380 ( .B1(n4850), .B2(keyinput112), .C1(n4849), .C2(keyinput96), 
        .A(n4848), .ZN(n4863) );
  AOI22_X1 U5381 ( .A1(n4853), .A2(keyinput127), .B1(n4852), .B2(keyinput118), 
        .ZN(n4851) );
  OAI221_X1 U5382 ( .B1(n4853), .B2(keyinput127), .C1(n4852), .C2(keyinput118), 
        .A(n4851), .ZN(n4862) );
  AOI22_X1 U5383 ( .A1(n4856), .A2(keyinput115), .B1(n4855), .B2(keyinput106), 
        .ZN(n4854) );
  OAI221_X1 U5384 ( .B1(n4856), .B2(keyinput115), .C1(n4855), .C2(keyinput106), 
        .A(n4854), .ZN(n4861) );
  AOI22_X1 U5385 ( .A1(n4859), .A2(keyinput102), .B1(keyinput94), .B2(n4858), 
        .ZN(n4857) );
  OAI221_X1 U5386 ( .B1(n4859), .B2(keyinput102), .C1(n4858), .C2(keyinput94), 
        .A(n4857), .ZN(n4860) );
  NOR4_X1 U5387 ( .A1(n4863), .A2(n4862), .A3(n4861), .A4(n4860), .ZN(n4864)
         );
  NAND4_X1 U5388 ( .A1(n4867), .A2(n4866), .A3(n4865), .A4(n4864), .ZN(n4934)
         );
  AOI22_X1 U5389 ( .A1(n2415), .A2(keyinput98), .B1(n4869), .B2(keyinput91), 
        .ZN(n4868) );
  OAI221_X1 U5390 ( .B1(n2415), .B2(keyinput98), .C1(n4869), .C2(keyinput91), 
        .A(n4868), .ZN(n4874) );
  XNOR2_X1 U5391 ( .A(n4870), .B(keyinput71), .ZN(n4873) );
  XNOR2_X1 U5392 ( .A(n4871), .B(keyinput63), .ZN(n4872) );
  OR3_X1 U5393 ( .A1(n4874), .A2(n4873), .A3(n4872), .ZN(n4883) );
  AOI22_X1 U5394 ( .A1(n4877), .A2(keyinput87), .B1(keyinput86), .B2(n4876), 
        .ZN(n4875) );
  OAI221_X1 U5395 ( .B1(n4877), .B2(keyinput87), .C1(n4876), .C2(keyinput86), 
        .A(n4875), .ZN(n4882) );
  INV_X1 U5396 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4879) );
  AOI22_X1 U5397 ( .A1(n4880), .A2(keyinput75), .B1(keyinput70), .B2(n4879), 
        .ZN(n4878) );
  OAI221_X1 U5398 ( .B1(n4880), .B2(keyinput75), .C1(n4879), .C2(keyinput70), 
        .A(n4878), .ZN(n4881) );
  NOR3_X1 U5399 ( .A1(n4883), .A2(n4882), .A3(n4881), .ZN(n4932) );
  AOI22_X1 U5400 ( .A1(n4886), .A2(keyinput34), .B1(keyinput35), .B2(n4885), 
        .ZN(n4884) );
  OAI221_X1 U5401 ( .B1(n4886), .B2(keyinput34), .C1(n4885), .C2(keyinput35), 
        .A(n4884), .ZN(n4897) );
  AOI22_X1 U5402 ( .A1(n2512), .A2(keyinput42), .B1(keyinput47), .B2(n3915), 
        .ZN(n4887) );
  OAI221_X1 U5403 ( .B1(n2512), .B2(keyinput42), .C1(n3915), .C2(keyinput47), 
        .A(n4887), .ZN(n4896) );
  AOI22_X1 U5404 ( .A1(n4890), .A2(keyinput38), .B1(n4889), .B2(keyinput43), 
        .ZN(n4888) );
  OAI221_X1 U5405 ( .B1(n4890), .B2(keyinput38), .C1(n4889), .C2(keyinput43), 
        .A(n4888), .ZN(n4895) );
  INV_X1 U5406 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4891) );
  XOR2_X1 U5407 ( .A(n4891), .B(keyinput54), .Z(n4893) );
  XNOR2_X1 U5408 ( .A(IR_REG_18__SCAN_IN), .B(keyinput51), .ZN(n4892) );
  NAND2_X1 U5409 ( .A1(n4893), .A2(n4892), .ZN(n4894) );
  NOR4_X1 U5410 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4931)
         );
  INV_X1 U5411 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4900) );
  AOI22_X1 U5412 ( .A1(n4900), .A2(keyinput26), .B1(n4899), .B2(keyinput30), 
        .ZN(n4898) );
  OAI221_X1 U5413 ( .B1(n4900), .B2(keyinput26), .C1(n4899), .C2(keyinput30), 
        .A(n4898), .ZN(n4912) );
  AOI22_X1 U5414 ( .A1(n3435), .A2(keyinput14), .B1(n4902), .B2(keyinput15), 
        .ZN(n4901) );
  OAI221_X1 U5415 ( .B1(n3435), .B2(keyinput14), .C1(n4902), .C2(keyinput15), 
        .A(n4901), .ZN(n4911) );
  AOI22_X1 U5416 ( .A1(n4905), .A2(keyinput6), .B1(keyinput3), .B2(n4904), 
        .ZN(n4903) );
  OAI221_X1 U5417 ( .B1(n4905), .B2(keyinput6), .C1(n4904), .C2(keyinput3), 
        .A(n4903), .ZN(n4910) );
  INV_X1 U5418 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4908) );
  AOI22_X1 U5419 ( .A1(n4908), .A2(keyinput21), .B1(n4907), .B2(keyinput29), 
        .ZN(n4906) );
  OAI221_X1 U5420 ( .B1(n4908), .B2(keyinput21), .C1(n4907), .C2(keyinput29), 
        .A(n4906), .ZN(n4909) );
  NOR4_X1 U5421 ( .A1(n4912), .A2(n4911), .A3(n4910), .A4(n4909), .ZN(n4930)
         );
  AOI22_X1 U5422 ( .A1(n4915), .A2(keyinput13), .B1(keyinput17), .B2(n4914), 
        .ZN(n4913) );
  OAI221_X1 U5423 ( .B1(n4915), .B2(keyinput13), .C1(n4914), .C2(keyinput17), 
        .A(n4913), .ZN(n4928) );
  AOI22_X1 U5424 ( .A1(n4918), .A2(keyinput85), .B1(keyinput69), .B2(n4917), 
        .ZN(n4916) );
  OAI221_X1 U5425 ( .B1(n4918), .B2(keyinput85), .C1(n4917), .C2(keyinput69), 
        .A(n4916), .ZN(n4927) );
  INV_X1 U5426 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4921) );
  AOI22_X1 U5427 ( .A1(n4921), .A2(keyinput45), .B1(keyinput57), .B2(n4920), 
        .ZN(n4919) );
  OAI221_X1 U5428 ( .B1(n4921), .B2(keyinput45), .C1(n4920), .C2(keyinput57), 
        .A(n4919), .ZN(n4926) );
  INV_X1 U5429 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4924) );
  AOI22_X1 U5430 ( .A1(n4924), .A2(keyinput5), .B1(keyinput9), .B2(n4923), 
        .ZN(n4922) );
  OAI221_X1 U5431 ( .B1(n4924), .B2(keyinput5), .C1(n4923), .C2(keyinput9), 
        .A(n4922), .ZN(n4925) );
  NOR4_X1 U5432 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n4929)
         );
  NAND4_X1 U5433 ( .A1(n4932), .A2(n4931), .A3(n4930), .A4(n4929), .ZN(n4933)
         );
  NOR3_X1 U5434 ( .A1(n4935), .A2(n4934), .A3(n4933), .ZN(n4973) );
  OAI22_X1 U5435 ( .A1(ADDR_REG_11__SCAN_IN), .A2(keyinput50), .B1(keyinput58), 
        .B2(DATAO_REG_17__SCAN_IN), .ZN(n4936) );
  AOI221_X1 U5436 ( .B1(ADDR_REG_11__SCAN_IN), .B2(keyinput50), .C1(
        DATAO_REG_17__SCAN_IN), .C2(keyinput58), .A(n4936), .ZN(n4943) );
  OAI22_X1 U5437 ( .A1(REG2_REG_14__SCAN_IN), .A2(keyinput62), .B1(keyinput66), 
        .B2(REG1_REG_16__SCAN_IN), .ZN(n4937) );
  AOI221_X1 U5438 ( .B1(REG2_REG_14__SCAN_IN), .B2(keyinput62), .C1(
        REG1_REG_16__SCAN_IN), .C2(keyinput66), .A(n4937), .ZN(n4942) );
  OAI22_X1 U5439 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput10), .B1(keyinput18), 
        .B2(REG0_REG_28__SCAN_IN), .ZN(n4938) );
  AOI221_X1 U5440 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput10), .C1(
        REG0_REG_28__SCAN_IN), .C2(keyinput18), .A(n4938), .ZN(n4941) );
  OAI22_X1 U5441 ( .A1(REG1_REG_8__SCAN_IN), .A2(keyinput22), .B1(keyinput46), 
        .B2(REG0_REG_7__SCAN_IN), .ZN(n4939) );
  AOI221_X1 U5442 ( .B1(REG1_REG_8__SCAN_IN), .B2(keyinput22), .C1(
        REG0_REG_7__SCAN_IN), .C2(keyinput46), .A(n4939), .ZN(n4940) );
  NAND4_X1 U5443 ( .A1(n4943), .A2(n4942), .A3(n4941), .A4(n4940), .ZN(n4971)
         );
  OAI22_X1 U5444 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput126), .B1(keyinput122), 
        .B2(REG0_REG_21__SCAN_IN), .ZN(n4944) );
  AOI221_X1 U5445 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput126), .C1(
        REG0_REG_21__SCAN_IN), .C2(keyinput122), .A(n4944), .ZN(n4951) );
  OAI22_X1 U5446 ( .A1(REG1_REG_26__SCAN_IN), .A2(keyinput114), .B1(
        REG0_REG_12__SCAN_IN), .B2(keyinput110), .ZN(n4945) );
  AOI221_X1 U5447 ( .B1(REG1_REG_26__SCAN_IN), .B2(keyinput114), .C1(
        keyinput110), .C2(REG0_REG_12__SCAN_IN), .A(n4945), .ZN(n4950) );
  OAI22_X1 U5448 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput82), .B1(DATAI_11_), 
        .B2(keyinput74), .ZN(n4946) );
  AOI221_X1 U5449 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput82), .C1(keyinput74), 
        .C2(DATAI_11_), .A(n4946), .ZN(n4949) );
  OAI22_X1 U5450 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput90), .B1(
        REG2_REG_4__SCAN_IN), .B2(keyinput78), .ZN(n4947) );
  AOI221_X1 U5451 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput90), .C1(keyinput78), .C2(REG2_REG_4__SCAN_IN), .A(n4947), .ZN(n4948) );
  NAND4_X1 U5452 ( .A1(n4951), .A2(n4950), .A3(n4949), .A4(n4948), .ZN(n4970)
         );
  OAI22_X1 U5453 ( .A1(REG1_REG_23__SCAN_IN), .A2(keyinput64), .B1(keyinput123), .B2(DATAI_6_), .ZN(n4952) );
  AOI221_X1 U5454 ( .B1(REG1_REG_23__SCAN_IN), .B2(keyinput64), .C1(DATAI_6_), 
        .C2(keyinput123), .A(n4952), .ZN(n4959) );
  OAI22_X1 U5455 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput0), .B1(keyinput59), 
        .B2(IR_REG_20__SCAN_IN), .ZN(n4953) );
  AOI221_X1 U5456 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput0), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput59), .A(n4953), .ZN(n4958) );
  OAI22_X1 U5457 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput107), .B1(
        REG0_REG_26__SCAN_IN), .B2(keyinput119), .ZN(n4954) );
  AOI221_X1 U5458 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput107), .C1(keyinput119), 
        .C2(REG0_REG_26__SCAN_IN), .A(n4954), .ZN(n4957) );
  OAI22_X1 U5459 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput103), .B1(
        keyinput124), .B2(REG3_REG_3__SCAN_IN), .ZN(n4955) );
  AOI221_X1 U5460 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput103), .C1(
        REG3_REG_3__SCAN_IN), .C2(keyinput124), .A(n4955), .ZN(n4956) );
  NAND4_X1 U5461 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4969)
         );
  OAI22_X1 U5462 ( .A1(REG1_REG_27__SCAN_IN), .A2(keyinput99), .B1(keyinput79), 
        .B2(ADDR_REG_9__SCAN_IN), .ZN(n4960) );
  AOI221_X1 U5463 ( .B1(REG1_REG_27__SCAN_IN), .B2(keyinput99), .C1(
        ADDR_REG_9__SCAN_IN), .C2(keyinput79), .A(n4960), .ZN(n4967) );
  OAI22_X1 U5464 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput2), .B1(
        REG0_REG_23__SCAN_IN), .B2(keyinput83), .ZN(n4961) );
  AOI221_X1 U5465 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput2), .C1(keyinput83), 
        .C2(REG0_REG_23__SCAN_IN), .A(n4961), .ZN(n4966) );
  OAI22_X1 U5466 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput55), .B1(
        DATAO_REG_2__SCAN_IN), .B2(keyinput67), .ZN(n4962) );
  AOI221_X1 U5467 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput55), .C1(keyinput67), 
        .C2(DATAO_REG_2__SCAN_IN), .A(n4962), .ZN(n4965) );
  OAI22_X1 U5468 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput95), .B1(DATAI_1_), 
        .B2(keyinput39), .ZN(n4963) );
  AOI221_X1 U5469 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput95), .C1(keyinput39), 
        .C2(DATAI_1_), .A(n4963), .ZN(n4964) );
  NAND4_X1 U5470 ( .A1(n4967), .A2(n4966), .A3(n4965), .A4(n4964), .ZN(n4968)
         );
  NOR4_X1 U5471 ( .A1(n4971), .A2(n4970), .A3(n4969), .A4(n4968), .ZN(n4972)
         );
  NAND3_X1 U5472 ( .A1(n4974), .A2(n4973), .A3(n4972), .ZN(n4991) );
  AOI211_X1 U5473 ( .C1(n2238), .C2(n4977), .A(n4976), .B(n4975), .ZN(n4978)
         );
  AOI211_X1 U5474 ( .C1(n4980), .C2(ADDR_REG_15__SCAN_IN), .A(n4979), .B(n4978), .ZN(n4987) );
  AOI21_X1 U5475 ( .B1(n4983), .B2(n4982), .A(n4981), .ZN(n4984) );
  NAND2_X1 U5476 ( .A1(n4985), .A2(n4984), .ZN(n4986) );
  OAI211_X1 U5477 ( .C1(n4989), .C2(n4988), .A(n4987), .B(n4986), .ZN(n4990)
         );
  XNOR2_X1 U5478 ( .A(n4991), .B(n4990), .ZN(U3255) );
  CLKBUF_X1 U2460 ( .A(n2527), .Z(n2740) );
  CLKBUF_X1 U2476 ( .A(n2895), .Z(n3043) );
  INV_X2 U2491 ( .A(n3015), .ZN(n3019) );
endmodule

