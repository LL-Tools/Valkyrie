

module b21_C_gen_AntiSAT_k_256_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503;

  NAND2_X1 U4983 ( .A1(n9465), .A2(n6126), .ZN(n6175) );
  INV_X2 U4984 ( .A(n5347), .ZN(n5363) );
  INV_X1 U4985 ( .A(n8892), .ZN(n8886) );
  NAND2_X1 U4986 ( .A1(n9142), .A2(n9085), .ZN(n9127) );
  INV_X2 U4987 ( .A(n6782), .ZN(n5839) );
  INV_X1 U4988 ( .A(n5353), .ZN(n6509) );
  INV_X1 U4989 ( .A(n9659), .ZN(n9848) );
  INV_X1 U4990 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U4991 ( .A1(n9192), .A2(n9083), .ZN(n9175) );
  NAND2_X1 U4992 ( .A1(n5559), .A2(n9636), .ZN(n9533) );
  NAND2_X1 U4993 ( .A1(n4492), .A2(n5178), .ZN(n5932) );
  AND2_X1 U4994 ( .A1(n6135), .A2(n9461), .ZN(n4478) );
  OR2_X1 U4995 ( .A1(n4972), .A2(n4636), .ZN(n4479) );
  NOR2_X2 U4996 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5075) );
  NAND3_X2 U4997 ( .A1(n5075), .A2(n5277), .A3(n5168), .ZN(n5313) );
  XNOR2_X2 U4998 ( .A(n8585), .B(n5104), .ZN(n8678) );
  OAI21_X2 U4999 ( .B1(n5531), .B2(n5164), .A(n5163), .ZN(n5562) );
  AOI21_X2 U5000 ( .B1(n4893), .B2(n5161), .A(n5160), .ZN(n5531) );
  OAI22_X2 U5001 ( .A1(n9254), .A2(n9077), .B1(n9407), .B2(n9279), .ZN(n9245)
         );
  AOI21_X2 U5002 ( .B1(n9296), .B2(n9275), .A(n9269), .ZN(n9254) );
  OR2_X1 U5003 ( .A1(n8666), .A2(n5007), .ZN(n4814) );
  CLKBUF_X1 U5004 ( .A(n9830), .Z(n4481) );
  NAND2_X1 U5005 ( .A1(n4686), .A2(n5352), .ZN(n6926) );
  INV_X1 U5006 ( .A(n8705), .ZN(n4808) );
  NAND2_X1 U5007 ( .A1(n7144), .A2(n8447), .ZN(n5997) );
  NAND2_X2 U5008 ( .A1(n6884), .A2(n6885), .ZN(n6883) );
  NAND2_X1 U5009 ( .A1(n6641), .A2(n6642), .ZN(n6643) );
  NAND2_X1 U5010 ( .A1(n8360), .A2(n8363), .ZN(n7146) );
  AOI22_X1 U5011 ( .A1(n5885), .A2(n9668), .B1(n5265), .B2(n6807), .ZN(n5326)
         );
  INV_X1 U5012 ( .A(n9669), .ZN(n7149) );
  INV_X1 U5013 ( .A(n7257), .ZN(n5949) );
  INV_X1 U5014 ( .A(n6807), .ZN(n10312) );
  NAND2_X1 U5015 ( .A1(n6141), .A2(n10369), .ZN(n6689) );
  BUF_X2 U5016 ( .A(n5872), .Z(n4483) );
  AND2_X1 U5017 ( .A1(n5364), .A2(n8204), .ZN(n5872) );
  NAND2_X1 U5018 ( .A1(n5364), .A2(n6461), .ZN(n5347) );
  CLKBUF_X2 U5019 ( .A(n6168), .Z(n8509) );
  AND2_X2 U5020 ( .A1(n5211), .A2(n5210), .ZN(n5304) );
  NAND2_X1 U5021 ( .A1(n5209), .A2(n10077), .ZN(n5221) );
  NAND2_X2 U5023 ( .A1(n4916), .A2(n4917), .ZN(n8204) );
  NOR2_X2 U5024 ( .A1(n4764), .A2(n5313), .ZN(n5183) );
  AOI21_X1 U5025 ( .B1(n4754), .B2(n9626), .A(n9651), .ZN(n9628) );
  MUX2_X1 U5026 ( .A(n6037), .B(n6036), .S(n10334), .Z(n6039) );
  MUX2_X1 U5027 ( .A(n6037), .B(n6027), .S(n10341), .Z(n6031) );
  OR2_X1 U5028 ( .A1(n6061), .A2(n10334), .ZN(n4614) );
  NAND2_X1 U5029 ( .A1(n4805), .A2(n4809), .ZN(n8640) );
  OAI21_X1 U5030 ( .B1(n8325), .B2(n9654), .A(n4739), .ZN(n4681) );
  OR2_X1 U5031 ( .A1(n9785), .A2(n9784), .ZN(n9788) );
  INV_X1 U5032 ( .A(n8324), .ZN(n10046) );
  AOI21_X1 U5033 ( .B1(n5051), .B2(n5053), .A(n4527), .ZN(n5050) );
  OAI22_X1 U5034 ( .A1(n9175), .A2(n9184), .B1(n9380), .B2(n9206), .ZN(n9160)
         );
  NAND2_X1 U5035 ( .A1(n9617), .A2(n4690), .ZN(n9512) );
  OAI21_X1 U5036 ( .B1(n9850), .B2(n4914), .A(n4623), .ZN(n6010) );
  NAND2_X1 U5037 ( .A1(n4908), .A2(n4515), .ZN(n9850) );
  NAND2_X1 U5038 ( .A1(n8588), .A2(n8587), .ZN(n9374) );
  XNOR2_X1 U5039 ( .A(n5870), .B(n5869), .ZN(n10096) );
  NAND2_X1 U5040 ( .A1(n5768), .A2(n5767), .ZN(n9832) );
  OAI21_X1 U5041 ( .B1(n6006), .B2(n4619), .A(n4615), .ZN(n9904) );
  AOI21_X1 U5042 ( .B1(n4756), .B2(n7999), .A(n5550), .ZN(n4692) );
  OAI22_X1 U5043 ( .A1(n8117), .A2(n5972), .B1(n9956), .B2(n10165), .ZN(n9950)
         );
  NAND2_X1 U5044 ( .A1(n8549), .A2(n8548), .ZN(n9388) );
  NAND2_X1 U5045 ( .A1(n7522), .A2(n6406), .ZN(n8076) );
  NAND2_X1 U5046 ( .A1(n8535), .A2(n8534), .ZN(n9394) );
  OR2_X1 U5047 ( .A1(n9922), .A2(n9910), .ZN(n9908) );
  NAND2_X1 U5048 ( .A1(n7926), .A2(n7925), .ZN(n7950) );
  NAND2_X1 U5049 ( .A1(n7370), .A2(n4514), .ZN(n7926) );
  NAND2_X1 U5050 ( .A1(n7313), .A2(n5072), .ZN(n7370) );
  NAND2_X1 U5051 ( .A1(n8105), .A2(n8104), .ZN(n9420) );
  NAND2_X1 U5052 ( .A1(n7234), .A2(n7233), .ZN(n7313) );
  OAI21_X1 U5053 ( .B1(n5658), .B2(n5657), .A(n5656), .ZN(n5684) );
  NAND2_X1 U5054 ( .A1(n6926), .A2(n6927), .ZN(n6925) );
  NAND2_X1 U5055 ( .A1(n5188), .A2(n5187), .ZN(n9649) );
  NAND2_X1 U5056 ( .A1(n6392), .A2(n6391), .ZN(n9436) );
  NAND2_X1 U5057 ( .A1(n5484), .A2(n5483), .ZN(n7994) );
  AND2_X2 U5058 ( .A1(n7023), .A2(n10375), .ZN(n10357) );
  INV_X2 U5059 ( .A(n10161), .ZN(n10157) );
  INV_X1 U5060 ( .A(n5994), .ZN(n8446) );
  OAI21_X1 U5061 ( .B1(n5924), .B2(n6773), .A(n9926), .ZN(n9648) );
  OAI211_X1 U5062 ( .C1(n5347), .C2(n6465), .A(n5316), .B(n5315), .ZN(n9575)
         );
  NAND4_X1 U5063 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n8945)
         );
  NAND4_X1 U5064 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n9669)
         );
  NAND4_X1 U5065 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n9668)
         );
  OAI211_X1 U5066 ( .C1(n5347), .C2(n6470), .A(n5298), .B(n5297), .ZN(n6807)
         );
  OAI211_X1 U5067 ( .C1(n5347), .C2(n6463), .A(n5280), .B(n5279), .ZN(n9611)
         );
  NAND2_X1 U5068 ( .A1(n6119), .A2(n8932), .ZN(n8741) );
  INV_X4 U5069 ( .A(n4478), .ZN(n4480) );
  INV_X2 U5070 ( .A(n6214), .ZN(n8622) );
  BUF_X4 U5071 ( .A(n5872), .Z(n4482) );
  INV_X1 U5072 ( .A(n8926), .ZN(n8763) );
  NAND2_X1 U5073 ( .A1(n6168), .A2(n8204), .ZN(n6241) );
  INV_X1 U5074 ( .A(n6135), .ZN(n9465) );
  NAND2_X1 U5075 ( .A1(n7298), .A2(n8473), .ZN(n6909) );
  INV_X2 U5076 ( .A(n9297), .ZN(n10369) );
  NAND2_X1 U5077 ( .A1(n6122), .A2(n6123), .ZN(n6135) );
  XNOR2_X1 U5078 ( .A(n6117), .B(n6073), .ZN(n9297) );
  NAND2_X1 U5079 ( .A1(n5182), .A2(n5181), .ZN(n10207) );
  NAND2_X1 U5080 ( .A1(n5198), .A2(n5197), .ZN(n7938) );
  AND2_X1 U5081 ( .A1(n5203), .A2(n5229), .ZN(n8473) );
  MUX2_X1 U5082 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6121), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6122) );
  NAND2_X1 U5083 ( .A1(n6147), .A2(n6146), .ZN(n6535) );
  MUX2_X1 U5084 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5207), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5209) );
  MUX2_X1 U5085 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5177), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5178) );
  XNOR2_X1 U5086 ( .A(n5205), .B(n4712), .ZN(n7298) );
  XNOR2_X1 U5087 ( .A(n5206), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5210) );
  MUX2_X1 U5088 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6145), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6146) );
  NAND2_X1 U5089 ( .A1(n6151), .A2(n6150), .ZN(n6534) );
  MUX2_X1 U5090 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5180), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5182) );
  MUX2_X1 U5091 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5196), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5198) );
  MUX2_X1 U5092 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6149), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6151) );
  OR2_X1 U5093 ( .A1(n5195), .A2(n5508), .ZN(n5196) );
  NAND2_X1 U5094 ( .A1(n6088), .A2(n4986), .ZN(n6147) );
  CLKBUF_X1 U5095 ( .A(n5208), .Z(n10077) );
  NAND2_X1 U5096 ( .A1(n6123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6125) );
  AND2_X1 U5097 ( .A1(n4944), .A2(n5183), .ZN(n4596) );
  AND2_X1 U5098 ( .A1(n5088), .A2(n4595), .ZN(n4594) );
  NAND2_X1 U5099 ( .A1(n4858), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4916) );
  AND2_X1 U5100 ( .A1(n5175), .A2(n4945), .ZN(n4944) );
  AND2_X1 U5101 ( .A1(n5099), .A2(n4535), .ZN(n5088) );
  AND4_X1 U5102 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5532), .ZN(n5175)
         );
  OAI21_X2 U5103 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5106), .ZN(n4917) );
  XNOR2_X1 U5104 ( .A(n5258), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6466) );
  INV_X4 U5105 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X2 U5106 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5277) );
  NOR2_X1 U5107 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5097) );
  NOR2_X1 U5108 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6066) );
  NOR2_X1 U5109 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6065) );
  NOR2_X1 U5110 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6064) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6068) );
  INV_X1 U5112 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7778) );
  NOR2_X1 U5113 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5035) );
  INV_X1 U5114 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6347) );
  INV_X1 U5115 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6283) );
  INV_X1 U5116 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U5117 ( .A1(n4667), .A2(n8301), .ZN(n8312) );
  OR4_X1 U5118 ( .A1(n9845), .A2(n9862), .A3(n9877), .A4(n8463), .ZN(n8464) );
  AND2_X4 U5119 ( .A1(n5248), .A2(n5226), .ZN(n5265) );
  XNOR2_X2 U5120 ( .A(n5950), .B(n7257), .ZN(n5992) );
  BUF_X4 U5121 ( .A(n5304), .Z(n4484) );
  INV_X1 U5122 ( .A(n6214), .ZN(n4485) );
  NAND2_X2 U5123 ( .A1(n6168), .A2(n4903), .ZN(n6214) );
  AND2_X4 U5124 ( .A1(n5221), .A2(n5210), .ZN(n5287) );
  AND2_X1 U5125 ( .A1(n5221), .A2(n10083), .ZN(n4486) );
  AND2_X1 U5126 ( .A1(n5221), .A2(n10083), .ZN(n4487) );
  OR2_X1 U5127 ( .A1(n9413), .A2(n9296), .ZN(n8849) );
  NAND2_X1 U5128 ( .A1(n7984), .A2(n4757), .ZN(n4756) );
  NOR2_X1 U5129 ( .A1(n7998), .A2(n4758), .ZN(n4757) );
  INV_X1 U5130 ( .A(n5502), .ZN(n4758) );
  INV_X1 U5131 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U5132 ( .A1(n8818), .A2(n8892), .ZN(n4798) );
  AOI21_X1 U5133 ( .B1(n8289), .B2(n8442), .A(n8288), .ZN(n4672) );
  OAI21_X1 U5134 ( .B1(n4784), .B2(n8874), .A(n4782), .ZN(n4781) );
  INV_X1 U5135 ( .A(n9135), .ZN(n4782) );
  AND2_X1 U5136 ( .A1(n4789), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5137 ( .A1(n4790), .A2(n4786), .ZN(n4785) );
  NAND2_X1 U5138 ( .A1(n8878), .A2(n9092), .ZN(n4787) );
  AND2_X1 U5139 ( .A1(n8435), .A2(n8430), .ZN(n8326) );
  NOR2_X1 U5140 ( .A1(n10046), .A2(n9748), .ZN(n8472) );
  NAND2_X1 U5141 ( .A1(n5155), .A2(n5154), .ZN(n5503) );
  NAND2_X1 U5142 ( .A1(n5136), .A2(n5135), .ZN(n5139) );
  NAND2_X1 U5143 ( .A1(n5059), .A2(n5060), .ZN(n5056) );
  AOI21_X1 U5144 ( .B1(n9244), .B2(n5062), .A(n9079), .ZN(n5061) );
  INV_X1 U5145 ( .A(n5063), .ZN(n5062) );
  OR2_X1 U5146 ( .A1(n9429), .A2(n9310), .ZN(n8834) );
  AOI21_X1 U5147 ( .B1(n8014), .B2(n8823), .A(n8822), .ZN(n8015) );
  NAND2_X2 U5148 ( .A1(n6535), .A2(n6534), .ZN(n6168) );
  NAND2_X1 U5149 ( .A1(n6788), .A2(n8189), .ZN(n8774) );
  NAND2_X1 U5150 ( .A1(n6925), .A2(n4496), .ZN(n5081) );
  NAND2_X1 U5151 ( .A1(n4745), .A2(n4744), .ZN(n4750) );
  NOR2_X1 U5152 ( .A1(n6028), .A2(n9979), .ZN(n4740) );
  AND2_X1 U5153 ( .A1(n8318), .A2(n8333), .ZN(n8467) );
  NAND2_X1 U5154 ( .A1(n9831), .A2(n9819), .ZN(n9813) );
  INV_X1 U5155 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U5156 ( .A1(n4888), .A2(n4887), .ZN(n8195) );
  AOI21_X1 U5157 ( .B1(n4890), .B2(n4892), .A(n4553), .ZN(n4887) );
  NAND2_X1 U5158 ( .A1(n5637), .A2(n5636), .ZN(n5658) );
  INV_X1 U5159 ( .A(n5632), .ZN(n5633) );
  AOI21_X1 U5160 ( .B1(n4872), .B2(n4870), .A(n4869), .ZN(n4868) );
  INV_X1 U5161 ( .A(n5588), .ZN(n4869) );
  INV_X1 U5162 ( .A(n5560), .ZN(n4870) );
  AND2_X1 U5163 ( .A1(n5588), .A2(n5567), .ZN(n5586) );
  INV_X1 U5164 ( .A(n5530), .ZN(n5164) );
  INV_X1 U5165 ( .A(n5504), .ZN(n5160) );
  AND2_X1 U5166 ( .A1(n5503), .A2(n5505), .ZN(n5161) );
  NAND2_X1 U5167 ( .A1(n4894), .A2(n5032), .ZN(n4893) );
  INV_X1 U5168 ( .A(n6379), .ZN(n6371) );
  NAND2_X1 U5169 ( .A1(n8162), .A2(n8163), .ZN(n4823) );
  AND2_X1 U5170 ( .A1(n8707), .A2(n5005), .ZN(n5004) );
  NAND2_X1 U5171 ( .A1(n5006), .A2(n5008), .ZN(n5005) );
  INV_X1 U5172 ( .A(n5009), .ZN(n5006) );
  NAND2_X1 U5173 ( .A1(n8668), .A2(n5010), .ZN(n5008) );
  AOI21_X1 U5174 ( .B1(n4799), .B2(n8896), .A(n8895), .ZN(n8924) );
  NAND2_X1 U5175 ( .A1(n4801), .A2(n4800), .ZN(n4799) );
  AND2_X1 U5176 ( .A1(n8501), .A2(n8500), .ZN(n8724) );
  OR2_X1 U5177 ( .A1(n9153), .A2(n6194), .ZN(n8501) );
  AND3_X1 U5178 ( .A1(n8112), .A2(n8111), .A3(n8110), .ZN(n9296) );
  OR2_X1 U5179 ( .A1(n6661), .A2(n6660), .ZN(n4718) );
  OR2_X1 U5180 ( .A1(n8613), .A2(n6758), .ZN(n9103) );
  OR2_X1 U5181 ( .A1(n9358), .A2(n9099), .ZN(n9092) );
  OR2_X1 U5182 ( .A1(n9380), .A2(n8722), .ZN(n8751) );
  AND2_X1 U5183 ( .A1(n8751), .A2(n8871), .ZN(n9184) );
  OR2_X1 U5184 ( .A1(n9400), .A2(n9237), .ZN(n8853) );
  NAND2_X1 U5185 ( .A1(n4952), .A2(n4949), .ZN(n9257) );
  NOR2_X1 U5186 ( .A1(n4951), .A2(n4950), .ZN(n4949) );
  INV_X1 U5187 ( .A(n9258), .ZN(n4951) );
  OR2_X1 U5188 ( .A1(n9423), .A2(n9295), .ZN(n5100) );
  OR2_X1 U5189 ( .A1(n6364), .A2(n7348), .ZN(n6393) );
  AND2_X1 U5190 ( .A1(n8015), .A2(n9070), .ZN(n8055) );
  NAND2_X1 U5191 ( .A1(n7928), .A2(n7927), .ZN(n4983) );
  NAND2_X1 U5192 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  NAND2_X1 U5193 ( .A1(n8495), .A2(n8494), .ZN(n9369) );
  INV_X1 U5194 ( .A(n7046), .ZN(n10398) );
  XNOR2_X1 U5195 ( .A(n6113), .B(n4832), .ZN(n8926) );
  NAND2_X1 U5196 ( .A1(n6112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6113) );
  AND2_X1 U5197 ( .A1(n7999), .A2(n5550), .ZN(n4755) );
  NOR2_X1 U5198 ( .A1(n7489), .A2(n7490), .ZN(n9672) );
  OR2_X1 U5199 ( .A1(n9692), .A2(n9691), .ZN(n4849) );
  OR2_X1 U5200 ( .A1(n9692), .A2(n4847), .ZN(n4845) );
  OR2_X1 U5201 ( .A1(n9709), .A2(n9691), .ZN(n4847) );
  AOI21_X1 U5202 ( .B1(n9740), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9739), .ZN(
        n9741) );
  NAND2_X1 U5203 ( .A1(n9808), .A2(n9809), .ZN(n5987) );
  OR2_X1 U5204 ( .A1(n9990), .A2(n9828), .ZN(n9794) );
  NOR2_X1 U5205 ( .A1(n4525), .A2(n4941), .ZN(n4940) );
  INV_X1 U5206 ( .A(n5980), .ZN(n4941) );
  NAND2_X1 U5207 ( .A1(n4567), .A2(n4571), .ZN(n5970) );
  INV_X1 U5208 ( .A(n4572), .ZN(n4571) );
  OAI21_X1 U5209 ( .B1(n4920), .B2(n4490), .A(n5968), .ZN(n4572) );
  NAND2_X1 U5210 ( .A1(n8209), .A2(n8208), .ZN(n8324) );
  NOR2_X1 U5211 ( .A1(n5313), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5400) );
  XNOR2_X1 U5212 ( .A(n5122), .B(n7648), .ZN(n5310) );
  INV_X2 U5213 ( .A(n5364), .ZN(n6433) );
  INV_X1 U5214 ( .A(n9657), .ZN(n9812) );
  INV_X1 U5215 ( .A(n9658), .ZN(n9828) );
  NAND2_X1 U5216 ( .A1(n5232), .A2(n5088), .ZN(n5179) );
  NAND2_X1 U5217 ( .A1(n4657), .A2(n8453), .ZN(n8223) );
  NOR2_X1 U5218 ( .A1(n4792), .A2(n5039), .ZN(n4791) );
  OAI21_X1 U5219 ( .B1(n8823), .B2(n4798), .A(n4793), .ZN(n4792) );
  OR2_X1 U5220 ( .A1(n4797), .A2(n8821), .ZN(n4793) );
  NAND2_X1 U5221 ( .A1(n4797), .A2(n4798), .ZN(n4795) );
  OR2_X1 U5222 ( .A1(n8290), .A2(n4684), .ZN(n4668) );
  NOR2_X1 U5223 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  INV_X1 U5224 ( .A(n8297), .ZN(n4671) );
  NOR2_X1 U5225 ( .A1(n4787), .A2(n4778), .ZN(n4777) );
  MUX2_X1 U5226 ( .A(n8869), .B(n8868), .S(n8892), .Z(n8872) );
  NAND2_X1 U5227 ( .A1(n4860), .A2(n9653), .ZN(n8405) );
  INV_X1 U5228 ( .A(n5763), .ZN(n4879) );
  OAI22_X1 U5229 ( .A1(n8884), .A2(n8886), .B1(n8892), .B2(n8887), .ZN(n4803)
         );
  NAND2_X1 U5230 ( .A1(n8323), .A2(n8322), .ZN(n8325) );
  AND2_X1 U5231 ( .A1(n4878), .A2(n4884), .ZN(n4877) );
  NOR2_X1 U5232 ( .A1(n5818), .A2(n4885), .ZN(n4884) );
  NAND2_X1 U5233 ( .A1(n4881), .A2(n4879), .ZN(n4878) );
  INV_X1 U5234 ( .A(n5789), .ZN(n4885) );
  INV_X1 U5235 ( .A(n4881), .ZN(n4880) );
  NOR2_X1 U5236 ( .A1(n5153), .A2(n5030), .ZN(n5029) );
  INV_X1 U5237 ( .A(n5149), .ZN(n5030) );
  INV_X1 U5238 ( .A(n5458), .ZN(n5153) );
  NAND2_X1 U5239 ( .A1(n5340), .A2(n5341), .ZN(n5127) );
  INV_X1 U5240 ( .A(n4829), .ZN(n4828) );
  INV_X1 U5241 ( .A(n6312), .ZN(n4827) );
  NAND2_X1 U5242 ( .A1(n6689), .A2(n6143), .ZN(n6144) );
  AND2_X1 U5243 ( .A1(n6142), .A2(n8926), .ZN(n6143) );
  NAND2_X1 U5244 ( .A1(n4977), .A2(n4981), .ZN(n4976) );
  INV_X1 U5245 ( .A(n4507), .ZN(n4977) );
  NAND2_X1 U5246 ( .A1(n4979), .A2(n8887), .ZN(n4978) );
  OR2_X1 U5247 ( .A1(n9388), .A2(n9207), .ZN(n9080) );
  OR2_X1 U5248 ( .A1(n9436), .A2(n8937), .ZN(n8829) );
  AOI21_X1 U5249 ( .B1(n5043), .B2(n5041), .A(n4526), .ZN(n5040) );
  INV_X1 U5250 ( .A(n5043), .ZN(n5042) );
  OR2_X1 U5251 ( .A1(n7964), .A2(n7955), .ZN(n8817) );
  NAND2_X1 U5252 ( .A1(n4770), .A2(n4765), .ZN(n8797) );
  NOR2_X1 U5253 ( .A1(n7374), .A2(n4766), .ZN(n4765) );
  INV_X1 U5254 ( .A(n6303), .ZN(n4766) );
  AND2_X1 U5255 ( .A1(n10359), .A2(n8781), .ZN(n4647) );
  NAND2_X1 U5256 ( .A1(n6181), .A2(n10393), .ZN(n8776) );
  AND2_X1 U5257 ( .A1(n6084), .A2(n4994), .ZN(n4993) );
  INV_X1 U5258 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U5259 ( .A1(n4831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6111) );
  INV_X1 U5260 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6072) );
  INV_X1 U5261 ( .A(n6083), .ZN(n4836) );
  INV_X1 U5262 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U5263 ( .A1(n9595), .A2(n9597), .ZN(n4741) );
  XNOR2_X1 U5264 ( .A(n5319), .B(n5839), .ZN(n5324) );
  XNOR2_X1 U5265 ( .A(n5283), .B(n5839), .ZN(n5285) );
  NAND2_X1 U5266 ( .A1(n4695), .A2(n5549), .ZN(n4694) );
  INV_X1 U5267 ( .A(n7999), .ZN(n4695) );
  INV_X1 U5268 ( .A(n5221), .ZN(n5211) );
  AND2_X1 U5269 ( .A1(n4842), .A2(n4841), .ZN(n9671) );
  NAND2_X1 U5270 ( .A1(n7488), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4841) );
  INV_X1 U5271 ( .A(n5983), .ZN(n4578) );
  NOR2_X1 U5272 ( .A1(n9826), .A2(n4670), .ZN(n4625) );
  OR2_X1 U5273 ( .A1(n5573), .A2(n5572), .ZN(n5596) );
  NAND2_X1 U5274 ( .A1(n5218), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5573) );
  INV_X1 U5275 ( .A(n5541), .ZN(n5218) );
  INV_X1 U5276 ( .A(n5969), .ZN(n4939) );
  OR2_X1 U5277 ( .A1(n5486), .A2(n5485), .ZN(n5516) );
  NAND2_X1 U5278 ( .A1(n9546), .A2(n7010), .ZN(n8421) );
  NAND2_X1 U5279 ( .A1(n10321), .A2(n9667), .ZN(n8416) );
  NAND2_X1 U5280 ( .A1(n7149), .A2(n9611), .ZN(n5995) );
  NAND2_X1 U5281 ( .A1(n8361), .A2(n5995), .ZN(n5994) );
  NAND2_X1 U5282 ( .A1(n5097), .A2(n5916), .ZN(n4761) );
  NAND2_X1 U5283 ( .A1(n5686), .A2(n5685), .ZN(n5709) );
  AOI21_X1 U5284 ( .B1(n4871), .B2(n4864), .A(n4499), .ZN(n4863) );
  INV_X1 U5285 ( .A(n5586), .ZN(n4873) );
  OAI21_X1 U5286 ( .B1(n5029), .B2(n5031), .A(n5503), .ZN(n5028) );
  NAND2_X1 U5287 ( .A1(n5503), .A2(n5157), .ZN(n5479) );
  NAND2_X1 U5288 ( .A1(n5437), .A2(n5102), .ZN(n5150) );
  NAND2_X1 U5289 ( .A1(n5139), .A2(n5138), .ZN(n5398) );
  AND2_X1 U5290 ( .A1(n5133), .A2(n5126), .ZN(n5023) );
  INV_X1 U5291 ( .A(n5127), .ZN(n5018) );
  XNOR2_X1 U5292 ( .A(n5130), .B(SI_7_), .ZN(n5374) );
  XNOR2_X1 U5293 ( .A(n5128), .B(SI_6_), .ZN(n5362) );
  NAND2_X1 U5294 ( .A1(n5127), .A2(n5126), .ZN(n5361) );
  AND2_X1 U5295 ( .A1(n5121), .A2(n5117), .ZN(n4608) );
  INV_X1 U5296 ( .A(SI_4_), .ZN(n7648) );
  NAND2_X1 U5297 ( .A1(n6381), .A2(n4519), .ZN(n7522) );
  AND2_X1 U5298 ( .A1(n6405), .A2(n6385), .ZN(n5011) );
  NOR2_X1 U5299 ( .A1(n7183), .A2(n4830), .ZN(n4829) );
  INV_X1 U5300 ( .A(n6316), .ZN(n4830) );
  NAND2_X1 U5301 ( .A1(n8652), .A2(n8519), .ZN(n5015) );
  INV_X1 U5302 ( .A(n8687), .ZN(n5016) );
  NAND2_X1 U5303 ( .A1(n6951), .A2(n6312), .ZN(n7177) );
  NAND2_X1 U5304 ( .A1(n6130), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6353) );
  INV_X1 U5305 ( .A(n6338), .ZN(n6130) );
  NAND2_X1 U5306 ( .A1(n6753), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8172) );
  INV_X1 U5307 ( .A(n8107), .ZN(n6753) );
  NOR2_X1 U5308 ( .A1(n8164), .A2(n4822), .ZN(n4821) );
  INV_X1 U5309 ( .A(n8099), .ZN(n4822) );
  XNOR2_X1 U5310 ( .A(n8076), .B(n8077), .ZN(n8075) );
  AND2_X1 U5311 ( .A1(n8596), .A2(n8595), .ZN(n8723) );
  AND2_X1 U5312 ( .A1(n8584), .A2(n8583), .ZN(n8722) );
  AND2_X1 U5313 ( .A1(n8178), .A2(n8177), .ZN(n9076) );
  NOR2_X1 U5314 ( .A1(n6591), .A2(n4509), .ZN(n6582) );
  OR2_X1 U5315 ( .A1(n6582), .A2(n6581), .ZN(n4720) );
  AND2_X1 U5316 ( .A1(n4718), .A2(n4717), .ZN(n6731) );
  NAND2_X1 U5317 ( .A1(n6728), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4717) );
  OR2_X1 U5318 ( .A1(n6731), .A2(n6730), .ZN(n4716) );
  AND2_X1 U5319 ( .A1(n4716), .A2(n4715), .ZN(n6857) );
  NAND2_X1 U5320 ( .A1(n6860), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5321 ( .A1(n9012), .A2(n9013), .ZN(n9015) );
  NOR2_X1 U5322 ( .A1(n9015), .A2(n9014), .ZN(n9026) );
  AND2_X1 U5323 ( .A1(n9121), .A2(n5101), .ZN(n9094) );
  NAND2_X1 U5324 ( .A1(n4635), .A2(n4633), .ZN(n9115) );
  OR2_X1 U5325 ( .A1(n4479), .A2(n9183), .ZN(n4635) );
  INV_X1 U5326 ( .A(n4634), .ZN(n4633) );
  OAI21_X1 U5327 ( .B1(n4479), .B2(n4510), .A(n4970), .ZN(n4634) );
  AND2_X1 U5328 ( .A1(n8614), .A2(n9103), .ZN(n9113) );
  AND2_X1 U5329 ( .A1(n9116), .A2(n5052), .ZN(n5051) );
  OR2_X1 U5330 ( .A1(n9135), .A2(n5053), .ZN(n5052) );
  INV_X1 U5331 ( .A(n9087), .ZN(n5053) );
  OR2_X1 U5332 ( .A1(n9369), .A2(n9137), .ZN(n9085) );
  OR2_X1 U5333 ( .A1(n8589), .A2(n8671), .ZN(n8591) );
  NAND2_X1 U5334 ( .A1(n4637), .A2(n4638), .ZN(n9147) );
  NAND2_X1 U5335 ( .A1(n9147), .A2(n9148), .ZN(n9146) );
  NAND2_X1 U5336 ( .A1(n9383), .A2(n9082), .ZN(n9083) );
  NAND2_X1 U5337 ( .A1(n9241), .A2(n4963), .ZN(n4961) );
  AOI21_X1 U5338 ( .B1(n4963), .B2(n8915), .A(n8721), .ZN(n4962) );
  NAND2_X1 U5339 ( .A1(n4961), .A2(n4959), .ZN(n9200) );
  NOR2_X1 U5340 ( .A1(n4966), .A2(n4960), .ZN(n4959) );
  INV_X1 U5341 ( .A(n4962), .ZN(n4960) );
  INV_X1 U5342 ( .A(n5061), .ZN(n5060) );
  AOI21_X1 U5343 ( .B1(n5061), .B2(n5063), .A(n4522), .ZN(n5059) );
  OR2_X1 U5344 ( .A1(n8536), .A2(n8661), .ZN(n8550) );
  AND2_X1 U5345 ( .A1(n8529), .A2(n8528), .ZN(n9237) );
  NOR2_X1 U5346 ( .A1(n9234), .A2(n4964), .ZN(n4963) );
  INV_X1 U5347 ( .A(n8853), .ZN(n4964) );
  OR2_X1 U5348 ( .A1(n9241), .A2(n8915), .ZN(n4965) );
  AND2_X1 U5349 ( .A1(n8853), .A2(n8855), .ZN(n9244) );
  NAND2_X1 U5350 ( .A1(n9257), .A2(n8851), .ZN(n9241) );
  NAND2_X1 U5351 ( .A1(n9306), .A2(n4956), .ZN(n4952) );
  NOR2_X1 U5352 ( .A1(n4958), .A2(n4957), .ZN(n4956) );
  INV_X1 U5353 ( .A(n9277), .ZN(n4957) );
  OR2_X1 U5354 ( .A1(n4954), .A2(n8720), .ZN(n4950) );
  AND2_X1 U5355 ( .A1(n9277), .A2(n4955), .ZN(n4954) );
  INV_X1 U5356 ( .A(n8754), .ZN(n4955) );
  AND2_X1 U5357 ( .A1(n8848), .A2(n8851), .ZN(n9258) );
  OR2_X1 U5358 ( .A1(n9420), .A2(n9312), .ZN(n8754) );
  NAND2_X1 U5359 ( .A1(n9285), .A2(n8837), .ZN(n4958) );
  NOR2_X1 U5360 ( .A1(n9288), .A2(n9413), .ZN(n9271) );
  NAND2_X1 U5361 ( .A1(n5066), .A2(n4508), .ZN(n5065) );
  INV_X1 U5362 ( .A(n5068), .ZN(n5066) );
  AND2_X1 U5363 ( .A1(n8849), .A2(n8843), .ZN(n9277) );
  NOR2_X1 U5364 ( .A1(n9285), .A2(n5069), .ZN(n5068) );
  INV_X1 U5365 ( .A(n5100), .ZN(n5069) );
  NAND2_X1 U5366 ( .A1(n9329), .A2(n9074), .ZN(n9303) );
  OR2_X1 U5367 ( .A1(n6395), .A2(n6133), .ZN(n6420) );
  AOI21_X1 U5368 ( .B1(n9341), .B2(n8831), .A(n8719), .ZN(n9307) );
  OR2_X1 U5369 ( .A1(n8050), .A2(n9436), .ZN(n9333) );
  NAND2_X1 U5370 ( .A1(n8827), .A2(n8824), .ZN(n4969) );
  AND2_X1 U5371 ( .A1(n8829), .A2(n8828), .ZN(n8827) );
  NOR2_X1 U5372 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  AND4_X1 U5373 ( .A1(n6358), .A2(n6357), .A3(n6356), .A4(n6355), .ZN(n8017)
         );
  AND2_X1 U5374 ( .A1(n8818), .A2(n8819), .ZN(n8911) );
  AND4_X1 U5375 ( .A1(n6369), .A2(n6368), .A3(n6367), .A4(n6366), .ZN(n8012)
         );
  NAND2_X1 U5376 ( .A1(n4772), .A2(n4767), .ZN(n8809) );
  NOR2_X1 U5377 ( .A1(n7923), .A2(n4768), .ZN(n4767) );
  INV_X1 U5378 ( .A(n6321), .ZN(n4768) );
  NAND2_X1 U5379 ( .A1(n6506), .A2(n6262), .ZN(n4772) );
  INV_X1 U5380 ( .A(n6291), .ZN(n6129) );
  INV_X1 U5381 ( .A(n4641), .ZN(n4640) );
  OAI21_X1 U5382 ( .B1(n4643), .B2(n4642), .A(n7315), .ZN(n4641) );
  NAND2_X1 U5383 ( .A1(n6128), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6291) );
  INV_X1 U5384 ( .A(n6269), .ZN(n6128) );
  OAI21_X1 U5385 ( .B1(n8902), .B2(n5048), .A(n10355), .ZN(n5047) );
  NAND2_X1 U5386 ( .A1(n7038), .A2(n8902), .ZN(n7112) );
  AND4_X1 U5387 ( .A1(n6213), .A2(n6212), .A3(n6211), .A4(n6210), .ZN(n7110)
         );
  NAND2_X1 U5388 ( .A1(n8776), .A2(n8775), .ZN(n7132) );
  INV_X1 U5389 ( .A(n7132), .ZN(n8899) );
  OR2_X1 U5390 ( .A1(n6415), .A2(P2_U3152), .ZN(n8931) );
  INV_X1 U5391 ( .A(n9311), .ZN(n10362) );
  NOR2_X1 U5392 ( .A1(n9101), .A2(n10434), .ZN(n4653) );
  NAND2_X1 U5393 ( .A1(n8577), .A2(n8576), .ZN(n9380) );
  NOR2_X1 U5394 ( .A1(n9245), .A2(n9244), .ZN(n9405) );
  AND2_X1 U5395 ( .A1(n8063), .A2(n6093), .ZN(n10377) );
  AND2_X1 U5396 ( .A1(n4993), .A2(n5073), .ZN(n4986) );
  AND2_X1 U5397 ( .A1(n6120), .A2(n5074), .ZN(n5073) );
  INV_X1 U5398 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U5399 ( .A1(n6108), .A2(n6107), .ZN(n6110) );
  XNOR2_X1 U5400 ( .A(n6111), .B(n6076), .ZN(n6685) );
  INV_X1 U5401 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7083) );
  AOI21_X1 U5402 ( .B1(n9536), .B2(n5585), .A(n5084), .ZN(n5083) );
  INV_X1 U5403 ( .A(n9554), .ZN(n5084) );
  NAND2_X1 U5404 ( .A1(n5251), .A2(n4516), .ZN(n4743) );
  NAND2_X1 U5405 ( .A1(n9670), .A2(n5265), .ZN(n5253) );
  AND2_X1 U5406 ( .A1(n5501), .A2(n5477), .ZN(n5087) );
  NAND2_X1 U5407 ( .A1(n5081), .A2(n6994), .ZN(n5416) );
  OAI21_X1 U5408 ( .B1(n4703), .B2(n5433), .A(n4706), .ZN(n4699) );
  OR2_X1 U5409 ( .A1(n7469), .A2(n7470), .ZN(n4706) );
  NOR2_X1 U5410 ( .A1(n5082), .A2(n5080), .ZN(n5079) );
  NAND2_X1 U5411 ( .A1(n4710), .A2(n9526), .ZN(n4709) );
  INV_X1 U5412 ( .A(n9526), .ZN(n4711) );
  NAND2_X1 U5413 ( .A1(n5251), .A2(n5239), .ZN(n4742) );
  NOR2_X1 U5414 ( .A1(n5919), .A2(n8482), .ZN(n4895) );
  MUX2_X1 U5415 ( .A(n8477), .B(n8476), .S(n8475), .Z(n8478) );
  NAND2_X1 U5416 ( .A1(n4900), .A2(n4679), .ZN(n4678) );
  AND2_X1 U5417 ( .A1(n4898), .A2(n4896), .ZN(n4679) );
  NAND2_X1 U5418 ( .A1(n4487), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5243) );
  AND2_X1 U5419 ( .A1(n10261), .A2(n6704), .ZN(n10276) );
  NAND2_X1 U5420 ( .A1(n10264), .A2(n6713), .ZN(n10281) );
  AND2_X1 U5421 ( .A1(n5439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5440) );
  OR2_X1 U5422 ( .A1(n5438), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5439) );
  NOR2_X1 U5423 ( .A1(n10297), .A2(n4546), .ZN(n6717) );
  AOI21_X1 U5424 ( .B1(n7101), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7100), .ZN(
        n7105) );
  OR2_X1 U5425 ( .A1(n7105), .A2(n7104), .ZN(n4842) );
  XNOR2_X1 U5426 ( .A(n9671), .B(n9678), .ZN(n7489) );
  OR2_X1 U5427 ( .A1(n9709), .A2(n4848), .ZN(n4846) );
  XNOR2_X1 U5428 ( .A(n4629), .B(n8468), .ZN(n4911) );
  NAND2_X1 U5429 ( .A1(n4628), .A2(n4626), .ZN(n4629) );
  INV_X1 U5430 ( .A(n8467), .ZN(n9784) );
  INV_X1 U5431 ( .A(n9656), .ZN(n9799) );
  NOR2_X1 U5432 ( .A1(n5984), .A2(n4581), .ZN(n4580) );
  INV_X1 U5433 ( .A(n5981), .ZN(n4581) );
  NAND2_X1 U5434 ( .A1(n9850), .A2(n4625), .ZN(n9823) );
  NAND2_X1 U5435 ( .A1(n9863), .A2(n8443), .ZN(n4908) );
  NAND2_X1 U5436 ( .A1(n9870), .A2(n9877), .ZN(n4942) );
  NAND2_X1 U5437 ( .A1(n4906), .A2(n8445), .ZN(n4905) );
  NAND2_X1 U5438 ( .A1(n4589), .A2(n4588), .ZN(n9888) );
  AOI21_X1 U5439 ( .B1(n4494), .B2(n4592), .A(n4543), .ZN(n4588) );
  INV_X1 U5440 ( .A(n5976), .ZN(n4592) );
  NAND2_X1 U5441 ( .A1(n6007), .A2(n8398), .ZN(n9890) );
  AOI21_X1 U5442 ( .B1(n4618), .B2(n4617), .A(n4616), .ZN(n4615) );
  INV_X1 U5443 ( .A(n8275), .ZN(n4616) );
  INV_X1 U5444 ( .A(n4621), .ZN(n4617) );
  NOR2_X1 U5445 ( .A1(n8264), .A2(n4622), .ZN(n4621) );
  AND2_X1 U5446 ( .A1(n8268), .A2(n8269), .ZN(n9942) );
  NAND2_X1 U5447 ( .A1(n9950), .A2(n9954), .ZN(n4936) );
  NAND2_X1 U5448 ( .A1(n4603), .A2(n4601), .ZN(n9952) );
  AOI21_X1 U5449 ( .B1(n4604), .B2(n4607), .A(n4602), .ZN(n4601) );
  INV_X1 U5450 ( .A(n8389), .ZN(n4602) );
  INV_X1 U5451 ( .A(n8033), .ZN(n6005) );
  AND2_X1 U5452 ( .A1(n8458), .A2(n4921), .ZN(n4920) );
  NAND2_X1 U5453 ( .A1(n4530), .A2(n5967), .ZN(n4921) );
  AOI21_X1 U5454 ( .B1(n4584), .B2(n4586), .A(n7450), .ZN(n4582) );
  INV_X1 U5455 ( .A(n4585), .ZN(n4584) );
  OAI22_X1 U5456 ( .A1(n4505), .A2(n4586), .B1(n7361), .B2(n9663), .ZN(n4585)
         );
  AND2_X1 U5457 ( .A1(n8240), .A2(n8368), .ZN(n8452) );
  NAND2_X1 U5458 ( .A1(n7007), .A2(n5960), .ZN(n7072) );
  INV_X1 U5459 ( .A(n5354), .ZN(n5213) );
  NAND2_X1 U5460 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5334) );
  AND2_X1 U5461 ( .A1(n6903), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U5462 ( .A1(n5958), .A2(n5957), .ZN(n6828) );
  AND2_X1 U5463 ( .A1(n8420), .A2(n8416), .ZN(n6826) );
  INV_X1 U5464 ( .A(n10149), .ZN(n9959) );
  INV_X1 U5465 ( .A(n9957), .ZN(n10147) );
  AND2_X1 U5466 ( .A1(n9670), .A2(n6851), .ZN(n6784) );
  NAND2_X1 U5467 ( .A1(n6784), .A2(n5992), .ZN(n4566) );
  NAND2_X1 U5468 ( .A1(n9460), .A2(n5363), .ZN(n4861) );
  AND2_X1 U5469 ( .A1(n6020), .A2(n6051), .ZN(n9768) );
  NAND2_X1 U5470 ( .A1(n5826), .A2(n5825), .ZN(n9801) );
  NAND2_X1 U5471 ( .A1(n8493), .A2(n5363), .ZN(n5826) );
  NAND2_X1 U5472 ( .A1(n5665), .A2(n5664), .ZN(n9895) );
  NAND2_X1 U5473 ( .A1(n5593), .A2(n5592), .ZN(n10030) );
  OR2_X1 U5474 ( .A1(n5364), .A2(n5259), .ZN(n5260) );
  XNOR2_X1 U5475 ( .A(n8207), .B(n8206), .ZN(n9457) );
  NAND2_X1 U5476 ( .A1(n5850), .A2(n5849), .ZN(n5870) );
  AND2_X1 U5477 ( .A1(n5871), .A2(n5855), .ZN(n5869) );
  NAND2_X1 U5478 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5479 ( .A1(n5232), .A2(n5234), .ZN(n5204) );
  OAI21_X1 U5480 ( .B1(n5562), .B2(n5561), .A(n5560), .ZN(n5587) );
  OR2_X1 U5481 ( .A1(n5402), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5438) );
  AND2_X1 U5482 ( .A1(n5344), .A2(n5343), .ZN(n6629) );
  XNOR2_X1 U5483 ( .A(n5120), .B(n5119), .ZN(n5294) );
  INV_X1 U5484 ( .A(SI_3_), .ZN(n5119) );
  OAI21_X1 U5485 ( .B1(n4810), .B2(n4808), .A(n4502), .ZN(n4806) );
  AOI21_X1 U5486 ( .B1(n5004), .B2(n5007), .A(n4545), .ZN(n4810) );
  NOR2_X1 U5487 ( .A1(n4811), .A2(n4808), .ZN(n4807) );
  INV_X1 U5488 ( .A(n5004), .ZN(n4811) );
  AOI21_X1 U5489 ( .B1(n4818), .B2(n4820), .A(n4523), .ZN(n4816) );
  NAND2_X1 U5490 ( .A1(n8624), .A2(n8623), .ZN(n9358) );
  AOI21_X1 U5491 ( .B1(n4488), .B2(n5007), .A(n4497), .ZN(n4809) );
  NAND2_X1 U5492 ( .A1(n4485), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5493 ( .A1(n8522), .A2(n8521), .ZN(n9400) );
  AND4_X1 U5494 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n7134)
         );
  AND4_X1 U5495 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n9295)
         );
  INV_X1 U5496 ( .A(n8699), .ZN(n8717) );
  AOI21_X1 U5497 ( .B1(n8929), .B2(n8928), .A(n8934), .ZN(n4775) );
  AND2_X1 U5498 ( .A1(n8927), .A2(n8926), .ZN(n4776) );
  INV_X1 U5499 ( .A(n8724), .ZN(n9137) );
  OAI211_X1 U5500 ( .C1(n6465), .C2(n6241), .A(n6217), .B(n6216), .ZN(n7046)
         );
  INV_X1 U5501 ( .A(n6685), .ZN(n6141) );
  NAND2_X1 U5502 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  NAND2_X1 U5503 ( .A1(n5798), .A2(n5797), .ZN(n9990) );
  NAND2_X1 U5504 ( .A1(n5514), .A2(n5513), .ZN(n8250) );
  NAND2_X1 U5505 ( .A1(n5719), .A2(n5718), .ZN(n10003) );
  NAND2_X1 U5506 ( .A1(n5836), .A2(n5835), .ZN(n9657) );
  OR2_X1 U5507 ( .A1(n9527), .A2(n5831), .ZN(n5808) );
  AOI21_X1 U5508 ( .B1(n9694), .B2(n9689), .A(n9688), .ZN(n9692) );
  OAI21_X1 U5509 ( .B1(n9742), .B2(n10288), .A(n10254), .ZN(n4857) );
  OR2_X1 U5510 ( .A1(n9743), .A2(n10288), .ZN(n4855) );
  XNOR2_X1 U5511 ( .A(n6050), .B(n8468), .ZN(n9759) );
  AOI21_X1 U5512 ( .B1(n4925), .B2(n4924), .A(n4521), .ZN(n4923) );
  NAND2_X1 U5513 ( .A1(n4927), .A2(n4925), .ZN(n6040) );
  NAND2_X1 U5514 ( .A1(n4927), .A2(n4929), .ZN(n5990) );
  NAND2_X1 U5515 ( .A1(n6777), .A2(n9926), .ZN(n10161) );
  NAND2_X1 U5516 ( .A1(n6061), .A2(n10344), .ZN(n4598) );
  AOI21_X1 U5517 ( .B1(n9759), .B2(n10332), .A(n4599), .ZN(n6061) );
  NAND2_X1 U5518 ( .A1(n4600), .A2(n4909), .ZN(n4599) );
  INV_X1 U5519 ( .A(n9760), .ZN(n4909) );
  INV_X1 U5520 ( .A(n9765), .ZN(n4600) );
  MUX2_X1 U5521 ( .A(n8756), .B(n8755), .S(n8886), .Z(n8785) );
  NAND2_X1 U5522 ( .A1(n4682), .A2(n5997), .ZN(n8216) );
  AND2_X1 U5523 ( .A1(n4683), .A2(n4684), .ZN(n4682) );
  AND2_X1 U5524 ( .A1(n8800), .A2(n8803), .ZN(n8808) );
  MUX2_X1 U5525 ( .A(n8799), .B(n8798), .S(n8886), .Z(n8800) );
  AND2_X1 U5526 ( .A1(n8797), .A2(n8809), .ZN(n8798) );
  AND2_X1 U5527 ( .A1(n4489), .A2(n8248), .ZN(n4664) );
  AND2_X1 U5528 ( .A1(n9942), .A2(n8266), .ZN(n4665) );
  NAND2_X1 U5529 ( .A1(n4796), .A2(n4517), .ZN(n8832) );
  INV_X1 U5530 ( .A(n8267), .ZN(n4666) );
  NAND2_X1 U5531 ( .A1(n4528), .A2(n4489), .ZN(n4663) );
  INV_X1 U5532 ( .A(n8871), .ZN(n4786) );
  MUX2_X1 U5533 ( .A(n8862), .B(n8861), .S(n8886), .Z(n8866) );
  OAI211_X1 U5534 ( .C1(n4672), .C2(n8328), .A(n4669), .B(n4668), .ZN(n4667)
         );
  NOR2_X1 U5535 ( .A1(n4781), .A2(n4783), .ZN(n4778) );
  AND2_X1 U5536 ( .A1(n4788), .A2(n4790), .ZN(n4783) );
  INV_X1 U5537 ( .A(n4781), .ZN(n4780) );
  NOR2_X1 U5538 ( .A1(n9135), .A2(n8743), .ZN(n4973) );
  NOR2_X1 U5539 ( .A1(n8911), .A2(n5044), .ZN(n5043) );
  INV_X1 U5540 ( .A(n7951), .ZN(n5044) );
  AND2_X1 U5541 ( .A1(n5078), .A2(n9519), .ZN(n5077) );
  NAND2_X1 U5542 ( .A1(n9587), .A2(n9585), .ZN(n5078) );
  NOR2_X1 U5543 ( .A1(n9649), .A2(n9497), .ZN(n4730) );
  OAI21_X1 U5544 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8201) );
  INV_X1 U5545 ( .A(n5871), .ZN(n4892) );
  INV_X1 U5546 ( .A(n4891), .ZN(n4890) );
  OAI21_X1 U5547 ( .B1(n5869), .B2(n4892), .A(n6041), .ZN(n4891) );
  INV_X1 U5548 ( .A(n4868), .ZN(n4865) );
  INV_X1 U5549 ( .A(n5479), .ZN(n5033) );
  NAND2_X1 U5550 ( .A1(n5141), .A2(n7598), .ZN(n5144) );
  INV_X1 U5551 ( .A(SI_14_), .ZN(n7612) );
  INV_X1 U5552 ( .A(SI_11_), .ZN(n7610) );
  INV_X1 U5553 ( .A(SI_9_), .ZN(n7598) );
  NAND2_X1 U5554 ( .A1(n7440), .A2(n7438), .ZN(n6379) );
  INV_X1 U5555 ( .A(n8667), .ZN(n5010) );
  OAI21_X1 U5556 ( .B1(n8885), .B2(n4804), .A(n4802), .ZN(n4801) );
  INV_X1 U5557 ( .A(n8884), .ZN(n4804) );
  INV_X1 U5558 ( .A(n4803), .ZN(n4802) );
  AND2_X1 U5559 ( .A1(n4507), .A2(n8888), .ZN(n4800) );
  OR2_X1 U5560 ( .A1(n8742), .A2(n6141), .ZN(n8892) );
  NAND2_X1 U5561 ( .A1(n8132), .A2(n4713), .ZN(n8982) );
  NAND2_X1 U5562 ( .A1(n7500), .A2(n7501), .ZN(n4713) );
  NOR2_X1 U5563 ( .A1(n9354), .A2(n4998), .ZN(n4997) );
  INV_X1 U5564 ( .A(n4999), .ZN(n4998) );
  OR2_X1 U5565 ( .A1(n9354), .A2(n9118), .ZN(n8884) );
  INV_X1 U5566 ( .A(n4638), .ZN(n4636) );
  INV_X1 U5567 ( .A(n4973), .ZN(n4972) );
  AOI21_X1 U5568 ( .B1(n4973), .B2(n9143), .A(n4971), .ZN(n4970) );
  INV_X1 U5569 ( .A(n8877), .ZN(n4971) );
  NOR2_X1 U5570 ( .A1(n9358), .A2(n9363), .ZN(n4999) );
  NAND2_X1 U5571 ( .A1(n9164), .A2(n8744), .ZN(n4638) );
  OR2_X1 U5572 ( .A1(n9369), .A2(n8724), .ZN(n8745) );
  AND2_X1 U5573 ( .A1(n9074), .A2(n4508), .ZN(n5067) );
  INV_X1 U5574 ( .A(n8792), .ZN(n4642) );
  NOR2_X1 U5575 ( .A1(n7233), .A2(n4644), .ZN(n4643) );
  INV_X1 U5576 ( .A(n8791), .ZN(n4644) );
  INV_X1 U5577 ( .A(n7111), .ZN(n5048) );
  AND2_X1 U5578 ( .A1(n5002), .A2(n10406), .ZN(n5001) );
  NOR2_X1 U5579 ( .A1(n7027), .A2(n7046), .ZN(n5002) );
  AND2_X1 U5580 ( .A1(n9332), .A2(n9423), .ZN(n9320) );
  OR2_X1 U5581 ( .A1(n8902), .A2(n7115), .ZN(n4648) );
  NOR2_X1 U5582 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4833) );
  INV_X1 U5583 ( .A(n9509), .ZN(n4689) );
  INV_X1 U5584 ( .A(n5784), .ZN(n4710) );
  NOR4_X1 U5585 ( .A1(n8472), .A2(n8471), .A3(n8470), .A4(n8469), .ZN(n8474)
         );
  OAI22_X1 U5586 ( .A1(n8327), .A2(n4739), .B1(n8472), .B2(n8430), .ZN(n4897)
         );
  NAND2_X1 U5587 ( .A1(n4681), .A2(n4680), .ZN(n8329) );
  NAND2_X1 U5588 ( .A1(n8338), .A2(n8328), .ZN(n4680) );
  INV_X1 U5589 ( .A(n8334), .ZN(n4627) );
  OR2_X1 U5590 ( .A1(n9979), .A2(n9799), .ZN(n8318) );
  OR2_X1 U5591 ( .A1(n6028), .A2(n9786), .ZN(n8331) );
  NOR2_X1 U5592 ( .A1(n8467), .A2(n4933), .ZN(n4932) );
  INV_X1 U5593 ( .A(n5988), .ZN(n4933) );
  INV_X1 U5594 ( .A(n5801), .ZN(n5799) );
  OR2_X1 U5595 ( .A1(n5770), .A2(n5769), .ZN(n5801) );
  NAND2_X1 U5596 ( .A1(n4735), .A2(n9861), .ZN(n4734) );
  AOI21_X1 U5597 ( .B1(n8284), .B2(n4907), .A(n8444), .ZN(n4906) );
  NOR2_X1 U5598 ( .A1(n10009), .A2(n9895), .ZN(n4735) );
  NAND2_X1 U5599 ( .A1(n4591), .A2(n5976), .ZN(n4590) );
  AOI21_X1 U5600 ( .B1(n9931), .B2(n5976), .A(n4520), .ZN(n4943) );
  INV_X1 U5601 ( .A(n5974), .ZN(n4591) );
  NOR2_X1 U5602 ( .A1(n4549), .A2(n4935), .ZN(n4934) );
  INV_X1 U5603 ( .A(n5973), .ZN(n4935) );
  NAND2_X1 U5604 ( .A1(n5217), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5541) );
  INV_X1 U5605 ( .A(n5539), .ZN(n5217) );
  NOR2_X1 U5606 ( .A1(n4490), .A2(n4569), .ZN(n4568) );
  INV_X1 U5607 ( .A(n5967), .ZN(n4569) );
  OR2_X1 U5608 ( .A1(n9497), .A2(n9645), .ZN(n8386) );
  AND2_X1 U5609 ( .A1(n6005), .A2(n8238), .ZN(n4912) );
  NAND2_X1 U5610 ( .A1(n10125), .A2(n10124), .ZN(n6004) );
  OR2_X1 U5611 ( .A1(n5516), .A2(n5515), .ZN(n5539) );
  INV_X1 U5612 ( .A(n5464), .ZN(n5216) );
  OR2_X1 U5613 ( .A1(n5446), .A2(n7473), .ZN(n5464) );
  AND2_X1 U5614 ( .A1(n8222), .A2(n8360), .ZN(n4683) );
  INV_X1 U5615 ( .A(n9815), .ZN(n9831) );
  NAND2_X1 U5616 ( .A1(n10122), .A2(n4730), .ZN(n9961) );
  INV_X1 U5617 ( .A(n7298), .ZN(n8480) );
  XNOR2_X1 U5618 ( .A(n8201), .B(n8200), .ZN(n8198) );
  NAND2_X1 U5619 ( .A1(n4876), .A2(n4874), .ZN(n5848) );
  AOI21_X1 U5620 ( .B1(n4877), .B2(n4880), .A(n4875), .ZN(n4874) );
  INV_X1 U5621 ( .A(n5817), .ZN(n4875) );
  NOR2_X1 U5622 ( .A1(n5790), .A2(n4882), .ZN(n4881) );
  INV_X1 U5623 ( .A(n5765), .ZN(n4882) );
  OAI21_X1 U5624 ( .B1(n5709), .B2(n4901), .A(n5712), .ZN(n5740) );
  INV_X1 U5625 ( .A(n5710), .ZN(n4901) );
  INV_X1 U5626 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5201) );
  AND2_X1 U5627 ( .A1(n5685), .A2(n5663), .ZN(n5683) );
  INV_X1 U5628 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5532) );
  XNOR2_X1 U5629 ( .A(n5162), .B(n7612), .ZN(n5530) );
  XNOR2_X1 U5630 ( .A(n5151), .B(n7610), .ZN(n5458) );
  NAND2_X1 U5631 ( .A1(n5146), .A2(n7828), .ZN(n5149) );
  OAI211_X1 U5632 ( .C1(n5127), .C2(n5022), .A(n5019), .B(n5024), .ZN(n5140)
         );
  INV_X1 U5633 ( .A(n5398), .ZN(n5024) );
  OR2_X1 U5634 ( .A1(n5022), .A2(n5023), .ZN(n5019) );
  INV_X1 U5635 ( .A(SI_5_), .ZN(n7656) );
  INV_X1 U5636 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5114) );
  INV_X1 U5637 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4859) );
  OR2_X1 U5638 ( .A1(n6379), .A2(n7436), .ZN(n6380) );
  OR2_X1 U5639 ( .A1(n8550), .A2(n8694), .ZN(n8564) );
  INV_X1 U5640 ( .A(n4819), .ZN(n4818) );
  OAI21_X1 U5641 ( .B1(n4821), .B2(n4820), .A(n8503), .ZN(n4819) );
  INV_X1 U5642 ( .A(n4823), .ZN(n4820) );
  OR2_X1 U5644 ( .A1(n7110), .A2(n8625), .ZN(n6239) );
  OR2_X1 U5645 ( .A1(n8653), .A2(n8652), .ZN(n8650) );
  XNOR2_X1 U5646 ( .A(n7442), .B(n8626), .ZN(n6382) );
  OR2_X1 U5647 ( .A1(n6322), .A2(n7815), .ZN(n6338) );
  AOI21_X1 U5648 ( .B1(n4827), .B2(n4829), .A(n4826), .ZN(n4825) );
  INV_X1 U5649 ( .A(n6332), .ZN(n4826) );
  NAND3_X1 U5650 ( .A1(n6191), .A2(n6173), .A3(n6883), .ZN(n6897) );
  INV_X1 U5651 ( .A(n6838), .ZN(n6191) );
  OR2_X1 U5652 ( .A1(n8087), .A2(n9009), .ZN(n8107) );
  OR2_X1 U5653 ( .A1(n8668), .A2(n5010), .ZN(n5009) );
  AOI22_X1 U5654 ( .A1(n4507), .A2(n8879), .B1(n4978), .B2(n4980), .ZN(n4975)
         );
  INV_X1 U5655 ( .A(n6175), .ZN(n8730) );
  NOR2_X1 U5656 ( .A1(n7274), .A2(n4552), .ZN(n8975) );
  NOR2_X1 U5657 ( .A1(n8975), .A2(n8976), .ZN(n8974) );
  NOR2_X1 U5658 ( .A1(n8974), .A2(n4721), .ZN(n7279) );
  AND2_X1 U5659 ( .A1(n8973), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5660 ( .A1(n7279), .A2(n7278), .ZN(n7343) );
  NAND2_X1 U5661 ( .A1(n7502), .A2(n4714), .ZN(n7504) );
  OR2_X1 U5662 ( .A1(n7503), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U5663 ( .A1(n7504), .A2(n7505), .ZN(n8132) );
  XNOR2_X1 U5664 ( .A(n8982), .B(n8983), .ZN(n8136) );
  NOR2_X1 U5665 ( .A1(n9026), .A2(n4562), .ZN(n9028) );
  NAND2_X1 U5666 ( .A1(n9028), .A2(n9029), .ZN(n9044) );
  AND2_X1 U5667 ( .A1(n9151), .A2(n4995), .ZN(n9062) );
  NOR2_X1 U5668 ( .A1(n9063), .A2(n4996), .ZN(n4995) );
  INV_X1 U5669 ( .A(n4997), .ZN(n4996) );
  NAND2_X1 U5670 ( .A1(n9115), .A2(n8725), .ZN(n9121) );
  NAND2_X1 U5671 ( .A1(n9151), .A2(n9086), .ZN(n9129) );
  INV_X1 U5672 ( .A(n8591), .ZN(n6757) );
  OR2_X1 U5673 ( .A1(n9374), .A2(n9186), .ZN(n9084) );
  INV_X1 U5674 ( .A(n8578), .ZN(n6756) );
  NOR2_X1 U5675 ( .A1(n9193), .A2(n9380), .ZN(n9176) );
  NOR2_X1 U5676 ( .A1(n9217), .A2(n5058), .ZN(n5057) );
  OAI21_X1 U5677 ( .B1(n9217), .B2(n5056), .A(n9080), .ZN(n5055) );
  INV_X1 U5678 ( .A(n5059), .ZN(n5058) );
  NOR2_X1 U5679 ( .A1(n9408), .A2(n9400), .ZN(n9224) );
  NAND2_X1 U5680 ( .A1(n9224), .A2(n9228), .ZN(n9225) );
  INV_X1 U5681 ( .A(n8523), .ZN(n6754) );
  AND2_X1 U5682 ( .A1(n8513), .A2(n8512), .ZN(n9263) );
  NAND2_X1 U5683 ( .A1(n6419), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8087) );
  INV_X1 U5684 ( .A(n6420), .ZN(n6419) );
  OAI21_X1 U5685 ( .B1(n8015), .B2(n4969), .A(n4967), .ZN(n9341) );
  INV_X1 U5686 ( .A(n4968), .ZN(n4967) );
  OAI21_X1 U5687 ( .B1(n4969), .B2(n9070), .A(n8829), .ZN(n4968) );
  AND2_X1 U5688 ( .A1(n9069), .A2(n5038), .ZN(n5037) );
  INV_X1 U5689 ( .A(n6393), .ZN(n6132) );
  NAND2_X1 U5690 ( .A1(n4991), .A2(n4987), .ZN(n8050) );
  AND2_X1 U5691 ( .A1(n4988), .A2(n4501), .ZN(n4987) );
  OAI21_X1 U5692 ( .B1(n7950), .B2(n5042), .A(n5040), .ZN(n9071) );
  NOR2_X1 U5693 ( .A1(n4990), .A2(n7964), .ZN(n8026) );
  NAND2_X1 U5694 ( .A1(n4992), .A2(n10435), .ZN(n4990) );
  AND2_X1 U5695 ( .A1(n8817), .A2(n8809), .ZN(n4982) );
  AND4_X1 U5696 ( .A1(n6344), .A2(n6343), .A3(n6342), .A4(n6341), .ZN(n7955)
         );
  AND2_X1 U5697 ( .A1(n8907), .A2(n7312), .ZN(n5072) );
  NAND2_X1 U5698 ( .A1(n7241), .A2(n8791), .ZN(n7243) );
  AND2_X1 U5699 ( .A1(n8794), .A2(n8792), .ZN(n8806) );
  AND4_X1 U5700 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n7310)
         );
  OR2_X1 U5701 ( .A1(n7199), .A2(n7332), .ZN(n7249) );
  AND4_X1 U5702 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6271), .ZN(n7194)
         );
  NAND2_X1 U5703 ( .A1(n8902), .A2(n4647), .ZN(n4645) );
  NAND2_X1 U5704 ( .A1(n5001), .A2(n7138), .ZN(n10366) );
  AND2_X1 U5705 ( .A1(n5002), .A2(n7138), .ZN(n10367) );
  AND4_X1 U5706 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n7120)
         );
  NAND2_X1 U5707 ( .A1(n7138), .A2(n7035), .ZN(n7042) );
  NAND2_X1 U5708 ( .A1(n4650), .A2(n8775), .ZN(n4649) );
  NAND2_X1 U5709 ( .A1(n9271), .A2(n9263), .ZN(n9408) );
  NAND2_X1 U5710 ( .A1(n6410), .A2(n6409), .ZN(n9429) );
  OR2_X1 U5711 ( .A1(n6091), .A2(n6090), .ZN(n6095) );
  NAND2_X1 U5712 ( .A1(n6074), .A2(n6073), .ZN(n6114) );
  AND2_X1 U5713 ( .A1(n6072), .A2(n7083), .ZN(n4835) );
  NAND2_X1 U5714 ( .A1(n4836), .A2(n6072), .ZN(n7082) );
  OR2_X1 U5715 ( .A1(n6285), .A2(n6284), .ZN(n6302) );
  AND2_X1 U5716 ( .A1(n6263), .A2(n6245), .ZN(n6572) );
  INV_X1 U5717 ( .A(n4692), .ZN(n9486) );
  OR2_X1 U5718 ( .A1(n5748), .A2(n5747), .ZN(n5770) );
  XNOR2_X1 U5719 ( .A(n5301), .B(n6782), .ZN(n5325) );
  NAND2_X1 U5720 ( .A1(n9616), .A2(n9619), .ZN(n4690) );
  NAND2_X1 U5721 ( .A1(n5214), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5406) );
  INV_X1 U5722 ( .A(n5382), .ZN(n5214) );
  AND2_X1 U5723 ( .A1(n9596), .A2(n5090), .ZN(n5089) );
  INV_X1 U5724 ( .A(n5760), .ZN(n5090) );
  AND2_X1 U5725 ( .A1(n5417), .A2(n5433), .ZN(n4705) );
  NAND2_X1 U5726 ( .A1(n7299), .A2(n7302), .ZN(n5417) );
  NAND2_X1 U5727 ( .A1(n5416), .A2(n5080), .ZN(n7300) );
  OR2_X1 U5728 ( .A1(n5406), .A2(n7303), .ZN(n5423) );
  NAND2_X1 U5729 ( .A1(n5215), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5446) );
  INV_X1 U5730 ( .A(n5423), .ZN(n5215) );
  NAND2_X1 U5731 ( .A1(n5644), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5667) );
  INV_X1 U5732 ( .A(n5646), .ZN(n5644) );
  NAND2_X1 U5733 ( .A1(n5690), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5722) );
  INV_X1 U5734 ( .A(n5692), .ZN(n5690) );
  INV_X1 U5735 ( .A(n6651), .ZN(n4753) );
  NAND2_X1 U5736 ( .A1(n4747), .A2(n4746), .ZN(n4751) );
  INV_X1 U5737 ( .A(n5285), .ZN(n4746) );
  NAND2_X1 U5738 ( .A1(n5284), .A2(n5285), .ZN(n5286) );
  NAND2_X1 U5739 ( .A1(n5631), .A2(n5630), .ZN(n9617) );
  INV_X1 U5740 ( .A(n4697), .ZN(n4696) );
  OAI21_X1 U5741 ( .B1(n4756), .B2(n5550), .A(n4693), .ZN(n4697) );
  AND2_X1 U5742 ( .A1(n4694), .A2(n5556), .ZN(n4693) );
  INV_X1 U5743 ( .A(n5302), .ZN(n5928) );
  NAND2_X1 U5744 ( .A1(n6613), .A2(n6612), .ZN(n6611) );
  OAI21_X1 U5745 ( .B1(n6466), .B2(n7256), .A(n4564), .ZN(n6607) );
  NAND2_X1 U5746 ( .A1(n6466), .A2(n7256), .ZN(n4564) );
  OR2_X1 U5747 ( .A1(n6442), .A2(n6441), .ZN(n4851) );
  NOR2_X1 U5748 ( .A1(n10233), .A2(n10232), .ZN(n10235) );
  AND2_X1 U5749 ( .A1(n10249), .A2(n10250), .ZN(n10247) );
  NOR2_X1 U5750 ( .A1(n10247), .A2(n4839), .ZN(n6635) );
  NOR2_X1 U5751 ( .A1(n10253), .A2(n4840), .ZN(n4839) );
  INV_X1 U5752 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U5753 ( .A1(n6635), .A2(n6634), .ZN(n6711) );
  AND2_X1 U5754 ( .A1(n6702), .A2(n6703), .ZN(n10262) );
  NAND2_X1 U5755 ( .A1(n6711), .A2(n4838), .ZN(n10266) );
  OR2_X1 U5756 ( .A1(n6712), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4838) );
  NAND2_X1 U5757 ( .A1(n10266), .A2(n10265), .ZN(n10264) );
  INV_X1 U5758 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7303) );
  INV_X1 U5759 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U5760 ( .A1(n10275), .A2(n4563), .ZN(n10294) );
  OR2_X1 U5761 ( .A1(n10290), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U5762 ( .A1(n10294), .A2(n10295), .ZN(n10293) );
  NAND2_X1 U5763 ( .A1(n6717), .A2(n6718), .ZN(n6875) );
  OAI21_X1 U5764 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6876), .A(n6875), .ZN(
        n6877) );
  AOI21_X1 U5765 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9687) );
  INV_X1 U5766 ( .A(n4932), .ZN(n4924) );
  NAND2_X1 U5767 ( .A1(n5827), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5878) );
  INV_X1 U5768 ( .A(n5829), .ZN(n5827) );
  INV_X1 U5769 ( .A(n4930), .ZN(n4929) );
  OAI22_X1 U5770 ( .A1(n8467), .A2(n4931), .B1(n9979), .B2(n9656), .ZN(n4930)
         );
  NAND2_X1 U5771 ( .A1(n5989), .A2(n5988), .ZN(n4931) );
  INV_X1 U5772 ( .A(n4624), .ZN(n4623) );
  OAI21_X1 U5773 ( .B1(n4625), .B2(n4914), .A(n8353), .ZN(n4624) );
  OAI21_X1 U5774 ( .B1(n5982), .B2(n4577), .A(n4574), .ZN(n9808) );
  AOI21_X1 U5775 ( .B1(n4576), .B2(n4575), .A(n4498), .ZN(n4574) );
  INV_X1 U5776 ( .A(n4580), .ZN(n4575) );
  NOR3_X1 U5777 ( .A1(n9908), .A2(n4734), .A3(n9998), .ZN(n9830) );
  NOR2_X1 U5778 ( .A1(n9908), .A2(n9895), .ZN(n9894) );
  NOR2_X1 U5779 ( .A1(n9908), .A2(n4733), .ZN(n9871) );
  INV_X1 U5780 ( .A(n4735), .ZN(n4733) );
  AND2_X1 U5781 ( .A1(n8276), .A2(n8398), .ZN(n9903) );
  NAND2_X1 U5782 ( .A1(n5594), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5619) );
  OR2_X1 U5783 ( .A1(n5619), .A2(n5618), .ZN(n5646) );
  NAND2_X1 U5784 ( .A1(n5975), .A2(n5974), .ZN(n9932) );
  AND2_X1 U5785 ( .A1(n10122), .A2(n4726), .ZN(n9938) );
  NOR2_X1 U5786 ( .A1(n10030), .A2(n4728), .ZN(n4726) );
  AND2_X1 U5787 ( .A1(n9951), .A2(n8389), .ZN(n8261) );
  AOI21_X1 U5788 ( .B1(n4912), .B2(n4606), .A(n4605), .ZN(n4604) );
  INV_X1 U5789 ( .A(n8386), .ZN(n4605) );
  INV_X1 U5790 ( .A(n4912), .ZN(n4607) );
  NAND2_X1 U5791 ( .A1(n4937), .A2(n5971), .ZN(n8117) );
  NOR2_X1 U5792 ( .A1(n4524), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U5793 ( .A1(n6004), .A2(n8238), .ZN(n8034) );
  NAND2_X1 U5794 ( .A1(n6004), .A2(n4912), .ZN(n8036) );
  NOR2_X1 U5795 ( .A1(n10141), .A2(n7994), .ZN(n10120) );
  AND2_X1 U5796 ( .A1(n10120), .A2(n10171), .ZN(n10122) );
  NAND2_X1 U5797 ( .A1(n4725), .A2(n4724), .ZN(n10141) );
  OR2_X1 U5798 ( .A1(n4587), .A2(n5964), .ZN(n4586) );
  INV_X1 U5799 ( .A(n5963), .ZN(n4587) );
  NOR2_X1 U5800 ( .A1(n7362), .A2(n7361), .ZN(n7448) );
  NAND2_X1 U5801 ( .A1(n7070), .A2(n5961), .ZN(n7400) );
  AOI21_X1 U5802 ( .B1(n6822), .B2(n6000), .A(n5999), .ZN(n7067) );
  AND2_X1 U5803 ( .A1(n8219), .A2(n5959), .ZN(n4918) );
  NAND2_X1 U5804 ( .A1(n5212), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5354) );
  NOR2_X1 U5805 ( .A1(n7154), .A2(n9575), .ZN(n6911) );
  NAND2_X1 U5806 ( .A1(n5997), .A2(n4683), .ZN(n8213) );
  NAND2_X1 U5807 ( .A1(n5952), .A2(n5994), .ZN(n6964) );
  INV_X1 U5808 ( .A(n9668), .ZN(n6965) );
  NOR2_X1 U5809 ( .A1(n5949), .A2(n6851), .ZN(n6970) );
  NAND2_X1 U5810 ( .A1(n6002), .A2(n8370), .ZN(n10146) );
  NAND2_X1 U5811 ( .A1(n4632), .A2(n4630), .ZN(n7010) );
  NAND2_X1 U5812 ( .A1(n6474), .A2(n5363), .ZN(n4632) );
  NOR2_X1 U5813 ( .A1(n4513), .A2(n4631), .ZN(n4630) );
  NOR2_X1 U5814 ( .A1(n5364), .A2(n10253), .ZN(n4631) );
  AND2_X1 U5815 ( .A1(n4915), .A2(n4537), .ZN(n10321) );
  OR2_X1 U5816 ( .A1(n6472), .A2(n5347), .ZN(n4915) );
  OR2_X1 U5817 ( .A1(n6960), .A2(n8480), .ZN(n10313) );
  OR2_X1 U5818 ( .A1(n6960), .A2(n6848), .ZN(n10329) );
  OR2_X1 U5819 ( .A1(n8328), .A2(n8480), .ZN(n10102) );
  AND2_X1 U5820 ( .A1(n5899), .A2(n5898), .ZN(n6482) );
  INV_X1 U5821 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4593) );
  XNOR2_X1 U5822 ( .A(n8198), .B(SI_30_), .ZN(n9460) );
  XNOR2_X1 U5823 ( .A(n8195), .B(n6047), .ZN(n9464) );
  XNOR2_X1 U5824 ( .A(n5848), .B(n5847), .ZN(n8493) );
  XNOR2_X1 U5825 ( .A(n5819), .B(n5818), .ZN(n8586) );
  NAND2_X1 U5826 ( .A1(n4886), .A2(n5789), .ZN(n5819) );
  NAND2_X1 U5827 ( .A1(n4883), .A2(n4881), .ZN(n4886) );
  NOR2_X1 U5828 ( .A1(n4761), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4760) );
  INV_X1 U5829 ( .A(n4761), .ZN(n4759) );
  NAND2_X1 U5830 ( .A1(n4883), .A2(n5765), .ZN(n5791) );
  AND2_X1 U5831 ( .A1(n5765), .A2(n5744), .ZN(n5763) );
  INV_X1 U5832 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U5833 ( .A1(n4866), .A2(n4868), .ZN(n5613) );
  NAND2_X1 U5834 ( .A1(n4867), .A2(n4872), .ZN(n4866) );
  INV_X1 U5835 ( .A(n5562), .ZN(n4867) );
  XNOR2_X1 U5836 ( .A(n5507), .B(n5506), .ZN(n6670) );
  INV_X1 U5837 ( .A(n5028), .ZN(n5027) );
  NAND2_X1 U5838 ( .A1(n4894), .A2(n5152), .ZN(n5480) );
  XNOR2_X1 U5839 ( .A(n5457), .B(n5458), .ZN(n6499) );
  NAND2_X1 U5840 ( .A1(n5150), .A2(n5149), .ZN(n5457) );
  XNOR2_X1 U5841 ( .A(n5437), .B(n5102), .ZN(n6506) );
  OAI21_X1 U5842 ( .B1(n5018), .B2(n5021), .A(n5020), .ZN(n5025) );
  INV_X1 U5843 ( .A(n5023), .ZN(n5021) );
  NAND2_X1 U5844 ( .A1(n5361), .A2(n4902), .ZN(n5373) );
  INV_X1 U5845 ( .A(n5362), .ZN(n4902) );
  XNOR2_X1 U5846 ( .A(n5361), .B(n5362), .ZN(n6474) );
  NAND2_X1 U5847 ( .A1(n5124), .A2(n5123), .ZN(n5340) );
  XNOR2_X1 U5848 ( .A(n5125), .B(n7656), .ZN(n5341) );
  INV_X1 U5849 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5168) );
  OR3_X1 U5850 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n5295) );
  AND2_X1 U5851 ( .A1(n6279), .A2(n6261), .ZN(n4834) );
  NAND2_X1 U5852 ( .A1(n6936), .A2(n6261), .ZN(n6815) );
  NAND2_X1 U5853 ( .A1(n6386), .A2(n6385), .ZN(n7524) );
  AND2_X1 U5854 ( .A1(n6381), .A2(n6380), .ZN(n6386) );
  XNOR2_X1 U5855 ( .A(n8572), .B(n8573), .ZN(n8642) );
  NAND2_X1 U5856 ( .A1(n7177), .A2(n6316), .ZN(n7184) );
  AND2_X1 U5857 ( .A1(n6840), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8630) );
  INV_X1 U5858 ( .A(n5014), .ZN(n5013) );
  OAI21_X1 U5859 ( .B1(n8687), .B2(n5015), .A(n8532), .ZN(n5014) );
  NAND2_X1 U5860 ( .A1(n8080), .A2(n8079), .ZN(n8083) );
  NAND2_X1 U5861 ( .A1(n8100), .A2(n8099), .ZN(n8165) );
  XNOR2_X1 U5862 ( .A(n6239), .B(n6237), .ZN(n6983) );
  NAND2_X1 U5863 ( .A1(n4770), .A2(n6303), .ZN(n7460) );
  INV_X1 U5864 ( .A(n8945), .ZN(n8183) );
  NAND2_X1 U5865 ( .A1(n8650), .A2(n8519), .ZN(n8688) );
  XNOR2_X1 U5866 ( .A(n6382), .B(n6383), .ZN(n7440) );
  NAND2_X1 U5867 ( .A1(n6883), .A2(n6173), .ZN(n6839) );
  NAND2_X1 U5868 ( .A1(n8100), .A2(n4821), .ZN(n4817) );
  NAND2_X1 U5869 ( .A1(n8170), .A2(n8169), .ZN(n9413) );
  NAND2_X1 U5870 ( .A1(n4814), .A2(n5004), .ZN(n8706) );
  NAND2_X1 U5871 ( .A1(n5003), .A2(n5008), .ZN(n8708) );
  NAND2_X1 U5872 ( .A1(n8666), .A2(n5009), .ZN(n5003) );
  INV_X1 U5873 ( .A(n8714), .ZN(n8696) );
  INV_X1 U5874 ( .A(n8630), .ZN(n8710) );
  INV_X1 U5875 ( .A(n8723), .ZN(n9186) );
  OR2_X1 U5876 ( .A1(n6521), .A2(n10380), .ZN(n8936) );
  INV_X1 U5877 ( .A(n4720), .ZN(n6580) );
  NOR2_X1 U5878 ( .A1(n6549), .A2(n6548), .ZN(n6566) );
  AND2_X1 U5879 ( .A1(n4720), .A2(n4719), .ZN(n6549) );
  NAND2_X1 U5880 ( .A1(n6556), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4719) );
  INV_X1 U5881 ( .A(n4718), .ZN(n6727) );
  INV_X1 U5882 ( .A(n4716), .ZN(n6854) );
  AND2_X1 U5883 ( .A1(n6537), .A2(n6535), .ZN(n10347) );
  NAND2_X1 U5884 ( .A1(n8735), .A2(n8734), .ZN(n9350) );
  INV_X1 U5885 ( .A(n9111), .ZN(n9362) );
  OAI21_X1 U5886 ( .B1(n9127), .B2(n5053), .A(n5051), .ZN(n9109) );
  NAND2_X1 U5887 ( .A1(n9146), .A2(n8748), .ZN(n9134) );
  NAND2_X1 U5888 ( .A1(n9183), .A2(n8751), .ZN(n9165) );
  AND2_X1 U5889 ( .A1(n9219), .A2(n9218), .ZN(n9391) );
  OAI21_X1 U5890 ( .B1(n9245), .B2(n5060), .A(n5059), .ZN(n9212) );
  NAND2_X1 U5891 ( .A1(n4965), .A2(n8853), .ZN(n9235) );
  AND2_X1 U5892 ( .A1(n4965), .A2(n4963), .ZN(n9233) );
  NOR2_X1 U5893 ( .A1(n9405), .A2(n5063), .ZN(n9223) );
  NOR2_X1 U5894 ( .A1(n4948), .A2(n4950), .ZN(n9259) );
  INV_X1 U5895 ( .A(n4952), .ZN(n4948) );
  INV_X1 U5896 ( .A(n9263), .ZN(n9407) );
  OAI21_X1 U5897 ( .B1(n4953), .B2(n4958), .A(n8754), .ZN(n9276) );
  INV_X1 U5898 ( .A(n9306), .ZN(n4953) );
  NAND2_X1 U5899 ( .A1(n9303), .A2(n5100), .ZN(n9284) );
  NAND2_X1 U5900 ( .A1(n8068), .A2(n8067), .ZN(n9324) );
  OR2_X1 U5901 ( .A1(n8055), .A2(n4969), .ZN(n8718) );
  NAND2_X1 U5902 ( .A1(n5045), .A2(n7951), .ZN(n8011) );
  NAND2_X1 U5903 ( .A1(n7950), .A2(n8897), .ZN(n5045) );
  NAND2_X1 U5904 ( .A1(n4983), .A2(n8809), .ZN(n7952) );
  NAND2_X1 U5905 ( .A1(n7112), .A2(n7111), .ZN(n10356) );
  NAND2_X1 U5906 ( .A1(n6688), .A2(n8765), .ZN(n7131) );
  NAND2_X1 U5907 ( .A1(n5071), .A2(n6792), .ZN(n7137) );
  INV_X1 U5908 ( .A(n9325), .ZN(n9338) );
  AND2_X1 U5909 ( .A1(n9328), .A2(n7034), .ZN(n9349) );
  NOR2_X1 U5910 ( .A1(n9356), .A2(n4653), .ZN(n4652) );
  INV_X2 U5911 ( .A(n10442), .ZN(n10444) );
  NAND2_X1 U5912 ( .A1(n10379), .A2(n10378), .ZN(n10383) );
  AND2_X1 U5913 ( .A1(n4986), .A2(n4985), .ZN(n4984) );
  INV_X1 U5914 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4985) );
  INV_X1 U5915 ( .A(n6126), .ZN(n9461) );
  NAND2_X1 U5916 ( .A1(n6110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6078) );
  INV_X1 U5917 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6507) );
  INV_X1 U5918 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6498) );
  INV_X1 U5919 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6490) );
  NOR2_X1 U5920 ( .A1(n6184), .A2(n4722), .ZN(n8960) );
  OAI22_X1 U5921 ( .A1(n6182), .A2(n4723), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        P2_IR_REG_2__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5922 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4723) );
  NOR2_X1 U5923 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6182) );
  AOI21_X1 U5924 ( .B1(n4491), .B2(n4711), .A(n4550), .ZN(n4708) );
  AOI21_X1 U5925 ( .B1(n9998), .B2(n5265), .A(n5759), .ZN(n9502) );
  XNOR2_X1 U5926 ( .A(n5325), .B(n5326), .ZN(n6806) );
  NAND2_X1 U5927 ( .A1(n5643), .A2(n5642), .ZN(n9910) );
  NAND2_X1 U5928 ( .A1(n4685), .A2(n5352), .ZN(n4687) );
  INV_X1 U5929 ( .A(n4686), .ZN(n4685) );
  INV_X1 U5930 ( .A(n10321), .ZN(n9545) );
  NAND2_X1 U5931 ( .A1(n9534), .A2(n5585), .ZN(n9553) );
  INV_X1 U5932 ( .A(n4699), .ZN(n4698) );
  NAND2_X1 U5933 ( .A1(n7299), .A2(n4518), .ZN(n4701) );
  CLKBUF_X1 U5934 ( .A(n9648), .Z(n9612) );
  NAND2_X1 U5935 ( .A1(n5617), .A2(n5616), .ZN(n10025) );
  OR2_X1 U5936 ( .A1(n5940), .A2(n10208), .ZN(n9578) );
  NAND2_X1 U5937 ( .A1(n5086), .A2(n5816), .ZN(n4754) );
  NAND2_X1 U5938 ( .A1(n9525), .A2(n9526), .ZN(n5086) );
  INV_X1 U5939 ( .A(n9578), .ZN(n9640) );
  OAI211_X1 U5940 ( .C1(n4678), .C2(n5105), .A(n8484), .B(n4677), .ZN(n4676)
         );
  NAND2_X1 U5941 ( .A1(n4678), .A2(n4495), .ZN(n4677) );
  NAND2_X1 U5942 ( .A1(n5248), .A2(n5918), .ZN(n8486) );
  NAND2_X1 U5943 ( .A1(n5288), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U5944 ( .A1(n5288), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5241) );
  INV_X1 U5945 ( .A(n4851), .ZN(n6627) );
  NAND2_X1 U5946 ( .A1(n4851), .A2(n4850), .ZN(n10219) );
  NAND2_X1 U5947 ( .A1(n6628), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4850) );
  OAI22_X1 U5948 ( .A1(n10219), .A2(n10220), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n10222), .ZN(n10242) );
  AND2_X1 U5949 ( .A1(n5443), .A2(n5459), .ZN(n10304) );
  NOR2_X1 U5950 ( .A1(n10279), .A2(n4843), .ZN(n10299) );
  AND2_X1 U5951 ( .A1(n10290), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4843) );
  NOR2_X1 U5952 ( .A1(n10299), .A2(n10298), .ZN(n10297) );
  INV_X1 U5953 ( .A(n4842), .ZN(n7487) );
  NOR2_X1 U5954 ( .A1(n9680), .A2(n10170), .ZN(n9693) );
  AND2_X1 U5955 ( .A1(n4849), .A2(n4848), .ZN(n9710) );
  NAND2_X1 U5956 ( .A1(n4845), .A2(n4846), .ZN(n9727) );
  AND2_X1 U5957 ( .A1(n4845), .A2(n4844), .ZN(n9731) );
  AND2_X1 U5958 ( .A1(n4846), .A2(n4560), .ZN(n4844) );
  NOR2_X1 U5959 ( .A1(n9755), .A2(n4738), .ZN(n4736) );
  NAND2_X1 U5960 ( .A1(n4910), .A2(n6058), .ZN(n9765) );
  NAND2_X1 U5961 ( .A1(n4911), .A2(n10152), .ZN(n4910) );
  OAI22_X1 U5962 ( .A1(n9786), .A2(n9957), .B1(n9749), .B2(n8408), .ZN(n6057)
         );
  NAND2_X1 U5963 ( .A1(n4928), .A2(n5988), .ZN(n9777) );
  NAND2_X1 U5964 ( .A1(n9823), .A2(n4913), .ZN(n9795) );
  NAND2_X1 U5965 ( .A1(n9823), .A2(n8297), .ZN(n9810) );
  NAND2_X1 U5966 ( .A1(n4579), .A2(n5983), .ZN(n9822) );
  NAND2_X1 U5967 ( .A1(n5982), .A2(n4580), .ZN(n4579) );
  NAND2_X1 U5968 ( .A1(n9850), .A2(n8295), .ZN(n9825) );
  NAND2_X1 U5969 ( .A1(n4908), .A2(n8442), .ZN(n9846) );
  NAND2_X1 U5970 ( .A1(n5982), .A2(n5981), .ZN(n9839) );
  NAND2_X1 U5971 ( .A1(n4942), .A2(n5980), .ZN(n9855) );
  NAND2_X1 U5972 ( .A1(n9890), .A2(n8284), .ZN(n9879) );
  OR2_X1 U5973 ( .A1(n9932), .A2(n9931), .ZN(n10024) );
  NAND2_X1 U5974 ( .A1(n4620), .A2(n8269), .ZN(n9918) );
  NAND2_X1 U5975 ( .A1(n6006), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U5976 ( .A1(n6006), .A2(n8391), .ZN(n9943) );
  NAND2_X1 U5977 ( .A1(n4936), .A2(n5973), .ZN(n9937) );
  NAND2_X1 U5978 ( .A1(n5970), .A2(n5969), .ZN(n8032) );
  AOI21_X1 U5979 ( .B1(n4573), .B2(n4920), .A(n4490), .ZN(n4570) );
  NAND2_X1 U5980 ( .A1(n10138), .A2(n5967), .ZN(n4573) );
  NAND2_X1 U5981 ( .A1(n4919), .A2(n5967), .ZN(n7939) );
  OR2_X1 U5982 ( .A1(n10138), .A2(n4530), .ZN(n4919) );
  NAND2_X1 U5983 ( .A1(n7398), .A2(n5963), .ZN(n7360) );
  NAND2_X1 U5984 ( .A1(n4565), .A2(n6826), .ZN(n6827) );
  INV_X1 U5985 ( .A(n5958), .ZN(n4565) );
  AND2_X1 U5986 ( .A1(n10161), .A2(n6850), .ZN(n10143) );
  OAI21_X1 U5987 ( .B1(n9776), .B2(n10036), .A(n6021), .ZN(n6022) );
  INV_X1 U5988 ( .A(n9801), .ZN(n10054) );
  NAND2_X1 U5989 ( .A1(n5872), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4673) );
  XNOR2_X1 U5990 ( .A(n6042), .B(n6041), .ZN(n10091) );
  NAND2_X1 U5991 ( .A1(n4889), .A2(n5871), .ZN(n6042) );
  XNOR2_X1 U5992 ( .A(n5764), .B(n5763), .ZN(n8561) );
  XNOR2_X1 U5993 ( .A(n5231), .B(n5230), .ZN(n7458) );
  INV_X1 U5994 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U5995 ( .A1(n5229), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  INV_X1 U5996 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7841) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7855) );
  AND2_X1 U5998 ( .A1(n5403), .A2(n5438), .ZN(n10272) );
  XNOR2_X1 U5999 ( .A(n5340), .B(n5341), .ZN(n6472) );
  NAND2_X1 U6000 ( .A1(n5293), .A2(n5294), .ZN(n4610) );
  OR2_X1 U6001 ( .A1(n5277), .A2(n5508), .ZN(n5278) );
  NOR2_X1 U6002 ( .A1(n7557), .A2(n10485), .ZN(n10484) );
  AOI21_X1 U6003 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10482), .ZN(n10481) );
  NOR2_X1 U6004 ( .A1(n10481), .A2(n10480), .ZN(n10479) );
  AND2_X1 U6005 ( .A1(n8621), .A2(n4551), .ZN(n4812) );
  AOI21_X1 U6006 ( .B1(n8666), .B2(n4807), .A(n4806), .ZN(n4813) );
  NAND2_X1 U6007 ( .A1(n4774), .A2(n4773), .ZN(P2_U3244) );
  AND2_X1 U6008 ( .A1(n4946), .A2(n8935), .ZN(n4773) );
  OAI21_X1 U6009 ( .B1(n8925), .B2(n4776), .A(n4775), .ZN(n4774) );
  AOI21_X1 U6010 ( .B1(n10306), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9746), .ZN(
        n4852) );
  OAI21_X1 U6011 ( .B1(n4493), .B2(n4857), .A(n8190), .ZN(n4856) );
  NAND2_X1 U6012 ( .A1(n4598), .A2(n4597), .ZN(n6060) );
  OR2_X1 U6013 ( .A1(n10344), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4597) );
  NOR2_X1 U6014 ( .A1(n4544), .A2(n4613), .ZN(n4612) );
  NOR2_X1 U6015 ( .A1(n10336), .A2(n6062), .ZN(n4613) );
  AND2_X1 U6016 ( .A1(n5004), .A2(n4545), .ZN(n4488) );
  AND2_X1 U6017 ( .A1(n8261), .A2(n8260), .ZN(n4489) );
  AND2_X1 U6018 ( .A1(n7994), .A2(n10150), .ZN(n4490) );
  AND4_X1 U6019 ( .A1(n4763), .A2(n4762), .A3(n5175), .A4(n4535), .ZN(n5189)
         );
  AND2_X1 U6020 ( .A1(n4529), .A2(n4709), .ZN(n4491) );
  NAND2_X1 U6021 ( .A1(n4594), .A2(n4596), .ZN(n4492) );
  AOI21_X1 U6022 ( .B1(n5561), .B2(n5560), .A(n4873), .ZN(n4872) );
  INV_X1 U6023 ( .A(n5415), .ZN(n5080) );
  AND2_X1 U6024 ( .A1(n9744), .A2(n10284), .ZN(n4493) );
  AND2_X1 U6025 ( .A1(n4943), .A2(n4590), .ZN(n4494) );
  OR2_X1 U6026 ( .A1(n9374), .A2(n8723), .ZN(n8744) );
  NAND2_X1 U6027 ( .A1(n6352), .A2(n6351), .ZN(n8010) );
  OR2_X1 U6028 ( .A1(n9586), .A2(n9587), .ZN(n9584) );
  AND2_X1 U6029 ( .A1(n8436), .A2(n4895), .ZN(n4495) );
  AND2_X1 U6030 ( .A1(n4559), .A2(n5371), .ZN(n4496) );
  NAND2_X1 U6031 ( .A1(n4861), .A2(n8197), .ZN(n9755) );
  INV_X1 U6032 ( .A(n9755), .ZN(n4860) );
  AND2_X1 U6033 ( .A1(n4545), .A2(n8611), .ZN(n4497) );
  AND2_X1 U6034 ( .A1(n10059), .A2(n9848), .ZN(n4498) );
  AND2_X1 U6035 ( .A1(n5611), .A2(SI_17_), .ZN(n4499) );
  NOR2_X1 U6036 ( .A1(n8010), .A2(n8141), .ZN(n4500) );
  AND2_X1 U6037 ( .A1(n4500), .A2(n4989), .ZN(n4501) );
  NOR2_X1 U6038 ( .A1(n7378), .A2(n7924), .ZN(n4992) );
  INV_X1 U6039 ( .A(n6683), .ZN(n4837) );
  OR3_X1 U6040 ( .A1(n8598), .A2(n8724), .A3(n8502), .ZN(n4502) );
  INV_X1 U6041 ( .A(n8897), .ZN(n5041) );
  NAND2_X1 U6042 ( .A1(n5478), .A2(n5477), .ZN(n7983) );
  NOR2_X1 U6043 ( .A1(n6418), .A2(n6118), .ZN(n8705) );
  NAND2_X1 U6044 ( .A1(n5462), .A2(n5461), .ZN(n10140) );
  INV_X1 U6045 ( .A(n10140), .ZN(n4724) );
  NAND2_X1 U6046 ( .A1(n4648), .A2(n4647), .ZN(n7117) );
  AND2_X1 U6047 ( .A1(n5352), .A2(n5092), .ZN(n9542) );
  NAND2_X1 U6048 ( .A1(n6336), .A2(n6335), .ZN(n7964) );
  AND2_X1 U6049 ( .A1(n4991), .A2(n4992), .ZN(n4503) );
  INV_X1 U6050 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6183) );
  INV_X1 U6051 ( .A(n6194), .ZN(n8556) );
  AND2_X1 U6052 ( .A1(n5221), .A2(n10083), .ZN(n5302) );
  AND2_X1 U6053 ( .A1(n5035), .A2(n5034), .ZN(n6184) );
  INV_X1 U6054 ( .A(n8189), .ZN(n6790) );
  AND2_X1 U6055 ( .A1(n6184), .A2(n6063), .ZN(n6200) );
  NAND2_X1 U6056 ( .A1(n10140), .A2(n7992), .ZN(n4504) );
  NAND4_X1 U6057 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n5950)
         );
  NAND2_X1 U6058 ( .A1(n6790), .A2(n6695), .ZN(n6688) );
  NAND4_X1 U6059 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n5955)
         );
  AND2_X1 U6060 ( .A1(n5962), .A2(n5961), .ZN(n4505) );
  OR2_X1 U6061 ( .A1(n5132), .A2(n5131), .ZN(n4506) );
  INV_X1 U6062 ( .A(n4914), .ZN(n4913) );
  NAND2_X1 U6063 ( .A1(n8302), .A2(n8297), .ZN(n4914) );
  NAND2_X1 U6064 ( .A1(n5560), .A2(n5167), .ZN(n5561) );
  OR2_X1 U6065 ( .A1(n9063), .A2(n8736), .ZN(n4507) );
  NAND2_X1 U6066 ( .A1(n5898), .A2(n5199), .ZN(n5248) );
  NAND2_X1 U6067 ( .A1(n8563), .A2(n8562), .ZN(n9383) );
  OR2_X1 U6068 ( .A1(n8010), .A2(n8017), .ZN(n8818) );
  INV_X1 U6069 ( .A(n10410), .ZN(n5000) );
  NAND2_X1 U6070 ( .A1(n9584), .A2(n9585), .ZN(n9518) );
  OR2_X1 U6071 ( .A1(n9420), .A2(n9278), .ZN(n4508) );
  NAND2_X1 U6072 ( .A1(n6071), .A2(n6200), .ZN(n6083) );
  AND2_X1 U6073 ( .A1(n6597), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U6074 ( .A1(n5017), .A2(n4506), .ZN(n5022) );
  NAND4_X1 U6075 ( .A1(n5243), .A2(n5241), .A3(n5242), .A4(n5240), .ZN(n9670)
         );
  AND2_X1 U6076 ( .A1(n8744), .A2(n8751), .ZN(n4510) );
  AND2_X1 U6077 ( .A1(n8825), .A2(n8824), .ZN(n9070) );
  INV_X1 U6078 ( .A(n9070), .ZN(n5039) );
  XOR2_X1 U6079 ( .A(n8337), .B(n8338), .Z(n8468) );
  AND4_X1 U6080 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n4511)
         );
  NAND2_X1 U6081 ( .A1(n5537), .A2(n5536), .ZN(n9497) );
  OR2_X1 U6082 ( .A1(n6241), .A2(n6467), .ZN(n4512) );
  OAI21_X1 U6083 ( .B1(n5785), .B2(n4711), .A(n4491), .ZN(n9627) );
  AND2_X1 U6084 ( .A1(n4483), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U6085 ( .A1(n5655), .A2(n4691), .ZN(n9586) );
  NAND2_X1 U6086 ( .A1(n9369), .A2(n8724), .ZN(n8748) );
  NAND2_X1 U6087 ( .A1(n8745), .A2(n8748), .ZN(n9143) );
  AND2_X1 U6088 ( .A1(n8909), .A2(n7369), .ZN(n4514) );
  OR2_X1 U6089 ( .A1(n9998), .A2(n9829), .ZN(n8295) );
  INV_X1 U6090 ( .A(n8295), .ZN(n4670) );
  NAND2_X1 U6091 ( .A1(n5075), .A2(n5277), .ZN(n5311) );
  AND2_X1 U6092 ( .A1(n6009), .A2(n8442), .ZN(n4515) );
  NAND2_X1 U6093 ( .A1(n5689), .A2(n5688), .ZN(n10009) );
  NAND2_X1 U6094 ( .A1(n5857), .A2(n5856), .ZN(n9979) );
  AND2_X1 U6095 ( .A1(n8860), .A2(n8863), .ZN(n9217) );
  INV_X1 U6096 ( .A(n9217), .ZN(n4966) );
  AND2_X1 U6097 ( .A1(n8331), .A2(n8334), .ZN(n8466) );
  INV_X1 U6098 ( .A(n9363), .ZN(n9086) );
  NAND2_X1 U6099 ( .A1(n8492), .A2(n8491), .ZN(n9363) );
  AND2_X1 U6100 ( .A1(n9670), .A2(n5239), .ZN(n4516) );
  NAND2_X1 U6101 ( .A1(n8727), .A2(n8726), .ZN(n9354) );
  INV_X1 U6102 ( .A(n6994), .ZN(n5082) );
  AND2_X1 U6103 ( .A1(n8826), .A2(n8827), .ZN(n4517) );
  INV_X1 U6104 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5916) );
  INV_X1 U6105 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4712) );
  AND2_X1 U6106 ( .A1(n4702), .A2(n7302), .ZN(n4518) );
  AND2_X1 U6107 ( .A1(n5011), .A2(n6380), .ZN(n4519) );
  NOR2_X1 U6108 ( .A1(n9910), .A2(n9920), .ZN(n4520) );
  NOR2_X1 U6109 ( .A1(n9786), .A2(n9772), .ZN(n4521) );
  NOR2_X1 U6110 ( .A1(n9228), .A2(n9078), .ZN(n4522) );
  INV_X1 U6111 ( .A(n5032), .ZN(n5031) );
  AND2_X1 U6112 ( .A1(n5152), .A2(n5033), .ZN(n5032) );
  AND2_X1 U6113 ( .A1(n8507), .A2(n8506), .ZN(n4523) );
  AND2_X1 U6114 ( .A1(n9497), .A2(n10126), .ZN(n4524) );
  AND2_X1 U6115 ( .A1(n10003), .A2(n9883), .ZN(n4525) );
  AND2_X1 U6116 ( .A1(n5175), .A2(n5183), .ZN(n5232) );
  INV_X1 U6117 ( .A(n4728), .ZN(n4727) );
  NAND2_X1 U6118 ( .A1(n4730), .A2(n4729), .ZN(n4728) );
  NOR2_X1 U6119 ( .A1(n8010), .A2(n8939), .ZN(n4526) );
  INV_X1 U6120 ( .A(n4738), .ZN(n4737) );
  NAND2_X1 U6121 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  AND2_X1 U6122 ( .A1(n8791), .A2(n8805), .ZN(n8904) );
  INV_X1 U6123 ( .A(n8874), .ZN(n4788) );
  AND2_X1 U6124 ( .A1(n9088), .A2(n9099), .ZN(n4527) );
  INV_X1 U6125 ( .A(n4619), .ZN(n4618) );
  NAND2_X1 U6126 ( .A1(n8272), .A2(n8269), .ZN(n4619) );
  NAND4_X1 U6127 ( .A1(n8257), .A2(n8256), .A3(n8386), .A4(n8255), .ZN(n4528)
         );
  INV_X1 U6128 ( .A(n4577), .ZN(n4576) );
  OR2_X1 U6129 ( .A1(n5985), .A2(n4578), .ZN(n4577) );
  AND2_X1 U6130 ( .A1(n8754), .A2(n8752), .ZN(n9285) );
  NAND2_X1 U6131 ( .A1(n8744), .A2(n8747), .ZN(n9164) );
  AND2_X1 U6132 ( .A1(n10046), .A2(n9748), .ZN(n8483) );
  INV_X1 U6133 ( .A(n4703), .ZN(n4702) );
  OR2_X1 U6134 ( .A1(n5456), .A2(n4704), .ZN(n4703) );
  AND2_X1 U6135 ( .A1(n5842), .A2(n5816), .ZN(n4529) );
  INV_X1 U6136 ( .A(n4872), .ZN(n4871) );
  OR2_X1 U6137 ( .A1(n10025), .A2(n9906), .ZN(n8272) );
  NOR2_X1 U6138 ( .A1(n10140), .A2(n9662), .ZN(n4530) );
  NAND2_X1 U6139 ( .A1(n5150), .A2(n5029), .ZN(n4894) );
  OR2_X1 U6140 ( .A1(n8820), .A2(n8892), .ZN(n4797) );
  AND2_X1 U6141 ( .A1(n8079), .A2(n8081), .ZN(n4531) );
  AND2_X1 U6142 ( .A1(n5039), .A2(n5040), .ZN(n4532) );
  AND2_X1 U6143 ( .A1(n5016), .A2(n8519), .ZN(n4533) );
  AND2_X1 U6144 ( .A1(n4833), .A2(n4832), .ZN(n4534) );
  AND2_X1 U6145 ( .A1(n5234), .A2(n4712), .ZN(n4535) );
  NOR2_X1 U6146 ( .A1(n4865), .A2(n5612), .ZN(n4864) );
  AND2_X1 U6147 ( .A1(n4504), .A2(n8370), .ZN(n4536) );
  AND2_X1 U6148 ( .A1(n5346), .A2(n5345), .ZN(n4537) );
  AND2_X1 U6149 ( .A1(n4665), .A2(n4664), .ZN(n4538) );
  AND2_X1 U6151 ( .A1(n4993), .A2(n6120), .ZN(n4539) );
  AND2_X1 U6152 ( .A1(n6008), .A2(n4905), .ZN(n4540) );
  AND2_X1 U6153 ( .A1(n4702), .A2(n5080), .ZN(n4541) );
  AND2_X1 U6154 ( .A1(n5679), .A2(n5680), .ZN(n9587) );
  INV_X1 U6155 ( .A(n4926), .ZN(n4925) );
  NAND2_X1 U6156 ( .A1(n4929), .A2(n6012), .ZN(n4926) );
  AND4_X1 U6158 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n7374)
         );
  INV_X1 U6159 ( .A(n7374), .ZN(n4769) );
  AND4_X1 U6160 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(n7923)
         );
  INV_X1 U6161 ( .A(n7923), .ZN(n4771) );
  NAND2_X1 U6162 ( .A1(n6088), .A2(n6084), .ZN(n6086) );
  AND2_X1 U6163 ( .A1(n10122), .A2(n8161), .ZN(n4542) );
  NAND2_X1 U6164 ( .A1(n8729), .A2(n8728), .ZN(n9063) );
  INV_X1 U6165 ( .A(n9063), .ZN(n4979) );
  NAND2_X1 U6166 ( .A1(n5874), .A2(n5873), .ZN(n6028) );
  INV_X1 U6167 ( .A(n8391), .ZN(n4622) );
  INV_X1 U6168 ( .A(n8398), .ZN(n4907) );
  NAND2_X1 U6169 ( .A1(n4817), .A2(n4823), .ZN(n8504) );
  NAND2_X1 U6170 ( .A1(n10024), .A2(n5976), .ZN(n9902) );
  INV_X1 U6171 ( .A(n4570), .ZN(n10119) );
  INV_X1 U6172 ( .A(n5288), .ZN(n5353) );
  AND2_X1 U6173 ( .A1(n9910), .A2(n9920), .ZN(n4543) );
  INV_X1 U6174 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U6175 ( .A1(n6049), .A2(n6048), .ZN(n8338) );
  INV_X1 U6176 ( .A(n8338), .ZN(n4739) );
  OR2_X1 U6177 ( .A1(n9533), .A2(n9536), .ZN(n9534) );
  NAND2_X1 U6178 ( .A1(n5085), .A2(n5083), .ZN(n9552) );
  NAND2_X1 U6179 ( .A1(n5776), .A2(n5775), .ZN(n9659) );
  AND2_X1 U6180 ( .A1(n8338), .A2(n7979), .ZN(n4544) );
  NAND2_X1 U6181 ( .A1(n10122), .A2(n4727), .ZN(n4731) );
  AND2_X1 U6182 ( .A1(n8633), .A2(n8610), .ZN(n4545) );
  AND2_X1 U6183 ( .A1(n10304), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4546) );
  INV_X1 U6184 ( .A(n5008), .ZN(n5007) );
  AND2_X1 U6185 ( .A1(n9303), .A2(n5068), .ZN(n4547) );
  AND2_X1 U6186 ( .A1(n4961), .A2(n4962), .ZN(n4548) );
  INV_X1 U6187 ( .A(n4732), .ZN(n9856) );
  NOR2_X1 U6188 ( .A1(n9908), .A2(n4734), .ZN(n4732) );
  AND2_X1 U6189 ( .A1(n10030), .A2(n9919), .ZN(n4549) );
  AND2_X1 U6190 ( .A1(n5846), .A2(n5845), .ZN(n4550) );
  OR2_X1 U6191 ( .A1(n9086), .A2(n8717), .ZN(n4551) );
  INV_X1 U6192 ( .A(n10124), .ZN(n4606) );
  NAND2_X1 U6193 ( .A1(n5571), .A2(n5570), .ZN(n9962) );
  INV_X1 U6194 ( .A(n9962), .ZN(n4729) );
  INV_X1 U6195 ( .A(n7458), .ZN(n5919) );
  NAND2_X1 U6196 ( .A1(n7177), .A2(n4829), .ZN(n7185) );
  NAND2_X1 U6197 ( .A1(n7241), .A2(n4643), .ZN(n7314) );
  NAND2_X1 U6198 ( .A1(n6925), .A2(n5371), .ZN(n6993) );
  OAI21_X1 U6199 ( .B1(n5046), .B2(n5047), .A(n7114), .ZN(n7193) );
  NAND2_X1 U6200 ( .A1(n7984), .A2(n5502), .ZN(n7997) );
  INV_X1 U6201 ( .A(n6142), .ZN(n6119) );
  NAND2_X1 U6202 ( .A1(n7448), .A2(n10105), .ZN(n10139) );
  INV_X1 U6203 ( .A(n10139), .ZN(n4725) );
  OAI21_X1 U6204 ( .B1(n7231), .B2(n8904), .A(n7232), .ZN(n7235) );
  NAND2_X1 U6205 ( .A1(n5081), .A2(n5079), .ZN(n7299) );
  NAND2_X1 U6206 ( .A1(n5189), .A2(n5097), .ZN(n5915) );
  AND2_X1 U6207 ( .A1(n7275), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U6208 ( .A1(n7070), .A2(n4505), .ZN(n7398) );
  NAND2_X1 U6209 ( .A1(n4705), .A2(n7300), .ZN(n7386) );
  AND2_X1 U6210 ( .A1(n6045), .A2(n6044), .ZN(n4553) );
  AND2_X1 U6211 ( .A1(n6407), .A2(n6390), .ZN(n8133) );
  NAND2_X1 U6212 ( .A1(n5091), .A2(n5351), .ZN(n5352) );
  AND2_X1 U6213 ( .A1(n7370), .A2(n7369), .ZN(n4554) );
  AND2_X1 U6214 ( .A1(n6828), .A2(n5959), .ZN(n4555) );
  AND2_X1 U6215 ( .A1(n7313), .A2(n7312), .ZN(n4556) );
  AND2_X1 U6216 ( .A1(n4648), .A2(n8781), .ZN(n4557) );
  INV_X1 U6217 ( .A(n8328), .ZN(n4684) );
  INV_X1 U6218 ( .A(n10128), .ZN(n10152) );
  AND3_X1 U6219 ( .A1(n4651), .A2(n6153), .A3(n4512), .ZN(n6695) );
  INV_X1 U6220 ( .A(n6695), .ZN(n6788) );
  NAND2_X1 U6221 ( .A1(n4772), .A2(n6321), .ZN(n7924) );
  INV_X1 U6222 ( .A(n7924), .ZN(n4989) );
  INV_X1 U6223 ( .A(n7964), .ZN(n4991) );
  NAND2_X1 U6224 ( .A1(n6643), .A2(n5255), .ZN(n6650) );
  AND2_X1 U6225 ( .A1(n8741), .A2(n8740), .ZN(n4558) );
  AND2_X1 U6226 ( .A1(n5249), .A2(n4743), .ZN(n6641) );
  NAND2_X1 U6227 ( .A1(n5393), .A2(n5394), .ZN(n4559) );
  INV_X1 U6228 ( .A(n4981), .ZN(n4980) );
  NAND2_X1 U6229 ( .A1(n8737), .A2(n8763), .ZN(n4981) );
  NAND2_X1 U6230 ( .A1(n9728), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4560) );
  NOR2_X1 U6231 ( .A1(n4558), .A2(n8934), .ZN(n4561) );
  INV_X1 U6232 ( .A(n5210), .ZN(n10083) );
  AND2_X1 U6233 ( .A1(n9027), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4562) );
  OR2_X1 U6234 ( .A1(n8486), .A2(n6023), .ZN(n9926) );
  NOR2_X2 U6235 ( .A1(n6777), .A2(n8190), .ZN(n9963) );
  OAI211_X1 U6236 ( .C1(n4611), .C2(n5294), .A(n4609), .B(n5310), .ZN(n5124)
         );
  INV_X1 U6237 ( .A(n4676), .ZN(n8490) );
  NAND2_X1 U6238 ( .A1(n8774), .A2(n6688), .ZN(n6686) );
  NOR2_X2 U6239 ( .A1(n9270), .A2(n9277), .ZN(n9269) );
  NAND2_X1 U6240 ( .A1(n9126), .A2(n9087), .ZN(n9110) );
  NAND2_X1 U6241 ( .A1(n4854), .A2(n9745), .ZN(n4853) );
  NOR2_X1 U6242 ( .A1(n6608), .A2(n6443), .ZN(n10200) );
  NOR2_X1 U6243 ( .A1(n7485), .A2(n7486), .ZN(n9677) );
  NOR2_X1 U6244 ( .A1(n6873), .A2(n6874), .ZN(n7096) );
  AOI21_X1 U6245 ( .B1(n9712), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9711), .ZN(
        n9714) );
  AOI21_X1 U6246 ( .B1(n9728), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9722), .ZN(
        n9723) );
  AOI21_X1 U6247 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6628), .A(n6620), .ZN(
        n10224) );
  NAND2_X1 U6248 ( .A1(n6625), .A2(n6624), .ZN(n6702) );
  OAI21_X1 U6249 ( .B1(n9744), .B2(n10296), .A(n4855), .ZN(n4854) );
  NAND2_X1 U6250 ( .A1(n5951), .A2(n4566), .ZN(n6962) );
  OAI21_X1 U6251 ( .B1(n5992), .B2(n6784), .A(n4566), .ZN(n7215) );
  NAND2_X1 U6252 ( .A1(n10138), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U6253 ( .A1(n4583), .A2(n4582), .ZN(n5966) );
  NAND2_X1 U6254 ( .A1(n7070), .A2(n4584), .ZN(n4583) );
  OAI21_X1 U6255 ( .B1(n7070), .B2(n4586), .A(n4584), .ZN(n7447) );
  NAND2_X1 U6256 ( .A1(n5975), .A2(n4494), .ZN(n4589) );
  NAND2_X1 U6257 ( .A1(n4596), .A2(n5088), .ZN(n5181) );
  NAND3_X1 U6258 ( .A1(n4594), .A2(n4596), .A3(n4593), .ZN(n5208) );
  NOR2_X1 U6259 ( .A1(n6959), .A2(n9670), .ZN(n6844) );
  NAND2_X1 U6260 ( .A1(n10125), .A2(n4604), .ZN(n4603) );
  OAI21_X1 U6261 ( .B1(n10125), .B2(n4607), .A(n4604), .ZN(n8118) );
  NAND2_X1 U6262 ( .A1(n5118), .A2(n4608), .ZN(n4609) );
  NAND2_X1 U6263 ( .A1(n5118), .A2(n5117), .ZN(n5293) );
  NAND2_X1 U6264 ( .A1(n4610), .A2(n5121), .ZN(n5309) );
  INV_X1 U6265 ( .A(n5121), .ZN(n4611) );
  NAND2_X1 U6266 ( .A1(n4614), .A2(n4612), .ZN(P1_U3520) );
  AOI21_X1 U6267 ( .B1(n6013), .B2(n9784), .A(n4627), .ZN(n4626) );
  NAND2_X1 U6268 ( .A1(n9785), .A2(n6013), .ZN(n4628) );
  NAND2_X1 U6269 ( .A1(n9788), .A2(n6013), .ZN(n6052) );
  NAND2_X1 U6270 ( .A1(n6002), .A2(n4536), .ZN(n7941) );
  NAND2_X1 U6271 ( .A1(n7941), .A2(n8381), .ZN(n6003) );
  NAND2_X1 U6272 ( .A1(n9183), .A2(n4510), .ZN(n4637) );
  OR2_X1 U6273 ( .A1(n7241), .A2(n4642), .ZN(n4639) );
  NAND2_X1 U6274 ( .A1(n4639), .A2(n4640), .ZN(n7928) );
  NAND3_X1 U6275 ( .A1(n4646), .A2(n8759), .A3(n4645), .ZN(n7116) );
  NAND2_X1 U6276 ( .A1(n7115), .A2(n4647), .ZN(n4646) );
  NAND2_X1 U6277 ( .A1(n8768), .A2(n4649), .ZN(n7039) );
  NAND4_X1 U6278 ( .A1(n6688), .A2(n8775), .A3(n8776), .A4(n8765), .ZN(n7129)
         );
  NAND3_X1 U6279 ( .A1(n6688), .A2(n8776), .A3(n8765), .ZN(n4650) );
  NAND3_X1 U6280 ( .A1(n9357), .A2(n5095), .A3(n4652), .ZN(n9441) );
  AND3_X2 U6281 ( .A1(n6071), .A2(n4511), .A3(n6200), .ZN(n6088) );
  NAND4_X1 U6282 ( .A1(n6071), .A2(n4511), .A3(n4993), .A4(n6200), .ZN(n6148)
         );
  NAND2_X1 U6283 ( .A1(n4656), .A2(n4654), .ZN(n8227) );
  INV_X1 U6284 ( .A(n4655), .ZN(n4654) );
  OAI21_X1 U6285 ( .B1(n8224), .B2(n8364), .A(n8413), .ZN(n4655) );
  NAND2_X1 U6286 ( .A1(n8223), .A2(n8421), .ZN(n4656) );
  NAND2_X1 U6287 ( .A1(n8218), .A2(n4684), .ZN(n4657) );
  NAND2_X1 U6288 ( .A1(n4659), .A2(n4658), .ZN(n8277) );
  OR2_X1 U6289 ( .A1(n4662), .A2(n4661), .ZN(n4658) );
  AND2_X1 U6290 ( .A1(n4660), .A2(n8271), .ZN(n4659) );
  NAND3_X1 U6291 ( .A1(n8249), .A2(n4538), .A3(n8247), .ZN(n4660) );
  INV_X1 U6292 ( .A(n4665), .ZN(n4661) );
  AND2_X1 U6293 ( .A1(n4666), .A2(n4663), .ZN(n4662) );
  AND2_X2 U6294 ( .A1(n4674), .A2(n4673), .ZN(n7257) );
  INV_X1 U6295 ( .A(n4675), .ZN(n4674) );
  OAI21_X1 U6296 ( .B1(n5347), .B2(n6467), .A(n5260), .ZN(n4675) );
  NAND2_X1 U6297 ( .A1(n5997), .A2(n8360), .ZN(n8214) );
  NAND2_X1 U6298 ( .A1(n5092), .A2(n9543), .ZN(n4686) );
  OAI21_X1 U6299 ( .B1(n9542), .B2(n9543), .A(n4687), .ZN(n9544) );
  NAND3_X1 U6300 ( .A1(n4690), .A2(n9617), .A3(n4689), .ZN(n4688) );
  NAND2_X1 U6301 ( .A1(n4688), .A2(n9510), .ZN(n4691) );
  NAND2_X1 U6302 ( .A1(n5555), .A2(n4696), .ZN(n9635) );
  NAND2_X1 U6303 ( .A1(n5416), .A2(n4541), .ZN(n4700) );
  NAND3_X1 U6304 ( .A1(n4701), .A2(n4700), .A3(n4698), .ZN(n7514) );
  NAND2_X1 U6305 ( .A1(n7386), .A2(n5436), .ZN(n7472) );
  INV_X1 U6306 ( .A(n5436), .ZN(n4704) );
  NAND2_X1 U6307 ( .A1(n5785), .A2(n4491), .ZN(n4707) );
  NAND2_X1 U6308 ( .A1(n4707), .A2(n4708), .ZN(n9480) );
  NAND2_X1 U6309 ( .A1(n5785), .A2(n5784), .ZN(n9525) );
  NAND2_X2 U6310 ( .A1(n5237), .A2(n6909), .ZN(n6782) );
  INV_X1 U6311 ( .A(n4731), .ZN(n9960) );
  AND2_X1 U6312 ( .A1(n9800), .A2(n4737), .ZN(n9754) );
  NAND2_X1 U6313 ( .A1(n9800), .A2(n4736), .ZN(n9747) );
  NAND2_X1 U6314 ( .A1(n9800), .A2(n4740), .ZN(n6051) );
  NAND2_X1 U6315 ( .A1(n9800), .A2(n9783), .ZN(n9778) );
  NAND2_X1 U6316 ( .A1(n4741), .A2(n9596), .ZN(n5761) );
  NAND2_X1 U6317 ( .A1(n5089), .A2(n4741), .ZN(n9501) );
  INV_X2 U6318 ( .A(n4742), .ZN(n5885) );
  NAND2_X1 U6319 ( .A1(n4752), .A2(n6651), .ZN(n4748) );
  NAND2_X1 U6320 ( .A1(n6650), .A2(n6653), .ZN(n4752) );
  NAND4_X1 U6321 ( .A1(n4748), .A2(n4751), .A3(n4750), .A4(n5286), .ZN(n9606)
         );
  INV_X1 U6322 ( .A(n6653), .ZN(n4744) );
  INV_X1 U6323 ( .A(n6650), .ZN(n4745) );
  INV_X1 U6324 ( .A(n5284), .ZN(n4747) );
  NAND2_X1 U6325 ( .A1(n4749), .A2(n4752), .ZN(n9605) );
  NAND2_X1 U6326 ( .A1(n4750), .A2(n4753), .ZN(n4749) );
  AND2_X1 U6327 ( .A1(n4751), .A2(n5286), .ZN(n9604) );
  NAND2_X1 U6328 ( .A1(n4756), .A2(n4755), .ZN(n9487) );
  AND2_X1 U6329 ( .A1(n5189), .A2(n4759), .ZN(n5195) );
  NAND2_X1 U6330 ( .A1(n5189), .A2(n4760), .ZN(n5197) );
  NAND4_X1 U6331 ( .A1(n5170), .A2(n5169), .A3(n5171), .A4(n7778), .ZN(n4764)
         );
  INV_X1 U6332 ( .A(n5313), .ZN(n4763) );
  INV_X1 U6333 ( .A(n4764), .ZN(n4762) );
  NAND2_X1 U6334 ( .A1(n6495), .A2(n6262), .ZN(n4770) );
  NAND2_X1 U6335 ( .A1(n8872), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U6336 ( .A1(n4779), .A2(n4777), .ZN(n8881) );
  INV_X1 U6337 ( .A(n8873), .ZN(n4789) );
  INV_X1 U6338 ( .A(n8870), .ZN(n4790) );
  NAND2_X1 U6339 ( .A1(n4794), .A2(n4791), .ZN(n4796) );
  NAND3_X1 U6340 ( .A1(n8816), .A2(n8815), .A3(n4795), .ZN(n4794) );
  NAND2_X1 U6341 ( .A1(n8666), .A2(n4488), .ZN(n4805) );
  OAI21_X1 U6342 ( .B1(n8640), .B2(n4813), .A(n4812), .ZN(P2_U3216) );
  NAND2_X1 U6343 ( .A1(n8100), .A2(n4818), .ZN(n4815) );
  NAND2_X1 U6344 ( .A1(n4815), .A2(n4816), .ZN(n8653) );
  OR2_X1 U6345 ( .A1(n6951), .A2(n4828), .ZN(n4824) );
  NAND2_X1 U6346 ( .A1(n4824), .A2(n4825), .ZN(n7290) );
  NAND2_X1 U6347 ( .A1(n6074), .A2(n4833), .ZN(n6112) );
  NAND2_X1 U6348 ( .A1(n6074), .A2(n4534), .ZN(n4831) );
  NAND2_X1 U6349 ( .A1(n6936), .A2(n4834), .ZN(n6816) );
  NAND2_X1 U6350 ( .A1(n6816), .A2(n6280), .ZN(n6301) );
  NAND2_X1 U6351 ( .A1(n4836), .A2(n4835), .ZN(n6116) );
  NOR2_X2 U6352 ( .A1(n6142), .A2(n4837), .ZN(n10411) );
  NAND2_X1 U6353 ( .A1(n6685), .A2(n8926), .ZN(n6142) );
  INV_X1 U6354 ( .A(n4849), .ZN(n9707) );
  NAND2_X1 U6355 ( .A1(n9712), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4848) );
  NAND3_X1 U6356 ( .A1(n4856), .A2(n4853), .A3(n4852), .ZN(P1_U3260) );
  NAND2_X1 U6357 ( .A1(n8704), .A2(n8560), .ZN(n8572) );
  NOR2_X1 U6358 ( .A1(n9731), .A2(n9730), .ZN(n9739) );
  NOR2_X1 U6359 ( .A1(n9675), .A2(n9676), .ZN(n9688) );
  INV_X4 U6360 ( .A(n8204), .ZN(n6461) );
  NAND2_X1 U6361 ( .A1(n5140), .A2(n5139), .ZN(n5418) );
  XNOR2_X2 U6362 ( .A(n5278), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U6363 ( .A1(n4859), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U6364 ( .A1(n5562), .A2(n4864), .ZN(n4862) );
  NAND2_X1 U6365 ( .A1(n4862), .A2(n4863), .ZN(n5634) );
  NAND2_X1 U6366 ( .A1(n5764), .A2(n4877), .ZN(n4876) );
  NAND2_X1 U6367 ( .A1(n5764), .A2(n5763), .ZN(n4883) );
  NAND2_X1 U6368 ( .A1(n5870), .A2(n4890), .ZN(n4888) );
  NAND2_X1 U6369 ( .A1(n5870), .A2(n5869), .ZN(n4889) );
  NAND2_X1 U6370 ( .A1(n4897), .A2(n8328), .ZN(n4896) );
  AOI21_X1 U6371 ( .B1(n4899), .B2(n4684), .A(n8483), .ZN(n4898) );
  OAI21_X1 U6372 ( .B1(n8327), .B2(n8337), .A(n8435), .ZN(n4899) );
  NAND2_X1 U6373 ( .A1(n8330), .A2(n8329), .ZN(n4900) );
  MUX2_X1 U6374 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6461), .Z(n5128) );
  MUX2_X1 U6375 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6461), .Z(n5151) );
  MUX2_X1 U6376 ( .A(n6673), .B(n6671), .S(n6461), .Z(n5158) );
  MUX2_X1 U6377 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4903), .Z(n5162) );
  MUX2_X1 U6378 ( .A(n6752), .B(n6750), .S(n4903), .Z(n5165) );
  MUX2_X1 U6379 ( .A(n5563), .B(n6765), .S(n4903), .Z(n5565) );
  MUX2_X1 U6380 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4903), .Z(n5611) );
  MUX2_X1 U6381 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4903), .Z(n5635) );
  MUX2_X1 U6382 ( .A(n8510), .B(n7841), .S(n4903), .Z(n5639) );
  MUX2_X1 U6383 ( .A(n5659), .B(n7852), .S(n4903), .Z(n5661) );
  MUX2_X1 U6384 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4903), .Z(n5711) );
  MUX2_X1 U6385 ( .A(n5713), .B(n7802), .S(n4903), .Z(n5715) );
  MUX2_X1 U6386 ( .A(n5741), .B(n7816), .S(n4903), .Z(n5742) );
  MUX2_X1 U6387 ( .A(n5766), .B(n7936), .S(n4903), .Z(n5787) );
  MUX2_X1 U6388 ( .A(n5792), .B(n8151), .S(n4903), .Z(n5794) );
  MUX2_X1 U6389 ( .A(n5820), .B(n8096), .S(n4903), .Z(n5822) );
  NAND2_X1 U6390 ( .A1(n6007), .A2(n4906), .ZN(n4904) );
  NAND2_X1 U6391 ( .A1(n4904), .A2(n4540), .ZN(n9881) );
  NAND3_X1 U6392 ( .A1(n4916), .A2(n4917), .A3(n5107), .ZN(n5246) );
  NAND2_X1 U6393 ( .A1(n4918), .A2(n6828), .ZN(n7007) );
  OR2_X1 U6394 ( .A1(n9793), .A2(n4926), .ZN(n4922) );
  OR2_X1 U6395 ( .A1(n9793), .A2(n5989), .ZN(n4928) );
  NAND2_X1 U6396 ( .A1(n4922), .A2(n4923), .ZN(n6050) );
  NAND2_X1 U6397 ( .A1(n9793), .A2(n4932), .ZN(n4927) );
  NAND2_X1 U6398 ( .A1(n4936), .A2(n4934), .ZN(n5975) );
  NAND2_X1 U6399 ( .A1(n5970), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U6400 ( .A1(n4942), .A2(n4940), .ZN(n5982) );
  NAND2_X1 U6401 ( .A1(n4947), .A2(n4561), .ZN(n4946) );
  XNOR2_X1 U6402 ( .A(n8739), .B(n10369), .ZN(n4947) );
  NAND2_X1 U6403 ( .A1(n9306), .A2(n8837), .ZN(n9292) );
  NAND2_X1 U6404 ( .A1(n4974), .A2(n4975), .ZN(n8738) );
  NAND2_X1 U6405 ( .A1(n9094), .A2(n4976), .ZN(n4974) );
  NAND2_X1 U6406 ( .A1(n4983), .A2(n4982), .ZN(n8014) );
  AND2_X2 U6407 ( .A1(n6126), .A2(n6135), .ZN(n6174) );
  NAND2_X1 U6408 ( .A1(n6088), .A2(n4984), .ZN(n6123) );
  INV_X1 U6409 ( .A(n7378), .ZN(n4988) );
  INV_X1 U6410 ( .A(n4992), .ZN(n7930) );
  NAND2_X1 U6411 ( .A1(n6088), .A2(n4539), .ZN(n6150) );
  NAND2_X1 U6412 ( .A1(n6150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6145) );
  AND2_X1 U6413 ( .A1(n9151), .A2(n4999), .ZN(n9112) );
  NAND2_X1 U6414 ( .A1(n9151), .A2(n4997), .ZN(n9100) );
  NAND3_X1 U6415 ( .A1(n5000), .A2(n5001), .A3(n7138), .ZN(n7199) );
  NAND2_X1 U6416 ( .A1(n8080), .A2(n4531), .ZN(n8100) );
  NAND2_X1 U6417 ( .A1(n8653), .A2(n4533), .ZN(n5012) );
  NAND2_X1 U6418 ( .A1(n5012), .A2(n5013), .ZN(n8659) );
  NAND2_X1 U6419 ( .A1(n5362), .A2(n5133), .ZN(n5017) );
  INV_X1 U6420 ( .A(n5022), .ZN(n5020) );
  INV_X1 U6421 ( .A(n5025), .ZN(n5397) );
  OR2_X1 U6422 ( .A1(n5150), .A2(n5031), .ZN(n5026) );
  NAND2_X1 U6423 ( .A1(n5026), .A2(n5027), .ZN(n5507) );
  INV_X1 U6424 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6425 ( .A1(n5036), .A2(n5037), .ZN(n9073) );
  NAND2_X1 U6426 ( .A1(n7950), .A2(n4532), .ZN(n5036) );
  NAND3_X1 U6427 ( .A1(n5039), .A2(n5040), .A3(n5042), .ZN(n5038) );
  NOR2_X1 U6428 ( .A1(n7038), .A2(n5048), .ZN(n5046) );
  NAND2_X1 U6429 ( .A1(n5049), .A2(n5050), .ZN(n9090) );
  NAND2_X1 U6430 ( .A1(n9127), .A2(n5051), .ZN(n5049) );
  NAND2_X1 U6431 ( .A1(n9127), .A2(n9135), .ZN(n9126) );
  AOI21_X1 U6432 ( .B1(n9245), .B2(n5057), .A(n5055), .ZN(n5054) );
  AND2_X1 U6433 ( .A1(n9400), .A2(n9261), .ZN(n5063) );
  NAND2_X1 U6434 ( .A1(n9329), .A2(n5067), .ZN(n5064) );
  NAND2_X1 U6435 ( .A1(n5064), .A2(n5065), .ZN(n9270) );
  NAND2_X1 U6436 ( .A1(n6789), .A2(n6788), .ZN(n5071) );
  NAND2_X1 U6437 ( .A1(n5070), .A2(n6793), .ZN(n6794) );
  NAND3_X1 U6438 ( .A1(n5071), .A2(n6792), .A3(n7132), .ZN(n5070) );
  NAND2_X1 U6439 ( .A1(n6794), .A2(n8901), .ZN(n7037) );
  INV_X1 U6440 ( .A(n7235), .ZN(n7234) );
  NAND2_X1 U6441 ( .A1(n6147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U6442 ( .A1(n5076), .A2(n5077), .ZN(n5708) );
  NAND2_X1 U6443 ( .A1(n9586), .A2(n9585), .ZN(n5076) );
  NAND2_X1 U6444 ( .A1(n9533), .A2(n5585), .ZN(n5085) );
  NAND2_X1 U6445 ( .A1(n5478), .A2(n5087), .ZN(n7984) );
  NAND2_X1 U6446 ( .A1(n9501), .A2(n9502), .ZN(n5762) );
  NAND2_X1 U6447 ( .A1(n5332), .A2(n5331), .ZN(n5091) );
  NAND3_X1 U6448 ( .A1(n5332), .A2(n5331), .A3(n5093), .ZN(n5092) );
  INV_X1 U6449 ( .A(n5351), .ZN(n5093) );
  NAND2_X1 U6450 ( .A1(n5417), .A2(n7300), .ZN(n7388) );
  NAND2_X1 U6451 ( .A1(n7039), .A2(n8757), .ZN(n7115) );
  AND2_X2 U6452 ( .A1(n10083), .A2(n5211), .ZN(n5288) );
  NAND2_X1 U6453 ( .A1(n6918), .A2(n6257), .ZN(n6936) );
  INV_X1 U6454 ( .A(n6022), .ZN(n6037) );
  OAI21_X1 U6455 ( .B1(n6461), .B2(n5114), .A(n5113), .ZN(n5116) );
  NAND2_X1 U6456 ( .A1(n6461), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6457 ( .A1(n6904), .A2(n8449), .ZN(n6903) );
  NAND2_X1 U6458 ( .A1(n4484), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6459 ( .A1(n5208), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5206) );
  NOR2_X1 U6460 ( .A1(n9480), .A2(n9477), .ZN(n5923) );
  OR2_X1 U6461 ( .A1(n9238), .A2(n8625), .ZN(n5094) );
  INV_X1 U6462 ( .A(n8806), .ZN(n7233) );
  AND3_X1 U6463 ( .A1(n8091), .A2(n8090), .A3(n8089), .ZN(n9312) );
  NAND2_X1 U6464 ( .A1(n5145), .A2(n5144), .ZN(n5437) );
  OR2_X1 U6465 ( .A1(n9355), .A2(n10436), .ZN(n5095) );
  OR2_X1 U6466 ( .A1(n8585), .A2(n5104), .ZN(n5096) );
  AND2_X1 U6467 ( .A1(n5943), .A2(n5920), .ZN(n5098) );
  AND4_X1 U6468 ( .A1(n5097), .A2(n5176), .A3(n7909), .A4(n5916), .ZN(n5099)
         );
  AND2_X1 U6469 ( .A1(n9091), .A2(n9092), .ZN(n5101) );
  AND2_X1 U6470 ( .A1(n8605), .A2(n8604), .ZN(n9119) );
  AND2_X1 U6471 ( .A1(n6119), .A2(n6417), .ZN(n9437) );
  INV_X1 U6472 ( .A(n10042), .ZN(n6029) );
  AND2_X1 U6473 ( .A1(n5149), .A2(n5148), .ZN(n5102) );
  INV_X1 U6474 ( .A(n4481), .ZN(n9840) );
  INV_X1 U6475 ( .A(n9358), .ZN(n9088) );
  AND2_X1 U6476 ( .A1(n5144), .A2(n5143), .ZN(n5103) );
  AND2_X1 U6477 ( .A1(n8571), .A2(n8570), .ZN(n9081) );
  INV_X1 U6478 ( .A(n9081), .ZN(n9082) );
  INV_X1 U6479 ( .A(n6028), .ZN(n9772) );
  XOR2_X1 U6480 ( .A(n9380), .B(n8599), .Z(n5104) );
  OR2_X1 U6481 ( .A1(n8191), .A2(n8476), .ZN(n5105) );
  NAND2_X1 U6482 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  INV_X1 U6483 ( .A(n5374), .ZN(n5131) );
  INV_X1 U6484 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6084) );
  INV_X1 U6485 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6073) );
  INV_X1 U6486 ( .A(SI_10_), .ZN(n7828) );
  INV_X1 U6487 ( .A(n8564), .ZN(n6755) );
  INV_X1 U6488 ( .A(n6353), .ZN(n6131) );
  OR2_X1 U6489 ( .A1(n8172), .A2(n8171), .ZN(n8523) );
  INV_X1 U6490 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6120) );
  INV_X1 U6491 ( .A(n7389), .ZN(n5433) );
  INV_X1 U6492 ( .A(n5736), .ZN(n5731) );
  INV_X1 U6493 ( .A(n5722), .ZN(n5720) );
  NAND2_X1 U6494 ( .A1(n5684), .A2(n5683), .ZN(n5686) );
  INV_X1 U6495 ( .A(n6814), .ZN(n6279) );
  NAND2_X1 U6496 ( .A1(n6755), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8578) );
  XNOR2_X1 U6497 ( .A(n8599), .B(n6788), .ZN(n6170) );
  NAND2_X1 U6498 ( .A1(n6131), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6364) );
  INV_X1 U6499 ( .A(n8084), .ZN(n8081) );
  INV_X1 U6500 ( .A(n8599), .ZN(n6304) );
  OR2_X1 U6501 ( .A1(n7020), .A2(n7018), .ZN(n6413) );
  NAND2_X1 U6502 ( .A1(n9086), .A2(n9119), .ZN(n9087) );
  NAND2_X1 U6503 ( .A1(n6756), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U6504 ( .A1(n6754), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U6505 ( .A1(n6132), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6395) );
  OR2_X1 U6506 ( .A1(n6305), .A2(n7176), .ZN(n6322) );
  NAND2_X1 U6507 ( .A1(n6129), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U6508 ( .A1(n6127), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6269) );
  INV_X1 U6509 ( .A(n9143), .ZN(n9148) );
  INV_X1 U6510 ( .A(n9324), .ZN(n9423) );
  INV_X1 U6511 ( .A(n9626), .ZN(n5842) );
  OR2_X1 U6512 ( .A1(n5878), .A2(n5877), .ZN(n5925) );
  NAND2_X1 U6513 ( .A1(n5799), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U6514 ( .A1(n5720), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5748) );
  INV_X1 U6515 ( .A(n5596), .ZN(n5594) );
  NAND2_X1 U6516 ( .A1(n5216), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5486) );
  OR2_X1 U6517 ( .A1(n10102), .A2(n8473), .ZN(n6023) );
  NAND2_X1 U6518 ( .A1(n4481), .A2(n10059), .ZN(n9815) );
  NAND2_X1 U6519 ( .A1(n7458), .A2(n8190), .ZN(n8328) );
  NAND2_X1 U6520 ( .A1(n5634), .A2(n5633), .ZN(n5637) );
  NAND2_X1 U6521 ( .A1(n5165), .A2(n7799), .ZN(n5560) );
  INV_X1 U6522 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5106) );
  INV_X1 U6523 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U6524 ( .A1(n6757), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8613) );
  INV_X1 U6525 ( .A(n7027), .ZN(n7035) );
  XNOR2_X1 U6526 ( .A(n6170), .B(n6172), .ZN(n6884) );
  INV_X1 U6527 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U6528 ( .A1(n6362), .A2(n6361), .ZN(n7442) );
  INV_X1 U6529 ( .A(n6174), .ZN(n6220) );
  INV_X1 U6530 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7815) );
  INV_X1 U6531 ( .A(n10349), .ZN(n8134) );
  OAI21_X1 U6532 ( .B1(n9094), .B2(n9093), .A(n10365), .ZN(n9098) );
  XNOR2_X1 U6533 ( .A(n9363), .B(n9119), .ZN(n9135) );
  INV_X1 U6534 ( .A(n9383), .ZN(n9199) );
  NAND2_X1 U6535 ( .A1(n8757), .A2(n8780), .ZN(n8901) );
  INV_X1 U6536 ( .A(n9437), .ZN(n10434) );
  INV_X1 U6537 ( .A(n9655), .ZN(n9786) );
  AND2_X1 U6538 ( .A1(n5891), .A2(n5892), .ZN(n9477) );
  OR2_X1 U6539 ( .A1(n5667), .A2(n5666), .ZN(n5692) );
  NAND2_X1 U6540 ( .A1(n5213), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5382) );
  OR2_X1 U6541 ( .A1(n6644), .A2(n8486), .ZN(n5924) );
  AND2_X1 U6542 ( .A1(n5879), .A2(n5925), .ZN(n9769) );
  AND2_X1 U6543 ( .A1(n8272), .A2(n8275), .ZN(n9931) );
  OR2_X1 U6544 ( .A1(n6769), .A2(n6768), .ZN(n6777) );
  INV_X1 U6545 ( .A(n10313), .ZN(n10032) );
  OR2_X1 U6546 ( .A1(n5932), .A2(n8191), .ZN(n9957) );
  AND2_X1 U6547 ( .A1(n6015), .A2(n8482), .ZN(n10128) );
  OR2_X1 U6548 ( .A1(n8486), .A2(n6024), .ZN(n6025) );
  AND2_X1 U6549 ( .A1(n5849), .A2(n5824), .ZN(n5847) );
  INV_X1 U6550 ( .A(n6787), .ZN(n10393) );
  AND2_X1 U6551 ( .A1(n8674), .A2(n10360), .ZN(n8714) );
  AOI21_X1 U6552 ( .B1(n9113), .B2(n8556), .A(n8618), .ZN(n9099) );
  AND4_X1 U6553 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n8937)
         );
  AND2_X1 U6554 ( .A1(n6529), .A2(n6528), .ZN(n10349) );
  INV_X1 U6555 ( .A(n9048), .ZN(n10350) );
  INV_X1 U6556 ( .A(n9309), .ZN(n10360) );
  INV_X1 U6557 ( .A(n8827), .ZN(n9068) );
  INV_X1 U6558 ( .A(n9321), .ZN(n9347) );
  AND2_X1 U6559 ( .A1(n10370), .A2(n7022), .ZN(n9325) );
  INV_X1 U6560 ( .A(n10411), .ZN(n10436) );
  INV_X1 U6561 ( .A(n10440), .ZN(n10426) );
  AND2_X1 U6562 ( .A1(n7313), .A2(n7236), .ZN(n10423) );
  NAND2_X1 U6563 ( .A1(n9313), .A2(n10418), .ZN(n10440) );
  OR2_X1 U6564 ( .A1(n10381), .A2(n6094), .ZN(n7020) );
  XNOR2_X1 U6565 ( .A(n6078), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7921) );
  AND2_X1 U6566 ( .A1(n6320), .A2(n6333), .ZN(n7275) );
  NOR2_X1 U6567 ( .A1(n5924), .A2(n5933), .ZN(n9607) );
  OR2_X1 U6568 ( .A1(n9629), .A2(n5831), .ZN(n5836) );
  INV_X1 U6569 ( .A(n4484), .ZN(n5831) );
  AOI21_X1 U6570 ( .B1(n10215), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6439), .ZN(
        n6442) );
  AND2_X1 U6571 ( .A1(n6017), .A2(n5932), .ZN(n10149) );
  AND2_X1 U6572 ( .A1(n5914), .A2(n6483), .ZN(n6026) );
  INV_X1 U6573 ( .A(n10329), .ZN(n10031) );
  AND2_X1 U6574 ( .A1(n5902), .A2(n5901), .ZN(n6488) );
  XNOR2_X1 U6575 ( .A(n5110), .B(n5109), .ZN(n5257) );
  INV_X1 U6576 ( .A(n9056), .ZN(n10351) );
  OR2_X1 U6577 ( .A1(n6426), .A2(n9311), .ZN(n8711) );
  INV_X1 U6578 ( .A(n9119), .ZN(n9149) );
  INV_X1 U6579 ( .A(n8722), .ZN(n9206) );
  AND4_X1 U6580 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n9310)
         );
  INV_X1 U6581 ( .A(n10347), .ZN(n7286) );
  OR2_X1 U6582 ( .A1(n7200), .A2(n10436), .ZN(n9321) );
  INV_X1 U6583 ( .A(n10455), .ZN(n10453) );
  AND2_X1 U6584 ( .A1(n10432), .A2(n10431), .ZN(n10452) );
  NAND2_X1 U6585 ( .A1(n6723), .A2(n7020), .ZN(n10442) );
  INV_X1 U6586 ( .A(n9607), .ZN(n9651) );
  NAND2_X1 U6587 ( .A1(n5863), .A2(n5862), .ZN(n9656) );
  INV_X1 U6588 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10218) );
  INV_X1 U6589 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10230) );
  INV_X1 U6590 ( .A(n10344), .ZN(n10341) );
  INV_X1 U6591 ( .A(n10336), .ZN(n10334) );
  INV_X1 U6592 ( .A(n10311), .ZN(n10309) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7832) );
  INV_X1 U6594 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7775) );
  NOR2_X1 U6595 ( .A1(n10487), .A2(n10486), .ZN(n10485) );
  NOR2_X1 U6596 ( .A1(n10484), .A2(n10483), .ZN(n10482) );
  AND2_X1 U6597 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5107) );
  AND2_X1 U6598 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6599 ( .A1(n8204), .A2(n5108), .ZN(n6166) );
  NAND2_X1 U6600 ( .A1(n5246), .A2(n6166), .ZN(n5110) );
  INV_X1 U6601 ( .A(SI_1_), .ZN(n5109) );
  MUX2_X1 U6602 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6461), .Z(n5256) );
  NAND2_X1 U6603 ( .A1(n5257), .A2(n5256), .ZN(n5112) );
  NAND2_X1 U6604 ( .A1(n5110), .A2(SI_1_), .ZN(n5111) );
  NAND2_X1 U6605 ( .A1(n5112), .A2(n5111), .ZN(n5275) );
  INV_X1 U6606 ( .A(SI_2_), .ZN(n5115) );
  XNOR2_X1 U6607 ( .A(n5116), .B(n5115), .ZN(n5276) );
  NAND2_X1 U6608 ( .A1(n5275), .A2(n5276), .ZN(n5118) );
  NAND2_X1 U6609 ( .A1(n5116), .A2(SI_2_), .ZN(n5117) );
  MUX2_X1 U6610 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6461), .Z(n5120) );
  NAND2_X1 U6611 ( .A1(n5120), .A2(SI_3_), .ZN(n5121) );
  MUX2_X1 U6612 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6461), .Z(n5122) );
  NAND2_X1 U6613 ( .A1(n5122), .A2(SI_4_), .ZN(n5123) );
  MUX2_X1 U6614 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6461), .Z(n5125) );
  NAND2_X1 U6615 ( .A1(n5125), .A2(SI_5_), .ZN(n5126) );
  NAND2_X1 U6616 ( .A1(n5128), .A2(SI_6_), .ZN(n5372) );
  MUX2_X1 U6617 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6461), .Z(n5130) );
  NAND2_X1 U6618 ( .A1(n5130), .A2(SI_7_), .ZN(n5129) );
  AND2_X1 U6619 ( .A1(n5372), .A2(n5129), .ZN(n5133) );
  INV_X1 U6620 ( .A(n5129), .ZN(n5132) );
  INV_X1 U6621 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5134) );
  MUX2_X1 U6622 ( .A(n6490), .B(n5134), .S(n6461), .Z(n5136) );
  INV_X1 U6623 ( .A(SI_8_), .ZN(n5135) );
  INV_X1 U6624 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6625 ( .A1(n5137), .A2(SI_8_), .ZN(n5138) );
  MUX2_X1 U6626 ( .A(n6498), .B(n7855), .S(n6461), .Z(n5141) );
  INV_X1 U6627 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6628 ( .A1(n5142), .A2(SI_9_), .ZN(n5143) );
  NAND2_X1 U6629 ( .A1(n5418), .A2(n5103), .ZN(n5145) );
  MUX2_X1 U6630 ( .A(n6507), .B(n7775), .S(n6461), .Z(n5146) );
  INV_X1 U6631 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6632 ( .A1(n5147), .A2(SI_10_), .ZN(n5148) );
  NAND2_X1 U6633 ( .A1(n5151), .A2(SI_11_), .ZN(n5152) );
  INV_X1 U6634 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6518) );
  MUX2_X1 U6635 ( .A(n6518), .B(n7832), .S(n6461), .Z(n5155) );
  INV_X1 U6636 ( .A(SI_12_), .ZN(n5154) );
  INV_X1 U6637 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6638 ( .A1(n5156), .A2(SI_12_), .ZN(n5157) );
  INV_X1 U6639 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6673) );
  INV_X1 U6640 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U6641 ( .A1(n5158), .A2(n7622), .ZN(n5505) );
  INV_X1 U6642 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U6643 ( .A1(n5159), .A2(SI_13_), .ZN(n5504) );
  NAND2_X1 U6644 ( .A1(n5162), .A2(SI_14_), .ZN(n5163) );
  INV_X1 U6645 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6752) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6750) );
  INV_X1 U6647 ( .A(SI_15_), .ZN(n7799) );
  INV_X1 U6648 ( .A(n5165), .ZN(n5166) );
  NAND2_X1 U6649 ( .A1(n5166), .A2(SI_15_), .ZN(n5167) );
  XNOR2_X1 U6650 ( .A(n5562), .B(n5561), .ZN(n6749) );
  NOR2_X1 U6651 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5171) );
  NOR2_X1 U6652 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5170) );
  NOR2_X1 U6653 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5169) );
  NOR2_X1 U6654 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5174) );
  NOR2_X1 U6655 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5173) );
  NOR2_X1 U6656 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5172) );
  NOR2_X1 U6657 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5176) );
  NAND2_X1 U6658 ( .A1(n5181), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6659 ( .A1(n5179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5180) );
  NAND2_X2 U6660 ( .A1(n5932), .A2(n10207), .ZN(n5364) );
  NAND2_X1 U6661 ( .A1(n6749), .A2(n5363), .ZN(n5188) );
  INV_X1 U6662 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5184) );
  AND2_X1 U6663 ( .A1(n5183), .A2(n5184), .ZN(n5509) );
  INV_X1 U6664 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6665 ( .A1(n5509), .A2(n5185), .ZN(n5568) );
  NAND2_X1 U6666 ( .A1(n5568), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U6667 ( .A1(n5533), .A2(n5532), .ZN(n5535) );
  NAND2_X1 U6668 ( .A1(n5535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5186) );
  XNOR2_X1 U6669 ( .A(n5186), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U6670 ( .A1(n4482), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6433), .B2(
        n9694), .ZN(n5187) );
  INV_X1 U6671 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6672 ( .A1(n5192), .A2(n5191), .ZN(n5194) );
  NAND2_X1 U6673 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U6674 ( .A(n5190), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5898) );
  OR2_X1 U6675 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  NAND2_X1 U6676 ( .A1(n5194), .A2(n5193), .ZN(n5895) );
  NOR2_X1 U6677 ( .A1(n5895), .A2(n7938), .ZN(n5199) );
  INV_X1 U6678 ( .A(n5189), .ZN(n5200) );
  NAND2_X1 U6679 ( .A1(n5200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6680 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  NAND2_X1 U6681 ( .A1(n5202), .A2(n5201), .ZN(n5229) );
  NAND2_X1 U6682 ( .A1(n5204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5205) );
  AND2_X4 U6683 ( .A1(n5248), .A2(n6909), .ZN(n5251) );
  NAND2_X1 U6684 ( .A1(n9649), .A2(n5251), .ZN(n5228) );
  NAND2_X1 U6685 ( .A1(n4492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6686 ( .A1(n6509), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6687 ( .A1(n5287), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5224) );
  INV_X1 U6688 ( .A(n5334), .ZN(n5212) );
  INV_X1 U6689 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5485) );
  INV_X1 U6690 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5515) );
  INV_X1 U6691 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6692 ( .A1(n5541), .A2(n5219), .ZN(n5220) );
  AND2_X1 U6693 ( .A1(n5573), .A2(n5220), .ZN(n9641) );
  NAND2_X1 U6694 ( .A1(n4484), .A2(n9641), .ZN(n5223) );
  NAND2_X1 U6695 ( .A1(n4487), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5222) );
  NAND4_X1 U6696 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(n9660)
         );
  INV_X1 U6697 ( .A(n6909), .ZN(n5226) );
  NAND2_X1 U6698 ( .A1(n9660), .A2(n5265), .ZN(n5227) );
  NAND2_X1 U6699 ( .A1(n5228), .A2(n5227), .ZN(n5238) );
  INV_X1 U6700 ( .A(n5232), .ZN(n5233) );
  NAND2_X1 U6701 ( .A1(n5233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5235) );
  MUX2_X1 U6702 ( .A(n5235), .B(P1_IR_REG_31__SCAN_IN), .S(n5234), .Z(n5236)
         );
  NAND2_X1 U6703 ( .A1(n5236), .A2(n5204), .ZN(n9745) );
  NAND2_X1 U6704 ( .A1(n5919), .A2(n9745), .ZN(n5237) );
  XNOR2_X1 U6705 ( .A(n5238), .B(n5839), .ZN(n5556) );
  AND2_X1 U6706 ( .A1(n7298), .A2(n9745), .ZN(n6848) );
  NAND2_X1 U6707 ( .A1(n7458), .A2(n6848), .ZN(n5239) );
  NAND2_X1 U6708 ( .A1(n5287), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5242) );
  INV_X1 U6709 ( .A(SI_0_), .ZN(n5245) );
  INV_X1 U6710 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5244) );
  OAI21_X1 U6711 ( .B1(n8204), .B2(n5245), .A(n5244), .ZN(n5247) );
  AND2_X1 U6712 ( .A1(n5247), .A2(n5246), .ZN(n10101) );
  MUX2_X1 U6713 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10101), .S(n5364), .Z(n6851)
         );
  INV_X1 U6714 ( .A(n5248), .ZN(n5250) );
  AOI22_X1 U6715 ( .A1(n5265), .A2(n6851), .B1(n5250), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U6716 ( .A1(n5251), .A2(n6851), .B1(n5250), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6717 ( .A1(n5253), .A2(n5252), .ZN(n6642) );
  INV_X1 U6718 ( .A(n6642), .ZN(n5254) );
  NAND2_X1 U6719 ( .A1(n5254), .A2(n6782), .ZN(n5255) );
  XNOR2_X1 U6720 ( .A(n5257), .B(n5256), .ZN(n6467) );
  NAND2_X1 U6721 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5258) );
  INV_X1 U6722 ( .A(n6466), .ZN(n5259) );
  NAND2_X1 U6723 ( .A1(n5251), .A2(n5949), .ZN(n5267) );
  NAND2_X1 U6724 ( .A1(n4486), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6725 ( .A1(n5304), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6726 ( .A1(n5287), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6727 ( .A1(n5950), .A2(n5265), .ZN(n5266) );
  XNOR2_X1 U6728 ( .A(n5268), .B(n5839), .ZN(n6653) );
  NAND2_X1 U6729 ( .A1(n5885), .A2(n5950), .ZN(n5270) );
  NAND2_X1 U6730 ( .A1(n5265), .A2(n5949), .ZN(n5269) );
  NAND2_X1 U6731 ( .A1(n5270), .A2(n5269), .ZN(n6651) );
  NAND2_X1 U6732 ( .A1(n5302), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6733 ( .A1(n5287), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6734 ( .A1(n5288), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6735 ( .A1(n4484), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6736 ( .A1(n9669), .A2(n5265), .ZN(n5282) );
  XNOR2_X1 U6737 ( .A(n5275), .B(n5276), .ZN(n6463) );
  NAND2_X1 U6738 ( .A1(n4482), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6739 ( .A1(n6433), .A2(n10215), .ZN(n5279) );
  NAND2_X1 U6740 ( .A1(n5251), .A2(n9611), .ZN(n5281) );
  NAND2_X1 U6741 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  AOI22_X1 U6742 ( .A1(n5885), .A2(n9669), .B1(n5265), .B2(n9611), .ZN(n5284)
         );
  NAND2_X1 U6743 ( .A1(n9606), .A2(n5286), .ZN(n6805) );
  NAND2_X1 U6744 ( .A1(n5287), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6745 ( .A1(n5288), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6746 ( .A1(n5302), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5290) );
  INV_X1 U6747 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U6748 ( .A1(n4484), .A2(n6435), .ZN(n5289) );
  NAND2_X1 U6749 ( .A1(n9668), .A2(n5265), .ZN(n5300) );
  XNOR2_X1 U6750 ( .A(n5293), .B(n5294), .ZN(n6470) );
  NAND2_X1 U6751 ( .A1(n4482), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6752 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5295), .ZN(n5296) );
  XNOR2_X1 U6753 ( .A(n5296), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U6754 ( .A1(n6433), .A2(n6628), .ZN(n5297) );
  NAND2_X1 U6755 ( .A1(n5251), .A2(n6807), .ZN(n5299) );
  NAND2_X1 U6756 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U6757 ( .A1(n5288), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6758 ( .A1(n5302), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5307) );
  INV_X1 U6759 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U6760 ( .A1(n6435), .A2(n9576), .ZN(n5303) );
  AND2_X1 U6761 ( .A1(n5303), .A2(n5334), .ZN(n9580) );
  NAND2_X1 U6762 ( .A1(n4484), .A2(n9580), .ZN(n5306) );
  NAND2_X1 U6763 ( .A1(n5287), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6764 ( .A1(n5955), .A2(n5265), .ZN(n5318) );
  XNOR2_X1 U6765 ( .A(n5309), .B(n5310), .ZN(n6465) );
  NAND2_X1 U6766 ( .A1(n4483), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6767 ( .A1(n5311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5312) );
  MUX2_X1 U6768 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5312), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5314) );
  AND2_X1 U6769 ( .A1(n5314), .A2(n5313), .ZN(n10222) );
  NAND2_X1 U6770 ( .A1(n6433), .A2(n10222), .ZN(n5315) );
  NAND2_X1 U6771 ( .A1(n5251), .A2(n9575), .ZN(n5317) );
  INV_X1 U6772 ( .A(n5324), .ZN(n5321) );
  AOI22_X1 U6773 ( .A1(n5885), .A2(n5955), .B1(n5265), .B2(n9575), .ZN(n5323)
         );
  INV_X1 U6774 ( .A(n5323), .ZN(n5320) );
  NAND2_X1 U6775 ( .A1(n5321), .A2(n5320), .ZN(n5329) );
  AND2_X1 U6776 ( .A1(n6806), .A2(n5329), .ZN(n5322) );
  NAND2_X1 U6777 ( .A1(n6805), .A2(n5322), .ZN(n5332) );
  XNOR2_X1 U6778 ( .A(n5324), .B(n5323), .ZN(n9571) );
  INV_X1 U6779 ( .A(n9571), .ZN(n5328) );
  INV_X1 U6780 ( .A(n5325), .ZN(n5327) );
  NAND2_X1 U6781 ( .A1(n5327), .A2(n5326), .ZN(n9569) );
  NAND2_X1 U6782 ( .A1(n5328), .A2(n9569), .ZN(n5330) );
  NAND2_X1 U6783 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  NAND2_X1 U6784 ( .A1(n5287), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6785 ( .A1(n5302), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5338) );
  INV_X1 U6786 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6787 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  AND2_X1 U6788 ( .A1(n5354), .A2(n5335), .ZN(n9548) );
  NAND2_X1 U6789 ( .A1(n4484), .A2(n9548), .ZN(n5337) );
  NAND2_X1 U6790 ( .A1(n5288), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5336) );
  NAND4_X1 U6791 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n9667)
         );
  NAND2_X1 U6792 ( .A1(n9667), .A2(n5265), .ZN(n5349) );
  NAND2_X1 U6793 ( .A1(n4483), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6794 ( .A1(n5313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5342) );
  MUX2_X1 U6795 ( .A(n5342), .B(P1_IR_REG_31__SCAN_IN), .S(n7778), .Z(n5344)
         );
  INV_X1 U6796 ( .A(n5400), .ZN(n5343) );
  NAND2_X1 U6797 ( .A1(n6433), .A2(n6629), .ZN(n5345) );
  NAND2_X1 U6798 ( .A1(n5251), .A2(n9545), .ZN(n5348) );
  NAND2_X1 U6799 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  XNOR2_X1 U6800 ( .A(n5350), .B(n5839), .ZN(n5351) );
  AOI22_X1 U6801 ( .A1(n5885), .A2(n9667), .B1(n5265), .B2(n9545), .ZN(n9543)
         );
  NAND2_X1 U6802 ( .A1(n6509), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6803 ( .A1(n5287), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5358) );
  INV_X1 U6804 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U6805 ( .A1(n5354), .A2(n6929), .ZN(n5355) );
  AND2_X1 U6806 ( .A1(n5382), .A2(n5355), .ZN(n7009) );
  NAND2_X1 U6807 ( .A1(n4484), .A2(n7009), .ZN(n5357) );
  NAND2_X1 U6808 ( .A1(n5302), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5356) );
  NAND4_X1 U6809 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n9666)
         );
  NAND2_X1 U6810 ( .A1(n9666), .A2(n5265), .ZN(n5366) );
  OR2_X1 U6811 ( .A1(n5400), .A2(n5508), .ZN(n5360) );
  INV_X1 U6812 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5376) );
  XNOR2_X1 U6813 ( .A(n5360), .B(n5376), .ZN(n10253) );
  NAND2_X1 U6814 ( .A1(n5251), .A2(n7010), .ZN(n5365) );
  NAND2_X1 U6815 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  XNOR2_X1 U6816 ( .A(n5367), .B(n6782), .ZN(n5368) );
  AOI22_X1 U6817 ( .A1(n5885), .A2(n9666), .B1(n5265), .B2(n7010), .ZN(n5369)
         );
  XNOR2_X1 U6818 ( .A(n5368), .B(n5369), .ZN(n6927) );
  INV_X1 U6819 ( .A(n5368), .ZN(n5370) );
  NAND2_X1 U6820 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6821 ( .A1(n5373), .A2(n5372), .ZN(n5375) );
  XNOR2_X1 U6822 ( .A(n5375), .B(n5374), .ZN(n6478) );
  NAND2_X1 U6823 ( .A1(n6478), .A2(n5363), .ZN(n5380) );
  NAND2_X1 U6824 ( .A1(n5400), .A2(n5376), .ZN(n5377) );
  NAND2_X1 U6825 ( .A1(n5377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U6826 ( .A(n5378), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6712) );
  AOI22_X1 U6827 ( .A1(n4483), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6433), .B2(
        n6712), .ZN(n5379) );
  NAND2_X1 U6828 ( .A1(n5380), .A2(n5379), .ZN(n7075) );
  NAND2_X1 U6829 ( .A1(n7075), .A2(n5251), .ZN(n5389) );
  NAND2_X1 U6830 ( .A1(n6509), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6831 ( .A1(n5287), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5386) );
  INV_X1 U6832 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6833 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  AND2_X1 U6834 ( .A1(n5406), .A2(n5383), .ZN(n7076) );
  NAND2_X1 U6835 ( .A1(n4484), .A2(n7076), .ZN(n5385) );
  NAND2_X1 U6836 ( .A1(n5302), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5384) );
  NAND4_X1 U6837 ( .A1(n5387), .A2(n5386), .A3(n5385), .A4(n5384), .ZN(n9665)
         );
  NAND2_X1 U6838 ( .A1(n9665), .A2(n5265), .ZN(n5388) );
  NAND2_X1 U6839 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  XNOR2_X1 U6840 ( .A(n5390), .B(n5839), .ZN(n5393) );
  NAND2_X1 U6841 ( .A1(n5885), .A2(n9665), .ZN(n5392) );
  NAND2_X1 U6842 ( .A1(n7075), .A2(n5265), .ZN(n5391) );
  AND2_X1 U6843 ( .A1(n5392), .A2(n5391), .ZN(n5394) );
  INV_X1 U6844 ( .A(n5393), .ZN(n5396) );
  INV_X1 U6845 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U6846 ( .A1(n5396), .A2(n5395), .ZN(n6994) );
  XNOR2_X1 U6847 ( .A(n5397), .B(n5398), .ZN(n6486) );
  NAND2_X1 U6848 ( .A1(n6486), .A2(n5363), .ZN(n5405) );
  NOR2_X1 U6849 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5399) );
  NAND2_X1 U6850 ( .A1(n5400), .A2(n5399), .ZN(n5402) );
  NAND2_X1 U6851 ( .A1(n5402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5401) );
  MUX2_X1 U6852 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5401), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5403) );
  AOI22_X1 U6853 ( .A1(n4482), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6433), .B2(
        n10272), .ZN(n5404) );
  NAND2_X1 U6854 ( .A1(n5405), .A2(n5404), .ZN(n7426) );
  NAND2_X1 U6855 ( .A1(n6509), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6856 ( .A1(n5287), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6857 ( .A1(n5406), .A2(n7303), .ZN(n5407) );
  AND2_X1 U6858 ( .A1(n5423), .A2(n5407), .ZN(n7409) );
  NAND2_X1 U6859 ( .A1(n4484), .A2(n7409), .ZN(n5409) );
  NAND2_X1 U6860 ( .A1(n5302), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5408) );
  NAND4_X1 U6861 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n9664)
         );
  AOI22_X1 U6862 ( .A1(n7426), .A2(n5265), .B1(n5885), .B2(n9664), .ZN(n5415)
         );
  NAND2_X1 U6863 ( .A1(n7426), .A2(n5251), .ZN(n5413) );
  NAND2_X1 U6864 ( .A1(n9664), .A2(n5265), .ZN(n5412) );
  NAND2_X1 U6865 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  XNOR2_X1 U6866 ( .A(n5414), .B(n6782), .ZN(n7302) );
  XNOR2_X1 U6867 ( .A(n5418), .B(n5103), .ZN(n6495) );
  NAND2_X1 U6868 ( .A1(n6495), .A2(n5363), .ZN(n5421) );
  NAND2_X1 U6869 ( .A1(n5438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5419) );
  XNOR2_X1 U6870 ( .A(n5419), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U6871 ( .A1(n4482), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6433), .B2(
        n10290), .ZN(n5420) );
  NAND2_X1 U6872 ( .A1(n5421), .A2(n5420), .ZN(n7361) );
  NAND2_X1 U6873 ( .A1(n7361), .A2(n5251), .ZN(n5430) );
  INV_X1 U6874 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6875 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  AND2_X1 U6876 ( .A1(n5446), .A2(n5424), .ZN(n7394) );
  NAND2_X1 U6877 ( .A1(n4484), .A2(n7394), .ZN(n5428) );
  NAND2_X1 U6878 ( .A1(n5287), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6879 ( .A1(n5302), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6880 ( .A1(n6509), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5425) );
  NAND4_X1 U6881 ( .A1(n5428), .A2(n5427), .A3(n5426), .A4(n5425), .ZN(n9663)
         );
  NAND2_X1 U6882 ( .A1(n9663), .A2(n5265), .ZN(n5429) );
  NAND2_X1 U6883 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  XNOR2_X1 U6884 ( .A(n5431), .B(n5839), .ZN(n5435) );
  AND2_X1 U6885 ( .A1(n5885), .A2(n9663), .ZN(n5432) );
  AOI21_X1 U6886 ( .B1(n7361), .B2(n5265), .A(n5432), .ZN(n5434) );
  XNOR2_X1 U6887 ( .A(n5435), .B(n5434), .ZN(n7389) );
  NAND2_X1 U6888 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  NAND2_X1 U6889 ( .A1(n6506), .A2(n5363), .ZN(n5445) );
  NAND2_X1 U6890 ( .A1(n5440), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5443) );
  INV_X1 U6891 ( .A(n5440), .ZN(n5442) );
  INV_X1 U6892 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6893 ( .A1(n5442), .A2(n5441), .ZN(n5459) );
  AOI22_X1 U6894 ( .A1(n4483), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6433), .B2(
        n10304), .ZN(n5444) );
  NAND2_X1 U6895 ( .A1(n5445), .A2(n5444), .ZN(n7474) );
  NAND2_X1 U6896 ( .A1(n7474), .A2(n5251), .ZN(n5453) );
  NAND2_X1 U6897 ( .A1(n6509), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6898 ( .A1(n5287), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6899 ( .A1(n5446), .A2(n7473), .ZN(n5447) );
  AND2_X1 U6900 ( .A1(n5464), .A2(n5447), .ZN(n7475) );
  NAND2_X1 U6901 ( .A1(n4484), .A2(n7475), .ZN(n5449) );
  NAND2_X1 U6902 ( .A1(n5302), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5448) );
  NAND4_X1 U6903 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n10148)
         );
  NAND2_X1 U6904 ( .A1(n10148), .A2(n5265), .ZN(n5452) );
  NAND2_X1 U6905 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  XNOR2_X1 U6906 ( .A(n5454), .B(n5839), .ZN(n7469) );
  AND2_X1 U6907 ( .A1(n5885), .A2(n10148), .ZN(n5455) );
  AOI21_X1 U6908 ( .B1(n7474), .B2(n5265), .A(n5455), .ZN(n7470) );
  AND2_X1 U6909 ( .A1(n7469), .A2(n7470), .ZN(n5456) );
  NAND2_X1 U6910 ( .A1(n6499), .A2(n5363), .ZN(n5462) );
  NAND2_X1 U6911 ( .A1(n5459), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U6912 ( .A(n5460), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U6913 ( .A1(n4483), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6433), .B2(
        n6876), .ZN(n5461) );
  NAND2_X1 U6914 ( .A1(n10140), .A2(n5251), .ZN(n5471) );
  NAND2_X1 U6915 ( .A1(n5287), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6916 ( .A1(n5302), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5468) );
  INV_X1 U6917 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6918 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  AND2_X1 U6919 ( .A1(n5486), .A2(n5465), .ZN(n10156) );
  NAND2_X1 U6920 ( .A1(n4484), .A2(n10156), .ZN(n5467) );
  NAND2_X1 U6921 ( .A1(n6509), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5466) );
  NAND4_X1 U6922 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n9662)
         );
  NAND2_X1 U6923 ( .A1(n9662), .A2(n5265), .ZN(n5470) );
  NAND2_X1 U6924 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  XNOR2_X1 U6925 ( .A(n5472), .B(n6782), .ZN(n5476) );
  AND2_X1 U6926 ( .A1(n5885), .A2(n9662), .ZN(n5473) );
  AOI21_X1 U6927 ( .B1(n10140), .B2(n5265), .A(n5473), .ZN(n5474) );
  XNOR2_X1 U6928 ( .A(n5476), .B(n5474), .ZN(n7515) );
  NAND2_X1 U6929 ( .A1(n7514), .A2(n7515), .ZN(n5478) );
  INV_X1 U6930 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U6931 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  XNOR2_X1 U6932 ( .A(n5480), .B(n5479), .ZN(n6516) );
  NAND2_X1 U6933 ( .A1(n6516), .A2(n5363), .ZN(n5484) );
  NOR2_X1 U6934 ( .A1(n5183), .A2(n5508), .ZN(n5481) );
  MUX2_X1 U6935 ( .A(n5508), .B(n5481), .S(P1_IR_REG_12__SCAN_IN), .Z(n5482)
         );
  OR2_X1 U6936 ( .A1(n5482), .A2(n5509), .ZN(n7097) );
  INV_X1 U6937 ( .A(n7097), .ZN(n7101) );
  AOI22_X1 U6938 ( .A1(n4483), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6433), .B2(
        n7101), .ZN(n5483) );
  NAND2_X1 U6939 ( .A1(n7994), .A2(n5251), .ZN(n5493) );
  NAND2_X1 U6940 ( .A1(n6509), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6941 ( .A1(n5287), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6942 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  AND2_X1 U6943 ( .A1(n5516), .A2(n5487), .ZN(n7989) );
  NAND2_X1 U6944 ( .A1(n4484), .A2(n7989), .ZN(n5489) );
  NAND2_X1 U6945 ( .A1(n5302), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5488) );
  NAND4_X1 U6946 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n10150)
         );
  NAND2_X1 U6947 ( .A1(n10150), .A2(n5265), .ZN(n5492) );
  NAND2_X1 U6948 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  XNOR2_X1 U6949 ( .A(n5494), .B(n5839), .ZN(n5496) );
  AND2_X1 U6950 ( .A1(n5885), .A2(n10150), .ZN(n5495) );
  AOI21_X1 U6951 ( .B1(n7994), .B2(n5265), .A(n5495), .ZN(n5497) );
  NAND2_X1 U6952 ( .A1(n5496), .A2(n5497), .ZN(n5502) );
  INV_X1 U6953 ( .A(n5496), .ZN(n5499) );
  INV_X1 U6954 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U6955 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  NAND2_X1 U6956 ( .A1(n5502), .A2(n5500), .ZN(n7986) );
  INV_X1 U6957 ( .A(n7986), .ZN(n5501) );
  AND2_X1 U6958 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  NAND2_X1 U6959 ( .A1(n6670), .A2(n5363), .ZN(n5514) );
  NOR2_X1 U6960 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  MUX2_X1 U6961 ( .A(n5508), .B(n5510), .S(P1_IR_REG_13__SCAN_IN), .Z(n5512)
         );
  INV_X1 U6962 ( .A(n5568), .ZN(n5511) );
  OR2_X1 U6963 ( .A1(n5512), .A2(n5511), .ZN(n7484) );
  INV_X1 U6964 ( .A(n7484), .ZN(n7488) );
  AOI22_X1 U6965 ( .A1(n4482), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6433), .B2(
        n7488), .ZN(n5513) );
  NAND2_X1 U6966 ( .A1(n8250), .A2(n5251), .ZN(n5523) );
  NAND2_X1 U6967 ( .A1(n6509), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U6968 ( .A1(n5287), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6969 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  AND2_X1 U6970 ( .A1(n5539), .A2(n5517), .ZN(n10132) );
  NAND2_X1 U6971 ( .A1(n4484), .A2(n10132), .ZN(n5519) );
  NAND2_X1 U6972 ( .A1(n5302), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5518) );
  NAND4_X1 U6973 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n9661)
         );
  NAND2_X1 U6974 ( .A1(n9661), .A2(n5265), .ZN(n5522) );
  NAND2_X1 U6975 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  XNOR2_X1 U6976 ( .A(n5524), .B(n5839), .ZN(n5526) );
  AND2_X1 U6977 ( .A1(n5885), .A2(n9661), .ZN(n5525) );
  AOI21_X1 U6978 ( .B1(n8250), .B2(n5265), .A(n5525), .ZN(n5527) );
  AND2_X1 U6979 ( .A1(n5526), .A2(n5527), .ZN(n7998) );
  INV_X1 U6980 ( .A(n5526), .ZN(n5529) );
  INV_X1 U6981 ( .A(n5527), .ZN(n5528) );
  NAND2_X1 U6982 ( .A1(n5529), .A2(n5528), .ZN(n7999) );
  XNOR2_X1 U6983 ( .A(n5531), .B(n5530), .ZN(n6674) );
  NAND2_X1 U6984 ( .A1(n6674), .A2(n5363), .ZN(n5537) );
  OR2_X1 U6985 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  AND2_X1 U6986 ( .A1(n5535), .A2(n5534), .ZN(n9674) );
  AOI22_X1 U6987 ( .A1(n4482), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6433), .B2(
        n9674), .ZN(n5536) );
  NAND2_X1 U6988 ( .A1(n9497), .A2(n5251), .ZN(n5547) );
  NAND2_X1 U6989 ( .A1(n5287), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6990 ( .A1(n6509), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5544) );
  INV_X1 U6991 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6992 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AND2_X1 U6993 ( .A1(n5541), .A2(n5540), .ZN(n9492) );
  NAND2_X1 U6994 ( .A1(n4484), .A2(n9492), .ZN(n5543) );
  NAND2_X1 U6995 ( .A1(n4487), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5542) );
  NAND4_X1 U6996 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5542), .ZN(n10126)
         );
  NAND2_X1 U6997 ( .A1(n10126), .A2(n5265), .ZN(n5546) );
  NAND2_X1 U6998 ( .A1(n5547), .A2(n5546), .ZN(n5548) );
  XNOR2_X1 U6999 ( .A(n5548), .B(n5839), .ZN(n5550) );
  INV_X1 U7000 ( .A(n5550), .ZN(n5549) );
  NAND2_X1 U7001 ( .A1(n9497), .A2(n5265), .ZN(n5552) );
  NAND2_X1 U7002 ( .A1(n5885), .A2(n10126), .ZN(n5551) );
  NAND2_X1 U7003 ( .A1(n5552), .A2(n5551), .ZN(n9489) );
  NAND2_X1 U7004 ( .A1(n9487), .A2(n9489), .ZN(n5555) );
  NAND2_X1 U7005 ( .A1(n9649), .A2(n5265), .ZN(n5554) );
  NAND2_X1 U7006 ( .A1(n5885), .A2(n9660), .ZN(n5553) );
  NAND2_X1 U7007 ( .A1(n5554), .A2(n5553), .ZN(n9638) );
  NAND2_X1 U7008 ( .A1(n9635), .A2(n9638), .ZN(n5559) );
  NAND2_X1 U7009 ( .A1(n5555), .A2(n9486), .ZN(n5558) );
  INV_X1 U7010 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U7011 ( .A1(n5558), .A2(n5557), .ZN(n9636) );
  INV_X1 U7012 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5563) );
  INV_X1 U7013 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6765) );
  INV_X1 U7014 ( .A(SI_16_), .ZN(n5564) );
  NAND2_X1 U7015 ( .A1(n5565), .A2(n5564), .ZN(n5588) );
  INV_X1 U7016 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7017 ( .A1(n5566), .A2(SI_16_), .ZN(n5567) );
  XNOR2_X1 U7018 ( .A(n5587), .B(n5586), .ZN(n8065) );
  NAND2_X1 U7019 ( .A1(n8065), .A2(n5363), .ZN(n5571) );
  OR3_X1 U7020 ( .A1(n5568), .A2(P1_IR_REG_14__SCAN_IN), .A3(
        P1_IR_REG_15__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7021 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5569) );
  XNOR2_X1 U7022 ( .A(n5569), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U7023 ( .A1(n4483), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6433), .B2(
        n9712), .ZN(n5570) );
  NAND2_X1 U7024 ( .A1(n9962), .A2(n5251), .ZN(n5580) );
  NAND2_X1 U7025 ( .A1(n5287), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7026 ( .A1(n4487), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5577) );
  INV_X1 U7027 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7028 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  AND2_X1 U7029 ( .A1(n5596), .A2(n5574), .ZN(n9964) );
  NAND2_X1 U7030 ( .A1(n4484), .A2(n9964), .ZN(n5576) );
  NAND2_X1 U7031 ( .A1(n6509), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5575) );
  NAND4_X1 U7032 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n9944)
         );
  NAND2_X1 U7033 ( .A1(n9944), .A2(n5265), .ZN(n5579) );
  NAND2_X1 U7034 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  XNOR2_X1 U7035 ( .A(n5581), .B(n5839), .ZN(n5584) );
  AND2_X1 U7036 ( .A1(n5885), .A2(n9944), .ZN(n5582) );
  AOI21_X1 U7037 ( .B1(n9962), .B2(n5265), .A(n5582), .ZN(n5583) );
  XNOR2_X1 U7038 ( .A(n5584), .B(n5583), .ZN(n9536) );
  NAND2_X1 U7039 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  INV_X1 U7040 ( .A(SI_17_), .ZN(n7576) );
  XNOR2_X1 U7041 ( .A(n5611), .B(n7576), .ZN(n5610) );
  XNOR2_X1 U7042 ( .A(n5613), .B(n5610), .ZN(n8101) );
  NAND2_X1 U7043 ( .A1(n8101), .A2(n5363), .ZN(n5593) );
  OAI21_X1 U7044 ( .B1(n5589), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  INV_X1 U7045 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U7046 ( .A1(n5590), .A2(n7659), .ZN(n5614) );
  OR2_X1 U7047 ( .A1(n5590), .A2(n7659), .ZN(n5591) );
  AND2_X1 U7048 ( .A1(n5614), .A2(n5591), .ZN(n9728) );
  AOI22_X1 U7049 ( .A1(n4482), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6433), .B2(
        n9728), .ZN(n5592) );
  NAND2_X1 U7050 ( .A1(n10030), .A2(n5251), .ZN(n5603) );
  INV_X1 U7051 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7052 ( .A1(n5596), .A2(n5595), .ZN(n5597) );
  NAND2_X1 U7053 ( .A1(n5619), .A2(n5597), .ZN(n9556) );
  NAND2_X1 U7054 ( .A1(n5287), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7055 ( .A1(n4487), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5598) );
  AND2_X1 U7056 ( .A1(n5599), .A2(n5598), .ZN(n5601) );
  NAND2_X1 U7057 ( .A1(n6509), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5600) );
  OAI211_X1 U7058 ( .C1(n9556), .C2(n5831), .A(n5601), .B(n5600), .ZN(n9919)
         );
  NAND2_X1 U7059 ( .A1(n9919), .A2(n5265), .ZN(n5602) );
  NAND2_X1 U7060 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  XNOR2_X1 U7061 ( .A(n5604), .B(n6782), .ZN(n5606) );
  AND2_X1 U7062 ( .A1(n5885), .A2(n9919), .ZN(n5605) );
  AOI21_X1 U7063 ( .B1(n10030), .B2(n5265), .A(n5605), .ZN(n5607) );
  XNOR2_X1 U7064 ( .A(n5606), .B(n5607), .ZN(n9554) );
  INV_X1 U7065 ( .A(n5606), .ZN(n5608) );
  NAND2_X1 U7066 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  NAND2_X1 U7067 ( .A1(n9552), .A2(n5609), .ZN(n5628) );
  INV_X1 U7068 ( .A(n5610), .ZN(n5612) );
  XNOR2_X1 U7069 ( .A(n5635), .B(SI_18_), .ZN(n5632) );
  XNOR2_X1 U7070 ( .A(n5634), .B(n5632), .ZN(n8166) );
  NAND2_X1 U7071 ( .A1(n8166), .A2(n5363), .ZN(n5617) );
  NAND2_X1 U7072 ( .A1(n5614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U7073 ( .A(n5615), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9740) );
  AOI22_X1 U7074 ( .A1(n4483), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6433), .B2(
        n9740), .ZN(n5616) );
  NAND2_X1 U7075 ( .A1(n10025), .A2(n5251), .ZN(n5624) );
  INV_X1 U7076 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7077 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  NAND2_X1 U7078 ( .A1(n5646), .A2(n5620), .ZN(n9927) );
  AOI22_X1 U7079 ( .A1(n4487), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n5287), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7080 ( .A1(n6509), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7081 ( .C1(n9927), .C2(n5831), .A(n5622), .B(n5621), .ZN(n9945)
         );
  NAND2_X1 U7082 ( .A1(n9945), .A2(n5265), .ZN(n5623) );
  NAND2_X1 U7083 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  XNOR2_X1 U7084 ( .A(n5625), .B(n5839), .ZN(n5629) );
  NAND2_X1 U7085 ( .A1(n5628), .A2(n5629), .ZN(n9616) );
  NAND2_X1 U7086 ( .A1(n10025), .A2(n5265), .ZN(n5627) );
  NAND2_X1 U7087 ( .A1(n9945), .A2(n5885), .ZN(n5626) );
  NAND2_X1 U7088 ( .A1(n5627), .A2(n5626), .ZN(n9619) );
  INV_X1 U7089 ( .A(n5628), .ZN(n5631) );
  INV_X1 U7090 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7091 ( .A1(n5635), .A2(SI_18_), .ZN(n5636) );
  INV_X1 U7092 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8510) );
  INV_X1 U7093 ( .A(SI_19_), .ZN(n5638) );
  NAND2_X1 U7094 ( .A1(n5639), .A2(n5638), .ZN(n5656) );
  INV_X1 U7095 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7096 ( .A1(n5640), .A2(SI_19_), .ZN(n5641) );
  NAND2_X1 U7097 ( .A1(n5656), .A2(n5641), .ZN(n5657) );
  XNOR2_X1 U7098 ( .A(n5658), .B(n5657), .ZN(n8508) );
  NAND2_X1 U7099 ( .A1(n8508), .A2(n5363), .ZN(n5643) );
  INV_X1 U7100 ( .A(n9745), .ZN(n8190) );
  AOI22_X1 U7101 ( .A1(n4483), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8190), .B2(
        n6433), .ZN(n5642) );
  NAND2_X1 U7102 ( .A1(n9910), .A2(n5251), .ZN(n5651) );
  INV_X1 U7103 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10021) );
  INV_X1 U7104 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7105 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U7106 ( .A1(n5667), .A2(n5647), .ZN(n9911) );
  OR2_X1 U7107 ( .A1(n9911), .A2(n5831), .ZN(n5649) );
  AOI22_X1 U7108 ( .A1(n5302), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n5287), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U7109 ( .C1(n5353), .C2(n10021), .A(n5649), .B(n5648), .ZN(n9920)
         );
  NAND2_X1 U7110 ( .A1(n9920), .A2(n5265), .ZN(n5650) );
  NAND2_X1 U7111 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  XNOR2_X1 U7112 ( .A(n5652), .B(n6782), .ZN(n9509) );
  NAND2_X1 U7113 ( .A1(n9910), .A2(n5265), .ZN(n5654) );
  NAND2_X1 U7114 ( .A1(n9920), .A2(n5885), .ZN(n5653) );
  NAND2_X1 U7115 ( .A1(n5654), .A2(n5653), .ZN(n9510) );
  NAND2_X1 U7116 ( .A1(n9512), .A2(n9509), .ZN(n5655) );
  INV_X1 U7117 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5659) );
  INV_X1 U7118 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7852) );
  INV_X1 U7119 ( .A(SI_20_), .ZN(n5660) );
  NAND2_X1 U7120 ( .A1(n5661), .A2(n5660), .ZN(n5685) );
  INV_X1 U7121 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7122 ( .A1(n5662), .A2(SI_20_), .ZN(n5663) );
  XNOR2_X1 U7123 ( .A(n5684), .B(n5683), .ZN(n8520) );
  NAND2_X1 U7124 ( .A1(n8520), .A2(n5363), .ZN(n5665) );
  NAND2_X1 U7125 ( .A1(n4482), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7126 ( .A1(n9895), .A2(n5251), .ZN(n5675) );
  INV_X1 U7127 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7128 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  AND2_X1 U7129 ( .A1(n5692), .A2(n5668), .ZN(n9896) );
  NAND2_X1 U7130 ( .A1(n9896), .A2(n4484), .ZN(n5673) );
  INV_X1 U7131 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U7132 ( .A1(n5287), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7133 ( .A1(n6509), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5669) );
  OAI211_X1 U7134 ( .C1(n5928), .C2(n10064), .A(n5670), .B(n5669), .ZN(n5671)
         );
  INV_X1 U7135 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U7136 ( .A1(n5673), .A2(n5672), .ZN(n9882) );
  NAND2_X1 U7137 ( .A1(n9882), .A2(n5265), .ZN(n5674) );
  NAND2_X1 U7138 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  XNOR2_X1 U7139 ( .A(n5676), .B(n6782), .ZN(n5679) );
  NAND2_X1 U7140 ( .A1(n9895), .A2(n5265), .ZN(n5678) );
  NAND2_X1 U7141 ( .A1(n9882), .A2(n5885), .ZN(n5677) );
  NAND2_X1 U7142 ( .A1(n5678), .A2(n5677), .ZN(n5680) );
  INV_X1 U7143 ( .A(n5679), .ZN(n5682) );
  INV_X1 U7144 ( .A(n5680), .ZN(n5681) );
  NAND2_X1 U7145 ( .A1(n5682), .A2(n5681), .ZN(n9585) );
  INV_X1 U7146 ( .A(SI_21_), .ZN(n5687) );
  XNOR2_X1 U7147 ( .A(n5711), .B(n5687), .ZN(n5710) );
  XNOR2_X1 U7148 ( .A(n5709), .B(n5710), .ZN(n8533) );
  NAND2_X1 U7149 ( .A1(n8533), .A2(n5363), .ZN(n5689) );
  NAND2_X1 U7150 ( .A1(n4482), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7151 ( .A1(n10009), .A2(n5251), .ZN(n5701) );
  INV_X1 U7152 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7153 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U7154 ( .A1(n5722), .A2(n5693), .ZN(n9873) );
  OR2_X1 U7155 ( .A1(n9873), .A2(n5831), .ZN(n5699) );
  INV_X1 U7156 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7157 ( .A1(n5287), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7158 ( .A1(n6509), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5694) );
  OAI211_X1 U7159 ( .C1(n5928), .C2(n5696), .A(n5695), .B(n5694), .ZN(n5697)
         );
  INV_X1 U7160 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U7161 ( .A1(n5699), .A2(n5698), .ZN(n9864) );
  NAND2_X1 U7162 ( .A1(n9864), .A2(n5265), .ZN(n5700) );
  NAND2_X1 U7163 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  XNOR2_X1 U7164 ( .A(n5702), .B(n6782), .ZN(n5704) );
  AND2_X1 U7165 ( .A1(n9864), .A2(n5885), .ZN(n5703) );
  AOI21_X1 U7166 ( .B1(n10009), .B2(n5265), .A(n5703), .ZN(n5705) );
  XNOR2_X1 U7167 ( .A(n5704), .B(n5705), .ZN(n9519) );
  INV_X1 U7168 ( .A(n5704), .ZN(n5706) );
  NAND2_X1 U7169 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  NAND2_X1 U7170 ( .A1(n5708), .A2(n5707), .ZN(n5737) );
  INV_X1 U7171 ( .A(n5737), .ZN(n5732) );
  NAND2_X1 U7172 ( .A1(n5711), .A2(SI_21_), .ZN(n5712) );
  INV_X1 U7173 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5713) );
  INV_X1 U7174 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7802) );
  INV_X1 U7175 ( .A(SI_22_), .ZN(n5714) );
  NAND2_X1 U7176 ( .A1(n5715), .A2(n5714), .ZN(n5738) );
  INV_X1 U7177 ( .A(n5715), .ZN(n5716) );
  NAND2_X1 U7178 ( .A1(n5716), .A2(SI_22_), .ZN(n5717) );
  NAND2_X1 U7179 ( .A1(n5738), .A2(n5717), .ZN(n5739) );
  XNOR2_X1 U7180 ( .A(n5740), .B(n5739), .ZN(n8547) );
  NAND2_X1 U7181 ( .A1(n8547), .A2(n5363), .ZN(n5719) );
  NAND2_X1 U7182 ( .A1(n4483), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5718) );
  INV_X1 U7183 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7184 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  NAND2_X1 U7185 ( .A1(n5748), .A2(n5723), .ZN(n9858) );
  OR2_X1 U7186 ( .A1(n9858), .A2(n5831), .ZN(n5729) );
  INV_X1 U7187 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7188 ( .A1(n5288), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7189 ( .A1(n5287), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5724) );
  OAI211_X1 U7190 ( .C1(n5726), .C2(n5928), .A(n5725), .B(n5724), .ZN(n5727)
         );
  INV_X1 U7191 ( .A(n5727), .ZN(n5728) );
  NAND2_X1 U7192 ( .A1(n5729), .A2(n5728), .ZN(n9883) );
  AND2_X1 U7193 ( .A1(n9883), .A2(n5885), .ZN(n5730) );
  AOI21_X1 U7194 ( .B1(n10003), .B2(n5265), .A(n5730), .ZN(n5736) );
  NAND2_X1 U7195 ( .A1(n5732), .A2(n5731), .ZN(n9595) );
  NAND2_X1 U7196 ( .A1(n10003), .A2(n5251), .ZN(n5734) );
  NAND2_X1 U7197 ( .A1(n9883), .A2(n5265), .ZN(n5733) );
  NAND2_X1 U7198 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  XNOR2_X1 U7199 ( .A(n5735), .B(n5839), .ZN(n9597) );
  NAND2_X1 U7200 ( .A1(n5737), .A2(n5736), .ZN(n9596) );
  OAI21_X2 U7201 ( .B1(n5740), .B2(n5739), .A(n5738), .ZN(n5764) );
  INV_X1 U7202 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5741) );
  INV_X1 U7203 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7816) );
  INV_X1 U7204 ( .A(SI_23_), .ZN(n7645) );
  NAND2_X1 U7205 ( .A1(n5742), .A2(n7645), .ZN(n5765) );
  INV_X1 U7206 ( .A(n5742), .ZN(n5743) );
  NAND2_X1 U7207 ( .A1(n5743), .A2(SI_23_), .ZN(n5744) );
  NAND2_X1 U7208 ( .A1(n8561), .A2(n5363), .ZN(n5746) );
  NAND2_X1 U7209 ( .A1(n4482), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5745) );
  NAND2_X2 U7210 ( .A1(n5746), .A2(n5745), .ZN(n9998) );
  NAND2_X1 U7211 ( .A1(n9998), .A2(n5251), .ZN(n5757) );
  INV_X1 U7212 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7213 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  NAND2_X1 U7214 ( .A1(n5770), .A2(n5749), .ZN(n9841) );
  OR2_X1 U7215 ( .A1(n9841), .A2(n5831), .ZN(n5755) );
  INV_X1 U7216 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7217 ( .A1(n5287), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7218 ( .A1(n6509), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5750) );
  OAI211_X1 U7219 ( .C1(n5928), .C2(n5752), .A(n5751), .B(n5750), .ZN(n5753)
         );
  INV_X1 U7220 ( .A(n5753), .ZN(n5754) );
  NAND2_X1 U7221 ( .A1(n5755), .A2(n5754), .ZN(n9865) );
  NAND2_X1 U7222 ( .A1(n9865), .A2(n5265), .ZN(n5756) );
  NAND2_X1 U7223 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  XNOR2_X1 U7224 ( .A(n5758), .B(n5839), .ZN(n5760) );
  AND2_X1 U7225 ( .A1(n9865), .A2(n5885), .ZN(n5759) );
  NAND2_X1 U7226 ( .A1(n5761), .A2(n5760), .ZN(n9500) );
  NAND2_X1 U7227 ( .A1(n5762), .A2(n9500), .ZN(n9562) );
  INV_X1 U7228 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5766) );
  INV_X1 U7229 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7936) );
  XNOR2_X1 U7230 ( .A(n5787), .B(SI_24_), .ZN(n5786) );
  XNOR2_X1 U7231 ( .A(n5791), .B(n5786), .ZN(n8575) );
  NAND2_X1 U7232 ( .A1(n8575), .A2(n5363), .ZN(n5768) );
  NAND2_X1 U7233 ( .A1(n4483), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7234 ( .A1(n9832), .A2(n5251), .ZN(n5778) );
  INV_X1 U7235 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7236 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  AND2_X1 U7237 ( .A1(n5801), .A2(n5771), .ZN(n9833) );
  NAND2_X1 U7238 ( .A1(n9833), .A2(n4484), .ZN(n5776) );
  INV_X1 U7239 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10057) );
  NAND2_X1 U7240 ( .A1(n5287), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7241 ( .A1(n5288), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5772) );
  OAI211_X1 U7242 ( .C1(n10057), .C2(n5928), .A(n5773), .B(n5772), .ZN(n5774)
         );
  INV_X1 U7243 ( .A(n5774), .ZN(n5775) );
  NAND2_X1 U7244 ( .A1(n9659), .A2(n5265), .ZN(n5777) );
  NAND2_X1 U7245 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  XNOR2_X1 U7246 ( .A(n5779), .B(n6782), .ZN(n5781) );
  AND2_X1 U7247 ( .A1(n9659), .A2(n5885), .ZN(n5780) );
  AOI21_X1 U7248 ( .B1(n9832), .B2(n5265), .A(n5780), .ZN(n5782) );
  XNOR2_X1 U7249 ( .A(n5781), .B(n5782), .ZN(n9563) );
  NAND2_X1 U7250 ( .A1(n9562), .A2(n9563), .ZN(n5785) );
  INV_X1 U7251 ( .A(n5781), .ZN(n5783) );
  NAND2_X1 U7252 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  INV_X1 U7253 ( .A(n5786), .ZN(n5790) );
  INV_X1 U7254 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7255 ( .A1(n5788), .A2(SI_24_), .ZN(n5789) );
  INV_X1 U7256 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5792) );
  INV_X1 U7257 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8151) );
  INV_X1 U7258 ( .A(SI_25_), .ZN(n5793) );
  NAND2_X1 U7259 ( .A1(n5794), .A2(n5793), .ZN(n5817) );
  INV_X1 U7260 ( .A(n5794), .ZN(n5795) );
  NAND2_X1 U7261 ( .A1(n5795), .A2(SI_25_), .ZN(n5796) );
  NAND2_X1 U7262 ( .A1(n5817), .A2(n5796), .ZN(n5818) );
  NAND2_X1 U7263 ( .A1(n8586), .A2(n5363), .ZN(n5798) );
  NAND2_X1 U7264 ( .A1(n4482), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7265 ( .A1(n9990), .A2(n5251), .ZN(n5810) );
  INV_X1 U7266 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7267 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U7268 ( .A1(n5829), .A2(n5802), .ZN(n9527) );
  INV_X1 U7269 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7270 ( .A1(n5287), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7271 ( .A1(n5288), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5803) );
  OAI211_X1 U7272 ( .C1(n5805), .C2(n5928), .A(n5804), .B(n5803), .ZN(n5806)
         );
  INV_X1 U7273 ( .A(n5806), .ZN(n5807) );
  NAND2_X1 U7274 ( .A1(n5808), .A2(n5807), .ZN(n9658) );
  NAND2_X1 U7275 ( .A1(n9658), .A2(n5265), .ZN(n5809) );
  NAND2_X1 U7276 ( .A1(n5810), .A2(n5809), .ZN(n5811) );
  XNOR2_X1 U7277 ( .A(n5811), .B(n6782), .ZN(n5813) );
  AND2_X1 U7278 ( .A1(n9658), .A2(n5885), .ZN(n5812) );
  AOI21_X1 U7279 ( .B1(n9990), .B2(n5265), .A(n5812), .ZN(n5814) );
  XNOR2_X1 U7280 ( .A(n5813), .B(n5814), .ZN(n9526) );
  INV_X1 U7281 ( .A(n5813), .ZN(n5815) );
  NAND2_X1 U7282 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  INV_X1 U7283 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5820) );
  INV_X1 U7284 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8096) );
  INV_X1 U7285 ( .A(SI_26_), .ZN(n5821) );
  NAND2_X1 U7286 ( .A1(n5822), .A2(n5821), .ZN(n5849) );
  INV_X1 U7287 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U7288 ( .A1(n5823), .A2(SI_26_), .ZN(n5824) );
  NAND2_X1 U7289 ( .A1(n4482), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7290 ( .A1(n9801), .A2(n5251), .ZN(n5838) );
  INV_X1 U7291 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U7292 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  NAND2_X1 U7293 ( .A1(n5878), .A2(n5830), .ZN(n9629) );
  INV_X1 U7294 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U7295 ( .A1(n6509), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7296 ( .A1(n5287), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5832) );
  OAI211_X1 U7297 ( .C1(n10052), .C2(n5928), .A(n5833), .B(n5832), .ZN(n5834)
         );
  INV_X1 U7298 ( .A(n5834), .ZN(n5835) );
  NAND2_X1 U7299 ( .A1(n9657), .A2(n5265), .ZN(n5837) );
  NAND2_X1 U7300 ( .A1(n5838), .A2(n5837), .ZN(n5840) );
  XNOR2_X1 U7301 ( .A(n5840), .B(n5839), .ZN(n5843) );
  AND2_X1 U7302 ( .A1(n9657), .A2(n5885), .ZN(n5841) );
  AOI21_X1 U7303 ( .B1(n9801), .B2(n5265), .A(n5841), .ZN(n5844) );
  XNOR2_X1 U7304 ( .A(n5843), .B(n5844), .ZN(n9626) );
  INV_X1 U7305 ( .A(n5843), .ZN(n5846) );
  INV_X1 U7306 ( .A(n5844), .ZN(n5845) );
  NAND2_X1 U7307 ( .A1(n5848), .A2(n5847), .ZN(n5850) );
  INV_X1 U7308 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5851) );
  INV_X1 U7309 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U7310 ( .A(n5851), .B(n10099), .S(n6461), .Z(n5853) );
  INV_X1 U7311 ( .A(SI_27_), .ZN(n5852) );
  NAND2_X1 U7312 ( .A1(n5853), .A2(n5852), .ZN(n5871) );
  INV_X1 U7313 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7314 ( .A1(n5854), .A2(SI_27_), .ZN(n5855) );
  NAND2_X1 U7315 ( .A1(n10096), .A2(n5363), .ZN(n5857) );
  NAND2_X1 U7316 ( .A1(n4483), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7317 ( .A1(n9979), .A2(n5251), .ZN(n5865) );
  XNOR2_X1 U7318 ( .A(n5878), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U7319 ( .A1(n9781), .A2(n4484), .ZN(n5863) );
  INV_X1 U7320 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7321 ( .A1(n5287), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7322 ( .A1(n5288), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5858) );
  OAI211_X1 U7323 ( .C1(n5860), .C2(n5928), .A(n5859), .B(n5858), .ZN(n5861)
         );
  INV_X1 U7324 ( .A(n5861), .ZN(n5862) );
  NAND2_X1 U7325 ( .A1(n9656), .A2(n5265), .ZN(n5864) );
  NAND2_X1 U7326 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  XNOR2_X1 U7327 ( .A(n5866), .B(n6782), .ZN(n5891) );
  NAND2_X1 U7328 ( .A1(n9979), .A2(n5265), .ZN(n5868) );
  NAND2_X1 U7329 ( .A1(n9656), .A2(n5885), .ZN(n5867) );
  NAND2_X1 U7330 ( .A1(n5868), .A2(n5867), .ZN(n5892) );
  INV_X1 U7331 ( .A(n5923), .ZN(n5921) );
  MUX2_X1 U7332 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6461), .Z(n6043) );
  INV_X1 U7333 ( .A(SI_28_), .ZN(n6044) );
  XNOR2_X1 U7334 ( .A(n6043), .B(n6044), .ZN(n6041) );
  NAND2_X1 U7335 ( .A1(n10091), .A2(n5363), .ZN(n5874) );
  NAND2_X1 U7336 ( .A1(n4483), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7337 ( .A1(n6028), .A2(n5265), .ZN(n5887) );
  INV_X1 U7338 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5876) );
  INV_X1 U7339 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5875) );
  OAI21_X1 U7340 ( .B1(n5878), .B2(n5876), .A(n5875), .ZN(n5879) );
  NAND2_X1 U7341 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5877) );
  NAND2_X1 U7342 ( .A1(n9769), .A2(n4484), .ZN(n5884) );
  INV_X1 U7343 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7344 ( .A1(n5287), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7345 ( .A1(n5288), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5880) );
  OAI211_X1 U7346 ( .C1(n6036), .C2(n5928), .A(n5881), .B(n5880), .ZN(n5882)
         );
  INV_X1 U7347 ( .A(n5882), .ZN(n5883) );
  NAND2_X1 U7348 ( .A1(n5884), .A2(n5883), .ZN(n9655) );
  NAND2_X1 U7349 ( .A1(n9655), .A2(n5885), .ZN(n5886) );
  NAND2_X1 U7350 ( .A1(n5887), .A2(n5886), .ZN(n5888) );
  XNOR2_X1 U7351 ( .A(n5888), .B(n6782), .ZN(n5890) );
  AOI22_X1 U7352 ( .A1(n6028), .A2(n5251), .B1(n5265), .B2(n9655), .ZN(n5889)
         );
  XNOR2_X1 U7353 ( .A(n5890), .B(n5889), .ZN(n5922) );
  INV_X1 U7354 ( .A(n5922), .ZN(n5943) );
  INV_X1 U7355 ( .A(n5891), .ZN(n5894) );
  INV_X1 U7356 ( .A(n5892), .ZN(n5893) );
  NAND2_X1 U7357 ( .A1(n5894), .A2(n5893), .ZN(n9476) );
  NAND3_X1 U7358 ( .A1(n5895), .A2(P1_B_REG_SCAN_IN), .A3(n7938), .ZN(n5897)
         );
  OR2_X1 U7359 ( .A1(n7938), .A2(P1_B_REG_SCAN_IN), .ZN(n5896) );
  AND2_X1 U7360 ( .A1(n5897), .A2(n5896), .ZN(n5899) );
  INV_X1 U7361 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7362 ( .A1(n6482), .A2(n5900), .ZN(n5902) );
  INV_X1 U7363 ( .A(n5898), .ZN(n8098) );
  NAND2_X1 U7364 ( .A1(n8098), .A2(n5895), .ZN(n5901) );
  NOR4_X1 U7365 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5906) );
  NOR4_X1 U7366 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5905) );
  NOR4_X1 U7367 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5904) );
  NOR4_X1 U7368 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5903) );
  NAND4_X1 U7369 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n5912)
         );
  NOR2_X1 U7370 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n5910) );
  NOR4_X1 U7371 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5909) );
  NOR4_X1 U7372 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5908) );
  NOR4_X1 U7373 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5907) );
  NAND4_X1 U7374 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n5911)
         );
  NOR2_X1 U7375 ( .A1(n5912), .A2(n5911), .ZN(n6032) );
  NAND2_X1 U7376 ( .A1(n6032), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7377 ( .A1(n6482), .A2(n5913), .ZN(n5914) );
  NAND2_X1 U7378 ( .A1(n8098), .A2(n7938), .ZN(n6483) );
  NAND2_X1 U7379 ( .A1(n6488), .A2(n6026), .ZN(n6644) );
  NAND2_X1 U7380 ( .A1(n5915), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U7381 ( .A(n5917), .B(n5916), .ZN(n6431) );
  AND2_X1 U7382 ( .A1(n6431), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5918) );
  INV_X1 U7383 ( .A(n8473), .ZN(n7356) );
  NAND2_X1 U7384 ( .A1(n7458), .A2(n7356), .ZN(n6960) );
  NAND2_X1 U7385 ( .A1(n5919), .A2(n8473), .ZN(n8191) );
  NAND2_X1 U7386 ( .A1(n10329), .A2(n8191), .ZN(n5933) );
  AND2_X1 U7387 ( .A1(n9476), .A2(n9607), .ZN(n5920) );
  NAND2_X1 U7388 ( .A1(n5921), .A2(n5098), .ZN(n5948) );
  NAND3_X1 U7389 ( .A1(n5923), .A2(n5922), .A3(n9607), .ZN(n5947) );
  OR2_X1 U7390 ( .A1(n6960), .A2(n7298), .ZN(n6773) );
  INV_X1 U7391 ( .A(n5925), .ZN(n9761) );
  INV_X1 U7392 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7393 ( .A1(n5287), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7394 ( .A1(n5288), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5926) );
  OAI211_X1 U7395 ( .C1(n5928), .C2(n6062), .A(n5927), .B(n5926), .ZN(n5929)
         );
  AOI21_X1 U7396 ( .B1(n9761), .B2(n4484), .A(n5929), .ZN(n8337) );
  NOR2_X1 U7397 ( .A1(n6909), .A2(n8190), .ZN(n5930) );
  NAND2_X1 U7398 ( .A1(n5919), .A2(n5930), .ZN(n8485) );
  OR2_X1 U7399 ( .A1(n8486), .A2(n8485), .ZN(n5931) );
  OR2_X1 U7400 ( .A1(n6644), .A2(n5931), .ZN(n5940) );
  INV_X1 U7401 ( .A(n5932), .ZN(n10208) );
  INV_X1 U7402 ( .A(n5933), .ZN(n5935) );
  OR2_X1 U7403 ( .A1(n8191), .A2(n6848), .ZN(n6766) );
  NAND3_X1 U7404 ( .A1(n5248), .A2(n6431), .A3(n6766), .ZN(n5934) );
  AOI21_X1 U7405 ( .B1(n6644), .B2(n5935), .A(n5934), .ZN(n5936) );
  OR2_X1 U7406 ( .A1(n5936), .A2(P1_U3084), .ZN(n5939) );
  AND2_X1 U7407 ( .A1(n6773), .A2(n8485), .ZN(n5937) );
  NOR2_X1 U7408 ( .A1(n8486), .A2(n5937), .ZN(n5938) );
  NAND2_X1 U7409 ( .A1(n6644), .A2(n5938), .ZN(n6647) );
  NAND2_X1 U7410 ( .A1(n5939), .A2(n6647), .ZN(n9642) );
  AOI22_X1 U7411 ( .A1(n9769), .A2(n9642), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5942) );
  NOR2_X2 U7412 ( .A1(n5940), .A2(n5932), .ZN(n9609) );
  NAND2_X1 U7413 ( .A1(n9656), .A2(n9609), .ZN(n5941) );
  OAI211_X1 U7414 ( .C1(n8337), .C2(n9578), .A(n5942), .B(n5941), .ZN(n5945)
         );
  NOR3_X1 U7415 ( .A1(n5943), .A2(n9651), .A3(n9476), .ZN(n5944) );
  AOI211_X1 U7416 ( .C1(n9612), .C2(n6028), .A(n5945), .B(n5944), .ZN(n5946)
         );
  NAND3_X1 U7417 ( .A1(n5948), .A2(n5947), .A3(n5946), .ZN(P1_U3218) );
  NAND2_X1 U7418 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  INV_X1 U7419 ( .A(n6962), .ZN(n5952) );
  INV_X1 U7420 ( .A(n9611), .ZN(n7061) );
  NAND2_X1 U7421 ( .A1(n9669), .A2(n7061), .ZN(n8361) );
  NAND2_X1 U7422 ( .A1(n7149), .A2(n7061), .ZN(n5953) );
  NAND2_X1 U7423 ( .A1(n6964), .A2(n5953), .ZN(n7147) );
  NAND2_X1 U7424 ( .A1(n6965), .A2(n6807), .ZN(n8360) );
  NAND2_X1 U7425 ( .A1(n9668), .A2(n10312), .ZN(n8363) );
  NAND2_X1 U7426 ( .A1(n7147), .A2(n7146), .ZN(n7145) );
  NAND2_X1 U7427 ( .A1(n6965), .A2(n10312), .ZN(n5954) );
  NAND2_X1 U7428 ( .A1(n7145), .A2(n5954), .ZN(n6904) );
  INV_X1 U7429 ( .A(n5955), .ZN(n7148) );
  NAND2_X1 U7430 ( .A1(n7148), .A2(n9575), .ZN(n8222) );
  INV_X1 U7431 ( .A(n9575), .ZN(n6914) );
  NAND2_X1 U7432 ( .A1(n5955), .A2(n6914), .ZN(n8415) );
  NAND2_X1 U7433 ( .A1(n8222), .A2(n8415), .ZN(n8449) );
  NAND2_X1 U7434 ( .A1(n7148), .A2(n6914), .ZN(n5956) );
  INV_X1 U7435 ( .A(n9667), .ZN(n9577) );
  NAND2_X1 U7436 ( .A1(n9577), .A2(n9545), .ZN(n8420) );
  INV_X1 U7437 ( .A(n6826), .ZN(n5957) );
  NAND2_X1 U7438 ( .A1(n9667), .A2(n9545), .ZN(n5959) );
  INV_X1 U7439 ( .A(n9666), .ZN(n9546) );
  INV_X1 U7440 ( .A(n7010), .ZN(n7263) );
  NAND2_X1 U7441 ( .A1(n9666), .A2(n7263), .ZN(n8220) );
  NAND2_X1 U7442 ( .A1(n8421), .A2(n8220), .ZN(n8219) );
  NAND2_X1 U7443 ( .A1(n9546), .A2(n7263), .ZN(n5960) );
  INV_X1 U7444 ( .A(n7075), .ZN(n7220) );
  NAND2_X1 U7445 ( .A1(n7220), .A2(n9665), .ZN(n8225) );
  INV_X1 U7446 ( .A(n9665), .ZN(n6931) );
  NAND2_X1 U7447 ( .A1(n6931), .A2(n7075), .ZN(n8369) );
  NAND2_X1 U7448 ( .A1(n8225), .A2(n8369), .ZN(n7071) );
  NAND2_X1 U7449 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  NAND2_X1 U7450 ( .A1(n7220), .A2(n6931), .ZN(n5961) );
  INV_X1 U7451 ( .A(n9664), .ZN(n7069) );
  OR2_X1 U7452 ( .A1(n7069), .A2(n7426), .ZN(n8240) );
  NAND2_X1 U7453 ( .A1(n7426), .A2(n7069), .ZN(n8368) );
  INV_X1 U7454 ( .A(n8452), .ZN(n5962) );
  NAND2_X1 U7455 ( .A1(n7426), .A2(n9664), .ZN(n5963) );
  AND2_X1 U7456 ( .A1(n7361), .A2(n9663), .ZN(n5964) );
  INV_X1 U7457 ( .A(n10148), .ZN(n7391) );
  OR2_X1 U7458 ( .A1(n7474), .A2(n7391), .ZN(n8245) );
  NAND2_X1 U7459 ( .A1(n7474), .A2(n7391), .ZN(n8236) );
  NAND2_X1 U7460 ( .A1(n8245), .A2(n8236), .ZN(n8456) );
  OR2_X1 U7461 ( .A1(n7474), .A2(n10148), .ZN(n5965) );
  NAND2_X1 U7462 ( .A1(n5966), .A2(n5965), .ZN(n10138) );
  NAND2_X1 U7463 ( .A1(n10140), .A2(n9662), .ZN(n5967) );
  INV_X1 U7464 ( .A(n10150), .ZN(n8006) );
  OR2_X1 U7465 ( .A1(n7994), .A2(n8006), .ZN(n8254) );
  NAND2_X1 U7466 ( .A1(n7994), .A2(n8006), .ZN(n8379) );
  NAND2_X1 U7467 ( .A1(n8254), .A2(n8379), .ZN(n8458) );
  OR2_X1 U7468 ( .A1(n8250), .A2(n9661), .ZN(n5968) );
  NAND2_X1 U7469 ( .A1(n8250), .A2(n9661), .ZN(n5969) );
  OR2_X1 U7470 ( .A1(n9497), .A2(n10126), .ZN(n5971) );
  NOR2_X1 U7471 ( .A1(n9649), .A2(n9660), .ZN(n5972) );
  INV_X1 U7472 ( .A(n9660), .ZN(n9956) );
  INV_X1 U7473 ( .A(n9649), .ZN(n10165) );
  INV_X1 U7474 ( .A(n9944), .ZN(n9558) );
  OR2_X1 U7475 ( .A1(n9962), .A2(n9558), .ZN(n8265) );
  NAND2_X1 U7476 ( .A1(n9962), .A2(n9558), .ZN(n8391) );
  NAND2_X1 U7477 ( .A1(n8265), .A2(n8391), .ZN(n9954) );
  NAND2_X1 U7478 ( .A1(n9962), .A2(n9944), .ZN(n5973) );
  OR2_X1 U7479 ( .A1(n10030), .A2(n9919), .ZN(n5974) );
  INV_X1 U7480 ( .A(n9945), .ZN(n9906) );
  NAND2_X1 U7481 ( .A1(n10025), .A2(n9906), .ZN(n8275) );
  NAND2_X1 U7482 ( .A1(n10025), .A2(n9945), .ZN(n5976) );
  OR2_X1 U7483 ( .A1(n9895), .A2(n9882), .ZN(n5977) );
  NAND2_X1 U7484 ( .A1(n9888), .A2(n5977), .ZN(n5979) );
  NAND2_X1 U7485 ( .A1(n9895), .A2(n9882), .ZN(n5978) );
  NAND2_X1 U7486 ( .A1(n5979), .A2(n5978), .ZN(n9870) );
  INV_X1 U7487 ( .A(n9864), .ZN(n9892) );
  OR2_X1 U7488 ( .A1(n10009), .A2(n9892), .ZN(n8280) );
  NAND2_X1 U7489 ( .A1(n10009), .A2(n9892), .ZN(n8285) );
  NAND2_X1 U7490 ( .A1(n8280), .A2(n8285), .ZN(n9877) );
  NAND2_X1 U7491 ( .A1(n10009), .A2(n9864), .ZN(n5980) );
  OR2_X1 U7492 ( .A1(n10003), .A2(n9883), .ZN(n5981) );
  NOR2_X1 U7493 ( .A1(n9998), .A2(n9865), .ZN(n5984) );
  NAND2_X1 U7494 ( .A1(n9998), .A2(n9865), .ZN(n5983) );
  AND2_X1 U7495 ( .A1(n9832), .A2(n9659), .ZN(n5985) );
  NAND2_X1 U7496 ( .A1(n9990), .A2(n9828), .ZN(n8302) );
  NAND2_X1 U7497 ( .A1(n9794), .A2(n8302), .ZN(n9809) );
  OR2_X1 U7498 ( .A1(n9990), .A2(n9658), .ZN(n5986) );
  NAND2_X1 U7499 ( .A1(n5987), .A2(n5986), .ZN(n9793) );
  NOR2_X1 U7500 ( .A1(n9801), .A2(n9657), .ZN(n5989) );
  NAND2_X1 U7501 ( .A1(n9801), .A2(n9657), .ZN(n5988) );
  NAND2_X1 U7502 ( .A1(n9979), .A2(n9799), .ZN(n8333) );
  NAND2_X1 U7503 ( .A1(n6028), .A2(n9786), .ZN(n8334) );
  NAND2_X1 U7504 ( .A1(n5990), .A2(n8466), .ZN(n5991) );
  NAND2_X1 U7505 ( .A1(n6040), .A2(n5991), .ZN(n9776) );
  NAND3_X1 U7506 ( .A1(n8485), .A2(n9745), .A3(n6782), .ZN(n10153) );
  NAND2_X1 U7507 ( .A1(n10153), .A2(n10102), .ZN(n10332) );
  INV_X1 U7508 ( .A(n10332), .ZN(n10036) );
  INV_X1 U7509 ( .A(n5992), .ZN(n6771) );
  INV_X1 U7510 ( .A(n6851), .ZN(n6959) );
  NAND2_X1 U7511 ( .A1(n6771), .A2(n6844), .ZN(n6770) );
  INV_X1 U7512 ( .A(n5950), .ZN(n8357) );
  NAND2_X1 U7513 ( .A1(n8357), .A2(n5949), .ZN(n5993) );
  NAND2_X1 U7514 ( .A1(n6770), .A2(n5993), .ZN(n6966) );
  NAND2_X1 U7515 ( .A1(n6966), .A2(n8446), .ZN(n5996) );
  NAND2_X1 U7516 ( .A1(n5996), .A2(n5995), .ZN(n7144) );
  INV_X1 U7517 ( .A(n7146), .ZN(n8447) );
  INV_X1 U7518 ( .A(n8222), .ZN(n8417) );
  NAND2_X1 U7519 ( .A1(n8213), .A2(n8415), .ZN(n6822) );
  AND2_X1 U7520 ( .A1(n8421), .A2(n8420), .ZN(n6000) );
  INV_X1 U7521 ( .A(n8416), .ZN(n5998) );
  NAND2_X1 U7522 ( .A1(n8421), .A2(n5998), .ZN(n8413) );
  NAND2_X1 U7523 ( .A1(n8413), .A2(n8220), .ZN(n5999) );
  INV_X1 U7524 ( .A(n7071), .ZN(n8451) );
  INV_X1 U7525 ( .A(n8369), .ZN(n8221) );
  AOI21_X1 U7526 ( .B1(n7067), .B2(n8451), .A(n8221), .ZN(n7401) );
  NAND2_X1 U7527 ( .A1(n7401), .A2(n8368), .ZN(n7357) );
  INV_X1 U7528 ( .A(n9663), .ZN(n7305) );
  OR2_X1 U7529 ( .A1(n7361), .A2(n7305), .ZN(n8244) );
  AND2_X1 U7530 ( .A1(n8244), .A2(n8240), .ZN(n8231) );
  NAND2_X1 U7531 ( .A1(n7357), .A2(n8231), .ZN(n6001) );
  NAND2_X1 U7532 ( .A1(n7361), .A2(n7305), .ZN(n8242) );
  NAND2_X1 U7533 ( .A1(n6001), .A2(n8242), .ZN(n7451) );
  INV_X1 U7534 ( .A(n8456), .ZN(n7450) );
  NAND2_X1 U7535 ( .A1(n7451), .A2(n7450), .ZN(n6002) );
  NAND2_X1 U7536 ( .A1(n8236), .A2(n8242), .ZN(n8232) );
  NAND2_X1 U7537 ( .A1(n8232), .A2(n8245), .ZN(n8370) );
  INV_X1 U7538 ( .A(n9662), .ZN(n7992) );
  OR2_X1 U7539 ( .A1(n10140), .A2(n7992), .ZN(n7940) );
  AND2_X1 U7540 ( .A1(n8254), .A2(n7940), .ZN(n8381) );
  NAND2_X1 U7541 ( .A1(n6003), .A2(n8379), .ZN(n10125) );
  XNOR2_X1 U7542 ( .A(n8250), .B(n9661), .ZN(n10124) );
  INV_X1 U7543 ( .A(n9661), .ZN(n9495) );
  NAND2_X1 U7544 ( .A1(n8250), .A2(n9495), .ZN(n8238) );
  INV_X1 U7545 ( .A(n10126), .ZN(n9645) );
  NAND2_X1 U7546 ( .A1(n9497), .A2(n9645), .ZN(n8258) );
  NAND2_X1 U7547 ( .A1(n8386), .A2(n8258), .ZN(n8033) );
  NAND2_X1 U7548 ( .A1(n9649), .A2(n9956), .ZN(n8389) );
  OR2_X1 U7549 ( .A1(n9649), .A2(n9956), .ZN(n9951) );
  AND2_X1 U7550 ( .A1(n8265), .A2(n9951), .ZN(n8394) );
  NAND2_X1 U7551 ( .A1(n9952), .A2(n8394), .ZN(n6006) );
  INV_X1 U7552 ( .A(n9919), .ZN(n9958) );
  AND2_X1 U7553 ( .A1(n10030), .A2(n9958), .ZN(n8264) );
  OR2_X1 U7554 ( .A1(n10030), .A2(n9958), .ZN(n8269) );
  INV_X1 U7555 ( .A(n9920), .ZN(n9893) );
  OR2_X1 U7556 ( .A1(n9910), .A2(n9893), .ZN(n8276) );
  NAND2_X1 U7557 ( .A1(n9910), .A2(n9893), .ZN(n8398) );
  NAND2_X1 U7558 ( .A1(n9904), .A2(n9903), .ZN(n6007) );
  INV_X1 U7559 ( .A(n9882), .ZN(n9907) );
  OR2_X1 U7560 ( .A1(n9895), .A2(n9907), .ZN(n8284) );
  NAND2_X1 U7561 ( .A1(n9895), .A2(n9907), .ZN(n9878) );
  INV_X1 U7562 ( .A(n9877), .ZN(n6008) );
  NAND2_X1 U7563 ( .A1(n9881), .A2(n8285), .ZN(n9863) );
  INV_X1 U7564 ( .A(n9883), .ZN(n9847) );
  OR2_X1 U7565 ( .A1(n10003), .A2(n9847), .ZN(n8443) );
  NAND2_X1 U7566 ( .A1(n10003), .A2(n9847), .ZN(n8442) );
  INV_X1 U7567 ( .A(n9865), .ZN(n9829) );
  NAND2_X1 U7568 ( .A1(n9998), .A2(n9829), .ZN(n8291) );
  NAND2_X1 U7569 ( .A1(n8295), .A2(n8291), .ZN(n9845) );
  INV_X1 U7570 ( .A(n9845), .ZN(n6009) );
  XNOR2_X1 U7571 ( .A(n9832), .B(n9848), .ZN(n9826) );
  NAND2_X1 U7572 ( .A1(n9832), .A2(n9848), .ZN(n8297) );
  INV_X1 U7573 ( .A(n8302), .ZN(n8309) );
  NAND2_X1 U7574 ( .A1(n9801), .A2(n9794), .ZN(n8308) );
  NAND2_X1 U7575 ( .A1(n9794), .A2(n9812), .ZN(n8304) );
  NAND2_X1 U7576 ( .A1(n8308), .A2(n8304), .ZN(n8353) );
  NAND2_X1 U7577 ( .A1(n9801), .A2(n9812), .ZN(n8441) );
  NAND2_X1 U7578 ( .A1(n6010), .A2(n8441), .ZN(n9785) );
  NAND2_X1 U7579 ( .A1(n9788), .A2(n8318), .ZN(n6011) );
  INV_X1 U7580 ( .A(n8466), .ZN(n6012) );
  NAND2_X1 U7581 ( .A1(n6011), .A2(n6012), .ZN(n6014) );
  INV_X1 U7582 ( .A(n8318), .ZN(n8426) );
  NOR2_X1 U7583 ( .A1(n6012), .A2(n8426), .ZN(n6013) );
  NAND2_X1 U7584 ( .A1(n6014), .A2(n6052), .ZN(n6016) );
  OR2_X1 U7585 ( .A1(n7458), .A2(n9745), .ZN(n6015) );
  NAND2_X1 U7586 ( .A1(n8473), .A2(n8480), .ZN(n8482) );
  NAND2_X1 U7587 ( .A1(n6016), .A2(n10152), .ZN(n6019) );
  INV_X1 U7588 ( .A(n8337), .ZN(n9654) );
  INV_X1 U7589 ( .A(n8191), .ZN(n6017) );
  AOI22_X1 U7590 ( .A1(n9654), .A2(n10149), .B1(n10147), .B2(n9656), .ZN(n6018) );
  NAND2_X1 U7591 ( .A1(n6019), .A2(n6018), .ZN(n9774) );
  INV_X1 U7592 ( .A(n9979), .ZN(n9783) );
  NAND2_X1 U7593 ( .A1(n6970), .A2(n7061), .ZN(n7153) );
  OR2_X1 U7594 ( .A1(n7153), .A2(n6807), .ZN(n7154) );
  AND2_X1 U7595 ( .A1(n6911), .A2(n10321), .ZN(n7008) );
  NAND2_X1 U7596 ( .A1(n7008), .A2(n7263), .ZN(n7074) );
  NOR2_X1 U7597 ( .A1(n7074), .A2(n7075), .ZN(n7073) );
  NAND2_X1 U7598 ( .A1(n7073), .A2(n7411), .ZN(n7362) );
  INV_X1 U7599 ( .A(n7474), .ZN(n10105) );
  INV_X1 U7600 ( .A(n8250), .ZN(n10171) );
  INV_X1 U7601 ( .A(n9497), .ZN(n8161) );
  INV_X1 U7602 ( .A(n10030), .ZN(n9941) );
  INV_X1 U7603 ( .A(n10025), .ZN(n9925) );
  NAND2_X1 U7604 ( .A1(n9938), .A2(n9925), .ZN(n9922) );
  INV_X1 U7605 ( .A(n10009), .ZN(n9876) );
  INV_X1 U7606 ( .A(n10003), .ZN(n9861) );
  INV_X1 U7607 ( .A(n9990), .ZN(n9819) );
  NOR2_X2 U7608 ( .A1(n9813), .A2(n9801), .ZN(n9800) );
  AOI21_X1 U7609 ( .B1(n9778), .B2(n6028), .A(n10313), .ZN(n6020) );
  NOR2_X1 U7610 ( .A1(n9774), .A2(n9768), .ZN(n6021) );
  INV_X1 U7611 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7612 ( .A1(n6023), .A2(n6766), .ZN(n6024) );
  NOR2_X1 U7613 ( .A1(n6488), .A2(n6025), .ZN(n6035) );
  AND2_X2 U7614 ( .A1(n6035), .A2(n6026), .ZN(n10344) );
  NAND2_X1 U7615 ( .A1(n10344), .A2(n10031), .ZN(n10042) );
  NAND2_X1 U7616 ( .A1(n6028), .A2(n6029), .ZN(n6030) );
  NAND2_X1 U7617 ( .A1(n6031), .A2(n6030), .ZN(P1_U3551) );
  INV_X1 U7618 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U7619 ( .A1(n6482), .A2(n6485), .ZN(n6034) );
  INV_X1 U7620 ( .A(n6032), .ZN(n6033) );
  AOI22_X1 U7621 ( .A1(n6034), .A2(n6483), .B1(n6482), .B2(n6033), .ZN(n6767)
         );
  AND2_X2 U7622 ( .A1(n6035), .A2(n6767), .ZN(n10336) );
  NAND2_X1 U7623 ( .A1(n10336), .A2(n10031), .ZN(n10076) );
  NAND2_X1 U7624 ( .A1(n6028), .A2(n7979), .ZN(n6038) );
  NAND2_X1 U7625 ( .A1(n6039), .A2(n6038), .ZN(P1_U3519) );
  INV_X1 U7626 ( .A(n6043), .ZN(n6045) );
  MUX2_X1 U7627 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8204), .Z(n8192) );
  INV_X1 U7628 ( .A(SI_29_), .ZN(n6046) );
  XNOR2_X1 U7629 ( .A(n8192), .B(n6046), .ZN(n6047) );
  NAND2_X1 U7630 ( .A1(n9464), .A2(n5363), .ZN(n6049) );
  NAND2_X1 U7631 ( .A1(n4482), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6048) );
  AOI211_X1 U7632 ( .C1(n8338), .C2(n6051), .A(n10313), .B(n9754), .ZN(n9760)
         );
  INV_X1 U7633 ( .A(P1_B_REG_SCAN_IN), .ZN(n6053) );
  OAI21_X1 U7634 ( .B1(n10207), .B2(n6053), .A(n10149), .ZN(n9749) );
  NAND2_X1 U7635 ( .A1(n6509), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7636 ( .A1(n5287), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7637 ( .A1(n4487), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6054) );
  AND3_X1 U7638 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n8408) );
  INV_X1 U7639 ( .A(n6057), .ZN(n6058) );
  NAND2_X1 U7640 ( .A1(n8338), .A2(n6029), .ZN(n6059) );
  NAND2_X1 U7641 ( .A1(n6060), .A2(n6059), .ZN(P1_U3552) );
  INV_X2 U7642 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U7643 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6067) );
  NAND4_X1 U7644 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n6070)
         );
  NAND4_X1 U7645 ( .A1(n6068), .A2(n6347), .A3(n6283), .A4(n6282), .ZN(n6069)
         );
  NOR2_X1 U7646 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  INV_X1 U7647 ( .A(n6116), .ZN(n6074) );
  INV_X1 U7648 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6075) );
  INV_X1 U7649 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7650 ( .A1(n6111), .A2(n6076), .ZN(n6077) );
  NAND2_X1 U7651 ( .A1(n6077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6108) );
  INV_X1 U7652 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6107) );
  NOR2_X1 U7653 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6082) );
  NOR2_X1 U7654 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6081) );
  NOR2_X1 U7655 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n6080) );
  NOR2_X1 U7656 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6079) );
  NAND2_X1 U7657 ( .A1(n6086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6085) );
  MUX2_X1 U7658 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6085), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6087) );
  AND2_X1 U7659 ( .A1(n6087), .A2(n6148), .ZN(n8063) );
  NOR2_X1 U7660 ( .A1(n7921), .A2(n8063), .ZN(n10381) );
  NOR2_X1 U7661 ( .A1(n6088), .A2(n6183), .ZN(n6089) );
  MUX2_X1 U7662 ( .A(n6183), .B(n6089), .S(P2_IR_REG_25__SCAN_IN), .Z(n6091)
         );
  INV_X1 U7663 ( .A(n6086), .ZN(n6090) );
  XOR2_X1 U7664 ( .A(n7921), .B(P2_B_REG_SCAN_IN), .Z(n6092) );
  NAND2_X1 U7665 ( .A1(n6095), .A2(n6092), .ZN(n6093) );
  INV_X1 U7666 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10382) );
  AND2_X1 U7667 ( .A1(n10377), .A2(n10382), .ZN(n6094) );
  INV_X1 U7668 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10384) );
  INV_X1 U7669 ( .A(n6095), .ZN(n8045) );
  NOR2_X1 U7670 ( .A1(n8045), .A2(n8063), .ZN(n10386) );
  AOI21_X1 U7671 ( .B1(n10377), .B2(n10384), .A(n10386), .ZN(n6679) );
  NOR4_X1 U7672 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6099) );
  NOR4_X1 U7673 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6098) );
  NOR4_X1 U7674 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6097) );
  NOR4_X1 U7675 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6096) );
  NAND4_X1 U7676 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n6105)
         );
  NOR2_X1 U7677 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n6103) );
  NOR4_X1 U7678 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6102) );
  NOR4_X1 U7679 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6101) );
  NOR4_X1 U7680 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6100) );
  NAND4_X1 U7681 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n6104)
         );
  OAI21_X1 U7682 ( .B1(n6105), .B2(n6104), .A(n10377), .ZN(n6678) );
  NAND2_X1 U7683 ( .A1(n6679), .A2(n6678), .ZN(n7018) );
  AND2_X1 U7684 ( .A1(n8045), .A2(n8063), .ZN(n6106) );
  NAND2_X1 U7685 ( .A1(n7921), .A2(n6106), .ZN(n6521) );
  OR2_X1 U7686 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  NAND2_X1 U7687 ( .A1(n6110), .A2(n6109), .ZN(n6492) );
  NAND2_X1 U7688 ( .A1(n6521), .A2(n6492), .ZN(n6415) );
  OR2_X1 U7689 ( .A1(n6413), .A2(n8931), .ZN(n6418) );
  NAND2_X1 U7690 ( .A1(n6114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U7691 ( .A(n6115), .B(n6075), .ZN(n6683) );
  NAND2_X1 U7692 ( .A1(n6116), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6117) );
  AND2_X1 U7693 ( .A1(n6683), .A2(n9297), .ZN(n8932) );
  INV_X1 U7694 ( .A(n8932), .ZN(n6417) );
  NAND2_X1 U7695 ( .A1(n6141), .A2(n8763), .ZN(n6491) );
  INV_X1 U7696 ( .A(n6491), .ZN(n6519) );
  OR2_X1 U7697 ( .A1(n9437), .A2(n6519), .ZN(n6118) );
  NAND2_X1 U7698 ( .A1(n8705), .A2(n8741), .ZN(n8502) );
  INV_X1 U7699 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6124) );
  XNOR2_X2 U7700 ( .A(n6125), .B(n6124), .ZN(n6126) );
  NAND2_X1 U7701 ( .A1(n4478), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6140) );
  INV_X1 U7702 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8135) );
  OR2_X1 U7703 ( .A1(n6175), .A2(n8135), .ZN(n6139) );
  NAND2_X2 U7704 ( .A1(n9461), .A2(n9465), .ZN(n6194) );
  NAND3_X1 U7705 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n6250) );
  INV_X1 U7706 ( .A(n6250), .ZN(n6127) );
  INV_X1 U7707 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7348) );
  INV_X1 U7708 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7709 ( .A1(n6395), .A2(n6133), .ZN(n6134) );
  NAND2_X1 U7710 ( .A1(n6420), .A2(n6134), .ZN(n9334) );
  OR2_X1 U7711 ( .A1(n6194), .A2(n9334), .ZN(n6138) );
  INV_X1 U7712 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7713 ( .A1(n6220), .A2(n6136), .ZN(n6137) );
  NOR2_X1 U7714 ( .A1(n8502), .A2(n9310), .ZN(n6412) );
  INV_X2 U7715 ( .A(n8741), .ZN(n8625) );
  NOR2_X1 U7716 ( .A1(n9310), .A2(n8625), .ZN(n8074) );
  NOR2_X1 U7717 ( .A1(n4808), .A2(n8074), .ZN(n6411) );
  NAND2_X1 U7718 ( .A1(n8763), .A2(n6683), .ZN(n7028) );
  NAND2_X4 U7719 ( .A1(n6144), .A2(n7028), .ZN(n8599) );
  NAND2_X1 U7720 ( .A1(n6148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6149) );
  INV_X2 U7721 ( .A(n6168), .ZN(n8066) );
  NAND2_X1 U7722 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6152) );
  XNOR2_X1 U7723 ( .A(n6152), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U7724 ( .A1(n8066), .A2(n8949), .ZN(n6153) );
  INV_X1 U7725 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6526) );
  OR2_X1 U7726 ( .A1(n6175), .A2(n6526), .ZN(n6157) );
  NAND2_X1 U7727 ( .A1(n6174), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6156) );
  INV_X1 U7728 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7052) );
  OR2_X1 U7729 ( .A1(n6194), .A2(n7052), .ZN(n6155) );
  INV_X1 U7730 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7051) );
  OR2_X1 U7731 ( .A1(n4480), .A2(n7051), .ZN(n6154) );
  AND4_X2 U7732 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n8189)
         );
  OR2_X1 U7733 ( .A1(n8189), .A2(n8625), .ZN(n6172) );
  NAND2_X1 U7734 ( .A1(n6174), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6163) );
  INV_X1 U7735 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10345) );
  OR2_X1 U7736 ( .A1(n6175), .A2(n10345), .ZN(n6162) );
  INV_X1 U7737 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6158) );
  OR2_X1 U7738 ( .A1(n4480), .A2(n6158), .ZN(n6161) );
  INV_X1 U7739 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6159) );
  OR2_X1 U7740 ( .A1(n6194), .A2(n6159), .ZN(n6160) );
  NAND2_X1 U7741 ( .A1(n8204), .A2(SI_0_), .ZN(n6165) );
  INV_X1 U7742 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7743 ( .A1(n6165), .A2(n6164), .ZN(n6167) );
  AND2_X1 U7744 ( .A1(n6167), .A2(n6166), .ZN(n9475) );
  MUX2_X1 U7745 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9475), .S(n8509), .Z(n10387)
         );
  NAND2_X1 U7746 ( .A1(n8945), .A2(n10387), .ZN(n7164) );
  INV_X1 U7747 ( .A(n7164), .ZN(n6791) );
  NAND2_X1 U7748 ( .A1(n6791), .A2(n8741), .ZN(n8184) );
  INV_X1 U7749 ( .A(n10387), .ZN(n8762) );
  NAND2_X1 U7750 ( .A1(n8762), .A2(n6304), .ZN(n6169) );
  AND2_X1 U7751 ( .A1(n8184), .A2(n6169), .ZN(n6885) );
  INV_X1 U7752 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7753 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  NAND2_X1 U7754 ( .A1(n6174), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6180) );
  OR2_X1 U7755 ( .A1(n6175), .A2(n10446), .ZN(n6179) );
  INV_X1 U7756 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6176) );
  OR2_X1 U7757 ( .A1(n6194), .A2(n6176), .ZN(n6178) );
  INV_X1 U7758 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7136) );
  OR2_X1 U7759 ( .A1(n4480), .A2(n7136), .ZN(n6177) );
  AND4_X2 U7760 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n6893)
         );
  INV_X1 U7761 ( .A(n6893), .ZN(n6181) );
  AND2_X1 U7762 ( .A1(n6181), .A2(n8741), .ZN(n6189) );
  INV_X1 U7763 ( .A(n6189), .ZN(n6187) );
  NAND2_X1 U7764 ( .A1(n8622), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7765 ( .A1(n8066), .A2(n8960), .ZN(n6185) );
  OAI211_X1 U7766 ( .C1(n6463), .C2(n6241), .A(n6186), .B(n6185), .ZN(n6787)
         );
  XNOR2_X1 U7767 ( .A(n8599), .B(n6787), .ZN(n6188) );
  INV_X1 U7768 ( .A(n6188), .ZN(n6894) );
  NAND2_X1 U7769 ( .A1(n6187), .A2(n6894), .ZN(n6190) );
  NAND2_X1 U7770 ( .A1(n6189), .A2(n6188), .ZN(n6192) );
  NAND2_X1 U7771 ( .A1(n6190), .A2(n6192), .ZN(n6838) );
  NAND2_X1 U7772 ( .A1(n6897), .A2(n6192), .ZN(n6208) );
  NAND2_X1 U7773 ( .A1(n6174), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6198) );
  INV_X1 U7774 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6193) );
  OR2_X1 U7775 ( .A1(n6175), .A2(n6193), .ZN(n6197) );
  OR2_X1 U7776 ( .A1(n6194), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6196) );
  INV_X1 U7777 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6551) );
  OR2_X1 U7778 ( .A1(n4480), .A2(n6551), .ZN(n6195) );
  NOR2_X1 U7779 ( .A1(n7134), .A2(n8625), .ZN(n6204) );
  NAND2_X1 U7780 ( .A1(n8622), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6203) );
  NOR2_X1 U7781 ( .A1(n6184), .A2(n6183), .ZN(n6199) );
  MUX2_X1 U7782 ( .A(n6183), .B(n6199), .S(P2_IR_REG_3__SCAN_IN), .Z(n6201) );
  NOR2_X1 U7783 ( .A1(n6201), .A2(n6200), .ZN(n6545) );
  NAND2_X1 U7784 ( .A1(n8066), .A2(n6545), .ZN(n6202) );
  OAI211_X1 U7785 ( .C1(n6470), .C2(n6241), .A(n6203), .B(n6202), .ZN(n7027)
         );
  XNOR2_X1 U7786 ( .A(n8599), .B(n7027), .ZN(n6984) );
  NAND2_X1 U7787 ( .A1(n6204), .A2(n6984), .ZN(n6218) );
  INV_X1 U7788 ( .A(n6204), .ZN(n6206) );
  INV_X1 U7789 ( .A(n6984), .ZN(n6205) );
  NAND2_X1 U7790 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  AND2_X1 U7791 ( .A1(n6218), .A2(n6207), .ZN(n6895) );
  NAND2_X1 U7792 ( .A1(n6208), .A2(n6895), .ZN(n6898) );
  NAND2_X1 U7793 ( .A1(n6174), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6213) );
  INV_X1 U7794 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6209) );
  OR2_X1 U7795 ( .A1(n6175), .A2(n6209), .ZN(n6212) );
  XNOR2_X1 U7796 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7041) );
  OR2_X1 U7797 ( .A1(n6194), .A2(n7041), .ZN(n6211) );
  INV_X1 U7798 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6555) );
  OR2_X1 U7799 ( .A1(n4480), .A2(n6555), .ZN(n6210) );
  NAND2_X1 U7800 ( .A1(n8622), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6217) );
  OR2_X1 U7801 ( .A1(n6200), .A2(n6183), .ZN(n6215) );
  XNOR2_X1 U7802 ( .A(n6215), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U7803 ( .A1(n8066), .A2(n6597), .ZN(n6216) );
  XNOR2_X1 U7804 ( .A(n8599), .B(n7046), .ZN(n6237) );
  AND2_X1 U7805 ( .A1(n6983), .A2(n6218), .ZN(n6219) );
  NAND2_X1 U7806 ( .A1(n6898), .A2(n6219), .ZN(n6982) );
  NAND2_X1 U7807 ( .A1(n6174), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6229) );
  INV_X1 U7808 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6221) );
  OR2_X1 U7809 ( .A1(n6175), .A2(n6221), .ZN(n6228) );
  INV_X1 U7810 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7811 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6222) );
  NAND2_X1 U7812 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  NAND2_X1 U7813 ( .A1(n6250), .A2(n6224), .ZN(n10376) );
  OR2_X1 U7814 ( .A1(n6194), .A2(n10376), .ZN(n6227) );
  INV_X1 U7815 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7816 ( .A1(n4480), .A2(n6225), .ZN(n6226) );
  NOR2_X1 U7817 ( .A1(n7120), .A2(n8625), .ZN(n6233) );
  INV_X1 U7818 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6460) );
  INV_X1 U7819 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7820 ( .A1(n6200), .A2(n6230), .ZN(n6285) );
  NAND2_X1 U7821 ( .A1(n6285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6242) );
  XNOR2_X1 U7822 ( .A(n6242), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6556) );
  INV_X1 U7823 ( .A(n6556), .ZN(n6590) );
  OAI22_X1 U7824 ( .A1(n6214), .A2(n6460), .B1(n8509), .B2(n6590), .ZN(n6231)
         );
  INV_X1 U7825 ( .A(n6231), .ZN(n6232) );
  OAI21_X1 U7826 ( .B1(n6472), .B2(n6241), .A(n6232), .ZN(n7113) );
  XNOR2_X1 U7827 ( .A(n7113), .B(n8599), .ZN(n6234) );
  NAND2_X1 U7828 ( .A1(n6233), .A2(n6234), .ZN(n6256) );
  INV_X1 U7829 ( .A(n6233), .ZN(n6235) );
  INV_X1 U7830 ( .A(n6234), .ZN(n6938) );
  NAND2_X1 U7831 ( .A1(n6235), .A2(n6938), .ZN(n6236) );
  AND2_X1 U7832 ( .A1(n6256), .A2(n6236), .ZN(n6919) );
  INV_X1 U7833 ( .A(n6237), .ZN(n6238) );
  NAND2_X1 U7834 ( .A1(n6239), .A2(n6238), .ZN(n6917) );
  AND2_X1 U7835 ( .A1(n6919), .A2(n6917), .ZN(n6240) );
  NAND2_X1 U7836 ( .A1(n6982), .A2(n6240), .ZN(n6918) );
  INV_X2 U7837 ( .A(n6241), .ZN(n6262) );
  NAND2_X1 U7838 ( .A1(n6474), .A2(n6262), .ZN(n6248) );
  INV_X1 U7839 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7840 ( .A1(n6242), .A2(n6282), .ZN(n6243) );
  NAND2_X1 U7841 ( .A1(n6243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7842 ( .A1(n6244), .A2(n6283), .ZN(n6263) );
  OR2_X1 U7843 ( .A1(n6244), .A2(n6283), .ZN(n6245) );
  INV_X1 U7844 ( .A(n6572), .ZN(n6565) );
  OAI22_X1 U7845 ( .A1(n6214), .A2(n6475), .B1(n8509), .B2(n6565), .ZN(n6246)
         );
  INV_X1 U7846 ( .A(n6246), .ZN(n6247) );
  NAND2_X1 U7847 ( .A1(n6248), .A2(n6247), .ZN(n10410) );
  XNOR2_X1 U7848 ( .A(n10410), .B(n8599), .ZN(n6258) );
  NAND2_X1 U7849 ( .A1(n6174), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6255) );
  INV_X1 U7850 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6249) );
  OR2_X1 U7851 ( .A1(n6175), .A2(n6249), .ZN(n6254) );
  INV_X1 U7852 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7123) );
  OR2_X1 U7853 ( .A1(n4480), .A2(n7123), .ZN(n6253) );
  INV_X1 U7854 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U7855 ( .A1(n6250), .A2(n7615), .ZN(n6251) );
  NAND2_X1 U7856 ( .A1(n6269), .A2(n6251), .ZN(n7125) );
  OR2_X1 U7857 ( .A1(n6194), .A2(n7125), .ZN(n6252) );
  NAND4_X1 U7858 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n10363)
         );
  NAND2_X1 U7859 ( .A1(n10363), .A2(n8741), .ZN(n6259) );
  XNOR2_X1 U7860 ( .A(n6258), .B(n6259), .ZN(n6937) );
  AND2_X1 U7861 ( .A1(n6937), .A2(n6256), .ZN(n6257) );
  INV_X1 U7862 ( .A(n6258), .ZN(n6260) );
  NAND2_X1 U7863 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  NAND2_X1 U7864 ( .A1(n6478), .A2(n6262), .ZN(n6267) );
  INV_X1 U7865 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U7866 ( .A1(n6263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6264) );
  INV_X1 U7867 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7868 ( .A(n6264), .B(n6281), .ZN(n6665) );
  OAI22_X1 U7869 ( .A1(n6214), .A2(n6481), .B1(n8509), .B2(n6665), .ZN(n6265)
         );
  INV_X1 U7870 ( .A(n6265), .ZN(n6266) );
  NAND2_X1 U7871 ( .A1(n6267), .A2(n6266), .ZN(n7332) );
  XNOR2_X1 U7872 ( .A(n7332), .B(n8599), .ZN(n6275) );
  NAND2_X1 U7873 ( .A1(n6174), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6274) );
  INV_X1 U7874 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6567) );
  OR2_X1 U7875 ( .A1(n6175), .A2(n6567), .ZN(n6273) );
  INV_X1 U7876 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7877 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  NAND2_X1 U7878 ( .A1(n6291), .A2(n6270), .ZN(n7202) );
  OR2_X1 U7879 ( .A1(n6194), .A2(n7202), .ZN(n6272) );
  INV_X1 U7880 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6575) );
  OR2_X1 U7881 ( .A1(n4480), .A2(n6575), .ZN(n6271) );
  NOR2_X1 U7882 ( .A1(n7194), .A2(n8625), .ZN(n6276) );
  NAND2_X1 U7883 ( .A1(n6275), .A2(n6276), .ZN(n6280) );
  INV_X1 U7884 ( .A(n6275), .ZN(n6950) );
  INV_X1 U7885 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U7886 ( .A1(n6950), .A2(n6277), .ZN(n6278) );
  NAND2_X1 U7887 ( .A1(n6280), .A2(n6278), .ZN(n6814) );
  NAND2_X1 U7888 ( .A1(n6486), .A2(n6262), .ZN(n6290) );
  NAND3_X1 U7889 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n6284) );
  NAND2_X1 U7890 ( .A1(n6302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  INV_X1 U7891 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6286) );
  XNOR2_X1 U7892 ( .A(n6287), .B(n6286), .ZN(n6735) );
  OAI22_X1 U7893 ( .A1(n6214), .A2(n6490), .B1(n8509), .B2(n6735), .ZN(n6288)
         );
  INV_X1 U7894 ( .A(n6288), .ZN(n6289) );
  NAND2_X1 U7895 ( .A1(n6290), .A2(n6289), .ZN(n7311) );
  XNOR2_X1 U7896 ( .A(n7311), .B(n8599), .ZN(n6297) );
  NAND2_X1 U7897 ( .A1(n6174), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6296) );
  INV_X1 U7898 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6659) );
  OR2_X1 U7899 ( .A1(n6175), .A2(n6659), .ZN(n6295) );
  INV_X1 U7900 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U7901 ( .A1(n6291), .A2(n7631), .ZN(n6292) );
  NAND2_X1 U7902 ( .A1(n6305), .A2(n6292), .ZN(n7247) );
  OR2_X1 U7903 ( .A1(n6194), .A2(n7247), .ZN(n6294) );
  INV_X1 U7904 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7248) );
  OR2_X1 U7905 ( .A1(n4480), .A2(n7248), .ZN(n6293) );
  NOR2_X1 U7906 ( .A1(n7310), .A2(n8625), .ZN(n6298) );
  NAND2_X1 U7907 ( .A1(n6297), .A2(n6298), .ZN(n6311) );
  INV_X1 U7908 ( .A(n6297), .ZN(n7168) );
  INV_X1 U7909 ( .A(n6298), .ZN(n6299) );
  NAND2_X1 U7910 ( .A1(n7168), .A2(n6299), .ZN(n6300) );
  AND2_X1 U7911 ( .A1(n6311), .A2(n6300), .ZN(n6948) );
  NAND2_X1 U7912 ( .A1(n6301), .A2(n6948), .ZN(n6951) );
  NOR2_X1 U7913 ( .A1(n6302), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6349) );
  OR2_X1 U7914 ( .A1(n6349), .A2(n6183), .ZN(n6317) );
  XNOR2_X1 U7915 ( .A(n6317), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7916 ( .A1(n8622), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8066), .B2(
        n6860), .ZN(n6303) );
  XNOR2_X1 U7917 ( .A(n7460), .B(n8626), .ZN(n6315) );
  NAND2_X1 U7918 ( .A1(n6174), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6310) );
  INV_X1 U7919 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6729) );
  OR2_X1 U7920 ( .A1(n6175), .A2(n6729), .ZN(n6309) );
  NAND2_X1 U7921 ( .A1(n6305), .A2(n7176), .ZN(n6306) );
  NAND2_X1 U7922 ( .A1(n6322), .A2(n6306), .ZN(n7323) );
  OR2_X1 U7923 ( .A1(n6194), .A2(n7323), .ZN(n6308) );
  INV_X1 U7924 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6736) );
  OR2_X1 U7925 ( .A1(n4480), .A2(n6736), .ZN(n6307) );
  NOR2_X1 U7926 ( .A1(n7374), .A2(n8625), .ZN(n6313) );
  XNOR2_X1 U7927 ( .A(n6315), .B(n6313), .ZN(n7181) );
  AND2_X1 U7928 ( .A1(n7181), .A2(n6311), .ZN(n6312) );
  INV_X1 U7929 ( .A(n6313), .ZN(n6314) );
  NAND2_X1 U7930 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U7931 ( .A1(n6317), .A2(n6347), .ZN(n6318) );
  NAND2_X1 U7932 ( .A1(n6318), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6319) );
  INV_X1 U7933 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6346) );
  OR2_X1 U7934 ( .A1(n6319), .A2(n6346), .ZN(n6320) );
  NAND2_X1 U7935 ( .A1(n6319), .A2(n6346), .ZN(n6333) );
  AOI22_X1 U7936 ( .A1(n8622), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8066), .B2(
        n7275), .ZN(n6321) );
  XNOR2_X1 U7937 ( .A(n7924), .B(n8599), .ZN(n6328) );
  NAND2_X1 U7938 ( .A1(n6174), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6327) );
  INV_X1 U7939 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6855) );
  OR2_X1 U7940 ( .A1(n6175), .A2(n6855), .ZN(n6326) );
  NAND2_X1 U7941 ( .A1(n6322), .A2(n7815), .ZN(n6323) );
  NAND2_X1 U7942 ( .A1(n6338), .A2(n6323), .ZN(n7380) );
  OR2_X1 U7943 ( .A1(n6194), .A2(n7380), .ZN(n6325) );
  INV_X1 U7944 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7381) );
  OR2_X1 U7945 ( .A1(n4480), .A2(n7381), .ZN(n6324) );
  NOR2_X1 U7946 ( .A1(n7923), .A2(n8625), .ZN(n6329) );
  NAND2_X1 U7947 ( .A1(n6328), .A2(n6329), .ZN(n6332) );
  INV_X1 U7948 ( .A(n6328), .ZN(n7288) );
  INV_X1 U7949 ( .A(n6329), .ZN(n6330) );
  NAND2_X1 U7950 ( .A1(n7288), .A2(n6330), .ZN(n6331) );
  NAND2_X1 U7951 ( .A1(n6332), .A2(n6331), .ZN(n7183) );
  NAND2_X1 U7952 ( .A1(n6499), .A2(n6262), .ZN(n6336) );
  NAND2_X1 U7953 ( .A1(n6333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6334) );
  XNOR2_X1 U7954 ( .A(n6334), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8973) );
  AOI22_X1 U7955 ( .A1(n8622), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8066), .B2(
        n8973), .ZN(n6335) );
  XNOR2_X1 U7956 ( .A(n7964), .B(n8626), .ZN(n6372) );
  NAND2_X1 U7957 ( .A1(n6174), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6344) );
  INV_X1 U7958 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7276) );
  OR2_X1 U7959 ( .A1(n6175), .A2(n7276), .ZN(n6343) );
  INV_X1 U7960 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7961 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  NAND2_X1 U7962 ( .A1(n6353), .A2(n6339), .ZN(n7965) );
  OR2_X1 U7963 ( .A1(n6194), .A2(n7965), .ZN(n6342) );
  INV_X1 U7964 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6340) );
  OR2_X1 U7965 ( .A1(n4480), .A2(n6340), .ZN(n6341) );
  NOR2_X1 U7966 ( .A1(n7955), .A2(n8625), .ZN(n6373) );
  XNOR2_X1 U7967 ( .A(n6372), .B(n6373), .ZN(n7289) );
  NAND2_X1 U7968 ( .A1(n6516), .A2(n6262), .ZN(n6352) );
  INV_X1 U7969 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6345) );
  AND3_X1 U7970 ( .A1(n6347), .A2(n6346), .A3(n6345), .ZN(n6348) );
  AND2_X1 U7971 ( .A1(n6349), .A2(n6348), .ZN(n6360) );
  OR2_X1 U7972 ( .A1(n6360), .A2(n6183), .ZN(n6350) );
  XNOR2_X1 U7973 ( .A(n6350), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7344) );
  AOI22_X1 U7974 ( .A1(n8622), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8066), .B2(
        n7344), .ZN(n6351) );
  XNOR2_X1 U7975 ( .A(n8010), .B(n8626), .ZN(n6375) );
  NAND2_X1 U7976 ( .A1(n6174), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6358) );
  INV_X1 U7977 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7277) );
  OR2_X1 U7978 ( .A1(n6175), .A2(n7277), .ZN(n6357) );
  INV_X1 U7979 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7958) );
  OR2_X1 U7980 ( .A1(n4480), .A2(n7958), .ZN(n6356) );
  INV_X1 U7981 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U7982 ( .A1(n6353), .A2(n7767), .ZN(n6354) );
  NAND2_X1 U7983 ( .A1(n6364), .A2(n6354), .ZN(n7957) );
  OR2_X1 U7984 ( .A1(n6194), .A2(n7957), .ZN(n6355) );
  OR2_X1 U7985 ( .A1(n8017), .A2(n8625), .ZN(n6376) );
  NAND2_X1 U7986 ( .A1(n6375), .A2(n6376), .ZN(n7438) );
  NAND2_X1 U7987 ( .A1(n6670), .A2(n6262), .ZN(n6362) );
  INV_X1 U7988 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7989 ( .A1(n6360), .A2(n6359), .ZN(n6746) );
  NAND2_X1 U7990 ( .A1(n6746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6387) );
  XNOR2_X1 U7991 ( .A(n6387), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7503) );
  AOI22_X1 U7992 ( .A1(n8622), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8066), .B2(
        n7503), .ZN(n6361) );
  NAND2_X1 U7993 ( .A1(n6174), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6369) );
  INV_X1 U7994 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6363) );
  OR2_X1 U7995 ( .A1(n6175), .A2(n6363), .ZN(n6368) );
  NAND2_X1 U7996 ( .A1(n6364), .A2(n7348), .ZN(n6365) );
  NAND2_X1 U7997 ( .A1(n6393), .A2(n6365), .ZN(n8022) );
  OR2_X1 U7998 ( .A1(n6194), .A2(n8022), .ZN(n6367) );
  INV_X1 U7999 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8023) );
  OR2_X1 U8000 ( .A1(n4480), .A2(n8023), .ZN(n6366) );
  NOR2_X1 U8001 ( .A1(n8012), .A2(n8625), .ZN(n6383) );
  AND2_X1 U8002 ( .A1(n7289), .A2(n6371), .ZN(n6370) );
  NAND2_X1 U8003 ( .A1(n7290), .A2(n6370), .ZN(n6381) );
  INV_X1 U8004 ( .A(n6372), .ZN(n6374) );
  NAND2_X1 U8005 ( .A1(n6374), .A2(n6373), .ZN(n7417) );
  INV_X1 U8006 ( .A(n6375), .ZN(n6378) );
  INV_X1 U8007 ( .A(n6376), .ZN(n6377) );
  NAND2_X1 U8008 ( .A1(n6378), .A2(n6377), .ZN(n7416) );
  AND2_X1 U8009 ( .A1(n7417), .A2(n7416), .ZN(n7436) );
  INV_X1 U8010 ( .A(n6382), .ZN(n6384) );
  NAND2_X1 U8011 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  NAND2_X1 U8012 ( .A1(n6674), .A2(n6262), .ZN(n6392) );
  INV_X1 U8013 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8014 ( .A1(n6387), .A2(n6744), .ZN(n6388) );
  NAND2_X1 U8015 ( .A1(n6388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6389) );
  INV_X1 U8016 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U8017 ( .A1(n6389), .A2(n6743), .ZN(n6407) );
  OR2_X1 U8018 ( .A1(n6389), .A2(n6743), .ZN(n6390) );
  AOI22_X1 U8019 ( .A1(n8622), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8133), .B2(
        n8066), .ZN(n6391) );
  XNOR2_X1 U8020 ( .A(n9436), .B(n8626), .ZN(n6400) );
  NAND2_X1 U8021 ( .A1(n6174), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6399) );
  INV_X1 U8022 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7501) );
  OR2_X1 U8023 ( .A1(n6175), .A2(n7501), .ZN(n6398) );
  INV_X1 U8024 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U8025 ( .A1(n6393), .A2(n7830), .ZN(n6394) );
  NAND2_X1 U8026 ( .A1(n6395), .A2(n6394), .ZN(n8059) );
  OR2_X1 U8027 ( .A1(n6194), .A2(n8059), .ZN(n6397) );
  INV_X1 U8028 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8051) );
  OR2_X1 U8029 ( .A1(n4480), .A2(n8051), .ZN(n6396) );
  OR2_X1 U8030 ( .A1(n8937), .A2(n8625), .ZN(n6401) );
  NAND2_X1 U8031 ( .A1(n6400), .A2(n6401), .ZN(n6406) );
  INV_X1 U8032 ( .A(n6400), .ZN(n6403) );
  INV_X1 U8033 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U8034 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  NAND2_X1 U8035 ( .A1(n6406), .A2(n6404), .ZN(n7525) );
  INV_X1 U8036 ( .A(n7525), .ZN(n6405) );
  NAND2_X1 U8037 ( .A1(n6749), .A2(n6262), .ZN(n6410) );
  NAND2_X1 U8038 ( .A1(n6407), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U8039 ( .A(n6408), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8994) );
  AOI22_X1 U8040 ( .A1(n8994), .A2(n8066), .B1(n8622), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6409) );
  XNOR2_X1 U8041 ( .A(n9429), .B(n8599), .ZN(n8077) );
  MUX2_X1 U8042 ( .A(n6412), .B(n6411), .S(n8075), .Z(n6430) );
  INV_X1 U8043 ( .A(n9429), .ZN(n9339) );
  AND2_X1 U8044 ( .A1(n6119), .A2(n4837), .ZN(n7022) );
  INV_X1 U8045 ( .A(n7022), .ZN(n10368) );
  NAND2_X1 U8046 ( .A1(n10411), .A2(n10369), .ZN(n6677) );
  OR2_X2 U8047 ( .A1(n8931), .A2(n6677), .ZN(n10375) );
  OAI21_X2 U8048 ( .B1(n6418), .B2(n10368), .A(n10375), .ZN(n8699) );
  NOR2_X1 U8049 ( .A1(n9339), .A2(n8717), .ZN(n6429) );
  NAND2_X1 U8050 ( .A1(n6413), .A2(n6677), .ZN(n6416) );
  NOR2_X1 U8051 ( .A1(n6491), .A2(n8932), .ZN(n6414) );
  NOR2_X1 U8052 ( .A1(n6415), .A2(n6414), .ZN(n7021) );
  NAND2_X1 U8053 ( .A1(n6416), .A2(n7021), .ZN(n6840) );
  OAI22_X1 U8054 ( .A1(n8710), .A2(n9334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6133), .ZN(n6428) );
  NOR2_X1 U8055 ( .A1(n6418), .A2(n6417), .ZN(n8674) );
  INV_X1 U8056 ( .A(n6535), .ZN(n6520) );
  NAND2_X1 U8057 ( .A1(n6519), .A2(n6520), .ZN(n9309) );
  NAND2_X1 U8058 ( .A1(n6174), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6425) );
  INV_X1 U8059 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U8060 ( .A1(n6420), .A2(n7667), .ZN(n6421) );
  NAND2_X1 U8061 ( .A1(n8087), .A2(n6421), .ZN(n9317) );
  OR2_X1 U8062 ( .A1(n9317), .A2(n6194), .ZN(n6424) );
  INV_X1 U8063 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8986) );
  OR2_X1 U8064 ( .A1(n6175), .A2(n8986), .ZN(n6423) );
  INV_X1 U8065 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9318) );
  OR2_X1 U8066 ( .A1(n4480), .A2(n9318), .ZN(n6422) );
  INV_X1 U8067 ( .A(n8674), .ZN(n6426) );
  NAND2_X1 U8068 ( .A1(n6519), .A2(n6535), .ZN(n9311) );
  OAI22_X1 U8069 ( .A1(n8696), .A2(n8937), .B1(n9295), .B2(n8711), .ZN(n6427)
         );
  OR4_X1 U8070 ( .A1(n6430), .A2(n6429), .A3(n6428), .A4(n6427), .ZN(P2_U3243)
         );
  INV_X1 U8071 ( .A(n6431), .ZN(n7531) );
  OR2_X1 U8072 ( .A1(n5248), .A2(n7531), .ZN(n6449) );
  OR2_X2 U8073 ( .A1(n6449), .A2(P1_U3084), .ZN(n10211) );
  INV_X1 U8074 ( .A(n10211), .ZN(P1_U4006) );
  NAND2_X1 U8075 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6492), .ZN(n10380) );
  INV_X2 U8076 ( .A(n8936), .ZN(P2_U3966) );
  OR2_X1 U8077 ( .A1(n7531), .A2(n8191), .ZN(n6432) );
  NAND2_X1 U8078 ( .A1(n6449), .A2(n6432), .ZN(n6452) );
  OR2_X1 U8079 ( .A1(n6452), .A2(n6433), .ZN(n6434) );
  NAND2_X1 U8080 ( .A1(n6434), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U8081 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6435), .ZN(n6808) );
  NAND2_X1 U8082 ( .A1(n10215), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6436) );
  OAI21_X1 U8083 ( .B1(n10215), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6436), .ZN(
        n10203) );
  INV_X1 U8084 ( .A(n10203), .ZN(n6438) );
  INV_X1 U8085 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6776) );
  MUX2_X1 U8086 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6776), .S(n6466), .Z(n6613)
         );
  AND2_X1 U8087 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6612) );
  NAND2_X1 U8088 ( .A1(n6466), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8089 ( .A1(n6611), .A2(n6437), .ZN(n10202) );
  NAND2_X1 U8090 ( .A1(n6438), .A2(n10202), .ZN(n10206) );
  INV_X1 U8091 ( .A(n10206), .ZN(n6439) );
  NAND2_X1 U8092 ( .A1(n6628), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6440) );
  OAI21_X1 U8093 ( .B1(n6628), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6440), .ZN(
        n6441) );
  OR2_X1 U8094 ( .A1(n5932), .A2(P1_U3084), .ZN(n10092) );
  OR2_X1 U8095 ( .A1(n6452), .A2(n10092), .ZN(n6446) );
  NOR2_X1 U8096 ( .A1(n6446), .A2(n10207), .ZN(n10284) );
  INV_X1 U8097 ( .A(n10284), .ZN(n10296) );
  AOI211_X1 U8098 ( .C1(n6442), .C2(n6441), .A(n6627), .B(n10296), .ZN(n6455)
         );
  INV_X1 U8099 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7256) );
  AND2_X1 U8100 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6606) );
  AND2_X1 U8101 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  AND2_X1 U8102 ( .A1(n6466), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8103 ( .A1(n10215), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6444) );
  OAI21_X1 U8104 ( .B1(n10215), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6444), .ZN(
        n10199) );
  NOR2_X1 U8105 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  AOI21_X1 U8106 ( .B1(n10215), .B2(P1_REG1_REG_2__SCAN_IN), .A(n10198), .ZN(
        n6448) );
  NAND2_X1 U8107 ( .A1(n6628), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6445) );
  OAI21_X1 U8108 ( .B1(n6628), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6445), .ZN(
        n6447) );
  NOR2_X1 U8109 ( .A1(n6448), .A2(n6447), .ZN(n6620) );
  INV_X1 U8110 ( .A(n6446), .ZN(n10192) );
  NAND2_X1 U8111 ( .A1(n10192), .A2(n10207), .ZN(n10288) );
  AOI211_X1 U8112 ( .C1(n6448), .C2(n6447), .A(n6620), .B(n10288), .ZN(n6454)
         );
  INV_X1 U8113 ( .A(n6449), .ZN(n6450) );
  NOR2_X2 U8114 ( .A1(P1_U3083), .A2(n6450), .ZN(n10306) );
  INV_X1 U8115 ( .A(n10306), .ZN(n10231) );
  INV_X1 U8116 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7538) );
  INV_X1 U8117 ( .A(n6628), .ZN(n6471) );
  INV_X1 U8118 ( .A(n10207), .ZN(n6451) );
  NAND2_X1 U8119 ( .A1(n6451), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10097) );
  NOR2_X1 U8120 ( .A1(n6452), .A2(n10097), .ZN(n10191) );
  NAND2_X1 U8121 ( .A1(n10191), .A2(n5932), .ZN(n10254) );
  OAI22_X1 U8122 ( .A1(n10231), .A2(n7538), .B1(n6471), .B2(n10254), .ZN(n6453) );
  OR4_X1 U8123 ( .A1(n6808), .A2(n6455), .A3(n6454), .A4(n6453), .ZN(P1_U3244)
         );
  NAND2_X1 U8124 ( .A1(n8204), .A2(P2_U3152), .ZN(n9463) );
  NOR2_X2 U8125 ( .A1(n8204), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9471) );
  AOI22_X1 U8126 ( .A1(n8960), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n9471), .ZN(n6456) );
  OAI21_X1 U8127 ( .B1(n6463), .B2(n9463), .A(n6456), .ZN(P2_U3356) );
  INV_X1 U8128 ( .A(n8949), .ZN(n6538) );
  CLKBUF_X1 U8129 ( .A(n9463), .Z(n9469) );
  INV_X1 U8130 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6457) );
  INV_X1 U8131 ( .A(n9471), .ZN(n7162) );
  OAI222_X1 U8132 ( .A1(P2_U3152), .A2(n6538), .B1(n9469), .B2(n6467), .C1(
        n6457), .C2(n7162), .ZN(P2_U3357) );
  INV_X1 U8133 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6458) );
  INV_X1 U8134 ( .A(n6545), .ZN(n6552) );
  OAI222_X1 U8135 ( .A1(n7162), .A2(n6458), .B1(n9469), .B2(n6470), .C1(
        P2_U3152), .C2(n6552), .ZN(P2_U3355) );
  INV_X1 U8136 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6459) );
  INV_X1 U8137 ( .A(n6597), .ZN(n6605) );
  OAI222_X1 U8138 ( .A1(n7162), .A2(n6459), .B1(n9469), .B2(n6465), .C1(
        P2_U3152), .C2(n6605), .ZN(P2_U3354) );
  OAI222_X1 U8139 ( .A1(n7162), .A2(n6460), .B1(n9469), .B2(n6472), .C1(
        P2_U3152), .C2(n6590), .ZN(P2_U3353) );
  NAND2_X1 U8140 ( .A1(n6461), .A2(P1_U3084), .ZN(n10081) );
  NAND2_X1 U8141 ( .A1(n8204), .A2(P1_U3084), .ZN(n10100) );
  INV_X1 U8142 ( .A(n10100), .ZN(n10079) );
  AOI22_X1 U8143 ( .A1(n10079), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n10215), 
        .B2(P1_STATE_REG_SCAN_IN), .ZN(n6462) );
  OAI21_X1 U8144 ( .B1(n6463), .B2(n10081), .A(n6462), .ZN(P1_U3351) );
  AOI22_X1 U8145 ( .A1(n10222), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10079), .ZN(n6464) );
  OAI21_X1 U8146 ( .B1(n6465), .B2(n10081), .A(n6464), .ZN(P1_U3349) );
  CLKBUF_X1 U8147 ( .A(n10100), .Z(n10086) );
  INV_X1 U8148 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6468) );
  OAI222_X1 U8149 ( .A1(n10086), .A2(n6468), .B1(n10081), .B2(n6467), .C1(
        n5259), .C2(P1_U3084), .ZN(P1_U3352) );
  INV_X1 U8150 ( .A(n10081), .ZN(n10095) );
  INV_X1 U8151 ( .A(n10095), .ZN(n10090) );
  INV_X1 U8152 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6469) );
  OAI222_X1 U8153 ( .A1(n6471), .A2(P1_U3084), .B1(n10090), .B2(n6470), .C1(
        n6469), .C2(n10100), .ZN(P1_U3350) );
  INV_X1 U8154 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6473) );
  INV_X1 U8155 ( .A(n6629), .ZN(n10239) );
  OAI222_X1 U8156 ( .A1(n10086), .A2(n6473), .B1(n10090), .B2(n6472), .C1(
        n10239), .C2(P1_U3084), .ZN(P1_U3348) );
  INV_X1 U8157 ( .A(n6474), .ZN(n6476) );
  OAI222_X1 U8158 ( .A1(n7162), .A2(n6475), .B1(n9469), .B2(n6476), .C1(
        P2_U3152), .C2(n6565), .ZN(P2_U3352) );
  INV_X1 U8159 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7833) );
  OAI222_X1 U8160 ( .A1(n10086), .A2(n7833), .B1(n10081), .B2(n6476), .C1(
        n10253), .C2(P1_U3084), .ZN(P1_U3347) );
  NAND2_X1 U8161 ( .A1(n8936), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n6477) );
  OAI21_X1 U8162 ( .B1(n8936), .B2(n9310), .A(n6477), .ZN(P2_U3567) );
  INV_X1 U8163 ( .A(n6712), .ZN(n6633) );
  INV_X1 U8164 ( .A(n6478), .ZN(n6480) );
  INV_X1 U8165 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6479) );
  OAI222_X1 U8166 ( .A1(n6633), .A2(P1_U3084), .B1(n10090), .B2(n6480), .C1(
        n6479), .C2(n10100), .ZN(P1_U3346) );
  OAI222_X1 U8167 ( .A1(n7162), .A2(n6481), .B1(n9469), .B2(n6480), .C1(
        P2_U3152), .C2(n6665), .ZN(P2_U3351) );
  NOR2_X1 U8168 ( .A1(n8486), .A2(n6482), .ZN(n10311) );
  NAND2_X1 U8169 ( .A1(n10311), .A2(n6483), .ZN(n6484) );
  OAI21_X1 U8170 ( .B1(n10311), .B2(n6485), .A(n6484), .ZN(P1_U3440) );
  INV_X1 U8171 ( .A(n6486), .ZN(n6489) );
  AOI22_X1 U8172 ( .A1(n10272), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10079), .ZN(n6487) );
  OAI21_X1 U8173 ( .B1(n6489), .B2(n10081), .A(n6487), .ZN(P1_U3345) );
  INV_X1 U8174 ( .A(n8486), .ZN(n6646) );
  NAND2_X1 U8175 ( .A1(n6488), .A2(n6646), .ZN(n6768) );
  OAI21_X1 U8176 ( .B1(n6646), .B2(n5900), .A(n6768), .ZN(P1_U3441) );
  OAI222_X1 U8177 ( .A1(n7162), .A2(n6490), .B1(n9469), .B2(n6489), .C1(
        P2_U3152), .C2(n6735), .ZN(P2_U3350) );
  OAI21_X1 U8178 ( .B1(n8931), .B2(n6491), .A(n8509), .ZN(n6494) );
  NOR2_X1 U8179 ( .A1(n6492), .A2(P2_U3152), .ZN(n8930) );
  INV_X1 U8180 ( .A(n8930), .ZN(n8934) );
  NAND2_X1 U8181 ( .A1(n8931), .A2(n8934), .ZN(n6493) );
  NAND2_X1 U8182 ( .A1(n6494), .A2(n6493), .ZN(n9056) );
  NOR2_X1 U8183 ( .A1(n10351), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8184 ( .A(n10290), .ZN(n6496) );
  INV_X1 U8185 ( .A(n6495), .ZN(n6497) );
  OAI222_X1 U8186 ( .A1(P1_U3084), .A2(n6496), .B1(n10081), .B2(n6497), .C1(
        n7855), .C2(n10100), .ZN(P1_U3344) );
  INV_X1 U8187 ( .A(n6860), .ZN(n6741) );
  OAI222_X1 U8188 ( .A1(n7162), .A2(n6498), .B1(n9469), .B2(n6497), .C1(n6741), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8189 ( .A(n6499), .ZN(n6515) );
  AOI22_X1 U8190 ( .A1(n8973), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9471), .ZN(n6500) );
  OAI21_X1 U8191 ( .B1(n6515), .B2(n9469), .A(n6500), .ZN(P2_U3347) );
  INV_X1 U8192 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U8193 ( .A1(n6174), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6504) );
  INV_X1 U8194 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6501) );
  OR2_X1 U8195 ( .A1(n6175), .A2(n6501), .ZN(n6503) );
  INV_X1 U8196 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9058) );
  OR2_X1 U8197 ( .A1(n4480), .A2(n9058), .ZN(n6502) );
  AND3_X1 U8198 ( .A1(n6504), .A2(n6503), .A3(n6502), .ZN(n8737) );
  INV_X1 U8199 ( .A(n8737), .ZN(n9059) );
  NAND2_X1 U8200 ( .A1(P2_U3966), .A2(n9059), .ZN(n6505) );
  OAI21_X1 U8201 ( .B1(P2_U3966), .B2(n7819), .A(n6505), .ZN(P2_U3583) );
  INV_X1 U8202 ( .A(n7275), .ZN(n6868) );
  INV_X1 U8203 ( .A(n6506), .ZN(n6508) );
  OAI222_X1 U8204 ( .A1(P2_U3152), .A2(n6868), .B1(n9469), .B2(n6508), .C1(
        n6507), .C2(n7162), .ZN(P2_U3348) );
  INV_X1 U8205 ( .A(n10304), .ZN(n6701) );
  OAI222_X1 U8206 ( .A1(P1_U3084), .A2(n6701), .B1(n10081), .B2(n6508), .C1(
        n7775), .C2(n10100), .ZN(P1_U3343) );
  INV_X1 U8207 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8208 ( .A1(n6509), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U8209 ( .A1(n5287), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U8210 ( .A1(n4487), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6510) );
  NAND3_X1 U8211 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(n9748) );
  NAND2_X1 U8212 ( .A1(P1_U4006), .A2(n9748), .ZN(n6513) );
  OAI21_X1 U8213 ( .B1(P1_U4006), .B2(n6514), .A(n6513), .ZN(P1_U3586) );
  INV_X1 U8214 ( .A(n6876), .ZN(n6872) );
  INV_X1 U8215 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7803) );
  OAI222_X1 U8216 ( .A1(P1_U3084), .A2(n6872), .B1(n10081), .B2(n6515), .C1(
        n7803), .C2(n10100), .ZN(P1_U3342) );
  INV_X1 U8217 ( .A(n6516), .ZN(n6517) );
  OAI222_X1 U8218 ( .A1(n10086), .A2(n7832), .B1(n10081), .B2(n6517), .C1(
        n7097), .C2(P1_U3084), .ZN(P1_U3341) );
  INV_X1 U8219 ( .A(n7344), .ZN(n7285) );
  OAI222_X1 U8220 ( .A1(n7162), .A2(n6518), .B1(n9469), .B2(n6517), .C1(
        P2_U3152), .C2(n7285), .ZN(P2_U3346) );
  OR2_X1 U8221 ( .A1(n8931), .A2(n6519), .ZN(n6524) );
  NAND2_X1 U8222 ( .A1(n6520), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9467) );
  OAI21_X1 U8223 ( .B1(n6521), .B2(n9467), .A(n8934), .ZN(n6522) );
  INV_X1 U8224 ( .A(n6522), .ZN(n6523) );
  NAND2_X1 U8225 ( .A1(n6524), .A2(n6523), .ZN(n6529) );
  NAND2_X1 U8226 ( .A1(n6529), .A2(n8509), .ZN(n6525) );
  NAND2_X1 U8227 ( .A1(n6525), .A2(n8936), .ZN(n6537) );
  INV_X1 U8228 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7669) );
  NOR2_X1 U8229 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7669), .ZN(n6533) );
  XOR2_X1 U8230 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8960), .Z(n8963) );
  MUX2_X1 U8231 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6526), .S(n8949), .Z(n8952)
         );
  AND2_X1 U8232 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8951) );
  NAND2_X1 U8233 ( .A1(n8952), .A2(n8951), .ZN(n8950) );
  OAI21_X1 U8234 ( .B1(n6526), .B2(n6538), .A(n8950), .ZN(n8962) );
  NAND2_X1 U8235 ( .A1(n8963), .A2(n8962), .ZN(n8961) );
  INV_X1 U8236 ( .A(n8961), .ZN(n6527) );
  AOI21_X1 U8237 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n8960), .A(n6527), .ZN(
        n6531) );
  XNOR2_X1 U8238 ( .A(n6545), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6530) );
  NOR2_X1 U8239 ( .A1(n6531), .A2(n6530), .ZN(n6544) );
  INV_X1 U8240 ( .A(n6534), .ZN(n9472) );
  NOR2_X1 U8241 ( .A1(n8066), .A2(n9472), .ZN(n6528) );
  AOI211_X1 U8242 ( .C1(n6531), .C2(n6530), .A(n6544), .B(n8134), .ZN(n6532)
         );
  AOI211_X1 U8243 ( .C1(n10351), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6533), .B(
        n6532), .ZN(n6543) );
  NOR2_X1 U8244 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  NAND2_X1 U8245 ( .A1(n6537), .A2(n6536), .ZN(n9048) );
  MUX2_X1 U8246 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7136), .S(n8960), .Z(n8959)
         );
  MUX2_X1 U8247 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7051), .S(n8949), .Z(n8947)
         );
  NAND3_X1 U8248 ( .A1(n8947), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n8946) );
  OAI21_X1 U8249 ( .B1(n7051), .B2(n6538), .A(n8946), .ZN(n8958) );
  NAND2_X1 U8250 ( .A1(n8959), .A2(n8958), .ZN(n8957) );
  NAND2_X1 U8251 ( .A1(n8960), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6539) );
  MUX2_X1 U8252 ( .A(n6551), .B(P2_REG2_REG_3__SCAN_IN), .S(n6545), .Z(n6540)
         );
  AOI21_X1 U8253 ( .B1(n8957), .B2(n6539), .A(n6540), .ZN(n6554) );
  INV_X1 U8254 ( .A(n6554), .ZN(n6600) );
  NAND3_X1 U8255 ( .A1(n6540), .A2(n8957), .A3(n6539), .ZN(n6541) );
  NAND3_X1 U8256 ( .A1(n10350), .A2(n6600), .A3(n6541), .ZN(n6542) );
  OAI211_X1 U8257 ( .C1(n7286), .C2(n6552), .A(n6543), .B(n6542), .ZN(P2_U3248) );
  NOR2_X1 U8258 ( .A1(n7615), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6940) );
  AOI21_X1 U8259 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6545), .A(n6544), .ZN(
        n6593) );
  XNOR2_X1 U8260 ( .A(n6597), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6592) );
  NOR2_X1 U8261 ( .A1(n6593), .A2(n6592), .ZN(n6591) );
  NAND2_X1 U8262 ( .A1(n6556), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U8263 ( .B1(n6556), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6546), .ZN(
        n6581) );
  NAND2_X1 U8264 ( .A1(n6572), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6547) );
  OAI21_X1 U8265 ( .B1(n6572), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6547), .ZN(
        n6548) );
  AOI211_X1 U8266 ( .C1(n6549), .C2(n6548), .A(n6566), .B(n8134), .ZN(n6550)
         );
  AOI211_X1 U8267 ( .C1(n10351), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6940), .B(
        n6550), .ZN(n6564) );
  NAND2_X1 U8268 ( .A1(n6556), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6559) );
  NOR2_X1 U8269 ( .A1(n6552), .A2(n6551), .ZN(n6596) );
  MUX2_X1 U8270 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6555), .S(n6597), .Z(n6553)
         );
  OAI21_X1 U8271 ( .B1(n6554), .B2(n6596), .A(n6553), .ZN(n6602) );
  OAI21_X1 U8272 ( .B1(n6555), .B2(n6605), .A(n6602), .ZN(n6586) );
  MUX2_X1 U8273 ( .A(n6225), .B(P2_REG2_REG_5__SCAN_IN), .S(n6556), .Z(n6585)
         );
  INV_X1 U8274 ( .A(n6585), .ZN(n6557) );
  NAND2_X1 U8275 ( .A1(n6586), .A2(n6557), .ZN(n6558) );
  NAND2_X1 U8276 ( .A1(n6559), .A2(n6558), .ZN(n6562) );
  MUX2_X1 U8277 ( .A(n7123), .B(P2_REG2_REG_6__SCAN_IN), .S(n6572), .Z(n6560)
         );
  INV_X1 U8278 ( .A(n6560), .ZN(n6561) );
  NAND2_X1 U8279 ( .A1(n6561), .A2(n6562), .ZN(n6573) );
  OAI211_X1 U8280 ( .C1(n6562), .C2(n6561), .A(n10350), .B(n6573), .ZN(n6563)
         );
  OAI211_X1 U8281 ( .C1(n7286), .C2(n6565), .A(n6564), .B(n6563), .ZN(P2_U3251) );
  NOR2_X1 U8282 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6268), .ZN(n6571) );
  AOI21_X1 U8283 ( .B1(n6572), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6566), .ZN(
        n6569) );
  MUX2_X1 U8284 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6567), .S(n6665), .Z(n6568)
         );
  NOR2_X1 U8285 ( .A1(n6569), .A2(n6568), .ZN(n6657) );
  AOI211_X1 U8286 ( .C1(n6569), .C2(n6568), .A(n6657), .B(n8134), .ZN(n6570)
         );
  AOI211_X1 U8287 ( .C1(n10351), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6571), .B(
        n6570), .ZN(n6579) );
  NAND2_X1 U8288 ( .A1(n6572), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8289 ( .A1(n6574), .A2(n6573), .ZN(n6577) );
  MUX2_X1 U8290 ( .A(n6575), .B(P2_REG2_REG_7__SCAN_IN), .S(n6665), .Z(n6576)
         );
  NAND2_X1 U8291 ( .A1(n6576), .A2(n6577), .ZN(n6664) );
  OAI211_X1 U8292 ( .C1(n6577), .C2(n6576), .A(n10350), .B(n6664), .ZN(n6578)
         );
  OAI211_X1 U8293 ( .C1(n7286), .C2(n6665), .A(n6579), .B(n6578), .ZN(P2_U3252) );
  NOR2_X1 U8294 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6223), .ZN(n6584) );
  AOI211_X1 U8295 ( .C1(n6582), .C2(n6581), .A(n8134), .B(n6580), .ZN(n6583)
         );
  AOI211_X1 U8296 ( .C1(n10351), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6584), .B(
        n6583), .ZN(n6589) );
  XNOR2_X1 U8297 ( .A(n6586), .B(n6585), .ZN(n6587) );
  NAND2_X1 U8298 ( .A1(n10350), .A2(n6587), .ZN(n6588) );
  OAI211_X1 U8299 ( .C1(n7286), .C2(n6590), .A(n6589), .B(n6588), .ZN(P2_U3250) );
  NAND2_X1 U8300 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6987) );
  INV_X1 U8301 ( .A(n6987), .ZN(n6595) );
  AOI211_X1 U8302 ( .C1(n6593), .C2(n6592), .A(n6591), .B(n8134), .ZN(n6594)
         );
  AOI211_X1 U8303 ( .C1(n10351), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6595), .B(
        n6594), .ZN(n6604) );
  INV_X1 U8304 ( .A(n6596), .ZN(n6599) );
  MUX2_X1 U8305 ( .A(n6555), .B(P2_REG2_REG_4__SCAN_IN), .S(n6597), .Z(n6598)
         );
  NAND3_X1 U8306 ( .A1(n6600), .A2(n6599), .A3(n6598), .ZN(n6601) );
  NAND3_X1 U8307 ( .A1(n10350), .A2(n6602), .A3(n6601), .ZN(n6603) );
  OAI211_X1 U8308 ( .C1(n7286), .C2(n6605), .A(n6604), .B(n6603), .ZN(P2_U3249) );
  INV_X1 U8309 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6619) );
  INV_X1 U8310 ( .A(n6606), .ZN(n6610) );
  INV_X1 U8311 ( .A(n6607), .ZN(n6609) );
  AOI211_X1 U8312 ( .C1(n6610), .C2(n6609), .A(n6608), .B(n10288), .ZN(n6617)
         );
  OAI211_X1 U8313 ( .C1(n6613), .C2(n6612), .A(n10284), .B(n6611), .ZN(n6614)
         );
  INV_X1 U8314 ( .A(n6614), .ZN(n6616) );
  INV_X1 U8315 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6775) );
  OAI22_X1 U8316 ( .A1(n10254), .A2(n5259), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6775), .ZN(n6615) );
  NOR3_X1 U8317 ( .A1(n6617), .A2(n6616), .A3(n6615), .ZN(n6618) );
  OAI21_X1 U8318 ( .B1(n10231), .B2(n6619), .A(n6618), .ZN(P1_U3242) );
  INV_X1 U8319 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6640) );
  INV_X1 U8320 ( .A(n10288), .ZN(n10302) );
  INV_X1 U8321 ( .A(n10253), .ZN(n6631) );
  XNOR2_X1 U8322 ( .A(n6631), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10257) );
  XNOR2_X1 U8323 ( .A(n10222), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10223) );
  INV_X1 U8324 ( .A(n10224), .ZN(n6621) );
  OAI22_X1 U8325 ( .A1(n10223), .A2(n6621), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n10222), .ZN(n10233) );
  NAND2_X1 U8326 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6629), .ZN(n6622) );
  OAI21_X1 U8327 ( .B1(n6629), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6622), .ZN(
        n10232) );
  AOI21_X1 U8328 ( .B1(n6629), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10235), .ZN(
        n6623) );
  INV_X1 U8329 ( .A(n6623), .ZN(n10256) );
  OAI22_X1 U8330 ( .A1(n10257), .A2(n10256), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6631), .ZN(n6625) );
  INV_X1 U8331 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7219) );
  AOI22_X1 U8332 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6712), .B1(n6633), .B2(
        n7219), .ZN(n6624) );
  OAI21_X1 U8333 ( .B1(n6625), .B2(n6624), .A(n6702), .ZN(n6637) );
  NOR2_X1 U8334 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6629), .ZN(n6626) );
  AOI21_X1 U8335 ( .B1(n6629), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6626), .ZN(
        n10243) );
  XNOR2_X1 U8336 ( .A(n10222), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U8337 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  OAI21_X1 U8338 ( .B1(n6629), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10241), .ZN(
        n6630) );
  INV_X1 U8339 ( .A(n6630), .ZN(n10249) );
  XNOR2_X1 U8340 ( .A(n10253), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10250) );
  INV_X1 U8341 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6632) );
  AOI22_X1 U8342 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6712), .B1(n6633), .B2(
        n6632), .ZN(n6634) );
  OAI21_X1 U8343 ( .B1(n6635), .B2(n6634), .A(n6711), .ZN(n6636) );
  AOI22_X1 U8344 ( .A1(n10302), .A2(n6637), .B1(n10284), .B2(n6636), .ZN(n6639) );
  INV_X1 U8345 ( .A(n10254), .ZN(n10305) );
  AND2_X1 U8346 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6996) );
  AOI21_X1 U8347 ( .B1(n10305), .B2(n6712), .A(n6996), .ZN(n6638) );
  OAI211_X1 U8348 ( .C1(n10231), .C2(n6640), .A(n6639), .B(n6638), .ZN(
        P1_U3248) );
  OAI21_X1 U8349 ( .B1(n6641), .B2(n6642), .A(n6643), .ZN(n10209) );
  AOI22_X1 U8350 ( .A1(n9607), .A2(n10209), .B1(n9648), .B2(n6851), .ZN(n6649)
         );
  NAND2_X1 U8351 ( .A1(n6644), .A2(n10329), .ZN(n6645) );
  NAND4_X1 U8352 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6766), .ZN(n9610)
         );
  AOI22_X1 U8353 ( .A1(n9640), .A2(n5950), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9610), .ZN(n6648) );
  NAND2_X1 U8354 ( .A1(n6649), .A2(n6648), .ZN(P1_U3230) );
  XNOR2_X1 U8355 ( .A(n6650), .B(n6651), .ZN(n6652) );
  XOR2_X1 U8356 ( .A(n6653), .B(n6652), .Z(n6656) );
  AOI22_X1 U8357 ( .A1(n9640), .A2(n9669), .B1(n9609), .B2(n9670), .ZN(n6655)
         );
  AOI22_X1 U8358 ( .A1(n9648), .A2(n5949), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9610), .ZN(n6654) );
  OAI211_X1 U8359 ( .C1(n6656), .C2(n9651), .A(n6655), .B(n6654), .ZN(P1_U3220) );
  NOR2_X1 U8360 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7631), .ZN(n6663) );
  INV_X1 U8361 ( .A(n6665), .ZN(n6658) );
  AOI21_X1 U8362 ( .B1(n6658), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6657), .ZN(
        n6661) );
  MUX2_X1 U8363 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6659), .S(n6735), .Z(n6660)
         );
  AOI211_X1 U8364 ( .C1(n6661), .C2(n6660), .A(n6727), .B(n8134), .ZN(n6662)
         );
  AOI211_X1 U8365 ( .C1(n10351), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6663), .B(
        n6662), .ZN(n6669) );
  OAI21_X1 U8366 ( .B1(n6665), .B2(n6575), .A(n6664), .ZN(n6667) );
  MUX2_X1 U8367 ( .A(n7248), .B(P2_REG2_REG_8__SCAN_IN), .S(n6735), .Z(n6666)
         );
  NAND2_X1 U8368 ( .A1(n6666), .A2(n6667), .ZN(n6734) );
  OAI211_X1 U8369 ( .C1(n6667), .C2(n6666), .A(n10350), .B(n6734), .ZN(n6668)
         );
  OAI211_X1 U8370 ( .C1(n7286), .C2(n6735), .A(n6669), .B(n6668), .ZN(P2_U3253) );
  INV_X1 U8371 ( .A(n6670), .ZN(n6672) );
  OAI222_X1 U8372 ( .A1(n10086), .A2(n6671), .B1(n10081), .B2(n6672), .C1(
        P1_U3084), .C2(n7484), .ZN(P1_U3340) );
  INV_X1 U8373 ( .A(n7503), .ZN(n7497) );
  OAI222_X1 U8374 ( .A1(n7162), .A2(n6673), .B1(n9463), .B2(n6672), .C1(n7497), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8375 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6675) );
  INV_X1 U8376 ( .A(n6674), .ZN(n6676) );
  INV_X1 U8377 ( .A(n8133), .ZN(n7500) );
  OAI222_X1 U8378 ( .A1(n7162), .A2(n6675), .B1(n9463), .B2(n6676), .C1(n7500), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8379 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7858) );
  INV_X1 U8380 ( .A(n9674), .ZN(n9678) );
  OAI222_X1 U8381 ( .A1(n10086), .A2(n7858), .B1(n10081), .B2(n6676), .C1(
        P1_U3084), .C2(n9678), .ZN(P1_U3339) );
  NAND4_X1 U8382 ( .A1(n6678), .A2(P2_STATE_REG_SCAN_IN), .A3(n7021), .A4(
        n6677), .ZN(n6680) );
  NOR2_X1 U8383 ( .A1(n6680), .A2(n6679), .ZN(n6723) );
  INV_X1 U8384 ( .A(n7020), .ZN(n6681) );
  AND2_X2 U8385 ( .A1(n6723), .A2(n6681), .ZN(n10455) );
  XNOR2_X1 U8386 ( .A(n6141), .B(n7028), .ZN(n6682) );
  NAND2_X1 U8387 ( .A1(n6682), .A2(n9297), .ZN(n9313) );
  AND2_X1 U8388 ( .A1(n6683), .A2(n10369), .ZN(n6684) );
  NAND2_X1 U8389 ( .A1(n6685), .A2(n6684), .ZN(n10418) );
  INV_X1 U8390 ( .A(n6686), .ZN(n8900) );
  NAND2_X1 U8391 ( .A1(n6686), .A2(n7164), .ZN(n6789) );
  INV_X1 U8392 ( .A(n6789), .ZN(n6687) );
  AOI21_X1 U8393 ( .B1(n8900), .B2(n6791), .A(n6687), .ZN(n7057) );
  NAND2_X1 U8394 ( .A1(n8183), .A2(n10387), .ZN(n6690) );
  NAND2_X1 U8395 ( .A1(n8774), .A2(n6690), .ZN(n8765) );
  INV_X1 U8396 ( .A(n8765), .ZN(n6692) );
  NAND2_X1 U8397 ( .A1(n8763), .A2(n4837), .ZN(n8740) );
  NAND2_X1 U8398 ( .A1(n6689), .A2(n8740), .ZN(n10365) );
  INV_X1 U8399 ( .A(n10365), .ZN(n9293) );
  NOR2_X1 U8400 ( .A1(n8900), .A2(n6690), .ZN(n6691) );
  AOI211_X1 U8401 ( .C1(n6692), .C2(n6688), .A(n9293), .B(n6691), .ZN(n6694)
         );
  OAI22_X1 U8402 ( .A1(n8183), .A2(n9309), .B1(n6893), .B2(n9311), .ZN(n6693)
         );
  NOR2_X1 U8403 ( .A1(n6694), .A2(n6693), .ZN(n7050) );
  NOR2_X1 U8404 ( .A1(n6788), .A2(n10387), .ZN(n7140) );
  INV_X1 U8405 ( .A(n7140), .ZN(n6697) );
  NAND2_X1 U8406 ( .A1(n10387), .A2(n6788), .ZN(n6696) );
  NAND2_X1 U8407 ( .A1(n6697), .A2(n6696), .ZN(n7053) );
  INV_X1 U8408 ( .A(n7053), .ZN(n6698) );
  AOI22_X1 U8409 ( .A1(n6698), .A2(n10411), .B1(n9437), .B2(n6788), .ZN(n6699)
         );
  OAI211_X1 U8410 ( .C1(n10426), .C2(n7057), .A(n7050), .B(n6699), .ZN(n6724)
         );
  NAND2_X1 U8411 ( .A1(n6724), .A2(n10455), .ZN(n6700) );
  OAI21_X1 U8412 ( .B1(n10455), .B2(n6526), .A(n6700), .ZN(P2_U3521) );
  INV_X1 U8413 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U8414 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6876), .B1(n6872), .B2(
        n10183), .ZN(n6707) );
  INV_X1 U8415 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U8416 ( .A1(n10304), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n10111), 
        .B2(n6701), .ZN(n10295) );
  INV_X1 U8417 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7432) );
  MUX2_X1 U8418 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7432), .S(n10272), .Z(n10263) );
  OR2_X1 U8419 ( .A1(n6712), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8420 ( .A1(n10263), .A2(n10262), .ZN(n10261) );
  NAND2_X1 U8421 ( .A1(n10272), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6704) );
  NOR2_X1 U8422 ( .A1(n10290), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6705) );
  AOI21_X1 U8423 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10290), .A(n6705), .ZN(
        n10277) );
  NAND2_X1 U8424 ( .A1(n10276), .A2(n10277), .ZN(n10275) );
  OAI21_X1 U8425 ( .B1(n10304), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10293), .ZN(
        n6706) );
  NAND2_X1 U8426 ( .A1(n6707), .A2(n6706), .ZN(n6870) );
  OAI21_X1 U8427 ( .B1(n6707), .B2(n6706), .A(n6870), .ZN(n6708) );
  INV_X1 U8428 ( .A(n6708), .ZN(n6722) );
  AND2_X1 U8429 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7516) );
  NOR2_X1 U8430 ( .A1(n10254), .A2(n6872), .ZN(n6709) );
  AOI211_X1 U8431 ( .C1(n10306), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7516), .B(
        n6709), .ZN(n6721) );
  NOR2_X1 U8432 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6876), .ZN(n6710) );
  AOI21_X1 U8433 ( .B1(n6876), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6710), .ZN(
        n6718) );
  INV_X1 U8434 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7406) );
  MUX2_X1 U8435 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7406), .S(n10272), .Z(n10265) );
  OR2_X1 U8436 ( .A1(n10272), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6713) );
  OR2_X1 U8437 ( .A1(n10290), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U8438 ( .A1(n10290), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U8439 ( .A1(n6715), .A2(n6714), .ZN(n10280) );
  NOR2_X1 U8440 ( .A1(n10281), .A2(n10280), .ZN(n10279) );
  NAND2_X1 U8441 ( .A1(n10304), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6716) );
  OAI21_X1 U8442 ( .B1(n10304), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6716), .ZN(
        n10298) );
  OAI21_X1 U8443 ( .B1(n6718), .B2(n6717), .A(n6875), .ZN(n6719) );
  NAND2_X1 U8444 ( .A1(n6719), .A2(n10284), .ZN(n6720) );
  OAI211_X1 U8445 ( .C1(n6722), .C2(n10288), .A(n6721), .B(n6720), .ZN(
        P1_U3252) );
  INV_X1 U8446 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6726) );
  NAND2_X1 U8447 ( .A1(n6724), .A2(n10444), .ZN(n6725) );
  OAI21_X1 U8448 ( .B1(n10444), .B2(n6726), .A(n6725), .ZN(P2_U3454) );
  AND2_X1 U8449 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6733) );
  INV_X1 U8450 ( .A(n6735), .ZN(n6728) );
  MUX2_X1 U8451 ( .A(n6729), .B(P2_REG1_REG_9__SCAN_IN), .S(n6860), .Z(n6730)
         );
  AOI211_X1 U8452 ( .C1(n6731), .C2(n6730), .A(n6854), .B(n8134), .ZN(n6732)
         );
  AOI211_X1 U8453 ( .C1(n10351), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6733), .B(
        n6732), .ZN(n6740) );
  OAI21_X1 U8454 ( .B1(n6735), .B2(n7248), .A(n6734), .ZN(n6738) );
  MUX2_X1 U8455 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6736), .S(n6860), .Z(n6737)
         );
  NAND2_X1 U8456 ( .A1(n6737), .A2(n6738), .ZN(n6861) );
  OAI211_X1 U8457 ( .C1(n6738), .C2(n6737), .A(n10350), .B(n6861), .ZN(n6739)
         );
  OAI211_X1 U8458 ( .C1(n7286), .C2(n6741), .A(n6740), .B(n6739), .ZN(P2_U3254) );
  INV_X1 U8459 ( .A(n8065), .ZN(n6764) );
  INV_X1 U8460 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6742) );
  NAND3_X1 U8461 ( .A1(n6744), .A2(n6743), .A3(n6742), .ZN(n6745) );
  OAI21_X1 U8462 ( .B1(n6746), .B2(n6745), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6747) );
  XNOR2_X1 U8463 ( .A(n6747), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9011) );
  AOI22_X1 U8464 ( .A1(n9011), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9471), .ZN(n6748) );
  OAI21_X1 U8465 ( .B1(n6764), .B2(n9469), .A(n6748), .ZN(P2_U3342) );
  INV_X1 U8466 ( .A(n6749), .ZN(n6751) );
  INV_X1 U8467 ( .A(n9694), .ZN(n9683) );
  OAI222_X1 U8468 ( .A1(n10100), .A2(n6750), .B1(n10081), .B2(n6751), .C1(
        n9683), .C2(P1_U3084), .ZN(P1_U3338) );
  INV_X1 U8469 ( .A(n8994), .ZN(n8983) );
  OAI222_X1 U8470 ( .A1(n7162), .A2(n6752), .B1(n9463), .B2(n6751), .C1(
        P2_U3152), .C2(n8983), .ZN(P2_U3343) );
  INV_X1 U8471 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9009) );
  INV_X1 U8472 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8171) );
  INV_X1 U8473 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8661) );
  INV_X1 U8474 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8694) );
  INV_X1 U8475 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U8476 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6758) );
  INV_X1 U8477 ( .A(n9103), .ZN(n6762) );
  INV_X1 U8478 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U8479 ( .A1(n8730), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U8480 ( .A1(n6174), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6759) );
  OAI211_X1 U8481 ( .C1(n4480), .C2(n9102), .A(n6760), .B(n6759), .ZN(n6761)
         );
  AOI21_X1 U8482 ( .B1(n6762), .B2(n8556), .A(n6761), .ZN(n9118) );
  NAND2_X1 U8483 ( .A1(n8936), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6763) );
  OAI21_X1 U8484 ( .B1(n9118), .B2(n8936), .A(n6763), .ZN(P2_U3581) );
  INV_X1 U8485 ( .A(n9712), .ZN(n9703) );
  OAI222_X1 U8486 ( .A1(n10100), .A2(n6765), .B1(n10090), .B2(n6764), .C1(
        P1_U3084), .C2(n9703), .ZN(P1_U3337) );
  NAND2_X1 U8487 ( .A1(n6767), .A2(n6766), .ZN(n6769) );
  OAI21_X1 U8488 ( .B1(n6771), .B2(n6844), .A(n6770), .ZN(n6772) );
  AOI222_X1 U8489 ( .A1(n10152), .A2(n6772), .B1(n9669), .B2(n10149), .C1(
        n9670), .C2(n10147), .ZN(n7214) );
  INV_X1 U8490 ( .A(n6773), .ZN(n6774) );
  NAND2_X1 U8491 ( .A1(n10161), .A2(n6774), .ZN(n10159) );
  INV_X1 U8492 ( .A(n10159), .ZN(n7011) );
  OAI22_X1 U8493 ( .A1(n10161), .A2(n6776), .B1(n6775), .B2(n9926), .ZN(n6781)
         );
  INV_X1 U8494 ( .A(n9963), .ZN(n7014) );
  NAND2_X1 U8495 ( .A1(n5949), .A2(n6851), .ZN(n6778) );
  NAND2_X1 U8496 ( .A1(n6778), .A2(n10032), .ZN(n6779) );
  OR2_X1 U8497 ( .A1(n6779), .A2(n6970), .ZN(n7213) );
  NOR2_X1 U8498 ( .A1(n7014), .A2(n7213), .ZN(n6780) );
  AOI211_X1 U8499 ( .C1(n7011), .C2(n5949), .A(n6781), .B(n6780), .ZN(n6786)
         );
  AND2_X1 U8500 ( .A1(n8485), .A2(n6782), .ZN(n6783) );
  NAND2_X1 U8501 ( .A1(n10161), .A2(n6783), .ZN(n9969) );
  OR2_X1 U8502 ( .A1(n9969), .A2(n7215), .ZN(n6785) );
  OAI211_X1 U8503 ( .C1(n10157), .C2(n7214), .A(n6786), .B(n6785), .ZN(
        P1_U3290) );
  NAND2_X1 U8504 ( .A1(n6893), .A2(n6787), .ZN(n8775) );
  NAND2_X1 U8505 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  NAND2_X1 U8506 ( .A1(n6893), .A2(n10393), .ZN(n6793) );
  NAND2_X1 U8507 ( .A1(n7134), .A2(n7027), .ZN(n8757) );
  INV_X1 U8508 ( .A(n7134), .ZN(n8944) );
  NAND2_X1 U8509 ( .A1(n8944), .A2(n7035), .ZN(n8780) );
  OAI21_X1 U8510 ( .B1(n6794), .B2(n8901), .A(n7037), .ZN(n7030) );
  INV_X1 U8511 ( .A(n7030), .ZN(n6800) );
  INV_X1 U8512 ( .A(n9313), .ZN(n7319) );
  OAI22_X1 U8513 ( .A1(n6893), .A2(n9309), .B1(n7110), .B2(n9311), .ZN(n6797)
         );
  INV_X1 U8514 ( .A(n8901), .ZN(n8768) );
  NAND3_X1 U8515 ( .A1(n7129), .A2(n8901), .A3(n8775), .ZN(n6795) );
  AOI21_X1 U8516 ( .B1(n7039), .B2(n6795), .A(n9293), .ZN(n6796) );
  AOI211_X1 U8517 ( .C1(n7030), .C2(n7319), .A(n6797), .B(n6796), .ZN(n7033)
         );
  AND2_X1 U8518 ( .A1(n7140), .A2(n10393), .ZN(n7138) );
  OAI211_X1 U8519 ( .C1(n7138), .C2(n7035), .A(n10411), .B(n7042), .ZN(n7024)
         );
  INV_X1 U8520 ( .A(n7024), .ZN(n6798) );
  AOI21_X1 U8521 ( .B1(n9437), .B2(n7027), .A(n6798), .ZN(n6799) );
  OAI211_X1 U8522 ( .C1(n6800), .C2(n10418), .A(n7033), .B(n6799), .ZN(n6802)
         );
  NAND2_X1 U8523 ( .A1(n6802), .A2(n10455), .ZN(n6801) );
  OAI21_X1 U8524 ( .B1(n10455), .B2(n6193), .A(n6801), .ZN(P2_U3523) );
  INV_X1 U8525 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8526 ( .A1(n6802), .A2(n10444), .ZN(n6803) );
  OAI21_X1 U8527 ( .B1(n10444), .B2(n6804), .A(n6803), .ZN(P2_U3460) );
  NAND2_X1 U8528 ( .A1(n6805), .A2(n6806), .ZN(n9570) );
  OAI21_X1 U8529 ( .B1(n6806), .B2(n6805), .A(n9570), .ZN(n6812) );
  INV_X1 U8530 ( .A(n9642), .ZN(n9622) );
  AOI22_X1 U8531 ( .A1(n6807), .A2(n9612), .B1(n9609), .B2(n9669), .ZN(n6810)
         );
  AOI21_X1 U8532 ( .B1(n9640), .B2(n5955), .A(n6808), .ZN(n6809) );
  OAI211_X1 U8533 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9622), .A(n6810), .B(
        n6809), .ZN(n6811) );
  AOI21_X1 U8534 ( .B1(n6812), .B2(n9607), .A(n6811), .ZN(n6813) );
  INV_X1 U8535 ( .A(n6813), .ZN(P1_U3216) );
  INV_X1 U8536 ( .A(n7332), .ZN(n7201) );
  AOI21_X1 U8537 ( .B1(n6815), .B2(n6814), .A(n4808), .ZN(n6817) );
  NAND2_X1 U8538 ( .A1(n6817), .A2(n6816), .ZN(n6821) );
  NOR2_X1 U8539 ( .A1(n8711), .A2(n7310), .ZN(n6819) );
  OAI22_X1 U8540 ( .A1(n8710), .A2(n7202), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6268), .ZN(n6818) );
  AOI211_X1 U8541 ( .C1(n8714), .C2(n10363), .A(n6819), .B(n6818), .ZN(n6820)
         );
  OAI211_X1 U8542 ( .C1(n7201), .C2(n8717), .A(n6821), .B(n6820), .ZN(P2_U3215) );
  NOR2_X1 U8543 ( .A1(n6822), .A2(n5957), .ZN(n7004) );
  AND2_X1 U8544 ( .A1(n6822), .A2(n5957), .ZN(n6823) );
  OAI21_X1 U8545 ( .B1(n7004), .B2(n6823), .A(n10152), .ZN(n6825) );
  AOI22_X1 U8546 ( .A1(n10149), .A2(n9666), .B1(n5955), .B2(n10147), .ZN(n6824) );
  AND2_X1 U8547 ( .A1(n6825), .A2(n6824), .ZN(n10325) );
  AND2_X1 U8548 ( .A1(n6828), .A2(n6827), .ZN(n10323) );
  INV_X1 U8549 ( .A(n9969), .ZN(n9933) );
  OAI21_X1 U8550 ( .B1(n6911), .B2(n10321), .A(n10032), .ZN(n6829) );
  OR2_X1 U8551 ( .A1(n6829), .A2(n7008), .ZN(n10320) );
  INV_X2 U8552 ( .A(n9926), .ZN(n10155) );
  AOI22_X1 U8553 ( .A1(n10157), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9548), .B2(
        n10155), .ZN(n6831) );
  NAND2_X1 U8554 ( .A1(n7011), .A2(n9545), .ZN(n6830) );
  OAI211_X1 U8555 ( .C1(n10320), .C2(n7014), .A(n6831), .B(n6830), .ZN(n6832)
         );
  AOI21_X1 U8556 ( .B1(n10323), .B2(n9933), .A(n6832), .ZN(n6833) );
  OAI21_X1 U8557 ( .B1(n10325), .B2(n10157), .A(n6833), .ZN(P1_U3286) );
  INV_X1 U8558 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7856) );
  INV_X1 U8559 ( .A(n8101), .ZN(n6836) );
  INV_X1 U8560 ( .A(n9728), .ZN(n9716) );
  OAI222_X1 U8561 ( .A1(n10086), .A2(n7856), .B1(n10090), .B2(n6836), .C1(
        P1_U3084), .C2(n9716), .ZN(P1_U3336) );
  NAND2_X1 U8562 ( .A1(n6083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6834) );
  MUX2_X1 U8563 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6834), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6835) );
  AND2_X1 U8564 ( .A1(n6835), .A2(n7082), .ZN(n9027) );
  INV_X1 U8565 ( .A(n9027), .ZN(n9006) );
  INV_X1 U8566 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8102) );
  OAI222_X1 U8567 ( .A1(P2_U3152), .A2(n9006), .B1(n9463), .B2(n6836), .C1(
        n8102), .C2(n7162), .ZN(P2_U3341) );
  INV_X1 U8568 ( .A(n6897), .ZN(n6837) );
  AOI211_X1 U8569 ( .C1(n6839), .C2(n6838), .A(n4808), .B(n6837), .ZN(n6843)
         );
  OR2_X1 U8570 ( .A1(n6840), .A2(P2_U3152), .ZN(n8186) );
  INV_X1 U8571 ( .A(n8186), .ZN(n6886) );
  OAI22_X1 U8572 ( .A1(n8717), .A2(n10393), .B1(n6886), .B2(n6176), .ZN(n6842)
         );
  OAI22_X1 U8573 ( .A1(n8696), .A2(n8189), .B1(n7134), .B2(n8711), .ZN(n6841)
         );
  OR3_X1 U8574 ( .A1(n6843), .A2(n6842), .A3(n6841), .ZN(P2_U3239) );
  AND2_X1 U8575 ( .A1(n9670), .A2(n6959), .ZN(n8355) );
  NOR2_X1 U8576 ( .A1(n6844), .A2(n8355), .ZN(n8448) );
  NAND2_X1 U8577 ( .A1(n8485), .A2(n6960), .ZN(n6845) );
  OR2_X1 U8578 ( .A1(n8448), .A2(n6845), .ZN(n6847) );
  NAND2_X1 U8579 ( .A1(n5950), .A2(n10149), .ZN(n6846) );
  AND2_X1 U8580 ( .A1(n6847), .A2(n6846), .ZN(n6958) );
  INV_X1 U8581 ( .A(n6848), .ZN(n6849) );
  NOR2_X1 U8582 ( .A1(n6960), .A2(n6849), .ZN(n6850) );
  OAI21_X1 U8583 ( .B1(n7011), .B2(n10143), .A(n6851), .ZN(n6853) );
  AOI22_X1 U8584 ( .A1(n10157), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10155), .ZN(n6852) );
  OAI211_X1 U8585 ( .C1(n10157), .C2(n6958), .A(n6853), .B(n6852), .ZN(
        P1_U3291) );
  NOR2_X1 U8586 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7815), .ZN(n6859) );
  MUX2_X1 U8587 ( .A(n6855), .B(P2_REG1_REG_10__SCAN_IN), .S(n7275), .Z(n6856)
         );
  NOR2_X1 U8588 ( .A1(n6857), .A2(n6856), .ZN(n7274) );
  AOI211_X1 U8589 ( .C1(n6857), .C2(n6856), .A(n7274), .B(n8134), .ZN(n6858)
         );
  AOI211_X1 U8590 ( .C1(n10351), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6859), .B(
        n6858), .ZN(n6867) );
  NAND2_X1 U8591 ( .A1(n6860), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6862) );
  NAND2_X1 U8592 ( .A1(n6862), .A2(n6861), .ZN(n6865) );
  MUX2_X1 U8593 ( .A(n7381), .B(P2_REG2_REG_10__SCAN_IN), .S(n7275), .Z(n6863)
         );
  INV_X1 U8594 ( .A(n6863), .ZN(n6864) );
  NAND2_X1 U8595 ( .A1(n6864), .A2(n6865), .ZN(n7267) );
  OAI211_X1 U8596 ( .C1(n6865), .C2(n6864), .A(n10350), .B(n7267), .ZN(n6866)
         );
  OAI211_X1 U8597 ( .C1(n7286), .C2(n6868), .A(n6867), .B(n6866), .ZN(P2_U3255) );
  INV_X1 U8598 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6869) );
  MUX2_X1 U8599 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6869), .S(n7097), .Z(n6874)
         );
  INV_X1 U8600 ( .A(n6870), .ZN(n6871) );
  AOI21_X1 U8601 ( .B1(n10183), .B2(n6872), .A(n6871), .ZN(n6873) );
  AOI21_X1 U8602 ( .B1(n6874), .B2(n6873), .A(n7096), .ZN(n6882) );
  NAND2_X1 U8603 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7987) );
  OAI21_X1 U8604 ( .B1(n10254), .B2(n7097), .A(n7987), .ZN(n6880) );
  XNOR2_X1 U8605 ( .A(n7101), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6878) );
  NOR2_X1 U8606 ( .A1(n6877), .A2(n6878), .ZN(n7100) );
  AOI211_X1 U8607 ( .C1(n6878), .C2(n6877), .A(n10296), .B(n7100), .ZN(n6879)
         );
  AOI211_X1 U8608 ( .C1(n10306), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6880), .B(
        n6879), .ZN(n6881) );
  OAI21_X1 U8609 ( .B1(n6882), .B2(n10288), .A(n6881), .ZN(P1_U3253) );
  OAI21_X1 U8610 ( .B1(n6885), .B2(n6884), .A(n6883), .ZN(n6889) );
  OAI22_X1 U8611 ( .A1(n8717), .A2(n6695), .B1(n6886), .B2(n7052), .ZN(n6888)
         );
  OAI22_X1 U8612 ( .A1(n8696), .A2(n8183), .B1(n6893), .B2(n8711), .ZN(n6887)
         );
  AOI211_X1 U8613 ( .C1(n8705), .C2(n6889), .A(n6888), .B(n6887), .ZN(n6890)
         );
  INV_X1 U8614 ( .A(n6890), .ZN(P2_U3224) );
  MUX2_X1 U8615 ( .A(P2_U3152), .B(n8630), .S(n7669), .Z(n6892) );
  OAI22_X1 U8616 ( .A1(n7035), .A2(n8717), .B1(n8711), .B2(n7110), .ZN(n6891)
         );
  AOI211_X1 U8617 ( .C1(n8714), .C2(n6181), .A(n6892), .B(n6891), .ZN(n6902)
         );
  NOR3_X1 U8618 ( .A1(n8502), .A2(n6894), .A3(n6893), .ZN(n6900) );
  INV_X1 U8619 ( .A(n6895), .ZN(n6896) );
  AOI21_X1 U8620 ( .B1(n6897), .B2(n6896), .A(n4808), .ZN(n6899) );
  OAI21_X1 U8621 ( .B1(n6900), .B2(n6899), .A(n6898), .ZN(n6901) );
  NAND2_X1 U8622 ( .A1(n6902), .A2(n6901), .ZN(P2_U3220) );
  INV_X1 U8623 ( .A(n10153), .ZN(n10131) );
  OAI21_X1 U8624 ( .B1(n6904), .B2(n8449), .A(n6903), .ZN(n7086) );
  OAI22_X1 U8625 ( .A1(n6965), .A2(n9957), .B1(n9577), .B2(n9959), .ZN(n6908)
         );
  INV_X1 U8626 ( .A(n8415), .ZN(n6905) );
  NOR2_X1 U8627 ( .A1(n8213), .A2(n6905), .ZN(n6906) );
  AOI211_X1 U8628 ( .C1(n8214), .C2(n8449), .A(n10128), .B(n6906), .ZN(n6907)
         );
  AOI211_X1 U8629 ( .C1(n10131), .C2(n7086), .A(n6908), .B(n6907), .ZN(n7089)
         );
  NOR2_X1 U8630 ( .A1(n6909), .A2(n9745), .ZN(n6910) );
  AND2_X1 U8631 ( .A1(n10161), .A2(n6910), .ZN(n10144) );
  INV_X1 U8632 ( .A(n7011), .ZN(n8122) );
  AOI21_X1 U8633 ( .B1(n9575), .B2(n7154), .A(n6911), .ZN(n7087) );
  NAND2_X1 U8634 ( .A1(n7087), .A2(n10143), .ZN(n6913) );
  AOI22_X1 U8635 ( .A1(n10157), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9580), .B2(
        n10155), .ZN(n6912) );
  OAI211_X1 U8636 ( .C1(n6914), .C2(n8122), .A(n6913), .B(n6912), .ZN(n6915)
         );
  AOI21_X1 U8637 ( .B1(n7086), .B2(n10144), .A(n6915), .ZN(n6916) );
  OAI21_X1 U8638 ( .B1(n7089), .B2(n10157), .A(n6916), .ZN(P1_U3287) );
  AND2_X1 U8639 ( .A1(n6982), .A2(n6917), .ZN(n6920) );
  OAI211_X1 U8640 ( .C1(n6920), .C2(n6919), .A(n6918), .B(n8705), .ZN(n6924)
         );
  INV_X1 U8641 ( .A(n7110), .ZN(n10361) );
  OAI22_X1 U8642 ( .A1(n8710), .A2(n10376), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6223), .ZN(n6922) );
  INV_X1 U8643 ( .A(n7113), .ZN(n10406) );
  INV_X1 U8644 ( .A(n10363), .ZN(n7197) );
  OAI22_X1 U8645 ( .A1(n10406), .A2(n8717), .B1(n8711), .B2(n7197), .ZN(n6921)
         );
  AOI211_X1 U8646 ( .C1(n8714), .C2(n10361), .A(n6922), .B(n6921), .ZN(n6923)
         );
  NAND2_X1 U8647 ( .A1(n6924), .A2(n6923), .ZN(P2_U3229) );
  OAI21_X1 U8648 ( .B1(n6927), .B2(n6926), .A(n6925), .ZN(n6928) );
  NAND2_X1 U8649 ( .A1(n6928), .A2(n9607), .ZN(n6935) );
  NAND2_X1 U8650 ( .A1(n9609), .A2(n9667), .ZN(n6930) );
  OR2_X1 U8651 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6929), .ZN(n10251) );
  OAI211_X1 U8652 ( .C1(n6931), .C2(n9578), .A(n6930), .B(n10251), .ZN(n6933)
         );
  INV_X1 U8653 ( .A(n9648), .ZN(n9634) );
  NOR2_X1 U8654 ( .A1(n9634), .A2(n7263), .ZN(n6932) );
  AOI211_X1 U8655 ( .C1(n7009), .C2(n9642), .A(n6933), .B(n6932), .ZN(n6934)
         );
  NAND2_X1 U8656 ( .A1(n6935), .A2(n6934), .ZN(P1_U3237) );
  OAI21_X1 U8657 ( .B1(n6937), .B2(n6918), .A(n6936), .ZN(n6946) );
  NOR3_X1 U8658 ( .A1(n8502), .A2(n6938), .A3(n6937), .ZN(n6939) );
  INV_X1 U8659 ( .A(n7120), .ZN(n8943) );
  OAI21_X1 U8660 ( .B1(n6939), .B2(n8714), .A(n8943), .ZN(n6944) );
  INV_X1 U8661 ( .A(n8711), .ZN(n8684) );
  INV_X1 U8662 ( .A(n7194), .ZN(n8942) );
  INV_X1 U8663 ( .A(n6940), .ZN(n6941) );
  OAI21_X1 U8664 ( .B1(n8710), .B2(n7125), .A(n6941), .ZN(n6942) );
  AOI21_X1 U8665 ( .B1(n8684), .B2(n8942), .A(n6942), .ZN(n6943) );
  OAI211_X1 U8666 ( .C1(n5000), .C2(n8717), .A(n6944), .B(n6943), .ZN(n6945)
         );
  AOI21_X1 U8667 ( .B1(n6946), .B2(n8705), .A(n6945), .ZN(n6947) );
  INV_X1 U8668 ( .A(n6947), .ZN(P2_U3241) );
  INV_X1 U8669 ( .A(n7311), .ZN(n10419) );
  INV_X1 U8670 ( .A(n6948), .ZN(n6949) );
  AOI21_X1 U8671 ( .B1(n6816), .B2(n6949), .A(n4808), .ZN(n6953) );
  NOR3_X1 U8672 ( .A1(n8502), .A2(n6950), .A3(n7194), .ZN(n6952) );
  OAI21_X1 U8673 ( .B1(n6953), .B2(n6952), .A(n6951), .ZN(n6957) );
  NOR2_X1 U8674 ( .A1(n8711), .A2(n7374), .ZN(n6955) );
  OAI22_X1 U8675 ( .A1(n8710), .A2(n7247), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7631), .ZN(n6954) );
  AOI211_X1 U8676 ( .C1(n8714), .C2(n8942), .A(n6955), .B(n6954), .ZN(n6956)
         );
  OAI211_X1 U8677 ( .C1(n10419), .C2(n8717), .A(n6957), .B(n6956), .ZN(
        P2_U3223) );
  INV_X1 U8678 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10194) );
  OAI21_X1 U8679 ( .B1(n6960), .B2(n6959), .A(n6958), .ZN(n6979) );
  NAND2_X1 U8680 ( .A1(n6979), .A2(n10344), .ZN(n6961) );
  OAI21_X1 U8681 ( .B1(n10344), .B2(n10194), .A(n6961), .ZN(P1_U3523) );
  INV_X1 U8682 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U8683 ( .A1(n6962), .A2(n8446), .ZN(n6963) );
  NAND2_X1 U8684 ( .A1(n6964), .A2(n6963), .ZN(n7065) );
  INV_X1 U8685 ( .A(n7065), .ZN(n6973) );
  OAI22_X1 U8686 ( .A1(n8357), .A2(n9957), .B1(n6965), .B2(n9959), .ZN(n6969)
         );
  INV_X1 U8687 ( .A(n6966), .ZN(n8359) );
  XNOR2_X1 U8688 ( .A(n8359), .B(n8446), .ZN(n6967) );
  NOR2_X1 U8689 ( .A1(n6967), .A2(n10128), .ZN(n6968) );
  AOI211_X1 U8690 ( .C1(n10131), .C2(n7065), .A(n6969), .B(n6968), .ZN(n7062)
         );
  OR2_X1 U8691 ( .A1(n6970), .A2(n7061), .ZN(n6971) );
  AND2_X1 U8692 ( .A1(n7153), .A2(n6971), .ZN(n7058) );
  AOI22_X1 U8693 ( .A1(n7058), .A2(n10032), .B1(n10031), .B2(n9611), .ZN(n6972) );
  OAI211_X1 U8694 ( .C1(n6973), .C2(n10102), .A(n7062), .B(n6972), .ZN(n6976)
         );
  NAND2_X1 U8695 ( .A1(n6976), .A2(n10344), .ZN(n6974) );
  OAI21_X1 U8696 ( .B1(n10344), .B2(n6975), .A(n6974), .ZN(P1_U3525) );
  INV_X1 U8697 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8698 ( .A1(n6976), .A2(n10336), .ZN(n6977) );
  OAI21_X1 U8699 ( .B1(n10336), .B2(n6978), .A(n6977), .ZN(P1_U3460) );
  INV_X1 U8700 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U8701 ( .A1(n6979), .A2(n10336), .ZN(n6980) );
  OAI21_X1 U8702 ( .B1(n10336), .B2(n6981), .A(n6980), .ZN(P1_U3454) );
  OAI21_X1 U8703 ( .B1(n6983), .B2(n6898), .A(n6982), .ZN(n6991) );
  INV_X1 U8704 ( .A(n8502), .ZN(n8700) );
  INV_X1 U8705 ( .A(n6983), .ZN(n6985) );
  NAND3_X1 U8706 ( .A1(n8700), .A2(n6985), .A3(n6984), .ZN(n6986) );
  AOI21_X1 U8707 ( .B1(n6986), .B2(n8696), .A(n7134), .ZN(n6990) );
  AOI22_X1 U8708 ( .A1(n8684), .A2(n8943), .B1(n7046), .B2(n8699), .ZN(n6988)
         );
  OAI211_X1 U8709 ( .C1(n7041), .C2(n8710), .A(n6988), .B(n6987), .ZN(n6989)
         );
  AOI211_X1 U8710 ( .C1(n8705), .C2(n6991), .A(n6990), .B(n6989), .ZN(n6992)
         );
  INV_X1 U8711 ( .A(n6992), .ZN(P2_U3232) );
  NAND2_X1 U8712 ( .A1(n4559), .A2(n6994), .ZN(n6995) );
  XNOR2_X1 U8713 ( .A(n6993), .B(n6995), .ZN(n7002) );
  NAND2_X1 U8714 ( .A1(n9609), .A2(n9666), .ZN(n6998) );
  INV_X1 U8715 ( .A(n6996), .ZN(n6997) );
  OAI211_X1 U8716 ( .C1(n7069), .C2(n9578), .A(n6998), .B(n6997), .ZN(n7000)
         );
  NOR2_X1 U8717 ( .A1(n9634), .A2(n7220), .ZN(n6999) );
  AOI211_X1 U8718 ( .C1(n7076), .C2(n9642), .A(n7000), .B(n6999), .ZN(n7001)
         );
  OAI21_X1 U8719 ( .B1(n7002), .B2(n9651), .A(n7001), .ZN(P1_U3211) );
  INV_X1 U8720 ( .A(n8420), .ZN(n7003) );
  NOR2_X1 U8721 ( .A1(n7004), .A2(n7003), .ZN(n7005) );
  XNOR2_X1 U8722 ( .A(n7005), .B(n8219), .ZN(n7006) );
  AOI222_X1 U8723 ( .A1(n10152), .A2(n7006), .B1(n9665), .B2(n10149), .C1(
        n9667), .C2(n10147), .ZN(n7226) );
  OAI21_X1 U8724 ( .B1(n4555), .B2(n8219), .A(n7007), .ZN(n7224) );
  OAI211_X1 U8725 ( .C1(n7008), .C2(n7263), .A(n10032), .B(n7074), .ZN(n7225)
         );
  AOI22_X1 U8726 ( .A1(n10157), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7009), .B2(
        n10155), .ZN(n7013) );
  NAND2_X1 U8727 ( .A1(n7011), .A2(n7010), .ZN(n7012) );
  OAI211_X1 U8728 ( .C1(n7225), .C2(n7014), .A(n7013), .B(n7012), .ZN(n7015)
         );
  AOI21_X1 U8729 ( .B1(n7224), .B2(n9933), .A(n7015), .ZN(n7016) );
  OAI21_X1 U8730 ( .B1(n7226), .B2(n10157), .A(n7016), .ZN(P1_U3285) );
  INV_X1 U8731 ( .A(n8166), .ZN(n7085) );
  AOI22_X1 U8732 ( .A1(n9740), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10079), .ZN(n7017) );
  OAI21_X1 U8733 ( .B1(n7085), .B2(n10081), .A(n7017), .ZN(P1_U3335) );
  INV_X1 U8734 ( .A(n7018), .ZN(n7019) );
  NAND4_X1 U8735 ( .A1(n7021), .A2(P2_STATE_REG_SCAN_IN), .A3(n7020), .A4(
        n7019), .ZN(n7023) );
  INV_X2 U8736 ( .A(n10357), .ZN(n10370) );
  NOR2_X1 U8737 ( .A1(n10370), .A2(n6551), .ZN(n7026) );
  OR2_X1 U8738 ( .A1(n7023), .A2(n10369), .ZN(n7200) );
  OAI22_X1 U8739 ( .A1(n7200), .A2(n7024), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10375), .ZN(n7025) );
  AOI211_X1 U8740 ( .C1(n9325), .C2(n7027), .A(n7026), .B(n7025), .ZN(n7032)
         );
  NOR2_X1 U8741 ( .A1(n7028), .A2(n9297), .ZN(n7029) );
  NAND2_X1 U8742 ( .A1(n10370), .A2(n7029), .ZN(n9328) );
  INV_X1 U8743 ( .A(n9328), .ZN(n7326) );
  NAND2_X1 U8744 ( .A1(n7030), .A2(n7326), .ZN(n7031) );
  OAI211_X1 U8745 ( .C1(n7033), .C2(n10357), .A(n7032), .B(n7031), .ZN(
        P2_U3293) );
  NAND2_X1 U8746 ( .A1(n10370), .A2(n7319), .ZN(n7034) );
  NAND2_X1 U8747 ( .A1(n7134), .A2(n7035), .ZN(n7036) );
  NAND2_X1 U8748 ( .A1(n7110), .A2(n7046), .ZN(n8758) );
  NAND2_X1 U8749 ( .A1(n10361), .A2(n10398), .ZN(n8781) );
  NAND2_X1 U8750 ( .A1(n8758), .A2(n8781), .ZN(n8902) );
  OAI21_X1 U8751 ( .B1(n7038), .B2(n8902), .A(n7112), .ZN(n10402) );
  INV_X1 U8752 ( .A(n10402), .ZN(n7049) );
  XNOR2_X1 U8753 ( .A(n7115), .B(n8902), .ZN(n7040) );
  OAI222_X1 U8754 ( .A1(n9309), .A2(n7134), .B1(n9311), .B2(n7120), .C1(n7040), 
        .C2(n9293), .ZN(n10400) );
  NAND2_X1 U8755 ( .A1(n10400), .A2(n10370), .ZN(n7048) );
  OAI22_X1 U8756 ( .A1(n10375), .A2(n7041), .B1(n6555), .B2(n10370), .ZN(n7045) );
  AND2_X1 U8757 ( .A1(n7042), .A2(n7046), .ZN(n7043) );
  OR2_X1 U8758 ( .A1(n7043), .A2(n10367), .ZN(n10399) );
  NOR2_X1 U8759 ( .A1(n10399), .A2(n9321), .ZN(n7044) );
  AOI211_X1 U8760 ( .C1(n9325), .C2(n7046), .A(n7045), .B(n7044), .ZN(n7047)
         );
  OAI211_X1 U8761 ( .C1(n9349), .C2(n7049), .A(n7048), .B(n7047), .ZN(P2_U3292) );
  MUX2_X1 U8762 ( .A(n7051), .B(n7050), .S(n10370), .Z(n7056) );
  OAI22_X1 U8763 ( .A1(n9321), .A2(n7053), .B1(n7052), .B2(n10375), .ZN(n7054)
         );
  AOI21_X1 U8764 ( .B1(n9325), .B2(n6788), .A(n7054), .ZN(n7055) );
  OAI211_X1 U8765 ( .C1(n9349), .C2(n7057), .A(n7056), .B(n7055), .ZN(P2_U3295) );
  AOI22_X1 U8766 ( .A1(n10157), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10155), .ZN(n7060) );
  NAND2_X1 U8767 ( .A1(n10143), .A2(n7058), .ZN(n7059) );
  OAI211_X1 U8768 ( .C1(n7061), .C2(n10159), .A(n7060), .B(n7059), .ZN(n7064)
         );
  NOR2_X1 U8769 ( .A1(n7062), .A2(n10157), .ZN(n7063) );
  AOI211_X1 U8770 ( .C1(n10144), .C2(n7065), .A(n7064), .B(n7063), .ZN(n7066)
         );
  INV_X1 U8771 ( .A(n7066), .ZN(P1_U3289) );
  XNOR2_X1 U8772 ( .A(n7067), .B(n7071), .ZN(n7068) );
  OAI222_X1 U8773 ( .A1(n9959), .A2(n7069), .B1(n9957), .B2(n9546), .C1(n10128), .C2(n7068), .ZN(n7207) );
  INV_X1 U8774 ( .A(n7207), .ZN(n7081) );
  OAI21_X1 U8775 ( .B1(n7072), .B2(n7071), .A(n7070), .ZN(n7209) );
  INV_X1 U8776 ( .A(n7073), .ZN(n7408) );
  AOI211_X1 U8777 ( .C1(n7075), .C2(n7074), .A(n10313), .B(n7073), .ZN(n7208)
         );
  NAND2_X1 U8778 ( .A1(n7208), .A2(n9963), .ZN(n7078) );
  AOI22_X1 U8779 ( .A1(n10157), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7076), .B2(
        n10155), .ZN(n7077) );
  OAI211_X1 U8780 ( .C1(n7220), .C2(n8122), .A(n7078), .B(n7077), .ZN(n7079)
         );
  AOI21_X1 U8781 ( .B1(n7209), .B2(n9933), .A(n7079), .ZN(n7080) );
  OAI21_X1 U8782 ( .B1(n7081), .B2(n10157), .A(n7080), .ZN(P1_U3284) );
  INV_X1 U8783 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U8784 ( .A1(n7082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7084) );
  XNOR2_X1 U8785 ( .A(n7084), .B(n7083), .ZN(n9042) );
  OAI222_X1 U8786 ( .A1(n7162), .A2(n8167), .B1(n9463), .B2(n7085), .C1(
        P2_U3152), .C2(n9042), .ZN(P2_U3340) );
  INV_X1 U8787 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7092) );
  INV_X1 U8788 ( .A(n7086), .ZN(n7090) );
  AOI22_X1 U8789 ( .A1(n7087), .A2(n10032), .B1(n10031), .B2(n9575), .ZN(n7088) );
  OAI211_X1 U8790 ( .C1(n7090), .C2(n10102), .A(n7089), .B(n7088), .ZN(n7093)
         );
  NAND2_X1 U8791 ( .A1(n7093), .A2(n10336), .ZN(n7091) );
  OAI21_X1 U8792 ( .B1(n10336), .B2(n7092), .A(n7091), .ZN(P1_U3466) );
  INV_X1 U8793 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U8794 ( .A1(n7093), .A2(n10344), .ZN(n7094) );
  OAI21_X1 U8795 ( .B1(n10344), .B2(n7095), .A(n7094), .ZN(P1_U3527) );
  INV_X1 U8796 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10177) );
  MUX2_X1 U8797 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10177), .S(n7484), .Z(n7099) );
  AOI21_X1 U8798 ( .B1(n6869), .B2(n7097), .A(n7096), .ZN(n7098) );
  NOR2_X1 U8799 ( .A1(n7098), .A2(n7099), .ZN(n7483) );
  AOI21_X1 U8800 ( .B1(n7099), .B2(n7098), .A(n7483), .ZN(n7109) );
  NAND2_X1 U8801 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8002) );
  OAI21_X1 U8802 ( .B1(n10254), .B2(n7484), .A(n8002), .ZN(n7107) );
  INV_X1 U8803 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7102) );
  MUX2_X1 U8804 ( .A(n7102), .B(P1_REG2_REG_13__SCAN_IN), .S(n7484), .Z(n7103)
         );
  INV_X1 U8805 ( .A(n7103), .ZN(n7104) );
  AOI211_X1 U8806 ( .C1(n7105), .C2(n7104), .A(n10296), .B(n7487), .ZN(n7106)
         );
  AOI211_X1 U8807 ( .C1(n10306), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7107), .B(
        n7106), .ZN(n7108) );
  OAI21_X1 U8808 ( .B1(n7109), .B2(n10288), .A(n7108), .ZN(P1_U3254) );
  NAND2_X1 U8809 ( .A1(n7110), .A2(n10398), .ZN(n7111) );
  NAND2_X1 U8810 ( .A1(n7120), .A2(n7113), .ZN(n8759) );
  NAND2_X1 U8811 ( .A1(n8943), .A2(n10406), .ZN(n8783) );
  NAND2_X1 U8812 ( .A1(n8759), .A2(n8783), .ZN(n10355) );
  NAND2_X1 U8813 ( .A1(n7120), .A2(n10406), .ZN(n7114) );
  NAND2_X1 U8814 ( .A1(n7197), .A2(n10410), .ZN(n8790) );
  NAND2_X1 U8815 ( .A1(n5000), .A2(n10363), .ZN(n8782) );
  AND2_X1 U8816 ( .A1(n8790), .A2(n8782), .ZN(n8905) );
  XNOR2_X1 U8817 ( .A(n7193), .B(n8905), .ZN(n10415) );
  INV_X1 U8818 ( .A(n10355), .ZN(n10359) );
  NAND2_X1 U8819 ( .A1(n7116), .A2(n8905), .ZN(n7240) );
  INV_X1 U8820 ( .A(n8905), .ZN(n7118) );
  NAND3_X1 U8821 ( .A1(n7117), .A2(n8759), .A3(n7118), .ZN(n7119) );
  NAND2_X1 U8822 ( .A1(n7240), .A2(n7119), .ZN(n7122) );
  OAI22_X1 U8823 ( .A1(n7120), .A2(n9309), .B1(n7194), .B2(n9311), .ZN(n7121)
         );
  AOI21_X1 U8824 ( .B1(n7122), .B2(n10365), .A(n7121), .ZN(n10414) );
  MUX2_X1 U8825 ( .A(n7123), .B(n10414), .S(n10370), .Z(n7128) );
  INV_X1 U8826 ( .A(n7199), .ZN(n7124) );
  AOI21_X1 U8827 ( .B1(n10410), .B2(n10366), .A(n7124), .ZN(n10412) );
  OAI22_X1 U8828 ( .A1(n9338), .A2(n5000), .B1(n10375), .B2(n7125), .ZN(n7126)
         );
  AOI21_X1 U8829 ( .B1(n10412), .B2(n9347), .A(n7126), .ZN(n7127) );
  OAI211_X1 U8830 ( .C1(n9349), .C2(n10415), .A(n7128), .B(n7127), .ZN(
        P2_U3290) );
  INV_X1 U8831 ( .A(n10375), .ZN(n9335) );
  INV_X1 U8832 ( .A(n7129), .ZN(n7130) );
  AOI21_X1 U8833 ( .B1(n7132), .B2(n7131), .A(n7130), .ZN(n7133) );
  OAI222_X1 U8834 ( .A1(n9309), .A2(n8189), .B1(n9311), .B2(n7134), .C1(n9293), 
        .C2(n7133), .ZN(n10394) );
  AOI21_X1 U8835 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n9335), .A(n10394), .ZN(
        n7135) );
  MUX2_X1 U8836 ( .A(n7136), .B(n7135), .S(n10370), .Z(n7143) );
  XNOR2_X1 U8837 ( .A(n7137), .B(n8899), .ZN(n10396) );
  INV_X1 U8838 ( .A(n9349), .ZN(n10358) );
  INV_X1 U8839 ( .A(n7138), .ZN(n7139) );
  OAI211_X1 U8840 ( .C1(n10393), .C2(n7140), .A(n7139), .B(n10411), .ZN(n10392) );
  OAI22_X1 U8841 ( .A1(n9338), .A2(n10393), .B1(n10392), .B2(n7200), .ZN(n7141) );
  AOI21_X1 U8842 ( .B1(n10396), .B2(n10358), .A(n7141), .ZN(n7142) );
  NAND2_X1 U8843 ( .A1(n7143), .A2(n7142), .ZN(P2_U3294) );
  XNOR2_X1 U8844 ( .A(n7144), .B(n7146), .ZN(n7152) );
  OAI21_X1 U8845 ( .B1(n7147), .B2(n7146), .A(n7145), .ZN(n10317) );
  OAI22_X1 U8846 ( .A1(n7149), .A2(n9957), .B1(n7148), .B2(n9959), .ZN(n7150)
         );
  AOI21_X1 U8847 ( .B1(n10317), .B2(n10131), .A(n7150), .ZN(n7151) );
  OAI21_X1 U8848 ( .B1(n10128), .B2(n7152), .A(n7151), .ZN(n10315) );
  INV_X1 U8849 ( .A(n10315), .ZN(n7161) );
  INV_X1 U8850 ( .A(n10143), .ZN(n8120) );
  INV_X1 U8851 ( .A(n7153), .ZN(n7155) );
  OAI21_X1 U8852 ( .B1(n7155), .B2(n10312), .A(n7154), .ZN(n10314) );
  NOR2_X1 U8853 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n9926), .ZN(n7157) );
  NOR2_X1 U8854 ( .A1(n8122), .A2(n10312), .ZN(n7156) );
  AOI211_X1 U8855 ( .C1(n10157), .C2(P1_REG2_REG_3__SCAN_IN), .A(n7157), .B(
        n7156), .ZN(n7158) );
  OAI21_X1 U8856 ( .B1(n8120), .B2(n10314), .A(n7158), .ZN(n7159) );
  AOI21_X1 U8857 ( .B1(n10144), .B2(n10317), .A(n7159), .ZN(n7160) );
  OAI21_X1 U8858 ( .B1(n10157), .B2(n7161), .A(n7160), .ZN(P1_U3288) );
  INV_X1 U8859 ( .A(n8508), .ZN(n7163) );
  OAI222_X1 U8860 ( .A1(n7162), .A2(n8510), .B1(n9469), .B2(n7163), .C1(n9297), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8861 ( .A1(P1_U3084), .A2(n9745), .B1(n10090), .B2(n7163), .C1(
        n7841), .C2(n10100), .ZN(P1_U3334) );
  OAI21_X1 U8862 ( .B1(n8945), .B2(n10387), .A(n7164), .ZN(n8898) );
  INV_X1 U8863 ( .A(n8898), .ZN(n10388) );
  AOI22_X1 U8864 ( .A1(n10388), .A2(n10365), .B1(n10362), .B2(n6790), .ZN(
        n10390) );
  OAI22_X1 U8865 ( .A1(n10390), .A2(n10357), .B1(n6159), .B2(n10375), .ZN(
        n7166) );
  AOI21_X1 U8866 ( .B1(n9338), .B2(n9321), .A(n8762), .ZN(n7165) );
  AOI211_X1 U8867 ( .C1(n10357), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7166), .B(
        n7165), .ZN(n7167) );
  OAI21_X1 U8868 ( .B1(n9349), .B2(n8898), .A(n7167), .ZN(P2_U3296) );
  INV_X1 U8869 ( .A(n6951), .ZN(n7170) );
  NOR3_X1 U8870 ( .A1(n8502), .A2(n7168), .A3(n7310), .ZN(n7169) );
  AOI21_X1 U8871 ( .B1(n7170), .B2(n8705), .A(n7169), .ZN(n7182) );
  OR2_X1 U8872 ( .A1(n7923), .A2(n9311), .ZN(n7172) );
  OR2_X1 U8873 ( .A1(n7310), .A2(n9309), .ZN(n7171) );
  NAND2_X1 U8874 ( .A1(n7172), .A2(n7171), .ZN(n7317) );
  NAND2_X1 U8875 ( .A1(n8674), .A2(n7317), .ZN(n7175) );
  INV_X1 U8876 ( .A(n7323), .ZN(n7173) );
  NAND2_X1 U8877 ( .A1(n8630), .A2(n7173), .ZN(n7174) );
  OAI211_X1 U8878 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7176), .A(n7175), .B(n7174), .ZN(n7179) );
  NOR2_X1 U8879 ( .A1(n7177), .A2(n4808), .ZN(n7178) );
  AOI211_X1 U8880 ( .C1(n7460), .C2(n8699), .A(n7179), .B(n7178), .ZN(n7180)
         );
  OAI21_X1 U8881 ( .B1(n7182), .B2(n7181), .A(n7180), .ZN(P2_U3233) );
  AOI21_X1 U8882 ( .B1(n7184), .B2(n7183), .A(n4808), .ZN(n7186) );
  NAND2_X1 U8883 ( .A1(n7186), .A2(n7185), .ZN(n7190) );
  NOR2_X1 U8884 ( .A1(n8711), .A2(n7955), .ZN(n7188) );
  OAI22_X1 U8885 ( .A1(n8710), .A2(n7380), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7815), .ZN(n7187) );
  AOI211_X1 U8886 ( .C1(n8714), .C2(n4769), .A(n7188), .B(n7187), .ZN(n7189)
         );
  OAI211_X1 U8887 ( .C1(n4989), .C2(n8717), .A(n7190), .B(n7189), .ZN(P2_U3219) );
  NOR2_X1 U8888 ( .A1(n10363), .A2(n10410), .ZN(n7192) );
  NAND2_X1 U8889 ( .A1(n10363), .A2(n10410), .ZN(n7191) );
  OAI21_X1 U8890 ( .B1(n7193), .B2(n7192), .A(n7191), .ZN(n7231) );
  OR2_X1 U8891 ( .A1(n7332), .A2(n7194), .ZN(n8791) );
  NAND2_X1 U8892 ( .A1(n7332), .A2(n7194), .ZN(n8805) );
  INV_X1 U8893 ( .A(n8904), .ZN(n7238) );
  XNOR2_X1 U8894 ( .A(n7231), .B(n7238), .ZN(n7334) );
  NAND2_X1 U8895 ( .A1(n7240), .A2(n8790), .ZN(n7195) );
  XNOR2_X1 U8896 ( .A(n7195), .B(n7238), .ZN(n7196) );
  OAI222_X1 U8897 ( .A1(n9309), .A2(n7197), .B1(n9311), .B2(n7310), .C1(n7196), 
        .C2(n9293), .ZN(n7330) );
  NAND2_X1 U8898 ( .A1(n7330), .A2(n10370), .ZN(n7206) );
  INV_X1 U8899 ( .A(n7249), .ZN(n7198) );
  AOI211_X1 U8900 ( .C1(n7332), .C2(n7199), .A(n10436), .B(n7198), .ZN(n7331)
         );
  INV_X1 U8901 ( .A(n7200), .ZN(n9182) );
  NOR2_X1 U8902 ( .A1(n9338), .A2(n7201), .ZN(n7204) );
  OAI22_X1 U8903 ( .A1(n10370), .A2(n6575), .B1(n7202), .B2(n10375), .ZN(n7203) );
  AOI211_X1 U8904 ( .C1(n7331), .C2(n9182), .A(n7204), .B(n7203), .ZN(n7205)
         );
  OAI211_X1 U8905 ( .C1(n9349), .C2(n7334), .A(n7206), .B(n7205), .ZN(P2_U3289) );
  AOI211_X1 U8906 ( .C1(n10332), .C2(n7209), .A(n7208), .B(n7207), .ZN(n7223)
         );
  INV_X1 U8907 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7210) );
  OAI22_X1 U8908 ( .A1(n10076), .A2(n7220), .B1(n10336), .B2(n7210), .ZN(n7211) );
  INV_X1 U8909 ( .A(n7211), .ZN(n7212) );
  OAI21_X1 U8910 ( .B1(n7223), .B2(n10334), .A(n7212), .ZN(P1_U3475) );
  OAI211_X1 U8911 ( .C1(n10036), .C2(n7215), .A(n7214), .B(n7213), .ZN(n7259)
         );
  INV_X1 U8912 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7216) );
  OAI22_X1 U8913 ( .A1(n10076), .A2(n7257), .B1(n10336), .B2(n7216), .ZN(n7217) );
  AOI21_X1 U8914 ( .B1(n7259), .B2(n10336), .A(n7217), .ZN(n7218) );
  INV_X1 U8915 ( .A(n7218), .ZN(P1_U3457) );
  OAI22_X1 U8916 ( .A1(n10042), .A2(n7220), .B1(n10344), .B2(n7219), .ZN(n7221) );
  INV_X1 U8917 ( .A(n7221), .ZN(n7222) );
  OAI21_X1 U8918 ( .B1(n7223), .B2(n10341), .A(n7222), .ZN(P1_U3530) );
  INV_X1 U8919 ( .A(n7224), .ZN(n7227) );
  OAI211_X1 U8920 ( .C1(n10036), .C2(n7227), .A(n7226), .B(n7225), .ZN(n7265)
         );
  INV_X1 U8921 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7228) );
  OAI22_X1 U8922 ( .A1(n10076), .A2(n7263), .B1(n10336), .B2(n7228), .ZN(n7229) );
  AOI21_X1 U8923 ( .B1(n7265), .B2(n10336), .A(n7229), .ZN(n7230) );
  INV_X1 U8924 ( .A(n7230), .ZN(P1_U3472) );
  OR2_X1 U8925 ( .A1(n7332), .A2(n8942), .ZN(n7232) );
  OR2_X1 U8926 ( .A1(n7311), .A2(n7310), .ZN(n8794) );
  NAND2_X1 U8927 ( .A1(n7311), .A2(n7310), .ZN(n8792) );
  NAND2_X1 U8928 ( .A1(n7235), .A2(n8806), .ZN(n7236) );
  INV_X1 U8929 ( .A(n10423), .ZN(n7255) );
  INV_X1 U8930 ( .A(n8790), .ZN(n7237) );
  NOR2_X1 U8931 ( .A1(n7238), .A2(n7237), .ZN(n7239) );
  NAND2_X1 U8932 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  INV_X1 U8933 ( .A(n7314), .ZN(n7242) );
  AOI21_X1 U8934 ( .B1(n7233), .B2(n7243), .A(n7242), .ZN(n7246) );
  NAND2_X1 U8935 ( .A1(n10423), .A2(n7319), .ZN(n7245) );
  AOI22_X1 U8936 ( .A1(n10360), .A2(n8942), .B1(n4769), .B2(n10362), .ZN(n7244) );
  OAI211_X1 U8937 ( .C1(n7246), .C2(n9293), .A(n7245), .B(n7244), .ZN(n10421)
         );
  NAND2_X1 U8938 ( .A1(n10421), .A2(n10370), .ZN(n7254) );
  OAI22_X1 U8939 ( .A1(n10370), .A2(n7248), .B1(n7247), .B2(n10375), .ZN(n7252) );
  AND2_X1 U8940 ( .A1(n7249), .A2(n7311), .ZN(n7250) );
  NOR2_X1 U8941 ( .A1(n7249), .A2(n7311), .ZN(n7320) );
  OR2_X1 U8942 ( .A1(n7250), .A2(n7320), .ZN(n10420) );
  NOR2_X1 U8943 ( .A1(n10420), .A2(n9321), .ZN(n7251) );
  AOI211_X1 U8944 ( .C1(n9325), .C2(n7311), .A(n7252), .B(n7251), .ZN(n7253)
         );
  OAI211_X1 U8945 ( .C1(n7255), .C2(n9328), .A(n7254), .B(n7253), .ZN(P2_U3288) );
  OAI22_X1 U8946 ( .A1(n10042), .A2(n7257), .B1(n10344), .B2(n7256), .ZN(n7258) );
  AOI21_X1 U8947 ( .B1(n7259), .B2(n10344), .A(n7258), .ZN(n7260) );
  INV_X1 U8948 ( .A(n7260), .ZN(P1_U3524) );
  INV_X1 U8949 ( .A(n8520), .ZN(n7297) );
  AOI22_X1 U8950 ( .A1(n4837), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n9471), .ZN(n7261) );
  OAI21_X1 U8951 ( .B1(n7297), .B2(n9463), .A(n7261), .ZN(P2_U3338) );
  INV_X1 U8952 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7262) );
  OAI22_X1 U8953 ( .A1(n10042), .A2(n7263), .B1(n10344), .B2(n7262), .ZN(n7264) );
  AOI21_X1 U8954 ( .B1(n7265), .B2(n10344), .A(n7264), .ZN(n7266) );
  INV_X1 U8955 ( .A(n7266), .ZN(P1_U3529) );
  NOR2_X1 U8956 ( .A1(n8973), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7270) );
  NAND2_X1 U8957 ( .A1(n7275), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U8958 ( .A1(n7268), .A2(n7267), .ZN(n8970) );
  MUX2_X1 U8959 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6340), .S(n8973), .Z(n7269)
         );
  INV_X1 U8960 ( .A(n7269), .ZN(n8969) );
  NOR2_X1 U8961 ( .A1(n8970), .A2(n8969), .ZN(n8968) );
  NOR2_X1 U8962 ( .A1(n7270), .A2(n8968), .ZN(n7273) );
  MUX2_X1 U8963 ( .A(n7958), .B(P2_REG2_REG_12__SCAN_IN), .S(n7344), .Z(n7271)
         );
  INV_X1 U8964 ( .A(n7271), .ZN(n7272) );
  NAND2_X1 U8965 ( .A1(n7272), .A2(n7273), .ZN(n7339) );
  OAI211_X1 U8966 ( .C1(n7273), .C2(n7272), .A(n10350), .B(n7339), .ZN(n7284)
         );
  MUX2_X1 U8967 ( .A(n7276), .B(P2_REG1_REG_11__SCAN_IN), .S(n8973), .Z(n8976)
         );
  MUX2_X1 U8968 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7277), .S(n7344), .Z(n7278)
         );
  OAI21_X1 U8969 ( .B1(n7279), .B2(n7278), .A(n7343), .ZN(n7282) );
  NOR2_X1 U8970 ( .A1(n7767), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7420) );
  INV_X1 U8971 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7280) );
  NOR2_X1 U8972 ( .A1(n9056), .A2(n7280), .ZN(n7281) );
  AOI211_X1 U8973 ( .C1(n10349), .C2(n7282), .A(n7420), .B(n7281), .ZN(n7283)
         );
  OAI211_X1 U8974 ( .C1(n7286), .C2(n7285), .A(n7284), .B(n7283), .ZN(P2_U3257) );
  INV_X1 U8975 ( .A(n7289), .ZN(n7287) );
  AOI21_X1 U8976 ( .B1(n7185), .B2(n7287), .A(n4808), .ZN(n7292) );
  NOR3_X1 U8977 ( .A1(n7288), .A2(n7923), .A3(n8502), .ZN(n7291) );
  NAND2_X1 U8978 ( .A1(n7290), .A2(n7289), .ZN(n7437) );
  OAI21_X1 U8979 ( .B1(n7292), .B2(n7291), .A(n7437), .ZN(n7296) );
  OAI22_X1 U8980 ( .A1(n8710), .A2(n7965), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6337), .ZN(n7294) );
  OAI22_X1 U8981 ( .A1(n8696), .A2(n7923), .B1(n8017), .B2(n8711), .ZN(n7293)
         );
  AOI211_X1 U8982 ( .C1(n7964), .C2(n8699), .A(n7294), .B(n7293), .ZN(n7295)
         );
  NAND2_X1 U8983 ( .A1(n7296), .A2(n7295), .ZN(P2_U3238) );
  OAI222_X1 U8984 ( .A1(n7298), .A2(P1_U3084), .B1(n10090), .B2(n7297), .C1(
        n7852), .C2(n10100), .ZN(P1_U3333) );
  NAND2_X1 U8985 ( .A1(n7299), .A2(n7300), .ZN(n7301) );
  XOR2_X1 U8986 ( .A(n7302), .B(n7301), .Z(n7309) );
  NAND2_X1 U8987 ( .A1(n9609), .A2(n9665), .ZN(n7304) );
  OR2_X1 U8988 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7303), .ZN(n10268) );
  OAI211_X1 U8989 ( .C1(n7305), .C2(n9578), .A(n7304), .B(n10268), .ZN(n7307)
         );
  INV_X1 U8990 ( .A(n7426), .ZN(n7411) );
  NOR2_X1 U8991 ( .A1(n9634), .A2(n7411), .ZN(n7306) );
  AOI211_X1 U8992 ( .C1(n7409), .C2(n9642), .A(n7307), .B(n7306), .ZN(n7308)
         );
  OAI21_X1 U8993 ( .B1(n7309), .B2(n9651), .A(n7308), .ZN(P1_U3219) );
  INV_X1 U8994 ( .A(n7310), .ZN(n8941) );
  NAND2_X1 U8995 ( .A1(n7311), .A2(n8941), .ZN(n7312) );
  NAND2_X1 U8996 ( .A1(n7460), .A2(n7374), .ZN(n8799) );
  NAND2_X1 U8997 ( .A1(n8797), .A2(n8799), .ZN(n8907) );
  OAI21_X1 U8998 ( .B1(n4556), .B2(n8907), .A(n7370), .ZN(n7459) );
  INV_X1 U8999 ( .A(n8907), .ZN(n7315) );
  NAND3_X1 U9000 ( .A1(n7314), .A2(n8907), .A3(n8792), .ZN(n7316) );
  AOI21_X1 U9001 ( .B1(n7928), .B2(n7316), .A(n9293), .ZN(n7318) );
  AOI211_X1 U9002 ( .C1(n7459), .C2(n7319), .A(n7318), .B(n7317), .ZN(n7463)
         );
  INV_X1 U9003 ( .A(n7320), .ZN(n7321) );
  INV_X1 U9004 ( .A(n7460), .ZN(n7322) );
  NAND2_X1 U9005 ( .A1(n7320), .A2(n7322), .ZN(n7378) );
  AOI21_X1 U9006 ( .B1(n7460), .B2(n7321), .A(n4988), .ZN(n7461) );
  NOR2_X1 U9007 ( .A1(n9338), .A2(n7322), .ZN(n7325) );
  OAI22_X1 U9008 ( .A1(n10370), .A2(n6736), .B1(n7323), .B2(n10375), .ZN(n7324) );
  AOI211_X1 U9009 ( .C1(n7461), .C2(n9347), .A(n7325), .B(n7324), .ZN(n7328)
         );
  NAND2_X1 U9010 ( .A1(n7459), .A2(n7326), .ZN(n7327) );
  OAI211_X1 U9011 ( .C1(n7463), .C2(n10357), .A(n7328), .B(n7327), .ZN(
        P2_U3287) );
  INV_X1 U9012 ( .A(n8533), .ZN(n7355) );
  AOI22_X1 U9013 ( .A1(n8763), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9471), .ZN(n7329) );
  OAI21_X1 U9014 ( .B1(n7355), .B2(n9463), .A(n7329), .ZN(P2_U3337) );
  AOI211_X1 U9015 ( .C1(n9437), .C2(n7332), .A(n7331), .B(n7330), .ZN(n7333)
         );
  OAI21_X1 U9016 ( .B1(n10426), .B2(n7334), .A(n7333), .ZN(n7336) );
  NAND2_X1 U9017 ( .A1(n7336), .A2(n10455), .ZN(n7335) );
  OAI21_X1 U9018 ( .B1(n10455), .B2(n6567), .A(n7335), .ZN(P2_U3527) );
  INV_X1 U9019 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U9020 ( .A1(n7336), .A2(n10444), .ZN(n7337) );
  OAI21_X1 U9021 ( .B1(n10444), .B2(n7338), .A(n7337), .ZN(P2_U3472) );
  NAND2_X1 U9022 ( .A1(n7344), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U9023 ( .A1(n7340), .A2(n7339), .ZN(n7342) );
  AOI22_X1 U9024 ( .A1(n7503), .A2(n8023), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7497), .ZN(n7341) );
  NOR2_X1 U9025 ( .A1(n7342), .A2(n7341), .ZN(n7496) );
  AOI21_X1 U9026 ( .B1(n7342), .B2(n7341), .A(n7496), .ZN(n7353) );
  AOI22_X1 U9027 ( .A1(n7503), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6363), .B2(
        n7497), .ZN(n7346) );
  OAI21_X1 U9028 ( .B1(n7344), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7343), .ZN(
        n7345) );
  NAND2_X1 U9029 ( .A1(n7346), .A2(n7345), .ZN(n7502) );
  OAI21_X1 U9030 ( .B1(n7346), .B2(n7345), .A(n7502), .ZN(n7347) );
  NAND2_X1 U9031 ( .A1(n7347), .A2(n10349), .ZN(n7352) );
  INV_X1 U9032 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7349) );
  OAI22_X1 U9033 ( .A1(n9056), .A2(n7349), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7348), .ZN(n7350) );
  AOI21_X1 U9034 ( .B1(n10347), .B2(n7503), .A(n7350), .ZN(n7351) );
  OAI211_X1 U9035 ( .C1(n7353), .C2(n9048), .A(n7352), .B(n7351), .ZN(P2_U3258) );
  INV_X1 U9036 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7354) );
  OAI222_X1 U9037 ( .A1(n7356), .A2(P1_U3084), .B1(n10090), .B2(n7355), .C1(
        n7354), .C2(n10100), .ZN(P1_U3332) );
  NAND2_X1 U9038 ( .A1(n7357), .A2(n8240), .ZN(n7358) );
  NAND2_X1 U9039 ( .A1(n8244), .A2(n8242), .ZN(n8455) );
  XNOR2_X1 U9040 ( .A(n7358), .B(n8455), .ZN(n7359) );
  AOI222_X1 U9041 ( .A1(n10152), .A2(n7359), .B1(n10148), .B2(n10149), .C1(
        n9664), .C2(n10147), .ZN(n10328) );
  XOR2_X1 U9042 ( .A(n7360), .B(n8455), .Z(n10333) );
  NAND2_X1 U9043 ( .A1(n10333), .A2(n9933), .ZN(n7368) );
  INV_X1 U9044 ( .A(n7361), .ZN(n10330) );
  INV_X1 U9045 ( .A(n7362), .ZN(n7407) );
  INV_X1 U9046 ( .A(n7448), .ZN(n7363) );
  OAI211_X1 U9047 ( .C1(n10330), .C2(n7407), .A(n7363), .B(n10032), .ZN(n10327) );
  INV_X1 U9048 ( .A(n10327), .ZN(n7366) );
  AOI22_X1 U9049 ( .A1(n10157), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7394), .B2(
        n10155), .ZN(n7364) );
  OAI21_X1 U9050 ( .B1(n10330), .B2(n10159), .A(n7364), .ZN(n7365) );
  AOI21_X1 U9051 ( .B1(n7366), .B2(n9963), .A(n7365), .ZN(n7367) );
  OAI211_X1 U9052 ( .C1(n10157), .C2(n10328), .A(n7368), .B(n7367), .ZN(
        P1_U3282) );
  OR2_X1 U9053 ( .A1(n7460), .A2(n4769), .ZN(n7369) );
  NAND2_X1 U9054 ( .A1(n7924), .A2(n7923), .ZN(n8803) );
  NAND2_X1 U9055 ( .A1(n8809), .A2(n8803), .ZN(n8909) );
  OAI21_X1 U9056 ( .B1(n4554), .B2(n8909), .A(n7926), .ZN(n10427) );
  NAND2_X1 U9057 ( .A1(n7928), .A2(n8799), .ZN(n7372) );
  INV_X1 U9058 ( .A(n8909), .ZN(n7371) );
  XNOR2_X1 U9059 ( .A(n7372), .B(n7371), .ZN(n7373) );
  NAND2_X1 U9060 ( .A1(n7373), .A2(n10365), .ZN(n7377) );
  OAI22_X1 U9061 ( .A1(n7955), .A2(n9311), .B1(n7374), .B2(n9309), .ZN(n7375)
         );
  INV_X1 U9062 ( .A(n7375), .ZN(n7376) );
  NAND2_X1 U9063 ( .A1(n7377), .A2(n7376), .ZN(n10430) );
  NAND2_X1 U9064 ( .A1(n7378), .A2(n7924), .ZN(n7379) );
  NAND2_X1 U9065 ( .A1(n7930), .A2(n7379), .ZN(n10428) );
  OAI22_X1 U9066 ( .A1(n10370), .A2(n7381), .B1(n7380), .B2(n10375), .ZN(n7382) );
  AOI21_X1 U9067 ( .B1(n9325), .B2(n7924), .A(n7382), .ZN(n7383) );
  OAI21_X1 U9068 ( .B1(n10428), .B2(n9321), .A(n7383), .ZN(n7384) );
  AOI21_X1 U9069 ( .B1(n10430), .B2(n10370), .A(n7384), .ZN(n7385) );
  OAI21_X1 U9070 ( .B1(n10427), .B2(n9349), .A(n7385), .ZN(P2_U3286) );
  INV_X1 U9071 ( .A(n7386), .ZN(n7387) );
  AOI21_X1 U9072 ( .B1(n7389), .B2(n7388), .A(n7387), .ZN(n7396) );
  NAND2_X1 U9073 ( .A1(n9609), .A2(n9664), .ZN(n7390) );
  NAND2_X1 U9074 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10285) );
  OAI211_X1 U9075 ( .C1(n7391), .C2(n9578), .A(n7390), .B(n10285), .ZN(n7393)
         );
  NOR2_X1 U9076 ( .A1(n9634), .A2(n10330), .ZN(n7392) );
  AOI211_X1 U9077 ( .C1(n7394), .C2(n9642), .A(n7393), .B(n7392), .ZN(n7395)
         );
  OAI21_X1 U9078 ( .B1(n7396), .B2(n9651), .A(n7395), .ZN(P1_U3229) );
  INV_X1 U9079 ( .A(n8547), .ZN(n7457) );
  AOI22_X1 U9080 ( .A1(n6141), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n9471), .ZN(n7397) );
  OAI21_X1 U9081 ( .B1(n7457), .B2(n9463), .A(n7397), .ZN(P2_U3336) );
  INV_X1 U9082 ( .A(n7398), .ZN(n7399) );
  AOI21_X1 U9083 ( .B1(n8452), .B2(n7400), .A(n7399), .ZN(n7405) );
  INV_X1 U9084 ( .A(n7405), .ZN(n7430) );
  INV_X1 U9085 ( .A(n10144), .ZN(n7415) );
  XNOR2_X1 U9086 ( .A(n7401), .B(n8452), .ZN(n7403) );
  AOI22_X1 U9087 ( .A1(n10147), .A2(n9665), .B1(n9663), .B2(n10149), .ZN(n7402) );
  OAI21_X1 U9088 ( .B1(n7403), .B2(n10128), .A(n7402), .ZN(n7404) );
  AOI21_X1 U9089 ( .B1(n7405), .B2(n10131), .A(n7404), .ZN(n7429) );
  MUX2_X1 U9090 ( .A(n7406), .B(n7429), .S(n10161), .Z(n7414) );
  AOI21_X1 U9091 ( .B1(n7426), .B2(n7408), .A(n7407), .ZN(n7427) );
  INV_X1 U9092 ( .A(n7409), .ZN(n7410) );
  OAI22_X1 U9093 ( .A1(n8122), .A2(n7411), .B1(n7410), .B2(n9926), .ZN(n7412)
         );
  AOI21_X1 U9094 ( .B1(n7427), .B2(n10143), .A(n7412), .ZN(n7413) );
  OAI211_X1 U9095 ( .C1(n7430), .C2(n7415), .A(n7414), .B(n7413), .ZN(P1_U3283) );
  NAND2_X1 U9096 ( .A1(n7438), .A2(n7416), .ZN(n7419) );
  NAND2_X1 U9097 ( .A1(n7437), .A2(n7417), .ZN(n7418) );
  XOR2_X1 U9098 ( .A(n7419), .B(n7418), .Z(n7425) );
  INV_X1 U9099 ( .A(n8012), .ZN(n8938) );
  INV_X1 U9100 ( .A(n7955), .ZN(n8940) );
  AOI22_X1 U9101 ( .A1(n8684), .A2(n8938), .B1(n8714), .B2(n8940), .ZN(n7422)
         );
  INV_X1 U9102 ( .A(n7420), .ZN(n7421) );
  OAI211_X1 U9103 ( .C1(n7957), .C2(n8710), .A(n7422), .B(n7421), .ZN(n7423)
         );
  AOI21_X1 U9104 ( .B1(n8010), .B2(n8699), .A(n7423), .ZN(n7424) );
  OAI21_X1 U9105 ( .B1(n7425), .B2(n4808), .A(n7424), .ZN(P2_U3226) );
  AOI22_X1 U9106 ( .A1(n7427), .A2(n10032), .B1(n10031), .B2(n7426), .ZN(n7428) );
  OAI211_X1 U9107 ( .C1(n10102), .C2(n7430), .A(n7429), .B(n7428), .ZN(n7433)
         );
  NAND2_X1 U9108 ( .A1(n7433), .A2(n10344), .ZN(n7431) );
  OAI21_X1 U9109 ( .B1(n10344), .B2(n7432), .A(n7431), .ZN(P1_U3531) );
  INV_X1 U9110 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9111 ( .A1(n7433), .A2(n10336), .ZN(n7434) );
  OAI21_X1 U9112 ( .B1(n10336), .B2(n7435), .A(n7434), .ZN(P1_U3478) );
  NAND2_X1 U9113 ( .A1(n7437), .A2(n7436), .ZN(n7439) );
  AND2_X1 U9114 ( .A1(n7439), .A2(n7438), .ZN(n7441) );
  XNOR2_X1 U9115 ( .A(n7441), .B(n7440), .ZN(n7446) );
  OAI22_X1 U9116 ( .A1(n8710), .A2(n8022), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7348), .ZN(n7444) );
  OAI22_X1 U9117 ( .A1(n8696), .A2(n8017), .B1(n8937), .B2(n8711), .ZN(n7443)
         );
  AOI211_X1 U9118 ( .C1(n8141), .C2(n8699), .A(n7444), .B(n7443), .ZN(n7445)
         );
  OAI21_X1 U9119 ( .B1(n7446), .B2(n4808), .A(n7445), .ZN(P2_U3236) );
  XNOR2_X1 U9120 ( .A(n7447), .B(n7450), .ZN(n10106) );
  OAI211_X1 U9121 ( .C1(n7448), .C2(n10105), .A(n10139), .B(n10032), .ZN(
        n10103) );
  INV_X1 U9122 ( .A(n10103), .ZN(n7455) );
  AOI22_X1 U9123 ( .A1(n10157), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7475), .B2(
        n10155), .ZN(n7449) );
  OAI21_X1 U9124 ( .B1(n10105), .B2(n10159), .A(n7449), .ZN(n7454) );
  XNOR2_X1 U9125 ( .A(n7451), .B(n7450), .ZN(n7452) );
  AOI222_X1 U9126 ( .A1(n10152), .A2(n7452), .B1(n9663), .B2(n10147), .C1(
        n9662), .C2(n10149), .ZN(n10104) );
  NOR2_X1 U9127 ( .A1(n10104), .A2(n10157), .ZN(n7453) );
  AOI211_X1 U9128 ( .C1(n7455), .C2(n9963), .A(n7454), .B(n7453), .ZN(n7456)
         );
  OAI21_X1 U9129 ( .B1(n9969), .B2(n10106), .A(n7456), .ZN(P1_U3281) );
  OAI222_X1 U9130 ( .A1(P1_U3084), .A2(n7458), .B1(n10090), .B2(n7457), .C1(
        n7802), .C2(n10100), .ZN(P1_U3331) );
  INV_X1 U9131 ( .A(n7459), .ZN(n7464) );
  AOI22_X1 U9132 ( .A1(n7461), .A2(n10411), .B1(n9437), .B2(n7460), .ZN(n7462)
         );
  OAI211_X1 U9133 ( .C1(n7464), .C2(n10418), .A(n7463), .B(n7462), .ZN(n7466)
         );
  NAND2_X1 U9134 ( .A1(n7466), .A2(n10455), .ZN(n7465) );
  OAI21_X1 U9135 ( .B1(n10455), .B2(n6729), .A(n7465), .ZN(P2_U3529) );
  INV_X1 U9136 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9137 ( .A1(n7466), .A2(n10444), .ZN(n7467) );
  OAI21_X1 U9138 ( .B1(n10444), .B2(n7468), .A(n7467), .ZN(P2_U3478) );
  XOR2_X1 U9139 ( .A(n7470), .B(n7469), .Z(n7471) );
  XNOR2_X1 U9140 ( .A(n7472), .B(n7471), .ZN(n7481) );
  NOR2_X1 U9141 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7473), .ZN(n10301) );
  AOI21_X1 U9142 ( .B1(n9640), .B2(n9662), .A(n10301), .ZN(n7479) );
  NAND2_X1 U9143 ( .A1(n7474), .A2(n9612), .ZN(n7478) );
  NAND2_X1 U9144 ( .A1(n9642), .A2(n7475), .ZN(n7477) );
  NAND2_X1 U9145 ( .A1(n9609), .A2(n9663), .ZN(n7476) );
  NAND4_X1 U9146 ( .A1(n7479), .A2(n7478), .A3(n7477), .A4(n7476), .ZN(n7480)
         );
  AOI21_X1 U9147 ( .B1(n7481), .B2(n9607), .A(n7480), .ZN(n7482) );
  INV_X1 U9148 ( .A(n7482), .ZN(P1_U3215) );
  INV_X1 U9149 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8159) );
  MUX2_X1 U9150 ( .A(n8159), .B(P1_REG1_REG_14__SCAN_IN), .S(n9674), .Z(n7486)
         );
  AOI21_X1 U9151 ( .B1(n10177), .B2(n7484), .A(n7483), .ZN(n7485) );
  AOI21_X1 U9152 ( .B1(n7486), .B2(n7485), .A(n9677), .ZN(n7495) );
  INV_X1 U9153 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7490) );
  AOI211_X1 U9154 ( .C1(n7490), .C2(n7489), .A(n10296), .B(n9672), .ZN(n7491)
         );
  INV_X1 U9155 ( .A(n7491), .ZN(n7494) );
  NAND2_X1 U9156 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9490) );
  OAI21_X1 U9157 ( .B1(n10254), .B2(n9678), .A(n9490), .ZN(n7492) );
  AOI21_X1 U9158 ( .B1(n10306), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7492), .ZN(
        n7493) );
  OAI211_X1 U9159 ( .C1(n7495), .C2(n10288), .A(n7494), .B(n7493), .ZN(
        P1_U3255) );
  AOI21_X1 U9160 ( .B1(n7497), .B2(n8023), .A(n7496), .ZN(n7499) );
  AOI22_X1 U9161 ( .A1(n8133), .A2(n8051), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7500), .ZN(n7498) );
  NOR2_X1 U9162 ( .A1(n7499), .A2(n7498), .ZN(n8127) );
  AOI21_X1 U9163 ( .B1(n7499), .B2(n7498), .A(n8127), .ZN(n7511) );
  AOI22_X1 U9164 ( .A1(n8133), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7501), .B2(
        n7500), .ZN(n7505) );
  OAI21_X1 U9165 ( .B1(n7505), .B2(n7504), .A(n8132), .ZN(n7509) );
  INV_X1 U9166 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U9167 ( .A1(n10347), .A2(n8133), .ZN(n7506) );
  NAND2_X1 U9168 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7526) );
  OAI211_X1 U9169 ( .C1(n7507), .C2(n9056), .A(n7506), .B(n7526), .ZN(n7508)
         );
  AOI21_X1 U9170 ( .B1(n7509), .B2(n10349), .A(n7508), .ZN(n7510) );
  OAI21_X1 U9171 ( .B1(n7511), .B2(n9048), .A(n7510), .ZN(P2_U3259) );
  INV_X1 U9172 ( .A(n8561), .ZN(n7513) );
  AOI21_X1 U9173 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9471), .A(n8930), .ZN(
        n7512) );
  OAI21_X1 U9174 ( .B1(n7513), .B2(n9463), .A(n7512), .ZN(P2_U3335) );
  XNOR2_X1 U9175 ( .A(n7514), .B(n7515), .ZN(n7521) );
  AOI21_X1 U9176 ( .B1(n9609), .B2(n10148), .A(n7516), .ZN(n7518) );
  NAND2_X1 U9177 ( .A1(n9642), .A2(n10156), .ZN(n7517) );
  OAI211_X1 U9178 ( .C1(n8006), .C2(n9578), .A(n7518), .B(n7517), .ZN(n7519)
         );
  AOI21_X1 U9179 ( .B1(n10140), .B2(n9648), .A(n7519), .ZN(n7520) );
  OAI21_X1 U9180 ( .B1(n7521), .B2(n9651), .A(n7520), .ZN(P1_U3234) );
  INV_X1 U9181 ( .A(n7522), .ZN(n7523) );
  AOI21_X1 U9182 ( .B1(n7525), .B2(n7524), .A(n7523), .ZN(n7530) );
  OAI21_X1 U9183 ( .B1(n8710), .B2(n8059), .A(n7526), .ZN(n7528) );
  OAI22_X1 U9184 ( .A1(n8696), .A2(n8012), .B1(n9310), .B2(n8711), .ZN(n7527)
         );
  AOI211_X1 U9185 ( .C1(n9436), .C2(n8699), .A(n7528), .B(n7527), .ZN(n7529)
         );
  OAI21_X1 U9186 ( .B1(n7530), .B2(n4808), .A(n7529), .ZN(P2_U3217) );
  NAND2_X1 U9187 ( .A1(n8561), .A2(n10095), .ZN(n7532) );
  NAND2_X1 U9188 ( .A1(n7531), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8489) );
  OAI211_X1 U9189 ( .C1(n7816), .C2(n10086), .A(n7532), .B(n8489), .ZN(
        P1_U3330) );
  INV_X1 U9190 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10496) );
  NOR2_X1 U9191 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7533) );
  AOI21_X1 U9192 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7533), .ZN(n10463) );
  NOR2_X1 U9193 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7534) );
  AOI21_X1 U9194 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7534), .ZN(n10466) );
  NOR2_X1 U9195 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7535) );
  AOI21_X1 U9196 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7535), .ZN(n10469) );
  NOR2_X1 U9197 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7536) );
  AOI21_X1 U9198 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7536), .ZN(n10472) );
  NOR2_X1 U9199 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7537) );
  AOI21_X1 U9200 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7537), .ZN(n10475) );
  NOR2_X1 U9201 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7544) );
  XOR2_X1 U9202 ( .A(n10230), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10503) );
  NAND2_X1 U9203 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7542) );
  XNOR2_X1 U9204 ( .A(n7538), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U9205 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7540) );
  XNOR2_X1 U9206 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n10218), .ZN(n10490) );
  AOI21_X1 U9207 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10456) );
  INV_X1 U9208 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10460) );
  NAND3_X1 U9209 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10458) );
  OAI21_X1 U9210 ( .B1(n10456), .B2(n10460), .A(n10458), .ZN(n10489) );
  NAND2_X1 U9211 ( .A1(n10490), .A2(n10489), .ZN(n7539) );
  NAND2_X1 U9212 ( .A1(n7540), .A2(n7539), .ZN(n10500) );
  NAND2_X1 U9213 ( .A1(n10501), .A2(n10500), .ZN(n7541) );
  NAND2_X1 U9214 ( .A1(n7542), .A2(n7541), .ZN(n10502) );
  NOR2_X1 U9215 ( .A1(n10503), .A2(n10502), .ZN(n7543) );
  NOR2_X1 U9216 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  NOR2_X1 U9217 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7545), .ZN(n10492) );
  AND2_X1 U9218 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7545), .ZN(n10491) );
  NOR2_X1 U9219 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10491), .ZN(n7546) );
  NOR2_X1 U9220 ( .A1(n10492), .A2(n7546), .ZN(n7547) );
  NAND2_X1 U9221 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7547), .ZN(n7549) );
  XOR2_X1 U9222 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7547), .Z(n10499) );
  NAND2_X1 U9223 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10499), .ZN(n7548) );
  NAND2_X1 U9224 ( .A1(n7549), .A2(n7548), .ZN(n7550) );
  NAND2_X1 U9225 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7550), .ZN(n7552) );
  XOR2_X1 U9226 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7550), .Z(n10488) );
  NAND2_X1 U9227 ( .A1(n10488), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U9228 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  NAND2_X1 U9229 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7553), .ZN(n7555) );
  XOR2_X1 U9230 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7553), .Z(n10498) );
  NAND2_X1 U9231 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10498), .ZN(n7554) );
  NAND2_X1 U9232 ( .A1(n7555), .A2(n7554), .ZN(n7556) );
  AND2_X1 U9233 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7556), .ZN(n7557) );
  XNOR2_X1 U9234 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7556), .ZN(n10487) );
  INV_X1 U9235 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U9236 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7558) );
  OAI21_X1 U9237 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7558), .ZN(n10483) );
  NAND2_X1 U9238 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7559) );
  OAI21_X1 U9239 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7559), .ZN(n10480) );
  AOI21_X1 U9240 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10479), .ZN(n10478) );
  NOR2_X1 U9241 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7560) );
  AOI21_X1 U9242 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7560), .ZN(n10477) );
  NAND2_X1 U9243 ( .A1(n10478), .A2(n10477), .ZN(n10476) );
  OAI21_X1 U9244 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10476), .ZN(n10474) );
  NAND2_X1 U9245 ( .A1(n10475), .A2(n10474), .ZN(n10473) );
  OAI21_X1 U9246 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10473), .ZN(n10471) );
  NAND2_X1 U9247 ( .A1(n10472), .A2(n10471), .ZN(n10470) );
  OAI21_X1 U9248 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10470), .ZN(n10468) );
  NAND2_X1 U9249 ( .A1(n10469), .A2(n10468), .ZN(n10467) );
  OAI21_X1 U9250 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10467), .ZN(n10465) );
  NAND2_X1 U9251 ( .A1(n10466), .A2(n10465), .ZN(n10464) );
  OAI21_X1 U9252 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10464), .ZN(n10462) );
  NAND2_X1 U9253 ( .A1(n10463), .A2(n10462), .ZN(n10461) );
  OAI21_X1 U9254 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10461), .ZN(n10495) );
  NOR2_X1 U9255 ( .A1(n10496), .A2(n10495), .ZN(n7561) );
  NAND2_X1 U9256 ( .A1(n10496), .A2(n10495), .ZN(n10494) );
  OAI21_X1 U9257 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7561), .A(n10494), .ZN(
        n7920) );
  OAI22_X1 U9258 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g104), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_g100), .ZN(n7562) );
  AOI221_X1 U9259 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g100), .C2(P1_IR_REG_9__SCAN_IN), .A(n7562), .ZN(n7569) );
  OAI22_X1 U9260 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_g83), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n7563) );
  AOI221_X1 U9261 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .C1(
        keyinput_g36), .C2(P2_REG3_REG_27__SCAN_IN), .A(n7563), .ZN(n7568) );
  OAI22_X1 U9262 ( .A1(SI_18_), .A2(keyinput_g14), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_g52), .ZN(n7564) );
  AOI221_X1 U9263 ( .B1(SI_18_), .B2(keyinput_g14), .C1(keyinput_g52), .C2(
        P2_REG3_REG_4__SCAN_IN), .A(n7564), .ZN(n7567) );
  OAI22_X1 U9264 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_g126), .B1(
        keyinput_g33), .B2(P2_RD_REG_SCAN_IN), .ZN(n7565) );
  AOI221_X1 U9265 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_g126), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n7565), .ZN(n7566) );
  NAND4_X1 U9266 ( .A1(n7569), .A2(n7568), .A3(n7567), .A4(n7566), .ZN(n7693)
         );
  OAI22_X1 U9267 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g105), .B1(
        keyinput_g85), .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7570) );
  AOI221_X1 U9268 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g105), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n7570), .ZN(n7596) );
  OAI22_X1 U9269 ( .A1(SI_22_), .A2(keyinput_g10), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n7571) );
  AOI221_X1 U9270 ( .B1(SI_22_), .B2(keyinput_g10), .C1(keyinput_g53), .C2(
        P2_REG3_REG_9__SCAN_IN), .A(n7571), .ZN(n7574) );
  OAI22_X1 U9271 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n7572) );
  AOI221_X1 U9272 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        keyinput_g41), .C2(P2_REG3_REG_19__SCAN_IN), .A(n7572), .ZN(n7573) );
  OAI211_X1 U9273 ( .C1(n7576), .C2(keyinput_g15), .A(n7574), .B(n7573), .ZN(
        n7575) );
  AOI21_X1 U9274 ( .B1(n7576), .B2(keyinput_g15), .A(n7575), .ZN(n7595) );
  AOI22_X1 U9275 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P1_IR_REG_18__SCAN_IN), 
        .B2(keyinput_g109), .ZN(n7577) );
  OAI221_X1 U9276 ( .B1(SI_31_), .B2(keyinput_g1), .C1(P1_IR_REG_18__SCAN_IN), 
        .C2(keyinput_g109), .A(n7577), .ZN(n7584) );
  AOI22_X1 U9277 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_g114), .ZN(n7578) );
  OAI221_X1 U9278 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_g114), .A(n7578), .ZN(n7583) );
  AOI22_X1 U9279 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_g124), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g101), .ZN(n7579) );
  OAI221_X1 U9280 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_g124), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g101), .A(n7579), .ZN(n7582) );
  AOI22_X1 U9281 ( .A1(SI_10_), .A2(keyinput_g22), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .ZN(n7580) );
  OAI221_X1 U9282 ( .B1(SI_10_), .B2(keyinput_g22), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_g78), .A(n7580), .ZN(n7581) );
  NOR4_X1 U9283 ( .A1(n7584), .A2(n7583), .A3(n7582), .A4(n7581), .ZN(n7594)
         );
  AOI22_X1 U9284 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_g122), .ZN(n7585) );
  OAI221_X1 U9285 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_g122), .A(n7585), .ZN(n7592) );
  AOI22_X1 U9286 ( .A1(SI_16_), .A2(keyinput_g16), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n7586) );
  OAI221_X1 U9287 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n7586), .ZN(n7591) );
  AOI22_X1 U9288 ( .A1(SI_27_), .A2(keyinput_g5), .B1(P1_IR_REG_2__SCAN_IN), 
        .B2(keyinput_g93), .ZN(n7587) );
  OAI221_X1 U9289 ( .B1(SI_27_), .B2(keyinput_g5), .C1(P1_IR_REG_2__SCAN_IN), 
        .C2(keyinput_g93), .A(n7587), .ZN(n7590) );
  AOI22_X1 U9290 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(SI_21_), .B2(keyinput_g11), .ZN(n7588) );
  OAI221_X1 U9291 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_21_), .C2(keyinput_g11), .A(n7588), .ZN(n7589) );
  NOR4_X1 U9292 ( .A1(n7592), .A2(n7591), .A3(n7590), .A4(n7589), .ZN(n7593)
         );
  NAND4_X1 U9293 ( .A1(n7596), .A2(n7595), .A3(n7594), .A4(n7593), .ZN(n7692)
         );
  INV_X1 U9294 ( .A(P2_B_REG_SCAN_IN), .ZN(n7599) );
  AOI22_X1 U9295 ( .A1(n7599), .A2(keyinput_g64), .B1(n7598), .B2(keyinput_g23), .ZN(n7597) );
  OAI221_X1 U9296 ( .B1(n7599), .B2(keyinput_g64), .C1(n7598), .C2(
        keyinput_g23), .A(n7597), .ZN(n7608) );
  INV_X1 U9297 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7601) );
  AOI22_X1 U9298 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_g89), .B1(n7601), 
        .B2(keyinput_g98), .ZN(n7600) );
  OAI221_X1 U9299 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .C1(n7601), .C2(keyinput_g98), .A(n7600), .ZN(n7607) );
  XNOR2_X1 U9300 ( .A(SI_30_), .B(keyinput_g2), .ZN(n7605) );
  XNOR2_X1 U9301 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_g99), .ZN(n7604) );
  XNOR2_X1 U9302 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g119), .ZN(n7603) );
  XNOR2_X1 U9303 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g112), .ZN(n7602) );
  NAND4_X1 U9304 ( .A1(n7605), .A2(n7604), .A3(n7603), .A4(n7602), .ZN(n7606)
         );
  NOR3_X1 U9305 ( .A1(n7608), .A2(n7607), .A3(n7606), .ZN(n7643) );
  AOI22_X1 U9306 ( .A1(n7610), .A2(keyinput_g21), .B1(keyinput_g49), .B2(n6223), .ZN(n7609) );
  OAI221_X1 U9307 ( .B1(n7610), .B2(keyinput_g21), .C1(n6223), .C2(
        keyinput_g49), .A(n7609), .ZN(n7619) );
  AOI22_X1 U9308 ( .A1(n7841), .A2(keyinput_g77), .B1(keyinput_g18), .B2(n7612), .ZN(n7611) );
  OAI221_X1 U9309 ( .B1(n7841), .B2(keyinput_g77), .C1(n7612), .C2(
        keyinput_g18), .A(n7611), .ZN(n7618) );
  INV_X1 U9310 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8709) );
  AOI22_X1 U9311 ( .A1(n8709), .A2(keyinput_g62), .B1(n7855), .B2(keyinput_g87), .ZN(n7613) );
  OAI221_X1 U9312 ( .B1(n8709), .B2(keyinput_g62), .C1(n7855), .C2(
        keyinput_g87), .A(n7613), .ZN(n7617) );
  AOI22_X1 U9313 ( .A1(n7348), .A2(keyinput_g56), .B1(keyinput_g61), .B2(n7615), .ZN(n7614) );
  OAI221_X1 U9314 ( .B1(n7348), .B2(keyinput_g56), .C1(n7615), .C2(
        keyinput_g61), .A(n7614), .ZN(n7616) );
  NOR4_X1 U9315 ( .A1(n7619), .A2(n7618), .A3(n7617), .A4(n7616), .ZN(n7642)
         );
  INV_X1 U9316 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U9317 ( .A1(n10310), .A2(keyinput_g125), .B1(keyinput_g58), .B2(
        n6337), .ZN(n7620) );
  OAI221_X1 U9318 ( .B1(n10310), .B2(keyinput_g125), .C1(n6337), .C2(
        keyinput_g58), .A(n7620), .ZN(n7629) );
  INV_X1 U9319 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10094) );
  INV_X1 U9320 ( .A(SI_13_), .ZN(n7622) );
  AOI22_X1 U9321 ( .A1(n10094), .A2(keyinput_g68), .B1(n7622), .B2(
        keyinput_g19), .ZN(n7621) );
  OAI221_X1 U9322 ( .B1(n10094), .B2(keyinput_g68), .C1(n7622), .C2(
        keyinput_g19), .A(n7621), .ZN(n7628) );
  AOI22_X1 U9323 ( .A1(n7936), .A2(keyinput_g72), .B1(keyinput_g73), .B2(n7816), .ZN(n7623) );
  OAI221_X1 U9324 ( .B1(n7936), .B2(keyinput_g72), .C1(n7816), .C2(
        keyinput_g73), .A(n7623), .ZN(n7627) );
  XNOR2_X1 U9325 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g117), .ZN(n7625) );
  XNOR2_X1 U9326 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_g55), .ZN(n7624)
         );
  NAND2_X1 U9327 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NOR4_X1 U9328 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n7641)
         );
  AOI22_X1 U9329 ( .A1(n7802), .A2(keyinput_g74), .B1(keyinput_g43), .B2(n7631), .ZN(n7630) );
  OAI221_X1 U9330 ( .B1(n7802), .B2(keyinput_g74), .C1(n7631), .C2(
        keyinput_g43), .A(n7630), .ZN(n7639) );
  XOR2_X1 U9331 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g92), .Z(n7638) );
  XOR2_X1 U9332 ( .A(SI_6_), .B(keyinput_g26), .Z(n7637) );
  XNOR2_X1 U9333 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g97), .ZN(n7635) );
  XNOR2_X1 U9334 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_g50), .ZN(n7634)
         );
  XNOR2_X1 U9335 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_g34), .ZN(n7633) );
  XNOR2_X1 U9336 ( .A(SI_3_), .B(keyinput_g29), .ZN(n7632) );
  NAND4_X1 U9337 ( .A1(n7635), .A2(n7634), .A3(n7633), .A4(n7632), .ZN(n7636)
         );
  NOR4_X1 U9338 ( .A1(n7639), .A2(n7638), .A3(n7637), .A4(n7636), .ZN(n7640)
         );
  NAND4_X1 U9339 ( .A1(n7643), .A2(n7642), .A3(n7641), .A4(n7640), .ZN(n7691)
         );
  AOI22_X1 U9340 ( .A1(n7645), .A2(keyinput_g9), .B1(keyinput_g76), .B2(n7852), 
        .ZN(n7644) );
  OAI221_X1 U9341 ( .B1(n7645), .B2(keyinput_g9), .C1(n7852), .C2(keyinput_g76), .A(n7644), .ZN(n7654) );
  INV_X1 U9342 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7800) );
  AOI22_X1 U9343 ( .A1(n7800), .A2(keyinput_g102), .B1(keyinput_g4), .B2(n6044), .ZN(n7646) );
  OAI221_X1 U9344 ( .B1(n7800), .B2(keyinput_g102), .C1(n6044), .C2(
        keyinput_g4), .A(n7646), .ZN(n7653) );
  INV_X1 U9345 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8681) );
  AOI22_X1 U9346 ( .A1(n7648), .A2(keyinput_g28), .B1(keyinput_g51), .B2(n8681), .ZN(n7647) );
  OAI221_X1 U9347 ( .B1(n7648), .B2(keyinput_g28), .C1(n8681), .C2(
        keyinput_g51), .A(n7647), .ZN(n7652) );
  XNOR2_X1 U9348 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g116), .ZN(n7650) );
  XNOR2_X1 U9349 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g103), .ZN(n7649) );
  NAND2_X1 U9350 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  NOR4_X1 U9351 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n7689)
         );
  AOI22_X1 U9352 ( .A1(n7656), .A2(keyinput_g27), .B1(keyinput_g39), .B2(n7815), .ZN(n7655) );
  OAI221_X1 U9353 ( .B1(n7656), .B2(keyinput_g27), .C1(n7815), .C2(
        keyinput_g39), .A(n7655), .ZN(n7665) );
  AOI22_X1 U9354 ( .A1(n6176), .A2(keyinput_g59), .B1(n8151), .B2(keyinput_g71), .ZN(n7657) );
  OAI221_X1 U9355 ( .B1(n6176), .B2(keyinput_g59), .C1(n8151), .C2(
        keyinput_g71), .A(n7657), .ZN(n7664) );
  INV_X1 U9356 ( .A(SI_24_), .ZN(n7777) );
  AOI22_X1 U9357 ( .A1(n7659), .A2(keyinput_g108), .B1(keyinput_g8), .B2(n7777), .ZN(n7658) );
  OAI221_X1 U9358 ( .B1(n7659), .B2(keyinput_g108), .C1(n7777), .C2(
        keyinput_g8), .A(n7658), .ZN(n7663) );
  XNOR2_X1 U9359 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g95), .ZN(n7661) );
  XNOR2_X1 U9360 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_g84), .ZN(n7660)
         );
  NAND2_X1 U9361 ( .A1(n7661), .A2(n7660), .ZN(n7662) );
  NOR4_X1 U9362 ( .A1(n7665), .A2(n7664), .A3(n7663), .A4(n7662), .ZN(n7688)
         );
  INV_X1 U9363 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10190) );
  AOI22_X1 U9364 ( .A1(n7667), .A2(keyinput_g48), .B1(keyinput_g0), .B2(n10190), .ZN(n7666) );
  OAI221_X1 U9365 ( .B1(n7667), .B2(keyinput_g48), .C1(n10190), .C2(
        keyinput_g0), .A(n7666), .ZN(n7676) );
  AOI22_X1 U9366 ( .A1(n7669), .A2(keyinput_g40), .B1(n8671), .B2(keyinput_g47), .ZN(n7668) );
  OAI221_X1 U9367 ( .B1(n7669), .B2(keyinput_g40), .C1(n8671), .C2(
        keyinput_g47), .A(n7668), .ZN(n7675) );
  XNOR2_X1 U9368 ( .A(SI_19_), .B(keyinput_g13), .ZN(n7673) );
  XNOR2_X1 U9369 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g111), .ZN(n7672) );
  XNOR2_X1 U9370 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_g121), .ZN(n7671) );
  XNOR2_X1 U9371 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n7670)
         );
  NAND4_X1 U9372 ( .A1(n7673), .A2(n7672), .A3(n7671), .A4(n7670), .ZN(n7674)
         );
  NOR3_X1 U9373 ( .A1(n7676), .A2(n7675), .A3(n7674), .ZN(n7687) );
  AOI22_X1 U9374 ( .A1(n6133), .A2(keyinput_g63), .B1(n7858), .B2(keyinput_g82), .ZN(n7677) );
  OAI221_X1 U9375 ( .B1(n6133), .B2(keyinput_g63), .C1(n7858), .C2(
        keyinput_g82), .A(n7677), .ZN(n7685) );
  INV_X1 U9376 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8645) );
  AOI22_X1 U9377 ( .A1(n10099), .A2(keyinput_g69), .B1(keyinput_g38), .B2(
        n8645), .ZN(n7678) );
  OAI221_X1 U9378 ( .B1(n10099), .B2(keyinput_g69), .C1(n8645), .C2(
        keyinput_g38), .A(n7678), .ZN(n7684) );
  XOR2_X1 U9379 ( .A(n7819), .B(keyinput_g65), .Z(n7682) );
  XNOR2_X1 U9380 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_g60), .ZN(n7681)
         );
  XNOR2_X1 U9381 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_g113), .ZN(n7680) );
  XNOR2_X1 U9382 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g106), .ZN(n7679) );
  NAND4_X1 U9383 ( .A1(n7682), .A2(n7681), .A3(n7680), .A4(n7679), .ZN(n7683)
         );
  NOR3_X1 U9384 ( .A1(n7685), .A2(n7684), .A3(n7683), .ZN(n7686) );
  NAND4_X1 U9385 ( .A1(n7689), .A2(n7688), .A3(n7687), .A4(n7686), .ZN(n7690)
         );
  NOR4_X1 U9386 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n7916)
         );
  OAI22_X1 U9387 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g94), .B1(SI_7_), 
        .B2(keyinput_g25), .ZN(n7694) );
  AOI221_X1 U9388 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g25), .C2(SI_7_), .A(n7694), .ZN(n7701) );
  OAI22_X1 U9389 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_g118), .B1(
        keyinput_g17), .B2(SI_15_), .ZN(n7695) );
  AOI221_X1 U9390 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_g118), .C1(SI_15_), .C2(keyinput_g17), .A(n7695), .ZN(n7700) );
  OAI22_X1 U9391 ( .A1(SI_2_), .A2(keyinput_g30), .B1(keyinput_g35), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n7696) );
  AOI221_X1 U9392 ( .B1(SI_2_), .B2(keyinput_g30), .C1(P2_REG3_REG_7__SCAN_IN), 
        .C2(keyinput_g35), .A(n7696), .ZN(n7699) );
  OAI22_X1 U9393 ( .A1(SI_12_), .A2(keyinput_g20), .B1(keyinput_g3), .B2(
        SI_29_), .ZN(n7697) );
  AOI221_X1 U9394 ( .B1(SI_12_), .B2(keyinput_g20), .C1(SI_29_), .C2(
        keyinput_g3), .A(n7697), .ZN(n7698) );
  NAND4_X1 U9395 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n7698), .ZN(n7729)
         );
  OAI22_X1 U9396 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n7702) );
  AOI221_X1 U9397 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g37), .C2(P2_REG3_REG_14__SCAN_IN), .A(n7702), .ZN(n7709) );
  OAI22_X1 U9398 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g96), .B1(
        keyinput_g91), .B2(P1_IR_REG_0__SCAN_IN), .ZN(n7703) );
  AOI221_X1 U9399 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g96), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_g91), .A(n7703), .ZN(n7708) );
  OAI22_X1 U9400 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g80), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n7704) );
  AOI221_X1 U9401 ( .B1(SI_25_), .B2(keyinput_g7), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_g80), .A(n7704), .ZN(n7707) );
  OAI22_X1 U9402 ( .A1(SI_20_), .A2(keyinput_g12), .B1(P1_IR_REG_29__SCAN_IN), 
        .B2(keyinput_g120), .ZN(n7705) );
  AOI221_X1 U9403 ( .B1(SI_20_), .B2(keyinput_g12), .C1(keyinput_g120), .C2(
        P1_IR_REG_29__SCAN_IN), .A(n7705), .ZN(n7706) );
  NAND4_X1 U9404 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .ZN(n7728)
         );
  OAI22_X1 U9405 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_g123), .B1(SI_8_), 
        .B2(keyinput_g24), .ZN(n7710) );
  AOI221_X1 U9406 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_g123), .C1(
        keyinput_g24), .C2(SI_8_), .A(n7710), .ZN(n7717) );
  OAI22_X1 U9407 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g127), .B1(
        keyinput_g46), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n7711) );
  AOI221_X1 U9408 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g127), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n7711), .ZN(n7716) );
  OAI22_X1 U9409 ( .A1(SI_26_), .A2(keyinput_g6), .B1(keyinput_g31), .B2(SI_1_), .ZN(n7712) );
  AOI221_X1 U9410 ( .B1(SI_26_), .B2(keyinput_g6), .C1(SI_1_), .C2(
        keyinput_g31), .A(n7712), .ZN(n7715) );
  OAI22_X1 U9411 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_g70), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .ZN(n7713) );
  AOI221_X1 U9412 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .C1(
        keyinput_g79), .C2(P2_DATAO_REG_17__SCAN_IN), .A(n7713), .ZN(n7714) );
  NAND4_X1 U9413 ( .A1(n7717), .A2(n7716), .A3(n7715), .A4(n7714), .ZN(n7727)
         );
  OAI22_X1 U9414 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .ZN(n7718) );
  AOI221_X1 U9415 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g90), .C2(P2_DATAO_REG_6__SCAN_IN), .A(n7718), .ZN(n7725) );
  OAI22_X1 U9416 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g44), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n7719) );
  AOI221_X1 U9417 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g110), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n7719), .ZN(n7724) );
  OAI22_X1 U9418 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g107), .B1(SI_0_), 
        .B2(keyinput_g32), .ZN(n7720) );
  AOI221_X1 U9419 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g107), .C1(
        keyinput_g32), .C2(SI_0_), .A(n7720), .ZN(n7723) );
  OAI22_X1 U9420 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_g66), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .ZN(n7721) );
  AOI221_X1 U9421 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .C1(
        keyinput_g67), .C2(P2_DATAO_REG_29__SCAN_IN), .A(n7721), .ZN(n7722) );
  NAND4_X1 U9422 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n7726)
         );
  NOR4_X1 U9423 ( .A1(n7729), .A2(n7728), .A3(n7727), .A4(n7726), .ZN(n7915)
         );
  XNOR2_X1 U9424 ( .A(n7909), .B(keyinput_g115), .ZN(n7914) );
  OAI22_X1 U9425 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_f33), .B1(SI_18_), 
        .B2(keyinput_f14), .ZN(n7730) );
  AOI221_X1 U9426 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .C1(
        keyinput_f14), .C2(SI_18_), .A(n7730), .ZN(n7737) );
  OAI22_X1 U9427 ( .A1(SI_9_), .A2(keyinput_f23), .B1(keyinput_f51), .B2(
        P2_REG3_REG_24__SCAN_IN), .ZN(n7731) );
  AOI221_X1 U9428 ( .B1(SI_9_), .B2(keyinput_f23), .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n7731), .ZN(n7736) );
  OAI22_X1 U9429 ( .A1(SI_25_), .A2(keyinput_f7), .B1(keyinput_f78), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7732) );
  AOI221_X1 U9430 ( .B1(SI_25_), .B2(keyinput_f7), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_f78), .A(n7732), .ZN(n7735) );
  OAI22_X1 U9431 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f99), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_f97), .ZN(n7733) );
  AOI221_X1 U9432 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f99), .C1(
        keyinput_f97), .C2(P1_IR_REG_6__SCAN_IN), .A(n7733), .ZN(n7734) );
  NAND4_X1 U9433 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), .ZN(n7872)
         );
  OAI22_X1 U9434 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f126), .B1(
        keyinput_f34), .B2(P2_STATE_REG_SCAN_IN), .ZN(n7738) );
  AOI221_X1 U9435 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f126), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n7738), .ZN(n7763) );
  OAI22_X1 U9436 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        SI_31_), .B2(keyinput_f1), .ZN(n7739) );
  AOI221_X1 U9437 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        keyinput_f1), .C2(SI_31_), .A(n7739), .ZN(n7742) );
  OAI22_X1 U9438 ( .A1(SI_17_), .A2(keyinput_f15), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(keyinput_f44), .ZN(n7740) );
  AOI221_X1 U9439 ( .B1(SI_17_), .B2(keyinput_f15), .C1(keyinput_f44), .C2(
        P2_REG3_REG_1__SCAN_IN), .A(n7740), .ZN(n7741) );
  OAI211_X1 U9440 ( .C1(n10099), .C2(keyinput_f69), .A(n7742), .B(n7741), .ZN(
        n7743) );
  AOI21_X1 U9441 ( .B1(n10099), .B2(keyinput_f69), .A(n7743), .ZN(n7762) );
  AOI22_X1 U9442 ( .A1(SI_20_), .A2(keyinput_f12), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n7744) );
  OAI221_X1 U9443 ( .B1(SI_20_), .B2(keyinput_f12), .C1(SI_26_), .C2(
        keyinput_f6), .A(n7744), .ZN(n7751) );
  AOI22_X1 U9444 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n7745) );
  OAI221_X1 U9445 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n7745), .ZN(n7750) );
  AOI22_X1 U9446 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput_f118), .ZN(n7746) );
  OAI221_X1 U9447 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_f118), .A(n7746), .ZN(n7749) );
  AOI22_X1 U9448 ( .A1(SI_8_), .A2(keyinput_f24), .B1(P1_IR_REG_9__SCAN_IN), 
        .B2(keyinput_f100), .ZN(n7747) );
  OAI221_X1 U9449 ( .B1(SI_8_), .B2(keyinput_f24), .C1(P1_IR_REG_9__SCAN_IN), 
        .C2(keyinput_f100), .A(n7747), .ZN(n7748) );
  NOR4_X1 U9450 ( .A1(n7751), .A2(n7750), .A3(n7749), .A4(n7748), .ZN(n7761)
         );
  AOI22_X1 U9451 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput_f124), .ZN(n7752) );
  OAI221_X1 U9452 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_f124), .A(n7752), .ZN(n7759) );
  AOI22_X1 U9453 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_f114), .ZN(n7753) );
  OAI221_X1 U9454 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_f114), .A(n7753), .ZN(n7758) );
  AOI22_X1 U9455 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_f113), .ZN(n7754) );
  OAI221_X1 U9456 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_f113), .A(n7754), .ZN(n7757) );
  AOI22_X1 U9457 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_B_REG_SCAN_IN), .B2(
        keyinput_f64), .ZN(n7755) );
  OAI221_X1 U9458 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P2_B_REG_SCAN_IN), .C2(
        keyinput_f64), .A(n7755), .ZN(n7756) );
  NOR4_X1 U9459 ( .A1(n7759), .A2(n7758), .A3(n7757), .A4(n7756), .ZN(n7760)
         );
  NAND4_X1 U9460 ( .A1(n7763), .A2(n7762), .A3(n7761), .A4(n7760), .ZN(n7871)
         );
  AOI22_X1 U9461 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput_f127), .ZN(n7764) );
  OAI221_X1 U9462 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput_f127), .A(n7764), .ZN(n7773) );
  AOI22_X1 U9463 ( .A1(SI_14_), .A2(keyinput_f18), .B1(P1_IR_REG_26__SCAN_IN), 
        .B2(keyinput_f117), .ZN(n7765) );
  OAI221_X1 U9464 ( .B1(SI_14_), .B2(keyinput_f18), .C1(P1_IR_REG_26__SCAN_IN), 
        .C2(keyinput_f117), .A(n7765), .ZN(n7772) );
  AOI22_X1 U9465 ( .A1(n6176), .A2(keyinput_f59), .B1(n7767), .B2(keyinput_f46), .ZN(n7766) );
  OAI221_X1 U9466 ( .B1(n6176), .B2(keyinput_f59), .C1(n7767), .C2(
        keyinput_f46), .A(n7766), .ZN(n7771) );
  INV_X1 U9467 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7769) );
  AOI22_X1 U9468 ( .A1(n7769), .A2(keyinput_f42), .B1(n7936), .B2(keyinput_f72), .ZN(n7768) );
  OAI221_X1 U9469 ( .B1(n7769), .B2(keyinput_f42), .C1(n7936), .C2(
        keyinput_f72), .A(n7768), .ZN(n7770) );
  NOR4_X1 U9470 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), .ZN(n7813)
         );
  AOI22_X1 U9471 ( .A1(n6046), .A2(keyinput_f3), .B1(n7775), .B2(keyinput_f86), 
        .ZN(n7774) );
  OAI221_X1 U9472 ( .B1(n6046), .B2(keyinput_f3), .C1(n7775), .C2(keyinput_f86), .A(n7774), .ZN(n7785) );
  AOI22_X1 U9473 ( .A1(n7778), .A2(keyinput_f96), .B1(keyinput_f8), .B2(n7777), 
        .ZN(n7776) );
  OAI221_X1 U9474 ( .B1(n7778), .B2(keyinput_f96), .C1(n7777), .C2(keyinput_f8), .A(n7776), .ZN(n7784) );
  XNOR2_X1 U9475 ( .A(SI_16_), .B(keyinput_f16), .ZN(n7782) );
  XNOR2_X1 U9476 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f95), .ZN(n7781) );
  XNOR2_X1 U9477 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_f121), .ZN(n7780) );
  XNOR2_X1 U9478 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n7779) );
  NAND4_X1 U9479 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n7783)
         );
  NOR3_X1 U9480 ( .A1(n7785), .A2(n7784), .A3(n7783), .ZN(n7812) );
  AOI22_X1 U9481 ( .A1(n8709), .A2(keyinput_f62), .B1(keyinput_f0), .B2(n10190), .ZN(n7786) );
  OAI221_X1 U9482 ( .B1(n8709), .B2(keyinput_f62), .C1(n10190), .C2(
        keyinput_f0), .A(n7786), .ZN(n7795) );
  INV_X1 U9483 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7788) );
  AOI22_X1 U9484 ( .A1(n8671), .A2(keyinput_f47), .B1(n7788), .B2(
        keyinput_f107), .ZN(n7787) );
  OAI221_X1 U9485 ( .B1(n8671), .B2(keyinput_f47), .C1(n7788), .C2(
        keyinput_f107), .A(n7787), .ZN(n7794) );
  INV_X1 U9486 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9024) );
  INV_X1 U9487 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U9488 ( .A1(n9024), .A2(keyinput_f60), .B1(keyinput_f67), .B2(
        n10087), .ZN(n7789) );
  OAI221_X1 U9489 ( .B1(n9024), .B2(keyinput_f60), .C1(n10087), .C2(
        keyinput_f67), .A(n7789), .ZN(n7793) );
  XNOR2_X1 U9490 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f105), .ZN(n7791) );
  XNOR2_X1 U9491 ( .A(SI_4_), .B(keyinput_f28), .ZN(n7790) );
  NAND2_X1 U9492 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  NOR4_X1 U9493 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n7811)
         );
  INV_X1 U9494 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7797) );
  AOI22_X1 U9495 ( .A1(n7797), .A2(keyinput_f94), .B1(keyinput_f56), .B2(n7348), .ZN(n7796) );
  OAI221_X1 U9496 ( .B1(n7797), .B2(keyinput_f94), .C1(n7348), .C2(
        keyinput_f56), .A(n7796), .ZN(n7809) );
  AOI22_X1 U9497 ( .A1(n7800), .A2(keyinput_f102), .B1(keyinput_f17), .B2(
        n7799), .ZN(n7798) );
  OAI221_X1 U9498 ( .B1(n7800), .B2(keyinput_f102), .C1(n7799), .C2(
        keyinput_f17), .A(n7798), .ZN(n7808) );
  AOI22_X1 U9499 ( .A1(n7803), .A2(keyinput_f85), .B1(n7802), .B2(keyinput_f74), .ZN(n7801) );
  OAI221_X1 U9500 ( .B1(n7803), .B2(keyinput_f85), .C1(n7802), .C2(
        keyinput_f74), .A(n7801), .ZN(n7807) );
  XNOR2_X1 U9501 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_f120), .ZN(n7805) );
  XNOR2_X1 U9502 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f110), .ZN(n7804) );
  NAND2_X1 U9503 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  NOR4_X1 U9504 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n7810)
         );
  NAND4_X1 U9505 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n7870)
         );
  AOI22_X1 U9506 ( .A1(n7816), .A2(keyinput_f73), .B1(keyinput_f39), .B2(n7815), .ZN(n7814) );
  OAI221_X1 U9507 ( .B1(n7816), .B2(keyinput_f73), .C1(n7815), .C2(
        keyinput_f39), .A(n7814), .ZN(n7826) );
  INV_X1 U9508 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7818) );
  INV_X1 U9509 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8689) );
  AOI22_X1 U9510 ( .A1(n7818), .A2(keyinput_f109), .B1(keyinput_f55), .B2(
        n8689), .ZN(n7817) );
  OAI221_X1 U9511 ( .B1(n7818), .B2(keyinput_f109), .C1(n8689), .C2(
        keyinput_f55), .A(n7817), .ZN(n7825) );
  XOR2_X1 U9512 ( .A(n7819), .B(keyinput_f65), .Z(n7823) );
  XNOR2_X1 U9513 ( .A(SI_12_), .B(keyinput_f20), .ZN(n7822) );
  XNOR2_X1 U9514 ( .A(SI_2_), .B(keyinput_f30), .ZN(n7821) );
  XNOR2_X1 U9515 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7820) );
  NAND4_X1 U9516 ( .A1(n7823), .A2(n7822), .A3(n7821), .A4(n7820), .ZN(n7824)
         );
  NOR3_X1 U9517 ( .A1(n7826), .A2(n7825), .A3(n7824), .ZN(n7868) );
  AOI22_X1 U9518 ( .A1(n10310), .A2(keyinput_f125), .B1(keyinput_f22), .B2(
        n7828), .ZN(n7827) );
  OAI221_X1 U9519 ( .B1(n10310), .B2(keyinput_f125), .C1(n7828), .C2(
        keyinput_f22), .A(n7827), .ZN(n7839) );
  INV_X1 U9520 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8612) );
  AOI22_X1 U9521 ( .A1(n8612), .A2(keyinput_f36), .B1(keyinput_f37), .B2(n7830), .ZN(n7829) );
  OAI221_X1 U9522 ( .B1(n8612), .B2(keyinput_f36), .C1(n7830), .C2(
        keyinput_f37), .A(n7829), .ZN(n7838) );
  AOI22_X1 U9523 ( .A1(n7833), .A2(keyinput_f90), .B1(n7832), .B2(keyinput_f84), .ZN(n7831) );
  OAI221_X1 U9524 ( .B1(n7833), .B2(keyinput_f90), .C1(n7832), .C2(
        keyinput_f84), .A(n7831), .ZN(n7837) );
  XNOR2_X1 U9525 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f116), .ZN(n7835) );
  XNOR2_X1 U9526 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_f88), .ZN(n7834)
         );
  NAND2_X1 U9527 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  NOR4_X1 U9528 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .ZN(n7867)
         );
  AOI22_X1 U9529 ( .A1(n7841), .A2(keyinput_f77), .B1(keyinput_f49), .B2(n6223), .ZN(n7840) );
  OAI221_X1 U9530 ( .B1(n7841), .B2(keyinput_f77), .C1(n6223), .C2(
        keyinput_f49), .A(n7840), .ZN(n7850) );
  AOI22_X1 U9531 ( .A1(n8151), .A2(keyinput_f71), .B1(keyinput_f54), .B2(n6159), .ZN(n7842) );
  OAI221_X1 U9532 ( .B1(n8151), .B2(keyinput_f71), .C1(n6159), .C2(
        keyinput_f54), .A(n7842), .ZN(n7849) );
  INV_X1 U9533 ( .A(SI_7_), .ZN(n7844) );
  AOI22_X1 U9534 ( .A1(n7844), .A2(keyinput_f25), .B1(keyinput_f38), .B2(n8645), .ZN(n7843) );
  OAI221_X1 U9535 ( .B1(n7844), .B2(keyinput_f25), .C1(n8645), .C2(
        keyinput_f38), .A(n7843), .ZN(n7848) );
  XNOR2_X1 U9536 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_f104), .ZN(n7846) );
  XNOR2_X1 U9537 ( .A(SI_19_), .B(keyinput_f13), .ZN(n7845) );
  NAND2_X1 U9538 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  NOR4_X1 U9539 ( .A1(n7850), .A2(n7849), .A3(n7848), .A4(n7847), .ZN(n7866)
         );
  INV_X1 U9540 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7853) );
  AOI22_X1 U9541 ( .A1(n7853), .A2(keyinput_f93), .B1(keyinput_f76), .B2(n7852), .ZN(n7851) );
  OAI221_X1 U9542 ( .B1(n7853), .B2(keyinput_f93), .C1(n7852), .C2(
        keyinput_f76), .A(n7851), .ZN(n7864) );
  AOI22_X1 U9543 ( .A1(n7856), .A2(keyinput_f79), .B1(keyinput_f87), .B2(n7855), .ZN(n7854) );
  OAI221_X1 U9544 ( .B1(n7856), .B2(keyinput_f79), .C1(n7855), .C2(
        keyinput_f87), .A(n7854), .ZN(n7863) );
  AOI22_X1 U9545 ( .A1(n7858), .A2(keyinput_f82), .B1(n8096), .B2(keyinput_f70), .ZN(n7857) );
  OAI221_X1 U9546 ( .B1(n7858), .B2(keyinput_f82), .C1(n8096), .C2(
        keyinput_f70), .A(n7857), .ZN(n7862) );
  XNOR2_X1 U9547 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f91), .ZN(n7860) );
  XNOR2_X1 U9548 ( .A(SI_3_), .B(keyinput_f29), .ZN(n7859) );
  NAND2_X1 U9549 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  NOR4_X1 U9550 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n7865)
         );
  NAND4_X1 U9551 ( .A1(n7868), .A2(n7867), .A3(n7866), .A4(n7865), .ZN(n7869)
         );
  NOR4_X1 U9552 ( .A1(n7872), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n7912)
         );
  OAI22_X1 U9553 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        keyinput_f35), .B2(P2_REG3_REG_7__SCAN_IN), .ZN(n7873) );
  AOI221_X1 U9554 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n7873), .ZN(n7880) );
  OAI22_X1 U9555 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_f106), .B1(
        keyinput_f58), .B2(P2_REG3_REG_11__SCAN_IN), .ZN(n7874) );
  AOI221_X1 U9556 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_f106), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n7874), .ZN(n7879) );
  OAI22_X1 U9557 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_f122), .B1(
        keyinput_f112), .B2(P1_IR_REG_21__SCAN_IN), .ZN(n7875) );
  AOI221_X1 U9558 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_f122), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_f112), .A(n7875), .ZN(n7878) );
  OAI22_X1 U9559 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n7876) );
  AOI221_X1 U9560 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        keyinput_f52), .C2(P2_REG3_REG_4__SCAN_IN), .A(n7876), .ZN(n7877) );
  NAND4_X1 U9561 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n7908)
         );
  OAI22_X1 U9562 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f111), .B1(
        keyinput_f81), .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7881) );
  AOI221_X1 U9563 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f111), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n7881), .ZN(n7888) );
  OAI22_X1 U9564 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f101), .B1(SI_23_), 
        .B2(keyinput_f9), .ZN(n7882) );
  AOI221_X1 U9565 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f9), .C2(SI_23_), .A(n7882), .ZN(n7887) );
  OAI22_X1 U9566 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f98), .B1(
        keyinput_f4), .B2(SI_28_), .ZN(n7883) );
  AOI221_X1 U9567 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f98), .C1(SI_28_), 
        .C2(keyinput_f4), .A(n7883), .ZN(n7886) );
  OAI22_X1 U9568 ( .A1(SI_21_), .A2(keyinput_f11), .B1(keyinput_f40), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7884) );
  AOI221_X1 U9569 ( .B1(SI_21_), .B2(keyinput_f11), .C1(P2_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n7884), .ZN(n7885) );
  NAND4_X1 U9570 ( .A1(n7888), .A2(n7887), .A3(n7886), .A4(n7885), .ZN(n7907)
         );
  OAI22_X1 U9571 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f108), .B1(
        keyinput_f21), .B2(SI_11_), .ZN(n7889) );
  AOI221_X1 U9572 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f108), .C1(SI_11_), .C2(keyinput_f21), .A(n7889), .ZN(n7896) );
  OAI22_X1 U9573 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_f123), .B1(
        keyinput_f48), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n7890) );
  AOI221_X1 U9574 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_f123), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n7890), .ZN(n7895) );
  OAI22_X1 U9575 ( .A1(SI_27_), .A2(keyinput_f5), .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .ZN(n7891) );
  AOI221_X1 U9576 ( .B1(SI_27_), .B2(keyinput_f5), .C1(keyinput_f66), .C2(
        P2_DATAO_REG_30__SCAN_IN), .A(n7891), .ZN(n7894) );
  OAI22_X1 U9577 ( .A1(SI_0_), .A2(keyinput_f32), .B1(keyinput_f45), .B2(
        P2_REG3_REG_21__SCAN_IN), .ZN(n7892) );
  AOI221_X1 U9578 ( .B1(SI_0_), .B2(keyinput_f32), .C1(P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n7892), .ZN(n7893) );
  NAND4_X1 U9579 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n7906)
         );
  OAI22_X1 U9580 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f103), .B1(SI_13_), 
        .B2(keyinput_f19), .ZN(n7897) );
  AOI221_X1 U9581 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f103), .C1(
        keyinput_f19), .C2(SI_13_), .A(n7897), .ZN(n7904) );
  OAI22_X1 U9582 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f92), .B1(
        keyinput_f83), .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7898) );
  AOI221_X1 U9583 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f92), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n7898), .ZN(n7903) );
  OAI22_X1 U9584 ( .A1(SI_22_), .A2(keyinput_f10), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n7899) );
  AOI221_X1 U9585 ( .B1(SI_22_), .B2(keyinput_f10), .C1(keyinput_f26), .C2(
        SI_6_), .A(n7899), .ZN(n7902) );
  OAI22_X1 U9586 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f119), .B1(SI_5_), 
        .B2(keyinput_f27), .ZN(n7900) );
  AOI221_X1 U9587 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f119), .C1(
        keyinput_f27), .C2(SI_5_), .A(n7900), .ZN(n7901) );
  NAND4_X1 U9588 ( .A1(n7904), .A2(n7903), .A3(n7902), .A4(n7901), .ZN(n7905)
         );
  NOR4_X1 U9589 ( .A1(n7908), .A2(n7907), .A3(n7906), .A4(n7905), .ZN(n7911)
         );
  XNOR2_X1 U9590 ( .A(n7909), .B(keyinput_f115), .ZN(n7910) );
  AOI21_X1 U9591 ( .B1(n7912), .B2(n7911), .A(n7910), .ZN(n7913) );
  AOI211_X1 U9592 ( .C1(n7916), .C2(n7915), .A(n7914), .B(n7913), .ZN(n7918)
         );
  XNOR2_X1 U9593 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7917) );
  XNOR2_X1 U9594 ( .A(n7918), .B(n7917), .ZN(n7919) );
  XNOR2_X1 U9595 ( .A(n7920), .B(n7919), .ZN(ADD_1071_U4) );
  INV_X1 U9596 ( .A(n8575), .ZN(n7937) );
  AOI22_X1 U9597 ( .A1(n7921), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9471), .ZN(n7922) );
  OAI21_X1 U9598 ( .B1(n7937), .B2(n9463), .A(n7922), .ZN(P2_U3334) );
  NAND2_X1 U9599 ( .A1(n7924), .A2(n4771), .ZN(n7925) );
  NAND2_X1 U9600 ( .A1(n7964), .A2(n7955), .ZN(n8804) );
  NAND2_X1 U9601 ( .A1(n8817), .A2(n8804), .ZN(n8897) );
  XNOR2_X1 U9602 ( .A(n7950), .B(n8897), .ZN(n7973) );
  INV_X1 U9603 ( .A(n8799), .ZN(n8801) );
  NOR2_X1 U9604 ( .A1(n8909), .A2(n8801), .ZN(n7927) );
  XNOR2_X1 U9605 ( .A(n7952), .B(n8897), .ZN(n7929) );
  INV_X1 U9606 ( .A(n8017), .ZN(n8939) );
  AOI222_X1 U9607 ( .A1(n10365), .A2(n7929), .B1(n4771), .B2(n10360), .C1(
        n8939), .C2(n10362), .ZN(n7968) );
  AOI21_X1 U9608 ( .B1(n7964), .B2(n7930), .A(n4503), .ZN(n7971) );
  AOI22_X1 U9609 ( .A1(n7971), .A2(n10411), .B1(n9437), .B2(n7964), .ZN(n7931)
         );
  OAI211_X1 U9610 ( .C1(n7973), .C2(n10426), .A(n7968), .B(n7931), .ZN(n7933)
         );
  NAND2_X1 U9611 ( .A1(n7933), .A2(n10455), .ZN(n7932) );
  OAI21_X1 U9612 ( .B1(n10455), .B2(n7276), .A(n7932), .ZN(P2_U3531) );
  INV_X1 U9613 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U9614 ( .A1(n7933), .A2(n10444), .ZN(n7934) );
  OAI21_X1 U9615 ( .B1(n10444), .B2(n7935), .A(n7934), .ZN(P2_U3484) );
  OAI222_X1 U9616 ( .A1(n7938), .A2(P1_U3084), .B1(n10090), .B2(n7937), .C1(
        n7936), .C2(n10100), .ZN(P1_U3329) );
  XOR2_X1 U9617 ( .A(n7939), .B(n8458), .Z(n7976) );
  INV_X1 U9618 ( .A(n7976), .ZN(n7949) );
  NAND2_X1 U9619 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  XOR2_X1 U9620 ( .A(n8458), .B(n7942), .Z(n7943) );
  OAI222_X1 U9621 ( .A1(n9959), .A2(n9495), .B1(n9957), .B2(n7992), .C1(n10128), .C2(n7943), .ZN(n7974) );
  INV_X1 U9622 ( .A(n7994), .ZN(n7946) );
  AOI211_X1 U9623 ( .C1(n7994), .C2(n10141), .A(n10313), .B(n10120), .ZN(n7975) );
  NAND2_X1 U9624 ( .A1(n7975), .A2(n9963), .ZN(n7945) );
  AOI22_X1 U9625 ( .A1(n10157), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7989), .B2(
        n10155), .ZN(n7944) );
  OAI211_X1 U9626 ( .C1(n7946), .C2(n10159), .A(n7945), .B(n7944), .ZN(n7947)
         );
  AOI21_X1 U9627 ( .B1(n7974), .B2(n10161), .A(n7947), .ZN(n7948) );
  OAI21_X1 U9628 ( .B1(n7949), .B2(n9969), .A(n7948), .ZN(P1_U3279) );
  NAND2_X1 U9629 ( .A1(n7964), .A2(n8940), .ZN(n7951) );
  NAND2_X1 U9630 ( .A1(n8010), .A2(n8017), .ZN(n8819) );
  XNOR2_X1 U9631 ( .A(n8011), .B(n8911), .ZN(n10441) );
  INV_X1 U9632 ( .A(n10441), .ZN(n7963) );
  NAND2_X1 U9633 ( .A1(n8014), .A2(n8804), .ZN(n7953) );
  XOR2_X1 U9634 ( .A(n8911), .B(n7953), .Z(n7954) );
  OAI222_X1 U9635 ( .A1(n9311), .A2(n8012), .B1(n9309), .B2(n7955), .C1(n7954), 
        .C2(n9293), .ZN(n10438) );
  INV_X1 U9636 ( .A(n8010), .ZN(n10435) );
  INV_X1 U9637 ( .A(n8026), .ZN(n7956) );
  OAI21_X1 U9638 ( .B1(n10435), .B2(n4503), .A(n7956), .ZN(n10437) );
  OAI22_X1 U9639 ( .A1(n10370), .A2(n7958), .B1(n7957), .B2(n10375), .ZN(n7959) );
  AOI21_X1 U9640 ( .B1(n8010), .B2(n9325), .A(n7959), .ZN(n7960) );
  OAI21_X1 U9641 ( .B1(n10437), .B2(n9321), .A(n7960), .ZN(n7961) );
  AOI21_X1 U9642 ( .B1(n10438), .B2(n10370), .A(n7961), .ZN(n7962) );
  OAI21_X1 U9643 ( .B1(n7963), .B2(n9349), .A(n7962), .ZN(P2_U3284) );
  INV_X1 U9644 ( .A(n7965), .ZN(n7966) );
  AOI22_X1 U9645 ( .A1(n10357), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7966), .B2(
        n9335), .ZN(n7967) );
  OAI21_X1 U9646 ( .B1(n4991), .B2(n9338), .A(n7967), .ZN(n7970) );
  NOR2_X1 U9647 ( .A1(n7968), .A2(n10357), .ZN(n7969) );
  AOI211_X1 U9648 ( .C1(n7971), .C2(n9347), .A(n7970), .B(n7969), .ZN(n7972)
         );
  OAI21_X1 U9649 ( .B1(n9349), .B2(n7973), .A(n7972), .ZN(P2_U3285) );
  AOI211_X1 U9650 ( .C1(n7976), .C2(n10332), .A(n7975), .B(n7974), .ZN(n7982)
         );
  INV_X1 U9651 ( .A(n10076), .ZN(n7979) );
  INV_X1 U9652 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7977) );
  NOR2_X1 U9653 ( .A1(n10336), .A2(n7977), .ZN(n7978) );
  AOI21_X1 U9654 ( .B1(n7994), .B2(n7979), .A(n7978), .ZN(n7980) );
  OAI21_X1 U9655 ( .B1(n7982), .B2(n10334), .A(n7980), .ZN(P1_U3490) );
  AOI22_X1 U9656 ( .A1(n7994), .A2(n6029), .B1(n10341), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7981) );
  OAI21_X1 U9657 ( .B1(n7982), .B2(n10341), .A(n7981), .ZN(P1_U3535) );
  INV_X1 U9658 ( .A(n7984), .ZN(n7985) );
  AOI21_X1 U9659 ( .B1(n7986), .B2(n7983), .A(n7985), .ZN(n7996) );
  INV_X1 U9660 ( .A(n9609), .ZN(n9646) );
  INV_X1 U9661 ( .A(n7987), .ZN(n7988) );
  AOI21_X1 U9662 ( .B1(n9640), .B2(n9661), .A(n7988), .ZN(n7991) );
  NAND2_X1 U9663 ( .A1(n9642), .A2(n7989), .ZN(n7990) );
  OAI211_X1 U9664 ( .C1(n9646), .C2(n7992), .A(n7991), .B(n7990), .ZN(n7993)
         );
  AOI21_X1 U9665 ( .B1(n7994), .B2(n9648), .A(n7993), .ZN(n7995) );
  OAI21_X1 U9666 ( .B1(n7996), .B2(n9651), .A(n7995), .ZN(P1_U3222) );
  INV_X1 U9667 ( .A(n7998), .ZN(n8000) );
  NAND2_X1 U9668 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  XNOR2_X1 U9669 ( .A(n7997), .B(n8001), .ZN(n8009) );
  INV_X1 U9670 ( .A(n8002), .ZN(n8003) );
  AOI21_X1 U9671 ( .B1(n9640), .B2(n10126), .A(n8003), .ZN(n8005) );
  NAND2_X1 U9672 ( .A1(n9642), .A2(n10132), .ZN(n8004) );
  OAI211_X1 U9673 ( .C1(n9646), .C2(n8006), .A(n8005), .B(n8004), .ZN(n8007)
         );
  AOI21_X1 U9674 ( .B1(n8250), .B2(n9612), .A(n8007), .ZN(n8008) );
  OAI21_X1 U9675 ( .B1(n8009), .B2(n9651), .A(n8008), .ZN(P1_U3232) );
  OR2_X1 U9676 ( .A1(n8141), .A2(n8012), .ZN(n8825) );
  NAND2_X1 U9677 ( .A1(n8141), .A2(n8012), .ZN(n8824) );
  OR2_X1 U9678 ( .A1(n9071), .A2(n9070), .ZN(n8047) );
  NAND2_X1 U9679 ( .A1(n9071), .A2(n9070), .ZN(n8013) );
  NAND2_X1 U9680 ( .A1(n8047), .A2(n8013), .ZN(n8144) );
  OR2_X1 U9681 ( .A1(n8144), .A2(n9313), .ZN(n8021) );
  AND2_X1 U9682 ( .A1(n8819), .A2(n8804), .ZN(n8823) );
  INV_X1 U9683 ( .A(n8818), .ZN(n8822) );
  NOR2_X1 U9684 ( .A1(n8015), .A2(n9070), .ZN(n8016) );
  OR2_X1 U9685 ( .A1(n8055), .A2(n8016), .ZN(n8019) );
  OAI22_X1 U9686 ( .A1(n8017), .A2(n9309), .B1(n8937), .B2(n9311), .ZN(n8018)
         );
  AOI21_X1 U9687 ( .B1(n8019), .B2(n10365), .A(n8018), .ZN(n8020) );
  NAND2_X1 U9688 ( .A1(n8021), .A2(n8020), .ZN(n8146) );
  OAI22_X1 U9689 ( .A1(n10370), .A2(n8023), .B1(n8022), .B2(n10375), .ZN(n8024) );
  AOI21_X1 U9690 ( .B1(n8141), .B2(n9325), .A(n8024), .ZN(n8029) );
  INV_X1 U9691 ( .A(n8141), .ZN(n8025) );
  OR2_X1 U9692 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  AND2_X1 U9693 ( .A1(n8050), .A2(n8027), .ZN(n8142) );
  NAND2_X1 U9694 ( .A1(n8142), .A2(n9347), .ZN(n8028) );
  OAI211_X1 U9695 ( .C1(n8144), .C2(n9328), .A(n8029), .B(n8028), .ZN(n8030)
         );
  AOI21_X1 U9696 ( .B1(n10370), .B2(n8146), .A(n8030), .ZN(n8031) );
  INV_X1 U9697 ( .A(n8031), .ZN(P2_U3283) );
  XNOR2_X1 U9698 ( .A(n8032), .B(n6005), .ZN(n8155) );
  INV_X1 U9699 ( .A(n8155), .ZN(n8044) );
  NAND2_X1 U9700 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  NAND3_X1 U9701 ( .A1(n8036), .A2(n10152), .A3(n8035), .ZN(n8038) );
  AOI22_X1 U9702 ( .A1(n10149), .A2(n9660), .B1(n9661), .B2(n10147), .ZN(n8037) );
  NAND2_X1 U9703 ( .A1(n8038), .A2(n8037), .ZN(n8153) );
  INV_X1 U9704 ( .A(n10122), .ZN(n8039) );
  AOI211_X1 U9705 ( .C1(n9497), .C2(n8039), .A(n10313), .B(n4542), .ZN(n8154)
         );
  NAND2_X1 U9706 ( .A1(n8154), .A2(n9963), .ZN(n8041) );
  AOI22_X1 U9707 ( .A1(n10157), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9492), .B2(
        n10155), .ZN(n8040) );
  OAI211_X1 U9708 ( .C1(n8161), .C2(n8122), .A(n8041), .B(n8040), .ZN(n8042)
         );
  AOI21_X1 U9709 ( .B1(n10161), .B2(n8153), .A(n8042), .ZN(n8043) );
  OAI21_X1 U9710 ( .B1(n8044), .B2(n9969), .A(n8043), .ZN(P1_U3277) );
  INV_X1 U9711 ( .A(n8586), .ZN(n8152) );
  AOI22_X1 U9712 ( .A1(n8045), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9471), .ZN(n8046) );
  OAI21_X1 U9713 ( .B1(n8152), .B2(n9463), .A(n8046), .ZN(P2_U3333) );
  NAND2_X1 U9714 ( .A1(n8141), .A2(n8938), .ZN(n9067) );
  NAND2_X1 U9715 ( .A1(n8047), .A2(n9067), .ZN(n8048) );
  NAND2_X1 U9716 ( .A1(n9436), .A2(n8937), .ZN(n8828) );
  XNOR2_X1 U9717 ( .A(n8048), .B(n9068), .ZN(n9439) );
  INV_X1 U9718 ( .A(n9333), .ZN(n8049) );
  AOI211_X1 U9719 ( .C1(n9436), .C2(n8050), .A(n10436), .B(n8049), .ZN(n9435)
         );
  INV_X1 U9720 ( .A(n9436), .ZN(n8052) );
  OAI22_X1 U9721 ( .A1(n8052), .A2(n9338), .B1(n10370), .B2(n8051), .ZN(n8053)
         );
  AOI21_X1 U9722 ( .B1(n9435), .B2(n9182), .A(n8053), .ZN(n8062) );
  INV_X1 U9723 ( .A(n8824), .ZN(n8054) );
  OAI211_X1 U9724 ( .C1(n8056), .C2(n8827), .A(n8718), .B(n10365), .ZN(n8058)
         );
  NAND2_X1 U9725 ( .A1(n8938), .A2(n10360), .ZN(n8057) );
  OAI211_X1 U9726 ( .C1(n9310), .C2(n9311), .A(n8058), .B(n8057), .ZN(n9434)
         );
  NOR2_X1 U9727 ( .A1(n10375), .A2(n8059), .ZN(n8060) );
  OAI21_X1 U9728 ( .B1(n9434), .B2(n8060), .A(n10370), .ZN(n8061) );
  OAI211_X1 U9729 ( .C1(n9439), .C2(n9349), .A(n8062), .B(n8061), .ZN(P2_U3282) );
  INV_X1 U9730 ( .A(n8493), .ZN(n8097) );
  AOI22_X1 U9731 ( .A1(n8063), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9471), .ZN(n8064) );
  OAI21_X1 U9732 ( .B1(n8097), .B2(n9463), .A(n8064), .ZN(P2_U3332) );
  NAND2_X1 U9733 ( .A1(n8065), .A2(n6262), .ZN(n8068) );
  AOI22_X1 U9734 ( .A1(n8622), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8066), .B2(
        n9011), .ZN(n8067) );
  XNOR2_X1 U9735 ( .A(n9324), .B(n8626), .ZN(n8069) );
  OR2_X1 U9736 ( .A1(n9295), .A2(n8625), .ZN(n8070) );
  NAND2_X1 U9737 ( .A1(n8069), .A2(n8070), .ZN(n8099) );
  INV_X1 U9738 ( .A(n8069), .ZN(n8072) );
  INV_X1 U9739 ( .A(n8070), .ZN(n8071) );
  NAND2_X1 U9740 ( .A1(n8072), .A2(n8071), .ZN(n8073) );
  NAND2_X1 U9741 ( .A1(n8099), .A2(n8073), .ZN(n8084) );
  NAND2_X1 U9742 ( .A1(n8075), .A2(n8074), .ZN(n8080) );
  INV_X1 U9743 ( .A(n8076), .ZN(n8078) );
  NAND2_X1 U9744 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  INV_X1 U9745 ( .A(n8100), .ZN(n8082) );
  AOI21_X1 U9746 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(n8095) );
  NAND2_X1 U9747 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8990) );
  OAI21_X1 U9748 ( .B1(n8710), .B2(n9317), .A(n8990), .ZN(n8093) );
  NAND2_X1 U9749 ( .A1(n8730), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8086) );
  NAND2_X1 U9750 ( .A1(n6174), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8085) );
  AND2_X1 U9751 ( .A1(n8086), .A2(n8085), .ZN(n8091) );
  NAND2_X1 U9752 ( .A1(n8087), .A2(n9009), .ZN(n8088) );
  AND2_X1 U9753 ( .A1(n8107), .A2(n8088), .ZN(n8106) );
  NAND2_X1 U9754 ( .A1(n8106), .A2(n8556), .ZN(n8090) );
  INV_X1 U9755 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9287) );
  OR2_X1 U9756 ( .A1(n4480), .A2(n9287), .ZN(n8089) );
  OAI22_X1 U9757 ( .A1(n8696), .A2(n9310), .B1(n9312), .B2(n8711), .ZN(n8092)
         );
  AOI211_X1 U9758 ( .C1(n9324), .C2(n8699), .A(n8093), .B(n8092), .ZN(n8094)
         );
  OAI21_X1 U9759 ( .B1(n8095), .B2(n4808), .A(n8094), .ZN(P2_U3228) );
  OAI222_X1 U9760 ( .A1(n8098), .A2(P1_U3084), .B1(n10090), .B2(n8097), .C1(
        n8096), .C2(n10086), .ZN(P1_U3327) );
  NAND2_X1 U9761 ( .A1(n8101), .A2(n6262), .ZN(n8105) );
  OAI22_X1 U9762 ( .A1(n6214), .A2(n8102), .B1(n8509), .B2(n9006), .ZN(n8103)
         );
  INV_X1 U9763 ( .A(n8103), .ZN(n8104) );
  XNOR2_X1 U9764 ( .A(n9420), .B(n8599), .ZN(n8162) );
  NOR2_X1 U9765 ( .A1(n9312), .A2(n8625), .ZN(n8163) );
  XNOR2_X1 U9766 ( .A(n8162), .B(n8163), .ZN(n8164) );
  XNOR2_X1 U9767 ( .A(n8165), .B(n8164), .ZN(n8116) );
  INV_X1 U9768 ( .A(n8106), .ZN(n9286) );
  OAI22_X1 U9769 ( .A1(n8710), .A2(n9286), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9009), .ZN(n8114) );
  NAND2_X1 U9770 ( .A1(n8107), .A2(n9024), .ZN(n8108) );
  NAND2_X1 U9771 ( .A1(n8172), .A2(n8108), .ZN(n9272) );
  OR2_X1 U9772 ( .A1(n9272), .A2(n6194), .ZN(n8112) );
  AOI22_X1 U9773 ( .A1(n6174), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n8730), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U9774 ( .A1(n4478), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8110) );
  OAI22_X1 U9775 ( .A1(n8696), .A2(n9295), .B1(n9296), .B2(n8711), .ZN(n8113)
         );
  AOI211_X1 U9776 ( .C1(n9420), .C2(n8699), .A(n8114), .B(n8113), .ZN(n8115)
         );
  OAI21_X1 U9777 ( .B1(n8116), .B2(n4808), .A(n8115), .ZN(P2_U3230) );
  INV_X1 U9778 ( .A(n8261), .ZN(n8461) );
  XNOR2_X1 U9779 ( .A(n8117), .B(n8461), .ZN(n10169) );
  INV_X1 U9780 ( .A(n10169), .ZN(n8126) );
  XNOR2_X1 U9781 ( .A(n8118), .B(n8261), .ZN(n8119) );
  OAI222_X1 U9782 ( .A1(n9959), .A2(n9558), .B1(n9957), .B2(n9645), .C1(n10128), .C2(n8119), .ZN(n10167) );
  OAI21_X1 U9783 ( .B1(n4542), .B2(n10165), .A(n9961), .ZN(n10166) );
  NOR2_X1 U9784 ( .A1(n10166), .A2(n8120), .ZN(n8124) );
  AOI22_X1 U9785 ( .A1(n10157), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9641), .B2(
        n10155), .ZN(n8121) );
  OAI21_X1 U9786 ( .B1(n10165), .B2(n8122), .A(n8121), .ZN(n8123) );
  AOI211_X1 U9787 ( .C1(n10167), .C2(n10161), .A(n8124), .B(n8123), .ZN(n8125)
         );
  OAI21_X1 U9788 ( .B1(n8126), .B2(n9969), .A(n8125), .ZN(P1_U3276) );
  NOR2_X1 U9789 ( .A1(n8133), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8128) );
  NOR2_X1 U9790 ( .A1(n8128), .A2(n8127), .ZN(n8993) );
  XNOR2_X1 U9791 ( .A(n8993), .B(n8994), .ZN(n8129) );
  NOR2_X1 U9792 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8129), .ZN(n8995) );
  AOI21_X1 U9793 ( .B1(n8129), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8995), .ZN(
        n8140) );
  INV_X1 U9794 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8131) );
  OR2_X1 U9795 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6133), .ZN(n8130) );
  OAI21_X1 U9796 ( .B1(n9056), .B2(n8131), .A(n8130), .ZN(n8138) );
  NOR2_X1 U9797 ( .A1(n8135), .A2(n8136), .ZN(n8984) );
  AOI211_X1 U9798 ( .C1(n8136), .C2(n8135), .A(n8984), .B(n8134), .ZN(n8137)
         );
  AOI211_X1 U9799 ( .C1(n10347), .C2(n8994), .A(n8138), .B(n8137), .ZN(n8139)
         );
  OAI21_X1 U9800 ( .B1(n8140), .B2(n9048), .A(n8139), .ZN(P2_U3260) );
  AOI22_X1 U9801 ( .A1(n8142), .A2(n10411), .B1(n9437), .B2(n8141), .ZN(n8143)
         );
  OAI21_X1 U9802 ( .B1(n8144), .B2(n10418), .A(n8143), .ZN(n8145) );
  NOR2_X1 U9803 ( .A1(n8146), .A2(n8145), .ZN(n8148) );
  MUX2_X1 U9804 ( .A(n6363), .B(n8148), .S(n10455), .Z(n8147) );
  INV_X1 U9805 ( .A(n8147), .ZN(P2_U3533) );
  INV_X1 U9806 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U9807 ( .A(n8149), .B(n8148), .S(n10444), .Z(n8150) );
  INV_X1 U9808 ( .A(n8150), .ZN(P2_U3490) );
  OAI222_X1 U9809 ( .A1(P1_U3084), .A2(n5895), .B1(n10090), .B2(n8152), .C1(
        n8151), .C2(n10086), .ZN(P1_U3328) );
  INV_X1 U9810 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8156) );
  AOI211_X1 U9811 ( .C1(n8155), .C2(n10332), .A(n8154), .B(n8153), .ZN(n8158)
         );
  MUX2_X1 U9812 ( .A(n8156), .B(n8158), .S(n10336), .Z(n8157) );
  OAI21_X1 U9813 ( .B1(n8161), .B2(n10076), .A(n8157), .ZN(P1_U3496) );
  MUX2_X1 U9814 ( .A(n8159), .B(n8158), .S(n10344), .Z(n8160) );
  OAI21_X1 U9815 ( .B1(n8161), .B2(n10042), .A(n8160), .ZN(P1_U3537) );
  NAND2_X1 U9816 ( .A1(n8166), .A2(n6262), .ZN(n8170) );
  OAI22_X1 U9817 ( .A1(n6214), .A2(n8167), .B1(n8509), .B2(n9042), .ZN(n8168)
         );
  INV_X1 U9818 ( .A(n8168), .ZN(n8169) );
  XNOR2_X1 U9819 ( .A(n9413), .B(n8626), .ZN(n8505) );
  NOR2_X1 U9820 ( .A1(n9296), .A2(n8625), .ZN(n8506) );
  XNOR2_X1 U9821 ( .A(n8505), .B(n8506), .ZN(n8503) );
  XNOR2_X1 U9822 ( .A(n8504), .B(n8503), .ZN(n8182) );
  OAI22_X1 U9823 ( .A1(n8710), .A2(n9272), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9024), .ZN(n8180) );
  NAND2_X1 U9824 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  AND2_X1 U9825 ( .A1(n8523), .A2(n8173), .ZN(n8654) );
  NAND2_X1 U9826 ( .A1(n8654), .A2(n8556), .ZN(n8178) );
  INV_X1 U9827 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U9828 ( .A1(n6174), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U9829 ( .A1(n8730), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8174) );
  OAI211_X1 U9830 ( .C1(n9256), .C2(n4480), .A(n8175), .B(n8174), .ZN(n8176)
         );
  INV_X1 U9831 ( .A(n8176), .ZN(n8177) );
  OAI22_X1 U9832 ( .A1(n8696), .A2(n9312), .B1(n9076), .B2(n8711), .ZN(n8179)
         );
  AOI211_X1 U9833 ( .C1(n9413), .C2(n8699), .A(n8180), .B(n8179), .ZN(n8181)
         );
  OAI21_X1 U9834 ( .B1(n8182), .B2(n4808), .A(n8181), .ZN(P2_U3240) );
  OAI22_X1 U9835 ( .A1(n8183), .A2(n8502), .B1(n4808), .B2(n8762), .ZN(n8185)
         );
  NAND2_X1 U9836 ( .A1(n8185), .A2(n8184), .ZN(n8188) );
  AOI22_X1 U9837 ( .A1(n8699), .A2(n10387), .B1(n8186), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n8187) );
  OAI211_X1 U9838 ( .C1(n8189), .C2(n8711), .A(n8188), .B(n8187), .ZN(P2_U3234) );
  NAND2_X1 U9839 ( .A1(n8190), .A2(n8480), .ZN(n8476) );
  NOR2_X1 U9840 ( .A1(n8192), .A2(SI_29_), .ZN(n8194) );
  NAND2_X1 U9841 ( .A1(n8192), .A2(SI_29_), .ZN(n8193) );
  MUX2_X1 U9842 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8204), .Z(n8200) );
  NAND2_X1 U9843 ( .A1(n4483), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U9844 ( .A1(n8405), .A2(n9748), .ZN(n8210) );
  INV_X1 U9845 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U9846 ( .A1(n8199), .A2(SI_30_), .ZN(n8203) );
  NAND2_X1 U9847 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  NAND2_X1 U9848 ( .A1(n8203), .A2(n8202), .ZN(n8207) );
  MUX2_X1 U9849 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8204), .Z(n8205) );
  XNOR2_X1 U9850 ( .A(n8205), .B(SI_31_), .ZN(n8206) );
  NAND2_X1 U9851 ( .A1(n9457), .A2(n5363), .ZN(n8209) );
  NAND2_X1 U9852 ( .A1(n4482), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U9853 ( .A1(n8210), .A2(n8324), .ZN(n8435) );
  INV_X1 U9854 ( .A(n8408), .ZN(n9653) );
  NAND2_X1 U9855 ( .A1(n9653), .A2(n9748), .ZN(n8211) );
  NAND2_X1 U9856 ( .A1(n9755), .A2(n8211), .ZN(n8430) );
  INV_X1 U9857 ( .A(n8326), .ZN(n8212) );
  AOI21_X1 U9858 ( .B1(n8328), .B2(n9654), .A(n8212), .ZN(n8330) );
  NAND3_X1 U9859 ( .A1(n8214), .A2(n8328), .A3(n8415), .ZN(n8215) );
  NAND2_X1 U9860 ( .A1(n8216), .A2(n8215), .ZN(n8224) );
  NAND2_X1 U9861 ( .A1(n8415), .A2(n8416), .ZN(n8217) );
  OAI21_X1 U9862 ( .B1(n8224), .B2(n8217), .A(n8420), .ZN(n8218) );
  INV_X1 U9863 ( .A(n8219), .ZN(n8453) );
  AND2_X1 U9864 ( .A1(n8225), .A2(n8220), .ZN(n8375) );
  AOI21_X1 U9865 ( .B1(n8223), .B2(n8375), .A(n8221), .ZN(n8229) );
  NAND3_X1 U9866 ( .A1(n8421), .A2(n8420), .A3(n8222), .ZN(n8364) );
  INV_X1 U9867 ( .A(n8225), .ZN(n8226) );
  AOI21_X1 U9868 ( .B1(n8227), .B2(n8369), .A(n8226), .ZN(n8228) );
  MUX2_X1 U9869 ( .A(n8229), .B(n8228), .S(n8328), .Z(n8241) );
  INV_X1 U9870 ( .A(n8368), .ZN(n8230) );
  NOR2_X1 U9871 ( .A1(n8232), .A2(n8230), .ZN(n8235) );
  OR2_X1 U9872 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  AND2_X1 U9873 ( .A1(n8233), .A2(n8245), .ZN(n8377) );
  NAND2_X1 U9874 ( .A1(n8254), .A2(n8377), .ZN(n8234) );
  AOI21_X1 U9875 ( .B1(n8241), .B2(n8235), .A(n8234), .ZN(n8237) );
  MUX2_X1 U9876 ( .A(n8237), .B(n8236), .S(n8328), .Z(n8249) );
  NAND2_X1 U9877 ( .A1(n8258), .A2(n8238), .ZN(n8387) );
  XNOR2_X1 U9878 ( .A(n10140), .B(n9662), .ZN(n10145) );
  NAND2_X1 U9879 ( .A1(n8379), .A2(n10145), .ZN(n8239) );
  NOR2_X1 U9880 ( .A1(n8387), .A2(n8239), .ZN(n8248) );
  NAND2_X1 U9881 ( .A1(n8241), .A2(n8240), .ZN(n8243) );
  NAND3_X1 U9882 ( .A1(n8243), .A2(n8242), .A3(n8368), .ZN(n8246) );
  NAND4_X1 U9883 ( .A1(n8246), .A2(n8328), .A3(n8245), .A4(n8244), .ZN(n8247)
         );
  INV_X1 U9884 ( .A(n8387), .ZN(n8253) );
  NAND2_X1 U9885 ( .A1(n8379), .A2(n8328), .ZN(n8251) );
  OR2_X1 U9886 ( .A1(n8250), .A2(n9495), .ZN(n8378) );
  OAI21_X1 U9887 ( .B1(n8381), .B2(n8251), .A(n8378), .ZN(n8252) );
  NAND2_X1 U9888 ( .A1(n8253), .A2(n8252), .ZN(n8257) );
  NAND2_X1 U9889 ( .A1(n8387), .A2(n4684), .ZN(n8256) );
  NAND2_X1 U9890 ( .A1(n8379), .A2(n4504), .ZN(n8376) );
  NAND3_X1 U9891 ( .A1(n8376), .A2(n4684), .A3(n8254), .ZN(n8255) );
  NAND2_X1 U9892 ( .A1(n8386), .A2(n8378), .ZN(n8259) );
  NAND3_X1 U9893 ( .A1(n8259), .A2(n4684), .A3(n8258), .ZN(n8260) );
  NAND2_X1 U9894 ( .A1(n8391), .A2(n8389), .ZN(n8263) );
  INV_X1 U9895 ( .A(n8394), .ZN(n8262) );
  MUX2_X1 U9896 ( .A(n8263), .B(n8262), .S(n8328), .Z(n8267) );
  INV_X1 U9897 ( .A(n8264), .ZN(n8268) );
  MUX2_X1 U9898 ( .A(n8265), .B(n8391), .S(n8328), .Z(n8266) );
  NAND2_X1 U9899 ( .A1(n8275), .A2(n8268), .ZN(n8392) );
  NAND2_X1 U9900 ( .A1(n8272), .A2(n8269), .ZN(n8343) );
  MUX2_X1 U9901 ( .A(n8392), .B(n8343), .S(n8328), .Z(n8270) );
  INV_X1 U9902 ( .A(n8270), .ZN(n8271) );
  AND2_X1 U9903 ( .A1(n8276), .A2(n8272), .ZN(n8274) );
  NAND2_X1 U9904 ( .A1(n9878), .A2(n8398), .ZN(n8273) );
  AOI21_X1 U9905 ( .B1(n8277), .B2(n8274), .A(n8273), .ZN(n8279) );
  AND2_X1 U9906 ( .A1(n8398), .A2(n8275), .ZN(n8344) );
  NAND2_X1 U9907 ( .A1(n8284), .A2(n8276), .ZN(n8345) );
  AOI21_X1 U9908 ( .B1(n8277), .B2(n8344), .A(n8345), .ZN(n8278) );
  MUX2_X1 U9909 ( .A(n8279), .B(n8278), .S(n8328), .Z(n8286) );
  AND2_X1 U9910 ( .A1(n8443), .A2(n8280), .ZN(n8342) );
  INV_X1 U9911 ( .A(n9878), .ZN(n8444) );
  NAND2_X1 U9912 ( .A1(n8280), .A2(n8444), .ZN(n8281) );
  AND2_X1 U9913 ( .A1(n8281), .A2(n8285), .ZN(n8282) );
  NAND2_X1 U9914 ( .A1(n8442), .A2(n8282), .ZN(n8399) );
  NAND2_X1 U9915 ( .A1(n8399), .A2(n8443), .ZN(n8352) );
  NAND2_X1 U9916 ( .A1(n8352), .A2(n8291), .ZN(n8283) );
  AOI21_X1 U9917 ( .B1(n8286), .B2(n8342), .A(n8283), .ZN(n8290) );
  INV_X1 U9918 ( .A(n8284), .ZN(n8445) );
  OAI21_X1 U9919 ( .B1(n8286), .B2(n8445), .A(n8285), .ZN(n8287) );
  NAND2_X1 U9920 ( .A1(n8287), .A2(n8342), .ZN(n8289) );
  OR2_X1 U9921 ( .A1(n9832), .A2(n9848), .ZN(n8296) );
  INV_X1 U9922 ( .A(n8296), .ZN(n8288) );
  INV_X1 U9923 ( .A(n8291), .ZN(n8292) );
  NAND2_X1 U9924 ( .A1(n8296), .A2(n8292), .ZN(n8293) );
  AND2_X1 U9925 ( .A1(n8293), .A2(n8297), .ZN(n8294) );
  NAND2_X1 U9926 ( .A1(n8294), .A2(n8302), .ZN(n8400) );
  NAND2_X1 U9927 ( .A1(n8296), .A2(n8295), .ZN(n8350) );
  NAND2_X1 U9928 ( .A1(n8350), .A2(n8297), .ZN(n8298) );
  NAND2_X1 U9929 ( .A1(n9794), .A2(n8298), .ZN(n8299) );
  MUX2_X1 U9930 ( .A(n8400), .B(n8299), .S(n8328), .Z(n8300) );
  INV_X1 U9931 ( .A(n8300), .ZN(n8301) );
  OAI22_X1 U9932 ( .A1(n8312), .A2(n9801), .B1(n4684), .B2(n8302), .ZN(n8303)
         );
  NAND2_X1 U9933 ( .A1(n8303), .A2(n9812), .ZN(n8307) );
  NAND2_X1 U9934 ( .A1(n8441), .A2(n8304), .ZN(n8305) );
  MUX2_X1 U9935 ( .A(n10054), .B(n8305), .S(n4684), .Z(n8306) );
  NAND2_X1 U9936 ( .A1(n8307), .A2(n8306), .ZN(n8317) );
  NAND2_X1 U9937 ( .A1(n8333), .A2(n8308), .ZN(n8311) );
  OAI21_X1 U9938 ( .B1(n9812), .B2(n8309), .A(n8318), .ZN(n8310) );
  MUX2_X1 U9939 ( .A(n8311), .B(n8310), .S(n8328), .Z(n8315) );
  INV_X1 U9940 ( .A(n8312), .ZN(n8313) );
  NAND2_X1 U9941 ( .A1(n8467), .A2(n8313), .ZN(n8314) );
  NAND2_X1 U9942 ( .A1(n8315), .A2(n8314), .ZN(n8316) );
  NAND2_X1 U9943 ( .A1(n8317), .A2(n8316), .ZN(n8320) );
  MUX2_X1 U9944 ( .A(n8333), .B(n8318), .S(n4684), .Z(n8319) );
  NAND2_X1 U9945 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  NAND2_X1 U9946 ( .A1(n8321), .A2(n8466), .ZN(n8323) );
  MUX2_X1 U9947 ( .A(n8334), .B(n8331), .S(n4684), .Z(n8322) );
  NAND2_X1 U9948 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  OR2_X1 U9949 ( .A1(n8338), .A2(n8337), .ZN(n8332) );
  NAND2_X1 U9950 ( .A1(n8332), .A2(n8331), .ZN(n8341) );
  OAI211_X1 U9951 ( .C1(n8426), .C2(n8441), .A(n8334), .B(n8333), .ZN(n8335)
         );
  INV_X1 U9952 ( .A(n8335), .ZN(n8336) );
  OR2_X1 U9953 ( .A1(n8341), .A2(n8336), .ZN(n8340) );
  NAND2_X1 U9954 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  NAND2_X1 U9955 ( .A1(n8340), .A2(n8339), .ZN(n8432) );
  INV_X1 U9956 ( .A(n8432), .ZN(n8407) );
  INV_X1 U9957 ( .A(n8341), .ZN(n8434) );
  INV_X1 U9958 ( .A(n8342), .ZN(n8349) );
  INV_X1 U9959 ( .A(n8344), .ZN(n8347) );
  INV_X1 U9960 ( .A(n8345), .ZN(n8346) );
  OAI21_X1 U9961 ( .B1(n4618), .B2(n8347), .A(n8346), .ZN(n8348) );
  OR2_X1 U9962 ( .A1(n8349), .A2(n8348), .ZN(n8351) );
  AOI21_X1 U9963 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8354) );
  OAI21_X1 U9964 ( .B1(n8354), .B2(n8400), .A(n8353), .ZN(n8427) );
  INV_X1 U9965 ( .A(n8427), .ZN(n8404) );
  INV_X1 U9966 ( .A(n8355), .ZN(n8356) );
  OAI211_X1 U9967 ( .C1(n8357), .C2(n5949), .A(n8473), .B(n8356), .ZN(n8358)
         );
  NAND3_X1 U9968 ( .A1(n8359), .A2(n5995), .A3(n8358), .ZN(n8362) );
  INV_X1 U9969 ( .A(n8360), .ZN(n8418) );
  AOI21_X1 U9970 ( .B1(n8362), .B2(n8361), .A(n8418), .ZN(n8367) );
  AND2_X1 U9971 ( .A1(n8415), .A2(n8363), .ZN(n8414) );
  INV_X1 U9972 ( .A(n8414), .ZN(n8366) );
  INV_X1 U9973 ( .A(n8364), .ZN(n8365) );
  OAI21_X1 U9974 ( .B1(n8367), .B2(n8366), .A(n8365), .ZN(n8374) );
  INV_X1 U9975 ( .A(n8392), .ZN(n8373) );
  NAND3_X1 U9976 ( .A1(n8370), .A2(n8369), .A3(n8368), .ZN(n8371) );
  NOR3_X1 U9977 ( .A1(n8387), .A2(n8376), .A3(n8371), .ZN(n8372) );
  AND4_X1 U9978 ( .A1(n8373), .A2(n8372), .A3(n8389), .A4(n8391), .ZN(n8397)
         );
  INV_X1 U9979 ( .A(n8397), .ZN(n8425) );
  AOI21_X1 U9980 ( .B1(n8413), .B2(n8374), .A(n8425), .ZN(n8402) );
  INV_X1 U9981 ( .A(n8375), .ZN(n8396) );
  INV_X1 U9982 ( .A(n8376), .ZN(n8385) );
  INV_X1 U9983 ( .A(n8377), .ZN(n8384) );
  INV_X1 U9984 ( .A(n8378), .ZN(n8383) );
  INV_X1 U9985 ( .A(n8379), .ZN(n8380) );
  NOR2_X1 U9986 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  AOI211_X1 U9987 ( .C1(n8385), .C2(n8384), .A(n8383), .B(n8382), .ZN(n8388)
         );
  OAI21_X1 U9988 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8390) );
  NAND2_X1 U9989 ( .A1(n8390), .A2(n8389), .ZN(n8393) );
  AOI211_X1 U9990 ( .C1(n8394), .C2(n8393), .A(n4622), .B(n8392), .ZN(n8395)
         );
  AOI21_X1 U9991 ( .B1(n8397), .B2(n8396), .A(n8395), .ZN(n8423) );
  INV_X1 U9992 ( .A(n8423), .ZN(n8401) );
  NOR3_X1 U9993 ( .A1(n8400), .A2(n4907), .A3(n8399), .ZN(n8429) );
  OAI21_X1 U9994 ( .B1(n8402), .B2(n8401), .A(n8429), .ZN(n8403) );
  NAND4_X1 U9995 ( .A1(n8434), .A2(n8467), .A3(n8404), .A4(n8403), .ZN(n8406)
         );
  INV_X1 U9996 ( .A(n8405), .ZN(n8470) );
  AOI21_X1 U9997 ( .B1(n8407), .B2(n8406), .A(n8470), .ZN(n8411) );
  INV_X1 U9998 ( .A(n8483), .ZN(n8436) );
  NAND2_X1 U9999 ( .A1(n9755), .A2(n8408), .ZN(n8409) );
  NAND2_X1 U10000 ( .A1(n8436), .A2(n8409), .ZN(n8471) );
  INV_X1 U10001 ( .A(n8472), .ZN(n8410) );
  OAI21_X1 U10002 ( .B1(n8411), .B2(n8471), .A(n8410), .ZN(n8412) );
  XNOR2_X1 U10003 ( .A(n8412), .B(n9745), .ZN(n8479) );
  NAND3_X1 U10004 ( .A1(n7144), .A2(n8414), .A3(n8413), .ZN(n8422) );
  OAI211_X1 U10005 ( .C1(n8418), .C2(n8417), .A(n8416), .B(n8415), .ZN(n8419)
         );
  NAND4_X1 U10006 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n8424)
         );
  OAI21_X1 U10007 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8428) );
  AOI211_X1 U10008 ( .C1(n8429), .C2(n8428), .A(n8427), .B(n8426), .ZN(n8433)
         );
  INV_X1 U10009 ( .A(n8430), .ZN(n8431) );
  AOI211_X1 U10010 ( .C1(n8434), .C2(n8433), .A(n8432), .B(n8431), .ZN(n8438)
         );
  INV_X1 U10011 ( .A(n8435), .ZN(n8437) );
  OAI211_X1 U10012 ( .C1(n8438), .C2(n8437), .A(n8473), .B(n8436), .ZN(n8439)
         );
  NAND3_X1 U10013 ( .A1(n8439), .A2(n8480), .A3(n9745), .ZN(n8477) );
  OR2_X1 U10014 ( .A1(n9801), .A2(n9812), .ZN(n8440) );
  NAND2_X1 U10015 ( .A1(n8441), .A2(n8440), .ZN(n9797) );
  NAND2_X1 U10016 ( .A1(n8443), .A2(n8442), .ZN(n9862) );
  NOR2_X1 U10017 ( .A1(n8445), .A2(n8444), .ZN(n9889) );
  INV_X1 U10018 ( .A(n9942), .ZN(n9936) );
  NAND3_X1 U10019 ( .A1(n8448), .A2(n8447), .A3(n8446), .ZN(n8450) );
  NOR4_X1 U10020 ( .A1(n8450), .A2(n5957), .A3(n5992), .A4(n8449), .ZN(n8454)
         );
  NAND4_X1 U10021 ( .A1(n8454), .A2(n8453), .A3(n8452), .A4(n8451), .ZN(n8457)
         );
  NOR4_X1 U10022 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n8459)
         );
  NAND4_X1 U10023 ( .A1(n6005), .A2(n8459), .A3(n10145), .A4(n10124), .ZN(
        n8460) );
  NOR4_X1 U10024 ( .A1(n9936), .A2(n8461), .A3(n9954), .A4(n8460), .ZN(n8462)
         );
  NAND4_X1 U10025 ( .A1(n9889), .A2(n9903), .A3(n9931), .A4(n8462), .ZN(n8463)
         );
  NOR4_X1 U10026 ( .A1(n9797), .A2(n9809), .A3(n9826), .A4(n8464), .ZN(n8465)
         );
  NAND4_X1 U10027 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n8469)
         );
  NOR2_X1 U10028 ( .A1(n8474), .A2(n8473), .ZN(n8475) );
  OAI21_X1 U10029 ( .B1(n8480), .B2(n8479), .A(n8478), .ZN(n8481) );
  INV_X1 U10030 ( .A(n8481), .ZN(n8484) );
  NOR4_X1 U10031 ( .A1(n8486), .A2(n5932), .A3(n10207), .A4(n8485), .ZN(n8488)
         );
  OAI21_X1 U10032 ( .B1(n8489), .B2(n5919), .A(P1_B_REG_SCAN_IN), .ZN(n8487)
         );
  OAI22_X1 U10033 ( .A1(n8490), .A2(n8489), .B1(n8488), .B2(n8487), .ZN(
        P1_U3240) );
  NAND2_X1 U10034 ( .A1(n10096), .A2(n6262), .ZN(n8492) );
  NAND2_X1 U10035 ( .A1(n4485), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10036 ( .A1(n8493), .A2(n6262), .ZN(n8495) );
  NAND2_X1 U10037 ( .A1(n8622), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8494) );
  XNOR2_X1 U10038 ( .A(n9369), .B(n8626), .ZN(n8598) );
  NAND2_X1 U10039 ( .A1(n8591), .A2(n8709), .ZN(n8496) );
  NAND2_X1 U10040 ( .A1(n8613), .A2(n8496), .ZN(n9153) );
  INV_X1 U10041 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U10042 ( .A1(n6174), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U10043 ( .A1(n8730), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U10044 ( .C1(n9154), .C2(n4480), .A(n8498), .B(n8497), .ZN(n8499)
         );
  INV_X1 U10045 ( .A(n8499), .ZN(n8500) );
  INV_X1 U10046 ( .A(n8505), .ZN(n8507) );
  NAND2_X1 U10047 ( .A1(n8508), .A2(n6262), .ZN(n8513) );
  OAI22_X1 U10048 ( .A1(n6214), .A2(n8510), .B1(n9297), .B2(n8509), .ZN(n8511)
         );
  INV_X1 U10049 ( .A(n8511), .ZN(n8512) );
  XNOR2_X1 U10050 ( .A(n9263), .B(n8599), .ZN(n8514) );
  OR2_X1 U10051 ( .A1(n9076), .A2(n8625), .ZN(n8515) );
  NAND2_X1 U10052 ( .A1(n8514), .A2(n8515), .ZN(n8519) );
  INV_X1 U10053 ( .A(n8514), .ZN(n8517) );
  INV_X1 U10054 ( .A(n8515), .ZN(n8516) );
  NAND2_X1 U10055 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  NAND2_X1 U10056 ( .A1(n8519), .A2(n8518), .ZN(n8652) );
  NAND2_X1 U10057 ( .A1(n8520), .A2(n6262), .ZN(n8522) );
  NAND2_X1 U10058 ( .A1(n8622), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8521) );
  XNOR2_X1 U10059 ( .A(n9400), .B(n8599), .ZN(n8531) );
  NAND2_X1 U10060 ( .A1(n8523), .A2(n8689), .ZN(n8524) );
  NAND2_X1 U10061 ( .A1(n8536), .A2(n8524), .ZN(n9248) );
  OR2_X1 U10062 ( .A1(n9248), .A2(n6194), .ZN(n8529) );
  INV_X1 U10063 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U10064 ( .A1(n8730), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10065 ( .A1(n6174), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8525) );
  OAI211_X1 U10066 ( .C1(n9249), .C2(n4480), .A(n8526), .B(n8525), .ZN(n8527)
         );
  INV_X1 U10067 ( .A(n8527), .ZN(n8528) );
  NOR2_X1 U10068 ( .A1(n9237), .A2(n8625), .ZN(n8530) );
  XNOR2_X1 U10069 ( .A(n8531), .B(n8530), .ZN(n8687) );
  NAND2_X1 U10070 ( .A1(n8531), .A2(n8530), .ZN(n8532) );
  NAND2_X1 U10071 ( .A1(n8533), .A2(n6262), .ZN(n8535) );
  NAND2_X1 U10072 ( .A1(n8622), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8534) );
  XNOR2_X1 U10073 ( .A(n9394), .B(n8599), .ZN(n8545) );
  NAND2_X1 U10074 ( .A1(n8536), .A2(n8661), .ZN(n8537) );
  NAND2_X1 U10075 ( .A1(n8550), .A2(n8537), .ZN(n9229) );
  OR2_X1 U10076 ( .A1(n9229), .A2(n6194), .ZN(n8542) );
  INV_X1 U10077 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U10078 ( .A1(n8730), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10079 ( .A1(n6174), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8538) );
  OAI211_X1 U10080 ( .C1(n4480), .C2(n9230), .A(n8539), .B(n8538), .ZN(n8540)
         );
  INV_X1 U10081 ( .A(n8540), .ZN(n8541) );
  NAND2_X1 U10082 ( .A1(n8542), .A2(n8541), .ZN(n9242) );
  NAND2_X1 U10083 ( .A1(n9242), .A2(n8741), .ZN(n8543) );
  XNOR2_X1 U10084 ( .A(n8545), .B(n8543), .ZN(n8660) );
  INV_X1 U10085 ( .A(n8543), .ZN(n8544) );
  AND2_X1 U10086 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  AOI21_X1 U10087 ( .B1(n8659), .B2(n8660), .A(n8546), .ZN(n8559) );
  NAND2_X1 U10088 ( .A1(n8547), .A2(n6262), .ZN(n8549) );
  NAND2_X1 U10089 ( .A1(n8622), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8548) );
  XOR2_X1 U10090 ( .A(n8599), .B(n9388), .Z(n8558) );
  XNOR2_X1 U10091 ( .A(n8559), .B(n8558), .ZN(n8701) );
  INV_X1 U10092 ( .A(n8701), .ZN(n8557) );
  NAND2_X1 U10093 ( .A1(n8550), .A2(n8694), .ZN(n8551) );
  AND2_X1 U10094 ( .A1(n8564), .A2(n8551), .ZN(n9214) );
  INV_X1 U10095 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10096 ( .A1(n6174), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10097 ( .A1(n8730), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8552) );
  OAI211_X1 U10098 ( .C1(n8554), .C2(n4480), .A(n8553), .B(n8552), .ZN(n8555)
         );
  AOI21_X1 U10099 ( .B1(n9214), .B2(n8556), .A(n8555), .ZN(n9238) );
  INV_X1 U10100 ( .A(n9238), .ZN(n9207) );
  NAND2_X1 U10101 ( .A1(n8557), .A2(n5094), .ZN(n8704) );
  NAND2_X1 U10102 ( .A1(n8559), .A2(n8558), .ZN(n8560) );
  NAND2_X1 U10103 ( .A1(n8561), .A2(n6262), .ZN(n8563) );
  NAND2_X1 U10104 ( .A1(n8622), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8562) );
  XNOR2_X1 U10105 ( .A(n9383), .B(n8599), .ZN(n8573) );
  NAND2_X1 U10106 ( .A1(n8564), .A2(n8645), .ZN(n8565) );
  NAND2_X1 U10107 ( .A1(n8578), .A2(n8565), .ZN(n9196) );
  OR2_X1 U10108 ( .A1(n9196), .A2(n6194), .ZN(n8571) );
  INV_X1 U10109 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10110 ( .A1(n8730), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10111 ( .A1(n6174), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8566) );
  OAI211_X1 U10112 ( .C1(n4480), .C2(n8568), .A(n8567), .B(n8566), .ZN(n8569)
         );
  INV_X1 U10113 ( .A(n8569), .ZN(n8570) );
  NOR2_X1 U10114 ( .A1(n9081), .A2(n8625), .ZN(n8641) );
  INV_X1 U10115 ( .A(n8572), .ZN(n8574) );
  AOI22_X2 U10116 ( .A1(n8642), .A2(n8641), .B1(n8574), .B2(n8573), .ZN(n8585)
         );
  NAND2_X1 U10117 ( .A1(n8575), .A2(n6262), .ZN(n8577) );
  NAND2_X1 U10118 ( .A1(n8622), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U10119 ( .A1(n8578), .A2(n8681), .ZN(n8579) );
  NAND2_X1 U10120 ( .A1(n8589), .A2(n8579), .ZN(n9179) );
  OR2_X1 U10121 ( .A1(n9179), .A2(n6194), .ZN(n8584) );
  INV_X1 U10122 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U10123 ( .A1(n6174), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10124 ( .A1(n8730), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8580) );
  OAI211_X1 U10125 ( .C1(n9178), .C2(n4480), .A(n8581), .B(n8580), .ZN(n8582)
         );
  INV_X1 U10126 ( .A(n8582), .ZN(n8583) );
  NAND2_X1 U10127 ( .A1(n9206), .A2(n8741), .ZN(n8677) );
  OAI21_X2 U10128 ( .B1(n8678), .B2(n8677), .A(n5096), .ZN(n8666) );
  NAND2_X1 U10129 ( .A1(n8586), .A2(n6262), .ZN(n8588) );
  NAND2_X1 U10130 ( .A1(n8622), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8587) );
  XNOR2_X1 U10131 ( .A(n9374), .B(n8599), .ZN(n8668) );
  NAND2_X1 U10132 ( .A1(n8589), .A2(n8671), .ZN(n8590) );
  AND2_X1 U10133 ( .A1(n8591), .A2(n8590), .ZN(n8670) );
  NAND2_X1 U10134 ( .A1(n8670), .A2(n8556), .ZN(n8596) );
  INV_X1 U10135 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U10136 ( .A1(n6174), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U10137 ( .A1(n8730), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8592) );
  OAI211_X1 U10138 ( .C1(n9162), .C2(n4480), .A(n8593), .B(n8592), .ZN(n8594)
         );
  INV_X1 U10139 ( .A(n8594), .ZN(n8595) );
  NAND2_X1 U10140 ( .A1(n9186), .A2(n8741), .ZN(n8667) );
  NAND2_X1 U10141 ( .A1(n9137), .A2(n8741), .ZN(n8597) );
  NOR2_X1 U10142 ( .A1(n8598), .A2(n8597), .ZN(n8611) );
  AOI21_X1 U10143 ( .B1(n8598), .B2(n8597), .A(n8611), .ZN(n8707) );
  XNOR2_X1 U10144 ( .A(n9363), .B(n8599), .ZN(n8606) );
  XNOR2_X1 U10145 ( .A(n8613), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U10146 ( .A1(n9132), .A2(n8556), .ZN(n8605) );
  INV_X1 U10147 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U10148 ( .A1(n6174), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10149 ( .A1(n8730), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8600) );
  OAI211_X1 U10150 ( .C1(n8602), .C2(n4480), .A(n8601), .B(n8600), .ZN(n8603)
         );
  INV_X1 U10151 ( .A(n8603), .ZN(n8604) );
  NOR2_X1 U10152 ( .A1(n9119), .A2(n8625), .ZN(n8607) );
  NAND2_X1 U10153 ( .A1(n8606), .A2(n8607), .ZN(n8633) );
  INV_X1 U10154 ( .A(n8606), .ZN(n8609) );
  INV_X1 U10155 ( .A(n8607), .ZN(n8608) );
  NAND2_X1 U10156 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  OAI22_X1 U10157 ( .A1(n8724), .A2(n8696), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8612), .ZN(n8620) );
  OAI21_X1 U10158 ( .B1(n8613), .B2(n8612), .A(n7769), .ZN(n8614) );
  INV_X1 U10159 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10160 ( .A1(n6174), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10161 ( .A1(n8730), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8615) );
  OAI211_X1 U10162 ( .C1(n8617), .C2(n4480), .A(n8616), .B(n8615), .ZN(n8618)
         );
  NOR2_X1 U10163 ( .A1(n9099), .A2(n8711), .ZN(n8619) );
  AOI211_X1 U10164 ( .C1(n8630), .C2(n9132), .A(n8620), .B(n8619), .ZN(n8621)
         );
  NAND2_X1 U10165 ( .A1(n10091), .A2(n6262), .ZN(n8624) );
  NAND2_X1 U10166 ( .A1(n8622), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8623) );
  OR2_X1 U10167 ( .A1(n9099), .A2(n8625), .ZN(n8627) );
  XNOR2_X1 U10168 ( .A(n8627), .B(n8626), .ZN(n8628) );
  XNOR2_X1 U10169 ( .A(n9358), .B(n8628), .ZN(n8629) );
  INV_X1 U10170 ( .A(n8629), .ZN(n8634) );
  NAND3_X1 U10171 ( .A1(n8634), .A2(n8705), .A3(n8633), .ZN(n8639) );
  NAND3_X1 U10172 ( .A1(n8640), .A2(n8705), .A3(n8629), .ZN(n8638) );
  NAND2_X1 U10173 ( .A1(n9149), .A2(n8714), .ZN(n8632) );
  AOI22_X1 U10174 ( .A1(n9113), .A2(n8630), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8631) );
  OAI211_X1 U10175 ( .C1(n9118), .C2(n8711), .A(n8632), .B(n8631), .ZN(n8636)
         );
  NOR3_X1 U10176 ( .A1(n8634), .A2(n8633), .A3(n4808), .ZN(n8635) );
  AOI211_X1 U10177 ( .C1(n9358), .C2(n8699), .A(n8636), .B(n8635), .ZN(n8637)
         );
  OAI211_X1 U10178 ( .C1(n8640), .C2(n8639), .A(n8638), .B(n8637), .ZN(
        P2_U3222) );
  NAND2_X1 U10179 ( .A1(n9082), .A2(n8700), .ZN(n8644) );
  OR2_X1 U10180 ( .A1(n8641), .A2(n4808), .ZN(n8643) );
  MUX2_X1 U10181 ( .A(n8644), .B(n8643), .S(n8642), .Z(n8649) );
  OAI22_X1 U10182 ( .A1(n9196), .A2(n8710), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8645), .ZN(n8647) );
  OAI22_X1 U10183 ( .A1(n8722), .A2(n8711), .B1(n9238), .B2(n8696), .ZN(n8646)
         );
  AOI211_X1 U10184 ( .C1(n9383), .C2(n8699), .A(n8647), .B(n8646), .ZN(n8648)
         );
  NAND2_X1 U10185 ( .A1(n8649), .A2(n8648), .ZN(P2_U3218) );
  INV_X1 U10186 ( .A(n8650), .ZN(n8651) );
  AOI21_X1 U10187 ( .B1(n8653), .B2(n8652), .A(n8651), .ZN(n8658) );
  INV_X1 U10188 ( .A(n8654), .ZN(n9255) );
  INV_X1 U10189 ( .A(n9237), .ZN(n9261) );
  INV_X1 U10190 ( .A(n9296), .ZN(n9260) );
  AOI22_X1 U10191 ( .A1(n8684), .A2(n9261), .B1(n8714), .B2(n9260), .ZN(n8655)
         );
  NAND2_X1 U10192 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9054) );
  OAI211_X1 U10193 ( .C1(n8710), .C2(n9255), .A(n8655), .B(n9054), .ZN(n8656)
         );
  AOI21_X1 U10194 ( .B1(n9407), .B2(n8699), .A(n8656), .ZN(n8657) );
  OAI21_X1 U10195 ( .B1(n8658), .B2(n4808), .A(n8657), .ZN(P2_U3221) );
  XNOR2_X1 U10196 ( .A(n8659), .B(n8660), .ZN(n8665) );
  OAI22_X1 U10197 ( .A1(n8710), .A2(n9229), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8661), .ZN(n8663) );
  OAI22_X1 U10198 ( .A1(n8696), .A2(n9237), .B1(n9238), .B2(n8711), .ZN(n8662)
         );
  AOI211_X1 U10199 ( .C1(n9394), .C2(n8699), .A(n8663), .B(n8662), .ZN(n8664)
         );
  OAI21_X1 U10200 ( .B1(n8665), .B2(n4808), .A(n8664), .ZN(P2_U3225) );
  XNOR2_X1 U10201 ( .A(n8668), .B(n8667), .ZN(n8669) );
  XNOR2_X1 U10202 ( .A(n8666), .B(n8669), .ZN(n8676) );
  OAI22_X1 U10203 ( .A1(n8724), .A2(n9311), .B1(n8722), .B2(n9309), .ZN(n9166)
         );
  INV_X1 U10204 ( .A(n8670), .ZN(n9163) );
  OAI22_X1 U10205 ( .A1(n9163), .A2(n8710), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8671), .ZN(n8673) );
  INV_X1 U10206 ( .A(n9374), .ZN(n9057) );
  NOR2_X1 U10207 ( .A1(n9057), .A2(n8717), .ZN(n8672) );
  AOI211_X1 U10208 ( .C1(n8674), .C2(n9166), .A(n8673), .B(n8672), .ZN(n8675)
         );
  OAI21_X1 U10209 ( .B1(n8676), .B2(n4808), .A(n8675), .ZN(P2_U3227) );
  INV_X1 U10210 ( .A(n9380), .ZN(n9177) );
  NAND2_X1 U10211 ( .A1(n8677), .A2(n8705), .ZN(n8680) );
  NAND2_X1 U10212 ( .A1(n9206), .A2(n8700), .ZN(n8679) );
  MUX2_X1 U10213 ( .A(n8680), .B(n8679), .S(n8678), .Z(n8686) );
  NOR2_X1 U10214 ( .A1(n9081), .A2(n8696), .ZN(n8683) );
  OAI22_X1 U10215 ( .A1(n9179), .A2(n8710), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8681), .ZN(n8682) );
  AOI211_X1 U10216 ( .C1(n9186), .C2(n8684), .A(n8683), .B(n8682), .ZN(n8685)
         );
  OAI211_X1 U10217 ( .C1(n9177), .C2(n8717), .A(n8686), .B(n8685), .ZN(
        P2_U3231) );
  XNOR2_X1 U10218 ( .A(n8688), .B(n8687), .ZN(n8693) );
  OAI22_X1 U10219 ( .A1(n8710), .A2(n9248), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8689), .ZN(n8691) );
  INV_X1 U10220 ( .A(n9242), .ZN(n9078) );
  OAI22_X1 U10221 ( .A1(n8696), .A2(n9076), .B1(n9078), .B2(n8711), .ZN(n8690)
         );
  AOI211_X1 U10222 ( .C1(n9400), .C2(n8699), .A(n8691), .B(n8690), .ZN(n8692)
         );
  OAI21_X1 U10223 ( .B1(n8693), .B2(n4808), .A(n8692), .ZN(P2_U3235) );
  INV_X1 U10224 ( .A(n9214), .ZN(n8695) );
  OAI22_X1 U10225 ( .A1(n8710), .A2(n8695), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8694), .ZN(n8698) );
  OAI22_X1 U10226 ( .A1(n9081), .A2(n8711), .B1(n9078), .B2(n8696), .ZN(n8697)
         );
  AOI211_X1 U10227 ( .C1(n9388), .C2(n8699), .A(n8698), .B(n8697), .ZN(n8703)
         );
  NAND3_X1 U10228 ( .A1(n8701), .A2(n8700), .A3(n9207), .ZN(n8702) );
  OAI211_X1 U10229 ( .C1(n8704), .C2(n4808), .A(n8703), .B(n8702), .ZN(
        P2_U3237) );
  INV_X1 U10230 ( .A(n9369), .ZN(n9155) );
  OAI211_X1 U10231 ( .C1(n8708), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8716)
         );
  OAI22_X1 U10232 ( .A1(n9153), .A2(n8710), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8709), .ZN(n8713) );
  NOR2_X1 U10233 ( .A1(n9119), .A2(n8711), .ZN(n8712) );
  AOI211_X1 U10234 ( .C1(n8714), .C2(n9186), .A(n8713), .B(n8712), .ZN(n8715)
         );
  OAI211_X1 U10235 ( .C1(n9155), .C2(n8717), .A(n8716), .B(n8715), .ZN(
        P2_U3242) );
  NAND2_X1 U10236 ( .A1(n9429), .A2(n9310), .ZN(n8833) );
  NAND2_X1 U10237 ( .A1(n8834), .A2(n8833), .ZN(n9340) );
  INV_X1 U10238 ( .A(n9340), .ZN(n8831) );
  INV_X1 U10239 ( .A(n8834), .ZN(n8719) );
  OR2_X1 U10240 ( .A1(n9324), .A2(n9295), .ZN(n8838) );
  NAND2_X1 U10241 ( .A1(n9324), .A2(n9295), .ZN(n8837) );
  NAND2_X1 U10242 ( .A1(n8838), .A2(n8837), .ZN(n9304) );
  INV_X1 U10243 ( .A(n9304), .ZN(n9308) );
  NAND2_X1 U10244 ( .A1(n9307), .A2(n9308), .ZN(n9306) );
  NAND2_X1 U10245 ( .A1(n9420), .A2(n9312), .ZN(n8752) );
  INV_X1 U10246 ( .A(n9285), .ZN(n9291) );
  NAND2_X1 U10247 ( .A1(n9413), .A2(n9296), .ZN(n8843) );
  INV_X1 U10248 ( .A(n8849), .ZN(n8720) );
  OR2_X1 U10249 ( .A1(n9407), .A2(n9076), .ZN(n8848) );
  NAND2_X1 U10250 ( .A1(n9407), .A2(n9076), .ZN(n8851) );
  NAND2_X1 U10251 ( .A1(n9400), .A2(n9237), .ZN(n8855) );
  INV_X1 U10252 ( .A(n9244), .ZN(n8915) );
  OR2_X1 U10253 ( .A1(n9394), .A2(n9078), .ZN(n8859) );
  NAND2_X1 U10254 ( .A1(n9394), .A2(n9078), .ZN(n8856) );
  NAND2_X1 U10255 ( .A1(n8859), .A2(n8856), .ZN(n9234) );
  INV_X1 U10256 ( .A(n8856), .ZN(n8721) );
  OR2_X1 U10257 ( .A1(n9388), .A2(n9238), .ZN(n8860) );
  NAND2_X1 U10258 ( .A1(n9388), .A2(n9238), .ZN(n8863) );
  OR2_X1 U10259 ( .A1(n9383), .A2(n9081), .ZN(n8865) );
  NAND2_X1 U10260 ( .A1(n9383), .A2(n9081), .ZN(n9185) );
  NAND2_X1 U10261 ( .A1(n8865), .A2(n9185), .ZN(n9201) );
  INV_X1 U10262 ( .A(n8860), .ZN(n9202) );
  NOR2_X1 U10263 ( .A1(n9201), .A2(n9202), .ZN(n8867) );
  NAND2_X1 U10264 ( .A1(n9200), .A2(n8867), .ZN(n9204) );
  NAND2_X1 U10265 ( .A1(n9380), .A2(n8722), .ZN(n8871) );
  NAND3_X1 U10266 ( .A1(n9204), .A2(n9184), .A3(n9185), .ZN(n9183) );
  NAND2_X1 U10267 ( .A1(n9374), .A2(n8723), .ZN(n8747) );
  INV_X1 U10268 ( .A(n9164), .ZN(n8918) );
  OR2_X1 U10269 ( .A1(n9363), .A2(n9119), .ZN(n8877) );
  NAND2_X1 U10270 ( .A1(n9358), .A2(n9099), .ZN(n8880) );
  NAND2_X1 U10271 ( .A1(n9092), .A2(n8880), .ZN(n9116) );
  INV_X1 U10272 ( .A(n9116), .ZN(n8725) );
  NAND2_X1 U10273 ( .A1(n9464), .A2(n6262), .ZN(n8727) );
  NAND2_X1 U10274 ( .A1(n4485), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U10275 ( .A1(n9354), .A2(n9118), .ZN(n8887) );
  NAND2_X1 U10276 ( .A1(n8884), .A2(n8887), .ZN(n9089) );
  INV_X1 U10277 ( .A(n9089), .ZN(n9091) );
  NAND2_X1 U10278 ( .A1(n9460), .A2(n6262), .ZN(n8729) );
  NAND2_X1 U10279 ( .A1(n8622), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8728) );
  INV_X1 U10280 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U10281 ( .A1(n8730), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U10282 ( .A1(n6174), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8731) );
  OAI211_X1 U10283 ( .C1(n4480), .C2(n8733), .A(n8732), .B(n8731), .ZN(n9095)
         );
  INV_X1 U10284 ( .A(n9095), .ZN(n8736) );
  NAND2_X1 U10285 ( .A1(n9457), .A2(n6262), .ZN(n8735) );
  NAND2_X1 U10286 ( .A1(n4485), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8734) );
  OR2_X1 U10287 ( .A1(n9350), .A2(n8737), .ZN(n8891) );
  NAND2_X1 U10288 ( .A1(n9063), .A2(n8736), .ZN(n8888) );
  NAND2_X1 U10289 ( .A1(n8891), .A2(n8888), .ZN(n8889) );
  NAND2_X1 U10290 ( .A1(n9350), .A2(n8737), .ZN(n8890) );
  OAI21_X1 U10291 ( .B1(n8738), .B2(n8889), .A(n8890), .ZN(n8739) );
  NAND2_X1 U10292 ( .A1(n8763), .A2(n10369), .ZN(n8742) );
  INV_X1 U10293 ( .A(n8748), .ZN(n8743) );
  AOI21_X1 U10294 ( .B1(n8745), .B2(n8744), .A(n8743), .ZN(n8750) );
  INV_X1 U10295 ( .A(n8745), .ZN(n8746) );
  AOI21_X1 U10296 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8749) );
  MUX2_X1 U10297 ( .A(n8750), .B(n8749), .S(n8892), .Z(n8874) );
  OAI211_X1 U10298 ( .C1(n8886), .C2(n8751), .A(n9148), .B(n8918), .ZN(n8873)
         );
  INV_X1 U10299 ( .A(n9201), .ZN(n8917) );
  AND2_X1 U10300 ( .A1(n8843), .A2(n8752), .ZN(n8753) );
  MUX2_X1 U10301 ( .A(n8754), .B(n8753), .S(n8886), .Z(n8842) );
  NAND2_X1 U10302 ( .A1(n8781), .A2(n8783), .ZN(n8756) );
  NAND2_X1 U10303 ( .A1(n8759), .A2(n8758), .ZN(n8755) );
  AND2_X1 U10304 ( .A1(n8758), .A2(n8757), .ZN(n8760) );
  OAI211_X1 U10305 ( .C1(n8785), .C2(n8760), .A(n8759), .B(n8790), .ZN(n8761)
         );
  NAND2_X1 U10306 ( .A1(n8761), .A2(n8892), .ZN(n8771) );
  INV_X1 U10307 ( .A(n8785), .ZN(n8769) );
  NAND2_X1 U10308 ( .A1(n8945), .A2(n8762), .ZN(n8772) );
  AND2_X1 U10309 ( .A1(n8772), .A2(n8763), .ZN(n8764) );
  OAI211_X1 U10310 ( .C1(n8765), .C2(n8764), .A(n8776), .B(n6688), .ZN(n8766)
         );
  NAND3_X1 U10311 ( .A1(n8766), .A2(n8775), .A3(n8892), .ZN(n8767) );
  NAND3_X1 U10312 ( .A1(n8769), .A2(n8768), .A3(n8767), .ZN(n8770) );
  NAND2_X1 U10313 ( .A1(n8771), .A2(n8770), .ZN(n8779) );
  NAND2_X1 U10314 ( .A1(n6688), .A2(n8772), .ZN(n8773) );
  NAND3_X1 U10315 ( .A1(n8775), .A2(n8774), .A3(n8773), .ZN(n8777) );
  NAND3_X1 U10316 ( .A1(n8777), .A2(n8886), .A3(n8776), .ZN(n8778) );
  NAND3_X1 U10317 ( .A1(n8779), .A2(n8782), .A3(n8778), .ZN(n8788) );
  AND2_X1 U10318 ( .A1(n8781), .A2(n8780), .ZN(n8784) );
  OAI211_X1 U10319 ( .C1(n8785), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8786)
         );
  NAND2_X1 U10320 ( .A1(n8786), .A2(n8886), .ZN(n8787) );
  NAND2_X1 U10321 ( .A1(n8788), .A2(n8787), .ZN(n8789) );
  OAI211_X1 U10322 ( .C1(n8790), .C2(n8892), .A(n8789), .B(n8904), .ZN(n8807)
         );
  NAND3_X1 U10323 ( .A1(n8807), .A2(n8806), .A3(n8791), .ZN(n8793) );
  NAND2_X1 U10324 ( .A1(n8793), .A2(n8792), .ZN(n8796) );
  NAND2_X1 U10325 ( .A1(n8797), .A2(n8794), .ZN(n8795) );
  MUX2_X1 U10326 ( .A(n8796), .B(n8795), .S(n8892), .Z(n8802) );
  OAI21_X1 U10327 ( .B1(n8802), .B2(n8801), .A(n8808), .ZN(n8816) );
  NAND2_X1 U10328 ( .A1(n8804), .A2(n8803), .ZN(n8813) );
  NAND3_X1 U10329 ( .A1(n8807), .A2(n8806), .A3(n8805), .ZN(n8811) );
  INV_X1 U10330 ( .A(n8808), .ZN(n8810) );
  OAI211_X1 U10331 ( .C1(n8811), .C2(n8810), .A(n8817), .B(n8809), .ZN(n8812)
         );
  MUX2_X1 U10332 ( .A(n8813), .B(n8812), .S(n8892), .Z(n8814) );
  INV_X1 U10333 ( .A(n8814), .ZN(n8815) );
  AND2_X1 U10334 ( .A1(n8818), .A2(n8817), .ZN(n8821) );
  INV_X1 U10335 ( .A(n8819), .ZN(n8820) );
  MUX2_X1 U10336 ( .A(n8825), .B(n8824), .S(n8886), .Z(n8826) );
  MUX2_X1 U10337 ( .A(n8829), .B(n8828), .S(n8892), .Z(n8830) );
  NAND3_X1 U10338 ( .A1(n8832), .A2(n8831), .A3(n8830), .ZN(n8836) );
  MUX2_X1 U10339 ( .A(n8834), .B(n8833), .S(n8886), .Z(n8835) );
  NAND3_X1 U10340 ( .A1(n8836), .A2(n9308), .A3(n8835), .ZN(n8840) );
  MUX2_X1 U10341 ( .A(n8838), .B(n8837), .S(n8892), .Z(n8839) );
  NAND3_X1 U10342 ( .A1(n8840), .A2(n9285), .A3(n8839), .ZN(n8841) );
  NAND3_X1 U10343 ( .A1(n8842), .A2(n8849), .A3(n8841), .ZN(n8850) );
  NAND2_X1 U10344 ( .A1(n8850), .A2(n8843), .ZN(n8844) );
  NAND2_X1 U10345 ( .A1(n8844), .A2(n8848), .ZN(n8845) );
  NAND3_X1 U10346 ( .A1(n8845), .A2(n8855), .A3(n8851), .ZN(n8846) );
  NAND3_X1 U10347 ( .A1(n8846), .A2(n8853), .A3(n8859), .ZN(n8847) );
  NAND3_X1 U10348 ( .A1(n8863), .A2(n8847), .A3(n8856), .ZN(n8862) );
  NAND3_X1 U10349 ( .A1(n8850), .A2(n8849), .A3(n8848), .ZN(n8852) );
  NAND2_X1 U10350 ( .A1(n8852), .A2(n8851), .ZN(n8854) );
  NAND2_X1 U10351 ( .A1(n8854), .A2(n8853), .ZN(n8857) );
  NAND3_X1 U10352 ( .A1(n8857), .A2(n8856), .A3(n8855), .ZN(n8858) );
  NAND3_X1 U10353 ( .A1(n8860), .A2(n8859), .A3(n8858), .ZN(n8861) );
  NAND3_X1 U10354 ( .A1(n8917), .A2(n8863), .A3(n8866), .ZN(n8864) );
  NAND3_X1 U10355 ( .A1(n9184), .A2(n8865), .A3(n8864), .ZN(n8869) );
  AND2_X1 U10356 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  AOI21_X1 U10357 ( .B1(n8871), .B2(n9185), .A(n8886), .ZN(n8870) );
  INV_X1 U10358 ( .A(n8880), .ZN(n8875) );
  AOI21_X1 U10359 ( .B1(n9119), .B2(n9363), .A(n8875), .ZN(n8876) );
  MUX2_X1 U10360 ( .A(n8877), .B(n8876), .S(n8892), .Z(n8878) );
  INV_X1 U10361 ( .A(n8887), .ZN(n8879) );
  AOI21_X1 U10362 ( .B1(n8881), .B2(n9099), .A(n8879), .ZN(n8883) );
  OAI211_X1 U10363 ( .C1(n8886), .C2(n9358), .A(n8881), .B(n8880), .ZN(n8882)
         );
  OAI21_X1 U10364 ( .B1(n8883), .B2(n8886), .A(n8882), .ZN(n8885) );
  INV_X1 U10365 ( .A(n8889), .ZN(n8922) );
  AND2_X1 U10366 ( .A1(n8890), .A2(n4507), .ZN(n8921) );
  MUX2_X1 U10367 ( .A(n8922), .B(n8921), .S(n8892), .Z(n8896) );
  INV_X1 U10368 ( .A(n8890), .ZN(n8894) );
  INV_X1 U10369 ( .A(n8891), .ZN(n8893) );
  MUX2_X1 U10370 ( .A(n8894), .B(n8893), .S(n8892), .Z(n8895) );
  INV_X1 U10371 ( .A(n8924), .ZN(n8929) );
  OAI21_X1 U10372 ( .B1(n4837), .B2(n6689), .A(n10436), .ZN(n8928) );
  NAND4_X1 U10373 ( .A1(n8900), .A2(n8899), .A3(n4837), .A4(n8898), .ZN(n8903)
         );
  NOR3_X1 U10374 ( .A1(n8903), .A2(n8902), .A3(n8901), .ZN(n8906) );
  NAND4_X1 U10375 ( .A1(n8906), .A2(n10359), .A3(n8905), .A4(n8904), .ZN(n8908) );
  NOR4_X1 U10376 ( .A1(n8909), .A2(n8908), .A3(n8907), .A4(n7233), .ZN(n8910)
         );
  NAND4_X1 U10377 ( .A1(n9070), .A2(n8911), .A3(n5041), .A4(n8910), .ZN(n8912)
         );
  NOR4_X1 U10378 ( .A1(n9304), .A2(n9340), .A3(n9068), .A4(n8912), .ZN(n8913)
         );
  NAND4_X1 U10379 ( .A1(n9258), .A2(n9277), .A3(n9285), .A4(n8913), .ZN(n8914)
         );
  NOR4_X1 U10380 ( .A1(n4966), .A2(n8915), .A3(n9234), .A4(n8914), .ZN(n8916)
         );
  NAND4_X1 U10381 ( .A1(n8918), .A2(n8917), .A3(n9184), .A4(n8916), .ZN(n8919)
         );
  NOR4_X1 U10382 ( .A1(n9116), .A2(n9135), .A3(n9143), .A4(n8919), .ZN(n8920)
         );
  NAND4_X1 U10383 ( .A1(n8922), .A2(n8921), .A3(n9091), .A4(n8920), .ZN(n8923)
         );
  XNOR2_X1 U10384 ( .A(n8923), .B(n10369), .ZN(n8927) );
  AOI21_X1 U10385 ( .B1(n8924), .B2(n6689), .A(n4837), .ZN(n8925) );
  INV_X1 U10386 ( .A(n8931), .ZN(n10378) );
  NAND4_X1 U10387 ( .A1(n10378), .A2(n9472), .A3(n8932), .A4(n10360), .ZN(
        n8933) );
  OAI211_X1 U10388 ( .C1(n6141), .C2(n8934), .A(n8933), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8935) );
  MUX2_X1 U10389 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9095), .S(P2_U3966), .Z(
        P2_U3582) );
  INV_X1 U10390 ( .A(n9099), .ZN(n9136) );
  MUX2_X1 U10391 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9136), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10392 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9149), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10393 ( .A(n9137), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8936), .Z(
        P2_U3578) );
  MUX2_X1 U10394 ( .A(n9186), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8936), .Z(
        P2_U3577) );
  MUX2_X1 U10395 ( .A(n9206), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8936), .Z(
        P2_U3576) );
  MUX2_X1 U10396 ( .A(n9082), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8936), .Z(
        P2_U3575) );
  MUX2_X1 U10397 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9207), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10398 ( .A(n9242), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8936), .Z(
        P2_U3573) );
  MUX2_X1 U10399 ( .A(n9261), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8936), .Z(
        P2_U3572) );
  INV_X1 U10400 ( .A(n9076), .ZN(n9279) );
  MUX2_X1 U10401 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9279), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10402 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9260), .S(P2_U3966), .Z(
        P2_U3570) );
  INV_X1 U10403 ( .A(n9312), .ZN(n9278) );
  MUX2_X1 U10404 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9278), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U10405 ( .A(n9295), .ZN(n9343) );
  MUX2_X1 U10406 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9343), .S(P2_U3966), .Z(
        P2_U3568) );
  INV_X1 U10407 ( .A(n8937), .ZN(n9342) );
  MUX2_X1 U10408 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9342), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10409 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8938), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10410 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8939), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10411 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8940), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10412 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n4771), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10413 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n4769), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10414 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8941), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10415 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8942), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10416 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n10363), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10417 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8943), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10418 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n10361), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10419 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8944), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10420 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6181), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10421 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6790), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10422 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8945), .S(P2_U3966), .Z(
        P2_U3552) );
  NOR2_X1 U10423 ( .A1(n5034), .A2(n6158), .ZN(n8948) );
  OAI211_X1 U10424 ( .C1(n8948), .C2(n8947), .A(n10350), .B(n8946), .ZN(n8956)
         );
  AOI22_X1 U10425 ( .A1(n10351), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8955) );
  NAND2_X1 U10426 ( .A1(n10347), .A2(n8949), .ZN(n8954) );
  OAI211_X1 U10427 ( .C1(n8952), .C2(n8951), .A(n10349), .B(n8950), .ZN(n8953)
         );
  NAND4_X1 U10428 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(
        P2_U3246) );
  OAI211_X1 U10429 ( .C1(n8959), .C2(n8958), .A(n10350), .B(n8957), .ZN(n8967)
         );
  AOI22_X1 U10430 ( .A1(n10351), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8966) );
  NAND2_X1 U10431 ( .A1(n10347), .A2(n8960), .ZN(n8965) );
  OAI211_X1 U10432 ( .C1(n8963), .C2(n8962), .A(n10349), .B(n8961), .ZN(n8964)
         );
  NAND4_X1 U10433 ( .A1(n8967), .A2(n8966), .A3(n8965), .A4(n8964), .ZN(
        P2_U3247) );
  AOI21_X1 U10434 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8971) );
  OR2_X1 U10435 ( .A1(n8971), .A2(n9048), .ZN(n8981) );
  NOR2_X1 U10436 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6337), .ZN(n8972) );
  AOI21_X1 U10437 ( .B1(n10351), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8972), .ZN(
        n8980) );
  NAND2_X1 U10438 ( .A1(n10347), .A2(n8973), .ZN(n8979) );
  AOI21_X1 U10439 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8977) );
  NAND2_X1 U10440 ( .A1(n10349), .A2(n8977), .ZN(n8978) );
  NAND4_X1 U10441 ( .A1(n8981), .A2(n8980), .A3(n8979), .A4(n8978), .ZN(
        P2_U3256) );
  NOR2_X1 U10442 ( .A1(n8983), .A2(n8982), .ZN(n8985) );
  NOR2_X1 U10443 ( .A1(n8985), .A2(n8984), .ZN(n8988) );
  XNOR2_X1 U10444 ( .A(n9011), .B(n8986), .ZN(n8987) );
  NAND2_X1 U10445 ( .A1(n8987), .A2(n8988), .ZN(n9012) );
  OAI21_X1 U10446 ( .B1(n8988), .B2(n8987), .A(n9012), .ZN(n8989) );
  NAND2_X1 U10447 ( .A1(n8989), .A2(n10349), .ZN(n9002) );
  INV_X1 U10448 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8991) );
  OAI21_X1 U10449 ( .B1(n9056), .B2(n8991), .A(n8990), .ZN(n8992) );
  AOI21_X1 U10450 ( .B1(n10347), .B2(n9011), .A(n8992), .ZN(n9001) );
  NOR2_X1 U10451 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  NOR2_X1 U10452 ( .A1(n8996), .A2(n8995), .ZN(n8999) );
  MUX2_X1 U10453 ( .A(n9318), .B(P2_REG2_REG_16__SCAN_IN), .S(n9011), .Z(n8997) );
  INV_X1 U10454 ( .A(n8997), .ZN(n8998) );
  NAND2_X1 U10455 ( .A1(n8998), .A2(n8999), .ZN(n9003) );
  OAI211_X1 U10456 ( .C1(n8999), .C2(n8998), .A(n10350), .B(n9003), .ZN(n9000)
         );
  NAND3_X1 U10457 ( .A1(n9002), .A2(n9001), .A3(n9000), .ZN(P2_U3261) );
  NAND2_X1 U10458 ( .A1(n9011), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U10459 ( .A1(n9004), .A2(n9003), .ZN(n9008) );
  NAND2_X1 U10460 ( .A1(n9027), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9022) );
  INV_X1 U10461 ( .A(n9022), .ZN(n9005) );
  AOI21_X1 U10462 ( .B1(n9287), .B2(n9006), .A(n9005), .ZN(n9007) );
  NAND2_X1 U10463 ( .A1(n9007), .A2(n9008), .ZN(n9021) );
  OAI211_X1 U10464 ( .C1(n9008), .C2(n9007), .A(n10350), .B(n9021), .ZN(n9020)
         );
  NOR2_X1 U10465 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9009), .ZN(n9010) );
  AOI21_X1 U10466 ( .B1(n10351), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9010), .ZN(
        n9019) );
  NAND2_X1 U10467 ( .A1(n10347), .A2(n9027), .ZN(n9018) );
  OR2_X1 U10468 ( .A1(n9011), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9013) );
  XNOR2_X1 U10469 ( .A(n9027), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9014) );
  AOI21_X1 U10470 ( .B1(n9015), .B2(n9014), .A(n9026), .ZN(n9016) );
  NAND2_X1 U10471 ( .A1(n10349), .A2(n9016), .ZN(n9017) );
  NAND4_X1 U10472 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(
        P2_U3262) );
  NAND2_X1 U10473 ( .A1(n9022), .A2(n9021), .ZN(n9037) );
  XNOR2_X1 U10474 ( .A(n9037), .B(n9042), .ZN(n9035) );
  XOR2_X1 U10475 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n9035), .Z(n9023) );
  NAND2_X1 U10476 ( .A1(n9023), .A2(n10350), .ZN(n9034) );
  NOR2_X1 U10477 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9024), .ZN(n9025) );
  AOI21_X1 U10478 ( .B1(n10351), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9025), .ZN(
        n9033) );
  INV_X1 U10479 ( .A(n9042), .ZN(n9036) );
  NAND2_X1 U10480 ( .A1(n10347), .A2(n9036), .ZN(n9032) );
  XNOR2_X1 U10481 ( .A(n9042), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9029) );
  OAI21_X1 U10482 ( .B1(n9029), .B2(n9028), .A(n9044), .ZN(n9030) );
  NAND2_X1 U10483 ( .A1(n10349), .A2(n9030), .ZN(n9031) );
  NAND4_X1 U10484 ( .A1(n9034), .A2(n9033), .A3(n9032), .A4(n9031), .ZN(
        P2_U3263) );
  NAND2_X1 U10485 ( .A1(n9035), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U10486 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NAND2_X1 U10487 ( .A1(n9039), .A2(n9038), .ZN(n9040) );
  XOR2_X1 U10488 ( .A(n9040), .B(P2_REG2_REG_19__SCAN_IN), .Z(n9049) );
  INV_X1 U10489 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U10490 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  NAND2_X1 U10491 ( .A1(n9044), .A2(n9043), .ZN(n9046) );
  INV_X1 U10492 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9045) );
  XNOR2_X1 U10493 ( .A(n9046), .B(n9045), .ZN(n9051) );
  INV_X1 U10494 ( .A(n9051), .ZN(n9047) );
  AOI22_X1 U10495 ( .A1(n9049), .A2(n10350), .B1(n9047), .B2(n10349), .ZN(
        n9053) );
  NOR2_X1 U10496 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  AOI211_X1 U10497 ( .C1(n10349), .C2(n9051), .A(n10347), .B(n9050), .ZN(n9052) );
  MUX2_X1 U10498 ( .A(n9053), .B(n9052), .S(n10369), .Z(n9055) );
  OAI211_X1 U10499 ( .C1(n5106), .C2(n9056), .A(n9055), .B(n9054), .ZN(
        P2_U3264) );
  INV_X1 U10500 ( .A(n9354), .ZN(n9101) );
  INV_X1 U10501 ( .A(n9394), .ZN(n9228) );
  NOR2_X1 U10502 ( .A1(n9333), .A2(n9429), .ZN(n9332) );
  INV_X1 U10503 ( .A(n9420), .ZN(n9075) );
  NAND2_X1 U10504 ( .A1(n9320), .A2(n9075), .ZN(n9288) );
  NOR2_X1 U10505 ( .A1(n9225), .A2(n9388), .ZN(n9213) );
  NAND2_X1 U10506 ( .A1(n9199), .A2(n9213), .ZN(n9193) );
  NAND2_X1 U10507 ( .A1(n9057), .A2(n9176), .ZN(n9168) );
  NOR2_X2 U10508 ( .A1(n9168), .A2(n9369), .ZN(n9151) );
  XOR2_X1 U10509 ( .A(n9350), .B(n9062), .Z(n9352) );
  NOR2_X1 U10510 ( .A1(n10370), .A2(n9058), .ZN(n9060) );
  AOI21_X1 U10511 ( .B1(n9472), .B2(P2_B_REG_SCAN_IN), .A(n9311), .ZN(n9096)
         );
  NAND2_X1 U10512 ( .A1(n9059), .A2(n9096), .ZN(n10113) );
  NOR2_X1 U10513 ( .A1(n10357), .A2(n10113), .ZN(n9064) );
  AOI211_X1 U10514 ( .C1(n9350), .C2(n9325), .A(n9060), .B(n9064), .ZN(n9061)
         );
  OAI21_X1 U10515 ( .B1(n9352), .B2(n9321), .A(n9061), .ZN(P2_U3265) );
  AOI21_X1 U10516 ( .B1(n9063), .B2(n9100), .A(n9062), .ZN(n10115) );
  NAND2_X1 U10517 ( .A1(n10115), .A2(n9347), .ZN(n9066) );
  AOI21_X1 U10518 ( .B1(n10357), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9064), .ZN(
        n9065) );
  OAI211_X1 U10519 ( .C1(n4979), .C2(n9338), .A(n9066), .B(n9065), .ZN(
        P2_U3266) );
  INV_X1 U10520 ( .A(n9413), .ZN(n9275) );
  AND2_X1 U10521 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  OR2_X1 U10522 ( .A1(n9436), .A2(n9342), .ZN(n9072) );
  NAND2_X1 U10523 ( .A1(n9073), .A2(n9072), .ZN(n9330) );
  NAND2_X1 U10524 ( .A1(n9330), .A2(n9340), .ZN(n9329) );
  NAND2_X1 U10525 ( .A1(n9339), .A2(n9310), .ZN(n9302) );
  AND2_X1 U10526 ( .A1(n9302), .A2(n9304), .ZN(n9074) );
  NOR2_X1 U10527 ( .A1(n9263), .A2(n9076), .ZN(n9077) );
  NOR2_X1 U10528 ( .A1(n9394), .A2(n9242), .ZN(n9079) );
  NAND2_X1 U10529 ( .A1(n5054), .A2(n9201), .ZN(n9192) );
  NAND2_X1 U10530 ( .A1(n9160), .A2(n9164), .ZN(n9159) );
  NAND2_X1 U10531 ( .A1(n9159), .A2(n9084), .ZN(n9144) );
  NAND2_X1 U10532 ( .A1(n9144), .A2(n9143), .ZN(n9142) );
  XNOR2_X1 U10533 ( .A(n9090), .B(n9089), .ZN(n9353) );
  INV_X1 U10534 ( .A(n9353), .ZN(n9108) );
  AOI21_X1 U10535 ( .B1(n9121), .B2(n9092), .A(n9091), .ZN(n9093) );
  NAND2_X1 U10536 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  OAI211_X1 U10537 ( .C1(n9099), .C2(n9309), .A(n9098), .B(n9097), .ZN(n9356)
         );
  OAI21_X1 U10538 ( .B1(n9112), .B2(n9101), .A(n9100), .ZN(n9355) );
  OAI22_X1 U10539 ( .A1(n9103), .A2(n10375), .B1(n9102), .B2(n10370), .ZN(
        n9104) );
  AOI21_X1 U10540 ( .B1(n9354), .B2(n9325), .A(n9104), .ZN(n9105) );
  OAI21_X1 U10541 ( .B1(n9355), .B2(n9321), .A(n9105), .ZN(n9106) );
  AOI21_X1 U10542 ( .B1(n9356), .B2(n10370), .A(n9106), .ZN(n9107) );
  OAI21_X1 U10543 ( .B1(n9108), .B2(n9349), .A(n9107), .ZN(P2_U3267) );
  OAI21_X1 U10544 ( .B1(n9110), .B2(n9116), .A(n9109), .ZN(n9111) );
  AOI21_X1 U10545 ( .B1(n9358), .B2(n9129), .A(n9112), .ZN(n9359) );
  AOI22_X1 U10546 ( .A1(n9113), .A2(n9335), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10357), .ZN(n9114) );
  OAI21_X1 U10547 ( .B1(n9088), .B2(n9338), .A(n9114), .ZN(n9124) );
  INV_X1 U10548 ( .A(n9115), .ZN(n9117) );
  AOI21_X1 U10549 ( .B1(n9117), .B2(n9116), .A(n9293), .ZN(n9122) );
  OAI22_X1 U10550 ( .A1(n9119), .A2(n9309), .B1(n9118), .B2(n9311), .ZN(n9120)
         );
  AOI21_X1 U10551 ( .B1(n9122), .B2(n9121), .A(n9120), .ZN(n9361) );
  NOR2_X1 U10552 ( .A1(n9361), .A2(n10357), .ZN(n9123) );
  AOI211_X1 U10553 ( .C1(n9359), .C2(n9347), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI21_X1 U10554 ( .B1(n9362), .B2(n9349), .A(n9125), .ZN(P2_U3268) );
  OAI21_X1 U10555 ( .B1(n9127), .B2(n9135), .A(n9126), .ZN(n9128) );
  INV_X1 U10556 ( .A(n9128), .ZN(n9367) );
  INV_X1 U10557 ( .A(n9151), .ZN(n9131) );
  INV_X1 U10558 ( .A(n9129), .ZN(n9130) );
  AOI21_X1 U10559 ( .B1(n9363), .B2(n9131), .A(n9130), .ZN(n9364) );
  AOI22_X1 U10560 ( .A1(n9132), .A2(n9335), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10357), .ZN(n9133) );
  OAI21_X1 U10561 ( .B1(n9086), .B2(n9338), .A(n9133), .ZN(n9140) );
  XOR2_X1 U10562 ( .A(n9135), .B(n9134), .Z(n9138) );
  AOI222_X1 U10563 ( .A1(n10365), .A2(n9138), .B1(n9137), .B2(n10360), .C1(
        n9136), .C2(n10362), .ZN(n9366) );
  NOR2_X1 U10564 ( .A1(n9366), .A2(n10357), .ZN(n9139) );
  AOI211_X1 U10565 ( .C1(n9364), .C2(n9347), .A(n9140), .B(n9139), .ZN(n9141)
         );
  OAI21_X1 U10566 ( .B1(n9367), .B2(n9349), .A(n9141), .ZN(P2_U3269) );
  OAI21_X1 U10567 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(n9145) );
  INV_X1 U10568 ( .A(n9145), .ZN(n9372) );
  OAI21_X1 U10569 ( .B1(n9148), .B2(n9147), .A(n9146), .ZN(n9150) );
  AOI222_X1 U10570 ( .A1(n10365), .A2(n9150), .B1(n9186), .B2(n10360), .C1(
        n9149), .C2(n10362), .ZN(n9371) );
  AOI211_X1 U10571 ( .C1(n9369), .C2(n9168), .A(n10436), .B(n9151), .ZN(n9368)
         );
  NAND2_X1 U10572 ( .A1(n9368), .A2(n9297), .ZN(n9152) );
  OAI211_X1 U10573 ( .C1(n10375), .C2(n9153), .A(n9371), .B(n9152), .ZN(n9157)
         );
  OAI22_X1 U10574 ( .A1(n9155), .A2(n9338), .B1(n10370), .B2(n9154), .ZN(n9156) );
  AOI21_X1 U10575 ( .B1(n9157), .B2(n10370), .A(n9156), .ZN(n9158) );
  OAI21_X1 U10576 ( .B1(n9372), .B2(n9349), .A(n9158), .ZN(P2_U3270) );
  OAI21_X1 U10577 ( .B1(n9160), .B2(n9164), .A(n9159), .ZN(n9161) );
  INV_X1 U10578 ( .A(n9161), .ZN(n9377) );
  OAI22_X1 U10579 ( .A1(n9163), .A2(n10375), .B1(n9162), .B2(n10370), .ZN(
        n9173) );
  XNOR2_X1 U10580 ( .A(n9165), .B(n9164), .ZN(n9167) );
  AOI21_X1 U10581 ( .B1(n9167), .B2(n10365), .A(n9166), .ZN(n9376) );
  INV_X1 U10582 ( .A(n9176), .ZN(n9170) );
  INV_X1 U10583 ( .A(n9168), .ZN(n9169) );
  AOI211_X1 U10584 ( .C1(n9374), .C2(n9170), .A(n10436), .B(n9169), .ZN(n9373)
         );
  NAND2_X1 U10585 ( .A1(n9373), .A2(n9297), .ZN(n9171) );
  AOI21_X1 U10586 ( .B1(n9376), .B2(n9171), .A(n10357), .ZN(n9172) );
  AOI211_X1 U10587 ( .C1(n9325), .C2(n9374), .A(n9173), .B(n9172), .ZN(n9174)
         );
  OAI21_X1 U10588 ( .B1(n9377), .B2(n9349), .A(n9174), .ZN(P2_U3271) );
  XOR2_X1 U10589 ( .A(n9184), .B(n9175), .Z(n9382) );
  AOI211_X1 U10590 ( .C1(n9380), .C2(n9193), .A(n10436), .B(n9176), .ZN(n9379)
         );
  NOR2_X1 U10591 ( .A1(n9177), .A2(n9338), .ZN(n9181) );
  OAI22_X1 U10592 ( .A1(n9179), .A2(n10375), .B1(n9178), .B2(n10370), .ZN(
        n9180) );
  AOI211_X1 U10593 ( .C1(n9379), .C2(n9182), .A(n9181), .B(n9180), .ZN(n9191)
         );
  NAND2_X1 U10594 ( .A1(n9183), .A2(n10365), .ZN(n9189) );
  AOI21_X1 U10595 ( .B1(n9204), .B2(n9185), .A(n9184), .ZN(n9188) );
  AOI22_X1 U10596 ( .A1(n9186), .A2(n10362), .B1(n10360), .B2(n9082), .ZN(
        n9187) );
  OAI21_X1 U10597 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(n9378) );
  NAND2_X1 U10598 ( .A1(n9378), .A2(n10370), .ZN(n9190) );
  OAI211_X1 U10599 ( .C1(n9382), .C2(n9349), .A(n9191), .B(n9190), .ZN(
        P2_U3272) );
  OAI21_X1 U10600 ( .B1(n5054), .B2(n9201), .A(n9192), .ZN(n9387) );
  INV_X1 U10601 ( .A(n9213), .ZN(n9195) );
  INV_X1 U10602 ( .A(n9193), .ZN(n9194) );
  AOI21_X1 U10603 ( .B1(n9383), .B2(n9195), .A(n9194), .ZN(n9384) );
  INV_X1 U10604 ( .A(n9196), .ZN(n9197) );
  AOI22_X1 U10605 ( .A1(n9197), .A2(n9335), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n10357), .ZN(n9198) );
  OAI21_X1 U10606 ( .B1(n9199), .B2(n9338), .A(n9198), .ZN(n9210) );
  INV_X1 U10607 ( .A(n9200), .ZN(n9203) );
  OAI21_X1 U10608 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9205) );
  NAND2_X1 U10609 ( .A1(n9205), .A2(n9204), .ZN(n9208) );
  AOI222_X1 U10610 ( .A1(n10365), .A2(n9208), .B1(n9207), .B2(n10360), .C1(
        n9206), .C2(n10362), .ZN(n9386) );
  NOR2_X1 U10611 ( .A1(n9386), .A2(n10357), .ZN(n9209) );
  AOI211_X1 U10612 ( .C1(n9384), .C2(n9347), .A(n9210), .B(n9209), .ZN(n9211)
         );
  OAI21_X1 U10613 ( .B1(n9387), .B2(n9349), .A(n9211), .ZN(P2_U3273) );
  XNOR2_X1 U10614 ( .A(n9212), .B(n4966), .ZN(n9392) );
  AOI21_X1 U10615 ( .B1(n9388), .B2(n9225), .A(n9213), .ZN(n9389) );
  INV_X1 U10616 ( .A(n9388), .ZN(n9216) );
  AOI22_X1 U10617 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n10357), .B1(n9214), 
        .B2(n9335), .ZN(n9215) );
  OAI21_X1 U10618 ( .B1(n9216), .B2(n9338), .A(n9215), .ZN(n9221) );
  OAI211_X1 U10619 ( .C1(n4548), .C2(n9217), .A(n9200), .B(n10365), .ZN(n9219)
         );
  AOI22_X1 U10620 ( .A1(n9082), .A2(n10362), .B1(n10360), .B2(n9242), .ZN(
        n9218) );
  NOR2_X1 U10621 ( .A1(n9391), .A2(n10357), .ZN(n9220) );
  AOI211_X1 U10622 ( .C1(n9389), .C2(n9347), .A(n9221), .B(n9220), .ZN(n9222)
         );
  OAI21_X1 U10623 ( .B1(n9392), .B2(n9349), .A(n9222), .ZN(P2_U3274) );
  XOR2_X1 U10624 ( .A(n9234), .B(n9223), .Z(n9398) );
  INV_X1 U10625 ( .A(n9224), .ZN(n9227) );
  INV_X1 U10626 ( .A(n9225), .ZN(n9226) );
  AOI21_X1 U10627 ( .B1(n9394), .B2(n9227), .A(n9226), .ZN(n9395) );
  NOR2_X1 U10628 ( .A1(n9228), .A2(n9338), .ZN(n9232) );
  OAI22_X1 U10629 ( .A1(n10370), .A2(n9230), .B1(n9229), .B2(n10375), .ZN(
        n9231) );
  AOI211_X1 U10630 ( .C1(n9395), .C2(n9347), .A(n9232), .B(n9231), .ZN(n9240)
         );
  AOI21_X1 U10631 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9236) );
  OAI222_X1 U10632 ( .A1(n9311), .A2(n9238), .B1(n9309), .B2(n9237), .C1(n9293), .C2(n9236), .ZN(n9393) );
  NAND2_X1 U10633 ( .A1(n9393), .A2(n10370), .ZN(n9239) );
  OAI211_X1 U10634 ( .C1(n9398), .C2(n9349), .A(n9240), .B(n9239), .ZN(
        P2_U3275) );
  XNOR2_X1 U10635 ( .A(n9241), .B(n9244), .ZN(n9243) );
  AOI222_X1 U10636 ( .A1(n10365), .A2(n9243), .B1(n9242), .B2(n10362), .C1(
        n9279), .C2(n10360), .ZN(n9403) );
  INV_X1 U10637 ( .A(n9405), .ZN(n9246) );
  NAND2_X1 U10638 ( .A1(n9245), .A2(n9244), .ZN(n9399) );
  NAND3_X1 U10639 ( .A1(n9246), .A2(n10358), .A3(n9399), .ZN(n9253) );
  XOR2_X1 U10640 ( .A(n9400), .B(n9408), .Z(n9401) );
  INV_X1 U10641 ( .A(n9400), .ZN(n9247) );
  NOR2_X1 U10642 ( .A1(n9247), .A2(n9338), .ZN(n9251) );
  OAI22_X1 U10643 ( .A1(n10370), .A2(n9249), .B1(n9248), .B2(n10375), .ZN(
        n9250) );
  AOI211_X1 U10644 ( .C1(n9401), .C2(n9347), .A(n9251), .B(n9250), .ZN(n9252)
         );
  OAI211_X1 U10645 ( .C1(n10357), .C2(n9403), .A(n9253), .B(n9252), .ZN(
        P2_U3276) );
  XOR2_X1 U10646 ( .A(n9258), .B(n9254), .Z(n9412) );
  OAI22_X1 U10647 ( .A1(n10370), .A2(n9256), .B1(n9255), .B2(n10375), .ZN(
        n9267) );
  OAI21_X1 U10648 ( .B1(n9259), .B2(n9258), .A(n9257), .ZN(n9262) );
  AOI222_X1 U10649 ( .A1(n10365), .A2(n9262), .B1(n9261), .B2(n10362), .C1(
        n9260), .C2(n10360), .ZN(n9411) );
  NOR2_X1 U10650 ( .A1(n9271), .A2(n9263), .ZN(n9406) );
  INV_X1 U10651 ( .A(n9406), .ZN(n9264) );
  NAND3_X1 U10652 ( .A1(n9264), .A2(n8625), .A3(n9408), .ZN(n9265) );
  AOI21_X1 U10653 ( .B1(n9411), .B2(n9265), .A(n10357), .ZN(n9266) );
  AOI211_X1 U10654 ( .C1(n9325), .C2(n9407), .A(n9267), .B(n9266), .ZN(n9268)
         );
  OAI21_X1 U10655 ( .B1(n9412), .B2(n9349), .A(n9268), .ZN(P2_U3277) );
  AOI21_X1 U10656 ( .B1(n9270), .B2(n9277), .A(n9269), .ZN(n9417) );
  AOI21_X1 U10657 ( .B1(n9413), .B2(n9288), .A(n9271), .ZN(n9414) );
  INV_X1 U10658 ( .A(n9272), .ZN(n9273) );
  AOI22_X1 U10659 ( .A1(n10357), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9273), 
        .B2(n9335), .ZN(n9274) );
  OAI21_X1 U10660 ( .B1(n9275), .B2(n9338), .A(n9274), .ZN(n9282) );
  XOR2_X1 U10661 ( .A(n9277), .B(n9276), .Z(n9280) );
  AOI222_X1 U10662 ( .A1(n10365), .A2(n9280), .B1(n9279), .B2(n10362), .C1(
        n9278), .C2(n10360), .ZN(n9416) );
  NOR2_X1 U10663 ( .A1(n9416), .A2(n10357), .ZN(n9281) );
  AOI211_X1 U10664 ( .C1(n9414), .C2(n9347), .A(n9282), .B(n9281), .ZN(n9283)
         );
  OAI21_X1 U10665 ( .B1(n9349), .B2(n9417), .A(n9283), .ZN(P2_U3278) );
  AOI21_X1 U10666 ( .B1(n9285), .B2(n9284), .A(n4547), .ZN(n9422) );
  OAI22_X1 U10667 ( .A1(n10370), .A2(n9287), .B1(n9286), .B2(n10375), .ZN(
        n9300) );
  INV_X1 U10668 ( .A(n9320), .ZN(n9290) );
  INV_X1 U10669 ( .A(n9288), .ZN(n9289) );
  AOI211_X1 U10670 ( .C1(n9420), .C2(n9290), .A(n10436), .B(n9289), .ZN(n9419)
         );
  XNOR2_X1 U10671 ( .A(n9292), .B(n9291), .ZN(n9294) );
  OAI222_X1 U10672 ( .A1(n9311), .A2(n9296), .B1(n9309), .B2(n9295), .C1(n9294), .C2(n9293), .ZN(n9418) );
  AOI21_X1 U10673 ( .B1(n9419), .B2(n9297), .A(n9418), .ZN(n9298) );
  NOR2_X1 U10674 ( .A1(n9298), .A2(n10357), .ZN(n9299) );
  AOI211_X1 U10675 ( .C1(n9325), .C2(n9420), .A(n9300), .B(n9299), .ZN(n9301)
         );
  OAI21_X1 U10676 ( .B1(n9349), .B2(n9422), .A(n9301), .ZN(P2_U3279) );
  AND2_X1 U10677 ( .A1(n9329), .A2(n9302), .ZN(n9305) );
  OAI21_X1 U10678 ( .B1(n9305), .B2(n9304), .A(n9303), .ZN(n9428) );
  OAI21_X1 U10679 ( .B1(n9308), .B2(n9307), .A(n9306), .ZN(n9316) );
  OAI22_X1 U10680 ( .A1(n9312), .A2(n9311), .B1(n9310), .B2(n9309), .ZN(n9315)
         );
  NOR2_X1 U10681 ( .A1(n9428), .A2(n9313), .ZN(n9314) );
  AOI211_X1 U10682 ( .C1(n10365), .C2(n9316), .A(n9315), .B(n9314), .ZN(n9427)
         );
  OR2_X1 U10683 ( .A1(n9427), .A2(n10357), .ZN(n9327) );
  OAI22_X1 U10684 ( .A1(n10370), .A2(n9318), .B1(n9317), .B2(n10375), .ZN(
        n9323) );
  NOR2_X1 U10685 ( .A1(n9332), .A2(n9423), .ZN(n9319) );
  OR2_X1 U10686 ( .A1(n9320), .A2(n9319), .ZN(n9424) );
  NOR2_X1 U10687 ( .A1(n9424), .A2(n9321), .ZN(n9322) );
  AOI211_X1 U10688 ( .C1(n9325), .C2(n9324), .A(n9323), .B(n9322), .ZN(n9326)
         );
  OAI211_X1 U10689 ( .C1(n9428), .C2(n9328), .A(n9327), .B(n9326), .ZN(
        P2_U3280) );
  OAI21_X1 U10690 ( .B1(n9330), .B2(n9340), .A(n9329), .ZN(n9331) );
  INV_X1 U10691 ( .A(n9331), .ZN(n9433) );
  AOI21_X1 U10692 ( .B1(n9429), .B2(n9333), .A(n9332), .ZN(n9430) );
  INV_X1 U10693 ( .A(n9334), .ZN(n9336) );
  AOI22_X1 U10694 ( .A1(n10357), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9336), 
        .B2(n9335), .ZN(n9337) );
  OAI21_X1 U10695 ( .B1(n9339), .B2(n9338), .A(n9337), .ZN(n9346) );
  XNOR2_X1 U10696 ( .A(n9341), .B(n9340), .ZN(n9344) );
  AOI222_X1 U10697 ( .A1(n10365), .A2(n9344), .B1(n9343), .B2(n10362), .C1(
        n9342), .C2(n10360), .ZN(n9432) );
  NOR2_X1 U10698 ( .A1(n9432), .A2(n10357), .ZN(n9345) );
  AOI211_X1 U10699 ( .C1(n9430), .C2(n9347), .A(n9346), .B(n9345), .ZN(n9348)
         );
  OAI21_X1 U10700 ( .B1(n9349), .B2(n9433), .A(n9348), .ZN(P2_U3281) );
  NAND2_X1 U10701 ( .A1(n9350), .A2(n9437), .ZN(n9351) );
  OAI211_X1 U10702 ( .C1(n9352), .C2(n10436), .A(n10113), .B(n9351), .ZN(n9440) );
  MUX2_X1 U10703 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9440), .S(n10455), .Z(
        P2_U3551) );
  NAND2_X1 U10704 ( .A1(n9353), .A2(n10440), .ZN(n9357) );
  MUX2_X1 U10705 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9441), .S(n10455), .Z(
        P2_U3549) );
  AOI22_X1 U10706 ( .A1(n9359), .A2(n10411), .B1(n9437), .B2(n9358), .ZN(n9360) );
  OAI211_X1 U10707 ( .C1(n9362), .C2(n10426), .A(n9361), .B(n9360), .ZN(n9442)
         );
  MUX2_X1 U10708 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9442), .S(n10455), .Z(
        P2_U3548) );
  AOI22_X1 U10709 ( .A1(n9364), .A2(n10411), .B1(n9437), .B2(n9363), .ZN(n9365) );
  OAI211_X1 U10710 ( .C1(n9367), .C2(n10426), .A(n9366), .B(n9365), .ZN(n9443)
         );
  MUX2_X1 U10711 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9443), .S(n10455), .Z(
        P2_U3547) );
  AOI21_X1 U10712 ( .B1(n9437), .B2(n9369), .A(n9368), .ZN(n9370) );
  OAI211_X1 U10713 ( .C1(n9372), .C2(n10426), .A(n9371), .B(n9370), .ZN(n9444)
         );
  MUX2_X1 U10714 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9444), .S(n10455), .Z(
        P2_U3546) );
  AOI21_X1 U10715 ( .B1(n9437), .B2(n9374), .A(n9373), .ZN(n9375) );
  OAI211_X1 U10716 ( .C1(n9377), .C2(n10426), .A(n9376), .B(n9375), .ZN(n9445)
         );
  MUX2_X1 U10717 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9445), .S(n10455), .Z(
        P2_U3545) );
  AOI211_X1 U10718 ( .C1(n9437), .C2(n9380), .A(n9379), .B(n9378), .ZN(n9381)
         );
  OAI21_X1 U10719 ( .B1(n9382), .B2(n10426), .A(n9381), .ZN(n9446) );
  MUX2_X1 U10720 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9446), .S(n10455), .Z(
        P2_U3544) );
  AOI22_X1 U10721 ( .A1(n9384), .A2(n10411), .B1(n9437), .B2(n9383), .ZN(n9385) );
  OAI211_X1 U10722 ( .C1(n9387), .C2(n10426), .A(n9386), .B(n9385), .ZN(n9447)
         );
  MUX2_X1 U10723 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9447), .S(n10455), .Z(
        P2_U3543) );
  AOI22_X1 U10724 ( .A1(n9389), .A2(n10411), .B1(n9437), .B2(n9388), .ZN(n9390) );
  OAI211_X1 U10725 ( .C1(n9392), .C2(n10426), .A(n9391), .B(n9390), .ZN(n9448)
         );
  MUX2_X1 U10726 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9448), .S(n10455), .Z(
        P2_U3542) );
  INV_X1 U10727 ( .A(n9393), .ZN(n9397) );
  AOI22_X1 U10728 ( .A1(n9395), .A2(n10411), .B1(n9437), .B2(n9394), .ZN(n9396) );
  OAI211_X1 U10729 ( .C1(n9398), .C2(n10426), .A(n9397), .B(n9396), .ZN(n9449)
         );
  MUX2_X1 U10730 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9449), .S(n10455), .Z(
        P2_U3541) );
  NAND2_X1 U10731 ( .A1(n9399), .A2(n10440), .ZN(n9404) );
  AOI22_X1 U10732 ( .A1(n9401), .A2(n10411), .B1(n9437), .B2(n9400), .ZN(n9402) );
  OAI211_X1 U10733 ( .C1(n9405), .C2(n9404), .A(n9403), .B(n9402), .ZN(n9450)
         );
  MUX2_X1 U10734 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9450), .S(n10455), .Z(
        P2_U3540) );
  NOR2_X1 U10735 ( .A1(n9406), .A2(n10436), .ZN(n9409) );
  AOI22_X1 U10736 ( .A1(n9409), .A2(n9408), .B1(n9437), .B2(n9407), .ZN(n9410)
         );
  OAI211_X1 U10737 ( .C1(n9412), .C2(n10426), .A(n9411), .B(n9410), .ZN(n9451)
         );
  MUX2_X1 U10738 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9451), .S(n10455), .Z(
        P2_U3539) );
  AOI22_X1 U10739 ( .A1(n9414), .A2(n10411), .B1(n9437), .B2(n9413), .ZN(n9415) );
  OAI211_X1 U10740 ( .C1(n9417), .C2(n10426), .A(n9416), .B(n9415), .ZN(n9452)
         );
  MUX2_X1 U10741 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9452), .S(n10455), .Z(
        P2_U3538) );
  AOI211_X1 U10742 ( .C1(n9437), .C2(n9420), .A(n9419), .B(n9418), .ZN(n9421)
         );
  OAI21_X1 U10743 ( .B1(n9422), .B2(n10426), .A(n9421), .ZN(n9453) );
  MUX2_X1 U10744 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9453), .S(n10455), .Z(
        P2_U3537) );
  OAI22_X1 U10745 ( .A1(n9424), .A2(n10436), .B1(n9423), .B2(n10434), .ZN(
        n9425) );
  INV_X1 U10746 ( .A(n9425), .ZN(n9426) );
  OAI211_X1 U10747 ( .C1(n10418), .C2(n9428), .A(n9427), .B(n9426), .ZN(n9454)
         );
  MUX2_X1 U10748 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9454), .S(n10455), .Z(
        P2_U3536) );
  AOI22_X1 U10749 ( .A1(n9430), .A2(n10411), .B1(n9437), .B2(n9429), .ZN(n9431) );
  OAI211_X1 U10750 ( .C1(n9433), .C2(n10426), .A(n9432), .B(n9431), .ZN(n9455)
         );
  MUX2_X1 U10751 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9455), .S(n10455), .Z(
        P2_U3535) );
  AOI211_X1 U10752 ( .C1(n9437), .C2(n9436), .A(n9435), .B(n9434), .ZN(n9438)
         );
  OAI21_X1 U10753 ( .B1(n10426), .B2(n9439), .A(n9438), .ZN(n9456) );
  MUX2_X1 U10754 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9456), .S(n10455), .Z(
        P2_U3534) );
  MUX2_X1 U10755 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9440), .S(n10444), .Z(
        P2_U3519) );
  MUX2_X1 U10756 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9441), .S(n10444), .Z(
        P2_U3517) );
  MUX2_X1 U10757 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9442), .S(n10444), .Z(
        P2_U3516) );
  MUX2_X1 U10758 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9443), .S(n10444), .Z(
        P2_U3515) );
  MUX2_X1 U10759 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9444), .S(n10444), .Z(
        P2_U3514) );
  MUX2_X1 U10760 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9445), .S(n10444), .Z(
        P2_U3513) );
  MUX2_X1 U10761 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9446), .S(n10444), .Z(
        P2_U3512) );
  MUX2_X1 U10762 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9447), .S(n10444), .Z(
        P2_U3511) );
  MUX2_X1 U10763 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9448), .S(n10444), .Z(
        P2_U3510) );
  MUX2_X1 U10764 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9449), .S(n10444), .Z(
        P2_U3509) );
  MUX2_X1 U10765 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9450), .S(n10444), .Z(
        P2_U3508) );
  MUX2_X1 U10766 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9451), .S(n10444), .Z(
        P2_U3507) );
  MUX2_X1 U10767 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9452), .S(n10444), .Z(
        P2_U3505) );
  MUX2_X1 U10768 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9453), .S(n10444), .Z(
        P2_U3502) );
  MUX2_X1 U10769 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9454), .S(n10444), .Z(
        P2_U3499) );
  MUX2_X1 U10770 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9455), .S(n10444), .Z(
        P2_U3496) );
  MUX2_X1 U10771 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9456), .S(n10444), .Z(
        P2_U3493) );
  INV_X1 U10772 ( .A(n9457), .ZN(n10082) );
  NOR4_X1 U10773 ( .A1(n6123), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6183), .A4(
        P2_U3152), .ZN(n9458) );
  AOI21_X1 U10774 ( .B1(n9471), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9458), .ZN(
        n9459) );
  OAI21_X1 U10775 ( .B1(n10082), .B2(n9463), .A(n9459), .ZN(P2_U3327) );
  INV_X1 U10776 ( .A(n9460), .ZN(n10084) );
  AOI22_X1 U10777 ( .A1(n9461), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9471), .ZN(n9462) );
  OAI21_X1 U10778 ( .B1(n10084), .B2(n9463), .A(n9462), .ZN(P2_U3328) );
  INV_X1 U10779 ( .A(n9464), .ZN(n10089) );
  AOI22_X1 U10780 ( .A1(n9465), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9471), .ZN(n9466) );
  OAI21_X1 U10781 ( .B1(n10089), .B2(n9469), .A(n9466), .ZN(P2_U3329) );
  INV_X1 U10782 ( .A(n10091), .ZN(n9470) );
  NAND2_X1 U10783 ( .A1(n9471), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9468) );
  OAI211_X1 U10784 ( .C1(n9470), .C2(n9469), .A(n9468), .B(n9467), .ZN(
        P2_U3330) );
  INV_X1 U10785 ( .A(n10096), .ZN(n9474) );
  AOI22_X1 U10786 ( .A1(n9472), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9471), .ZN(n9473) );
  OAI21_X1 U10787 ( .B1(n9474), .B2(n9463), .A(n9473), .ZN(P2_U3331) );
  MUX2_X1 U10788 ( .A(n9475), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10789 ( .A(n9476), .ZN(n9478) );
  NOR2_X1 U10790 ( .A1(n9478), .A2(n9477), .ZN(n9479) );
  XNOR2_X1 U10791 ( .A(n9480), .B(n9479), .ZN(n9485) );
  AOI22_X1 U10792 ( .A1(n9657), .A2(n9609), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9482) );
  NAND2_X1 U10793 ( .A1(n9781), .A2(n9642), .ZN(n9481) );
  OAI211_X1 U10794 ( .C1(n9786), .C2(n9578), .A(n9482), .B(n9481), .ZN(n9483)
         );
  AOI21_X1 U10795 ( .B1(n9979), .B2(n9612), .A(n9483), .ZN(n9484) );
  OAI21_X1 U10796 ( .B1(n9485), .B2(n9651), .A(n9484), .ZN(P1_U3212) );
  NAND2_X1 U10797 ( .A1(n9487), .A2(n9486), .ZN(n9488) );
  XOR2_X1 U10798 ( .A(n9489), .B(n9488), .Z(n9499) );
  INV_X1 U10799 ( .A(n9490), .ZN(n9491) );
  AOI21_X1 U10800 ( .B1(n9640), .B2(n9660), .A(n9491), .ZN(n9494) );
  NAND2_X1 U10801 ( .A1(n9642), .A2(n9492), .ZN(n9493) );
  OAI211_X1 U10802 ( .C1(n9646), .C2(n9495), .A(n9494), .B(n9493), .ZN(n9496)
         );
  AOI21_X1 U10803 ( .B1(n9497), .B2(n9648), .A(n9496), .ZN(n9498) );
  OAI21_X1 U10804 ( .B1(n9499), .B2(n9651), .A(n9498), .ZN(P1_U3213) );
  NAND2_X1 U10805 ( .A1(n9501), .A2(n9500), .ZN(n9503) );
  XNOR2_X1 U10806 ( .A(n9503), .B(n9502), .ZN(n9508) );
  NAND2_X1 U10807 ( .A1(n9659), .A2(n9640), .ZN(n9505) );
  AOI22_X1 U10808 ( .A1(n9883), .A2(n9609), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9504) );
  OAI211_X1 U10809 ( .C1(n9622), .C2(n9841), .A(n9505), .B(n9504), .ZN(n9506)
         );
  AOI21_X1 U10810 ( .B1(n9998), .B2(n9648), .A(n9506), .ZN(n9507) );
  OAI21_X1 U10811 ( .B1(n9508), .B2(n9651), .A(n9507), .ZN(P1_U3214) );
  XOR2_X1 U10812 ( .A(n9510), .B(n9509), .Z(n9511) );
  XNOR2_X1 U10813 ( .A(n9512), .B(n9511), .ZN(n9517) );
  NAND2_X1 U10814 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9736) );
  OAI21_X1 U10815 ( .B1(n9646), .B2(n9906), .A(n9736), .ZN(n9513) );
  AOI21_X1 U10816 ( .B1(n9640), .B2(n9882), .A(n9513), .ZN(n9514) );
  OAI21_X1 U10817 ( .B1(n9622), .B2(n9911), .A(n9514), .ZN(n9515) );
  AOI21_X1 U10818 ( .B1(n9910), .B2(n9612), .A(n9515), .ZN(n9516) );
  OAI21_X1 U10819 ( .B1(n9517), .B2(n9651), .A(n9516), .ZN(P1_U3217) );
  XOR2_X1 U10820 ( .A(n9519), .B(n9518), .Z(n9524) );
  AOI22_X1 U10821 ( .A1(n9883), .A2(n9640), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9521) );
  NAND2_X1 U10822 ( .A1(n9609), .A2(n9882), .ZN(n9520) );
  OAI211_X1 U10823 ( .C1(n9622), .C2(n9873), .A(n9521), .B(n9520), .ZN(n9522)
         );
  AOI21_X1 U10824 ( .B1(n10009), .B2(n9612), .A(n9522), .ZN(n9523) );
  OAI21_X1 U10825 ( .B1(n9524), .B2(n9651), .A(n9523), .ZN(P1_U3221) );
  XOR2_X1 U10826 ( .A(n9526), .B(n9525), .Z(n9532) );
  INV_X1 U10827 ( .A(n9527), .ZN(n9816) );
  AOI22_X1 U10828 ( .A1(n9816), .A2(n9642), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9529) );
  NAND2_X1 U10829 ( .A1(n9659), .A2(n9609), .ZN(n9528) );
  OAI211_X1 U10830 ( .C1(n9812), .C2(n9578), .A(n9529), .B(n9528), .ZN(n9530)
         );
  AOI21_X1 U10831 ( .B1(n9990), .B2(n9648), .A(n9530), .ZN(n9531) );
  OAI21_X1 U10832 ( .B1(n9532), .B2(n9651), .A(n9531), .ZN(P1_U3223) );
  INV_X1 U10833 ( .A(n9534), .ZN(n9535) );
  AOI21_X1 U10834 ( .B1(n9536), .B2(n9533), .A(n9535), .ZN(n9541) );
  AOI22_X1 U10835 ( .A1(n9609), .A2(n9660), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n9538) );
  NAND2_X1 U10836 ( .A1(n9642), .A2(n9964), .ZN(n9537) );
  OAI211_X1 U10837 ( .C1(n9958), .C2(n9578), .A(n9538), .B(n9537), .ZN(n9539)
         );
  AOI21_X1 U10838 ( .B1(n9962), .B2(n9612), .A(n9539), .ZN(n9540) );
  OAI21_X1 U10839 ( .B1(n9541), .B2(n9651), .A(n9540), .ZN(P1_U3224) );
  NAND2_X1 U10840 ( .A1(n9544), .A2(n9607), .ZN(n9551) );
  AOI22_X1 U10841 ( .A1(n9545), .A2(n9612), .B1(n9609), .B2(n5955), .ZN(n9550)
         );
  AND2_X1 U10842 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U10843 ( .A1(n9578), .A2(n9546), .ZN(n9547) );
  AOI211_X1 U10844 ( .C1(n9548), .C2(n9642), .A(n10236), .B(n9547), .ZN(n9549)
         );
  NAND3_X1 U10845 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(P1_U3225) );
  OAI21_X1 U10846 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9555) );
  NAND2_X1 U10847 ( .A1(n9555), .A2(n9607), .ZN(n9561) );
  INV_X1 U10848 ( .A(n9556), .ZN(n9939) );
  AOI22_X1 U10849 ( .A1(n9640), .A2(n9945), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n9557) );
  OAI21_X1 U10850 ( .B1(n9558), .B2(n9646), .A(n9557), .ZN(n9559) );
  AOI21_X1 U10851 ( .B1(n9939), .B2(n9642), .A(n9559), .ZN(n9560) );
  OAI211_X1 U10852 ( .C1(n9941), .C2(n9634), .A(n9561), .B(n9560), .ZN(
        P1_U3226) );
  XOR2_X1 U10853 ( .A(n9563), .B(n9562), .Z(n9568) );
  AOI22_X1 U10854 ( .A1(n9865), .A2(n9609), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9565) );
  NAND2_X1 U10855 ( .A1(n9833), .A2(n9642), .ZN(n9564) );
  OAI211_X1 U10856 ( .C1(n9828), .C2(n9578), .A(n9565), .B(n9564), .ZN(n9566)
         );
  AOI21_X1 U10857 ( .B1(n9832), .B2(n9612), .A(n9566), .ZN(n9567) );
  OAI21_X1 U10858 ( .B1(n9568), .B2(n9651), .A(n9567), .ZN(P1_U3227) );
  NAND2_X1 U10859 ( .A1(n9570), .A2(n9569), .ZN(n9572) );
  AOI21_X1 U10860 ( .B1(n9572), .B2(n9571), .A(n9651), .ZN(n9574) );
  OR2_X1 U10861 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  NAND2_X1 U10862 ( .A1(n9574), .A2(n9573), .ZN(n9583) );
  AOI22_X1 U10863 ( .A1(n9575), .A2(n9612), .B1(n9609), .B2(n9668), .ZN(n9582)
         );
  NOR2_X1 U10864 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9576), .ZN(n10226) );
  NOR2_X1 U10865 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  AOI211_X1 U10866 ( .C1(n9580), .C2(n9642), .A(n10226), .B(n9579), .ZN(n9581)
         );
  NAND3_X1 U10867 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(P1_U3228) );
  INV_X1 U10868 ( .A(n9895), .ZN(n10066) );
  INV_X1 U10869 ( .A(n9585), .ZN(n9589) );
  OAI21_X1 U10870 ( .B1(n9587), .B2(n9589), .A(n9586), .ZN(n9588) );
  OAI21_X1 U10871 ( .B1(n9584), .B2(n9589), .A(n9588), .ZN(n9590) );
  NAND2_X1 U10872 ( .A1(n9590), .A2(n9607), .ZN(n9594) );
  AOI22_X1 U10873 ( .A1(n9864), .A2(n9640), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9591) );
  OAI21_X1 U10874 ( .B1(n9893), .B2(n9646), .A(n9591), .ZN(n9592) );
  AOI21_X1 U10875 ( .B1(n9896), .B2(n9642), .A(n9592), .ZN(n9593) );
  OAI211_X1 U10876 ( .C1(n10066), .C2(n9634), .A(n9594), .B(n9593), .ZN(
        P1_U3231) );
  NAND2_X1 U10877 ( .A1(n9595), .A2(n9596), .ZN(n9598) );
  XNOR2_X1 U10878 ( .A(n9598), .B(n9597), .ZN(n9603) );
  NAND2_X1 U10879 ( .A1(n9865), .A2(n9640), .ZN(n9600) );
  AOI22_X1 U10880 ( .A1(n9864), .A2(n9609), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9599) );
  OAI211_X1 U10881 ( .C1(n9622), .C2(n9858), .A(n9600), .B(n9599), .ZN(n9601)
         );
  AOI21_X1 U10882 ( .B1(n10003), .B2(n9648), .A(n9601), .ZN(n9602) );
  OAI21_X1 U10883 ( .B1(n9603), .B2(n9651), .A(n9602), .ZN(P1_U3233) );
  OAI21_X1 U10884 ( .B1(n9604), .B2(n9605), .A(n9606), .ZN(n9608) );
  NAND2_X1 U10885 ( .A1(n9608), .A2(n9607), .ZN(n9615) );
  AOI22_X1 U10886 ( .A1(n9640), .A2(n9668), .B1(n9609), .B2(n5950), .ZN(n9614)
         );
  AOI22_X1 U10887 ( .A1(n9612), .A2(n9611), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9610), .ZN(n9613) );
  NAND3_X1 U10888 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(P1_U3235) );
  NAND2_X1 U10889 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  XOR2_X1 U10890 ( .A(n9619), .B(n9618), .Z(n9625) );
  NAND2_X1 U10891 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9725) );
  OAI21_X1 U10892 ( .B1(n9646), .B2(n9958), .A(n9725), .ZN(n9620) );
  AOI21_X1 U10893 ( .B1(n9640), .B2(n9920), .A(n9620), .ZN(n9621) );
  OAI21_X1 U10894 ( .B1(n9622), .B2(n9927), .A(n9621), .ZN(n9623) );
  AOI21_X1 U10895 ( .B1(n10025), .B2(n9648), .A(n9623), .ZN(n9624) );
  OAI21_X1 U10896 ( .B1(n9625), .B2(n9651), .A(n9624), .ZN(P1_U3236) );
  NAND2_X1 U10897 ( .A1(n9628), .A2(n9627), .ZN(n9633) );
  INV_X1 U10898 ( .A(n9629), .ZN(n9802) );
  AOI22_X1 U10899 ( .A1(n9802), .A2(n9642), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9630) );
  OAI21_X1 U10900 ( .B1(n9828), .B2(n9646), .A(n9630), .ZN(n9631) );
  AOI21_X1 U10901 ( .B1(n9640), .B2(n9656), .A(n9631), .ZN(n9632) );
  OAI211_X1 U10902 ( .C1(n10054), .C2(n9634), .A(n9633), .B(n9632), .ZN(
        P1_U3238) );
  NAND2_X1 U10903 ( .A1(n9635), .A2(n9636), .ZN(n9637) );
  XOR2_X1 U10904 ( .A(n9638), .B(n9637), .Z(n9652) );
  NAND2_X1 U10905 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9681) );
  INV_X1 U10906 ( .A(n9681), .ZN(n9639) );
  AOI21_X1 U10907 ( .B1(n9640), .B2(n9944), .A(n9639), .ZN(n9644) );
  NAND2_X1 U10908 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  OAI211_X1 U10909 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9647)
         );
  AOI21_X1 U10910 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(n9650) );
  OAI21_X1 U10911 ( .B1(n9652), .B2(n9651), .A(n9650), .ZN(P1_U3239) );
  MUX2_X1 U10912 ( .A(n9653), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10211), .Z(
        P1_U3585) );
  MUX2_X1 U10913 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9654), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10914 ( .A(n9655), .B(P1_DATAO_REG_28__SCAN_IN), .S(n10211), .Z(
        P1_U3583) );
  MUX2_X1 U10915 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9656), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10916 ( .A(n9657), .B(P1_DATAO_REG_26__SCAN_IN), .S(n10211), .Z(
        P1_U3581) );
  MUX2_X1 U10917 ( .A(n9658), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10211), .Z(
        P1_U3580) );
  MUX2_X1 U10918 ( .A(n9659), .B(P1_DATAO_REG_24__SCAN_IN), .S(n10211), .Z(
        P1_U3579) );
  MUX2_X1 U10919 ( .A(n9865), .B(P1_DATAO_REG_23__SCAN_IN), .S(n10211), .Z(
        P1_U3578) );
  MUX2_X1 U10920 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9883), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10921 ( .A(n9864), .B(P1_DATAO_REG_21__SCAN_IN), .S(n10211), .Z(
        P1_U3576) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9882), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10923 ( .A(n9920), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10211), .Z(
        P1_U3574) );
  MUX2_X1 U10924 ( .A(n9945), .B(P1_DATAO_REG_18__SCAN_IN), .S(n10211), .Z(
        P1_U3573) );
  MUX2_X1 U10925 ( .A(n9919), .B(P1_DATAO_REG_17__SCAN_IN), .S(n10211), .Z(
        P1_U3572) );
  MUX2_X1 U10926 ( .A(n9944), .B(P1_DATAO_REG_16__SCAN_IN), .S(n10211), .Z(
        P1_U3571) );
  MUX2_X1 U10927 ( .A(n9660), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10211), .Z(
        P1_U3570) );
  MUX2_X1 U10928 ( .A(n10126), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10211), .Z(
        P1_U3569) );
  MUX2_X1 U10929 ( .A(n9661), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10211), .Z(
        P1_U3568) );
  MUX2_X1 U10930 ( .A(n10150), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10211), .Z(
        P1_U3567) );
  MUX2_X1 U10931 ( .A(n9662), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10211), .Z(
        P1_U3566) );
  MUX2_X1 U10932 ( .A(n10148), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10211), .Z(
        P1_U3565) );
  MUX2_X1 U10933 ( .A(n9663), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10211), .Z(
        P1_U3564) );
  MUX2_X1 U10934 ( .A(n9664), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10211), .Z(
        P1_U3563) );
  MUX2_X1 U10935 ( .A(n9665), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10211), .Z(
        P1_U3562) );
  MUX2_X1 U10936 ( .A(n9666), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10211), .Z(
        P1_U3561) );
  MUX2_X1 U10937 ( .A(n9667), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10211), .Z(
        P1_U3560) );
  MUX2_X1 U10938 ( .A(n5955), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10211), .Z(
        P1_U3559) );
  MUX2_X1 U10939 ( .A(n9668), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10211), .Z(
        P1_U3558) );
  MUX2_X1 U10940 ( .A(n9669), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10211), .Z(
        P1_U3557) );
  MUX2_X1 U10941 ( .A(n5950), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10211), .Z(
        P1_U3556) );
  MUX2_X1 U10942 ( .A(n9670), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10211), .Z(
        P1_U3555) );
  INV_X1 U10943 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9676) );
  INV_X1 U10944 ( .A(n9671), .ZN(n9673) );
  XOR2_X1 U10945 ( .A(n9694), .B(n9687), .Z(n9675) );
  AOI211_X1 U10946 ( .C1(n9676), .C2(n9675), .A(n10296), .B(n9688), .ZN(n9686)
         );
  INV_X1 U10947 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10170) );
  AOI21_X1 U10948 ( .B1(n8159), .B2(n9678), .A(n9677), .ZN(n9695) );
  INV_X1 U10949 ( .A(n9695), .ZN(n9679) );
  XOR2_X1 U10950 ( .A(n9694), .B(n9679), .Z(n9680) );
  AOI211_X1 U10951 ( .C1(n10170), .C2(n9680), .A(n10288), .B(n9693), .ZN(n9685) );
  NAND2_X1 U10952 ( .A1(n10306), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9682) );
  OAI211_X1 U10953 ( .C1(n10254), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9684)
         );
  OR3_X1 U10954 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(P1_U3256) );
  INV_X1 U10955 ( .A(n9687), .ZN(n9689) );
  NAND2_X1 U10956 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9712), .ZN(n9690) );
  OAI21_X1 U10957 ( .B1(n9712), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9690), .ZN(
        n9691) );
  AOI211_X1 U10958 ( .C1(n9692), .C2(n9691), .A(n9707), .B(n10296), .ZN(n9706)
         );
  AOI21_X1 U10959 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9700) );
  INV_X1 U10960 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9696) );
  OR2_X1 U10961 ( .A1(n9712), .A2(n9696), .ZN(n9698) );
  NAND2_X1 U10962 ( .A1(n9712), .A2(n9696), .ZN(n9697) );
  AND2_X1 U10963 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  NOR2_X1 U10964 ( .A1(n9700), .A2(n9699), .ZN(n9711) );
  AOI211_X1 U10965 ( .C1(n9700), .C2(n9699), .A(n9711), .B(n10288), .ZN(n9705)
         );
  NAND2_X1 U10966 ( .A1(n10306), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9702) );
  NAND2_X1 U10967 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9701) );
  OAI211_X1 U10968 ( .C1(n10254), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9704)
         );
  OR3_X1 U10969 ( .A1(n9706), .A2(n9705), .A3(n9704), .ZN(P1_U3257) );
  INV_X1 U10970 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U10971 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9728), .ZN(n9708) );
  OAI21_X1 U10972 ( .B1(n9728), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9708), .ZN(
        n9709) );
  AOI211_X1 U10973 ( .C1(n9710), .C2(n9709), .A(n9727), .B(n10296), .ZN(n9719)
         );
  XNOR2_X1 U10974 ( .A(n9728), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9713) );
  NOR2_X1 U10975 ( .A1(n9714), .A2(n9713), .ZN(n9722) );
  AOI211_X1 U10976 ( .C1(n9714), .C2(n9713), .A(n9722), .B(n10288), .ZN(n9718)
         );
  NAND2_X1 U10977 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9715) );
  OAI21_X1 U10978 ( .B1(n10254), .B2(n9716), .A(n9715), .ZN(n9717) );
  NOR3_X1 U10979 ( .A1(n9719), .A2(n9718), .A3(n9717), .ZN(n9720) );
  OAI21_X1 U10980 ( .B1(n10231), .B2(n9721), .A(n9720), .ZN(P1_U3258) );
  XOR2_X1 U10981 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9740), .Z(n9724) );
  NAND2_X1 U10982 ( .A1(n9724), .A2(n9723), .ZN(n9737) );
  OAI21_X1 U10983 ( .B1(n9724), .B2(n9723), .A(n9737), .ZN(n9734) );
  INV_X1 U10984 ( .A(n9740), .ZN(n9726) );
  OAI21_X1 U10985 ( .B1(n10254), .B2(n9726), .A(n9725), .ZN(n9733) );
  NAND2_X1 U10986 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9740), .ZN(n9729) );
  OAI21_X1 U10987 ( .B1(n9740), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9729), .ZN(
        n9730) );
  AOI211_X1 U10988 ( .C1(n9731), .C2(n9730), .A(n9739), .B(n10296), .ZN(n9732)
         );
  AOI211_X1 U10989 ( .C1(n10302), .C2(n9734), .A(n9733), .B(n9732), .ZN(n9735)
         );
  OAI21_X1 U10990 ( .B1(n10231), .B2(n10496), .A(n9735), .ZN(P1_U3259) );
  INV_X1 U10991 ( .A(n9736), .ZN(n9746) );
  OAI21_X1 U10992 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9740), .A(n9737), .ZN(
        n9738) );
  XOR2_X1 U10993 ( .A(n9738), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9743) );
  INV_X1 U10994 ( .A(n9743), .ZN(n9742) );
  XOR2_X1 U10995 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9741), .Z(n9744) );
  XNOR2_X1 U10996 ( .A(n10046), .B(n9747), .ZN(n9971) );
  NAND2_X1 U10997 ( .A1(n9971), .A2(n10143), .ZN(n9753) );
  INV_X1 U10998 ( .A(n9748), .ZN(n9750) );
  NOR2_X1 U10999 ( .A1(n9750), .A2(n9749), .ZN(n9974) );
  INV_X1 U11000 ( .A(n9974), .ZN(n9751) );
  NOR2_X1 U11001 ( .A1(n10157), .A2(n9751), .ZN(n9756) );
  AOI21_X1 U11002 ( .B1(n10157), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9756), .ZN(
        n9752) );
  OAI211_X1 U11003 ( .C1(n10046), .C2(n10159), .A(n9753), .B(n9752), .ZN(
        P1_U3261) );
  XNOR2_X1 U11004 ( .A(n9755), .B(n9754), .ZN(n9975) );
  NAND2_X1 U11005 ( .A1(n9975), .A2(n10143), .ZN(n9758) );
  AOI21_X1 U11006 ( .B1(n10157), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9756), .ZN(
        n9757) );
  OAI211_X1 U11007 ( .C1(n4860), .C2(n10159), .A(n9758), .B(n9757), .ZN(
        P1_U3262) );
  INV_X1 U11008 ( .A(n9759), .ZN(n9767) );
  NAND2_X1 U11009 ( .A1(n9760), .A2(n9963), .ZN(n9763) );
  AOI22_X1 U11010 ( .A1(n9761), .A2(n10155), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10157), .ZN(n9762) );
  OAI211_X1 U11011 ( .C1(n4739), .C2(n10159), .A(n9763), .B(n9762), .ZN(n9764)
         );
  AOI21_X1 U11012 ( .B1(n9765), .B2(n10161), .A(n9764), .ZN(n9766) );
  OAI21_X1 U11013 ( .B1(n9767), .B2(n9969), .A(n9766), .ZN(P1_U3355) );
  NAND2_X1 U11014 ( .A1(n9768), .A2(n9963), .ZN(n9771) );
  AOI22_X1 U11015 ( .A1(n9769), .A2(n10155), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10157), .ZN(n9770) );
  OAI211_X1 U11016 ( .C1(n9772), .C2(n10159), .A(n9771), .B(n9770), .ZN(n9773)
         );
  AOI21_X1 U11017 ( .B1(n9774), .B2(n10161), .A(n9773), .ZN(n9775) );
  OAI21_X1 U11018 ( .B1(n9776), .B2(n9969), .A(n9775), .ZN(P1_U3263) );
  XNOR2_X1 U11019 ( .A(n9777), .B(n9784), .ZN(n9982) );
  INV_X1 U11020 ( .A(n9800), .ZN(n9780) );
  INV_X1 U11021 ( .A(n9778), .ZN(n9779) );
  AOI211_X1 U11022 ( .C1(n9979), .C2(n9780), .A(n10313), .B(n9779), .ZN(n9978)
         );
  AOI22_X1 U11023 ( .A1(n9781), .A2(n10155), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10157), .ZN(n9782) );
  OAI21_X1 U11024 ( .B1(n9783), .B2(n10159), .A(n9782), .ZN(n9791) );
  AOI21_X1 U11025 ( .B1(n9785), .B2(n9784), .A(n10128), .ZN(n9789) );
  OAI22_X1 U11026 ( .A1(n9786), .A2(n9959), .B1(n9812), .B2(n9957), .ZN(n9787)
         );
  AOI21_X1 U11027 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(n9981) );
  NOR2_X1 U11028 ( .A1(n9981), .A2(n10157), .ZN(n9790) );
  AOI211_X1 U11029 ( .C1(n9963), .C2(n9978), .A(n9791), .B(n9790), .ZN(n9792)
         );
  OAI21_X1 U11030 ( .B1(n9982), .B2(n9969), .A(n9792), .ZN(P1_U3264) );
  XNOR2_X1 U11031 ( .A(n9793), .B(n9797), .ZN(n9985) );
  INV_X1 U11032 ( .A(n9985), .ZN(n9807) );
  NAND2_X1 U11033 ( .A1(n9795), .A2(n9794), .ZN(n9796) );
  XOR2_X1 U11034 ( .A(n9797), .B(n9796), .Z(n9798) );
  OAI222_X1 U11035 ( .A1(n9957), .A2(n9828), .B1(n9959), .B2(n9799), .C1(
        n10128), .C2(n9798), .ZN(n9983) );
  AOI211_X1 U11036 ( .C1(n9801), .C2(n9813), .A(n10313), .B(n9800), .ZN(n9984)
         );
  NAND2_X1 U11037 ( .A1(n9984), .A2(n9963), .ZN(n9804) );
  AOI22_X1 U11038 ( .A1(n9802), .A2(n10155), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10157), .ZN(n9803) );
  OAI211_X1 U11039 ( .C1(n10054), .C2(n10159), .A(n9804), .B(n9803), .ZN(n9805) );
  AOI21_X1 U11040 ( .B1(n9983), .B2(n10161), .A(n9805), .ZN(n9806) );
  OAI21_X1 U11041 ( .B1(n9807), .B2(n9969), .A(n9806), .ZN(P1_U3265) );
  XOR2_X1 U11042 ( .A(n9808), .B(n9809), .Z(n9992) );
  XNOR2_X1 U11043 ( .A(n9810), .B(n9809), .ZN(n9811) );
  OAI222_X1 U11044 ( .A1(n9959), .A2(n9812), .B1(n9957), .B2(n9848), .C1(n9811), .C2(n10128), .ZN(n9988) );
  INV_X1 U11045 ( .A(n9813), .ZN(n9814) );
  AOI211_X1 U11046 ( .C1(n9990), .C2(n9815), .A(n10313), .B(n9814), .ZN(n9989)
         );
  NAND2_X1 U11047 ( .A1(n9989), .A2(n9963), .ZN(n9818) );
  AOI22_X1 U11048 ( .A1(n9816), .A2(n10155), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10157), .ZN(n9817) );
  OAI211_X1 U11049 ( .C1(n9819), .C2(n10159), .A(n9818), .B(n9817), .ZN(n9820)
         );
  AOI21_X1 U11050 ( .B1(n9988), .B2(n10161), .A(n9820), .ZN(n9821) );
  OAI21_X1 U11051 ( .B1(n9992), .B2(n9969), .A(n9821), .ZN(P1_U3266) );
  XOR2_X1 U11052 ( .A(n9822), .B(n9826), .Z(n9995) );
  INV_X1 U11053 ( .A(n9995), .ZN(n9838) );
  INV_X1 U11054 ( .A(n9823), .ZN(n9824) );
  AOI21_X1 U11055 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(n9827) );
  OAI222_X1 U11056 ( .A1(n9957), .A2(n9829), .B1(n9959), .B2(n9828), .C1(
        n10128), .C2(n9827), .ZN(n9993) );
  INV_X1 U11057 ( .A(n9832), .ZN(n10059) );
  AOI211_X1 U11058 ( .C1(n9832), .C2(n9840), .A(n10313), .B(n9831), .ZN(n9994)
         );
  NAND2_X1 U11059 ( .A1(n9994), .A2(n9963), .ZN(n9835) );
  AOI22_X1 U11060 ( .A1(n9833), .A2(n10155), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10157), .ZN(n9834) );
  OAI211_X1 U11061 ( .C1(n10059), .C2(n10159), .A(n9835), .B(n9834), .ZN(n9836) );
  AOI21_X1 U11062 ( .B1(n9993), .B2(n10161), .A(n9836), .ZN(n9837) );
  OAI21_X1 U11063 ( .B1(n9838), .B2(n9969), .A(n9837), .ZN(P1_U3267) );
  XOR2_X1 U11064 ( .A(n9845), .B(n9839), .Z(n10002) );
  AOI21_X1 U11065 ( .B1(n9998), .B2(n9856), .A(n4481), .ZN(n9999) );
  INV_X1 U11066 ( .A(n9998), .ZN(n9844) );
  INV_X1 U11067 ( .A(n9841), .ZN(n9842) );
  AOI22_X1 U11068 ( .A1(n9842), .A2(n10155), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10157), .ZN(n9843) );
  OAI21_X1 U11069 ( .B1(n9844), .B2(n10159), .A(n9843), .ZN(n9853) );
  AOI21_X1 U11070 ( .B1(n9846), .B2(n9845), .A(n10128), .ZN(n9851) );
  OAI22_X1 U11071 ( .A1(n9848), .A2(n9959), .B1(n9847), .B2(n9957), .ZN(n9849)
         );
  AOI21_X1 U11072 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n10001) );
  NOR2_X1 U11073 ( .A1(n10001), .A2(n10157), .ZN(n9852) );
  AOI211_X1 U11074 ( .C1(n9999), .C2(n10143), .A(n9853), .B(n9852), .ZN(n9854)
         );
  OAI21_X1 U11075 ( .B1(n10002), .B2(n9969), .A(n9854), .ZN(P1_U3268) );
  XNOR2_X1 U11076 ( .A(n9855), .B(n9862), .ZN(n10007) );
  INV_X1 U11077 ( .A(n9871), .ZN(n9857) );
  AOI21_X1 U11078 ( .B1(n10003), .B2(n9857), .A(n4732), .ZN(n10004) );
  INV_X1 U11079 ( .A(n9858), .ZN(n9859) );
  AOI22_X1 U11080 ( .A1(n9859), .A2(n10155), .B1(n10157), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9860) );
  OAI21_X1 U11081 ( .B1(n9861), .B2(n10159), .A(n9860), .ZN(n9868) );
  XOR2_X1 U11082 ( .A(n9863), .B(n9862), .Z(n9866) );
  AOI222_X1 U11083 ( .A1(n10152), .A2(n9866), .B1(n9865), .B2(n10149), .C1(
        n9864), .C2(n10147), .ZN(n10006) );
  NOR2_X1 U11084 ( .A1(n10006), .A2(n10157), .ZN(n9867) );
  AOI211_X1 U11085 ( .C1(n10004), .C2(n10143), .A(n9868), .B(n9867), .ZN(n9869) );
  OAI21_X1 U11086 ( .B1(n9969), .B2(n10007), .A(n9869), .ZN(P1_U3269) );
  XNOR2_X1 U11087 ( .A(n9870), .B(n9877), .ZN(n10012) );
  INV_X1 U11088 ( .A(n9894), .ZN(n9872) );
  AOI211_X1 U11089 ( .C1(n10009), .C2(n9872), .A(n10313), .B(n9871), .ZN(
        n10008) );
  INV_X1 U11090 ( .A(n9873), .ZN(n9874) );
  AOI22_X1 U11091 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n10157), .B1(n9874), 
        .B2(n10155), .ZN(n9875) );
  OAI21_X1 U11092 ( .B1(n9876), .B2(n10159), .A(n9875), .ZN(n9886) );
  NAND3_X1 U11093 ( .A1(n9879), .A2(n9878), .A3(n9877), .ZN(n9880) );
  NAND2_X1 U11094 ( .A1(n9881), .A2(n9880), .ZN(n9884) );
  AOI222_X1 U11095 ( .A1(n10152), .A2(n9884), .B1(n9883), .B2(n10149), .C1(
        n9882), .C2(n10147), .ZN(n10011) );
  NOR2_X1 U11096 ( .A1(n10011), .A2(n10157), .ZN(n9885) );
  AOI211_X1 U11097 ( .C1(n10008), .C2(n9963), .A(n9886), .B(n9885), .ZN(n9887)
         );
  OAI21_X1 U11098 ( .B1(n9969), .B2(n10012), .A(n9887), .ZN(P1_U3270) );
  XNOR2_X1 U11099 ( .A(n9888), .B(n9889), .ZN(n10015) );
  INV_X1 U11100 ( .A(n10015), .ZN(n9901) );
  XOR2_X1 U11101 ( .A(n9890), .B(n9889), .Z(n9891) );
  OAI222_X1 U11102 ( .A1(n9957), .A2(n9893), .B1(n9959), .B2(n9892), .C1(n9891), .C2(n10128), .ZN(n10013) );
  AOI211_X1 U11103 ( .C1(n9895), .C2(n9908), .A(n10313), .B(n9894), .ZN(n10014) );
  NAND2_X1 U11104 ( .A1(n10014), .A2(n9963), .ZN(n9898) );
  AOI22_X1 U11105 ( .A1(n10157), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9896), 
        .B2(n10155), .ZN(n9897) );
  OAI211_X1 U11106 ( .C1(n10066), .C2(n10159), .A(n9898), .B(n9897), .ZN(n9899) );
  AOI21_X1 U11107 ( .B1(n10013), .B2(n10161), .A(n9899), .ZN(n9900) );
  OAI21_X1 U11108 ( .B1(n9901), .B2(n9969), .A(n9900), .ZN(P1_U3271) );
  XNOR2_X1 U11109 ( .A(n9902), .B(n9903), .ZN(n10020) );
  INV_X1 U11110 ( .A(n10020), .ZN(n9917) );
  XOR2_X1 U11111 ( .A(n9904), .B(n9903), .Z(n9905) );
  OAI222_X1 U11112 ( .A1(n9959), .A2(n9907), .B1(n9957), .B2(n9906), .C1(n9905), .C2(n10128), .ZN(n10018) );
  INV_X1 U11113 ( .A(n9910), .ZN(n10070) );
  INV_X1 U11114 ( .A(n9908), .ZN(n9909) );
  AOI211_X1 U11115 ( .C1(n9910), .C2(n9922), .A(n10313), .B(n9909), .ZN(n10019) );
  NAND2_X1 U11116 ( .A1(n10019), .A2(n9963), .ZN(n9914) );
  INV_X1 U11117 ( .A(n9911), .ZN(n9912) );
  AOI22_X1 U11118 ( .A1(n10157), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9912), 
        .B2(n10155), .ZN(n9913) );
  OAI211_X1 U11119 ( .C1(n10070), .C2(n10159), .A(n9914), .B(n9913), .ZN(n9915) );
  AOI21_X1 U11120 ( .B1(n10018), .B2(n10161), .A(n9915), .ZN(n9916) );
  OAI21_X1 U11121 ( .B1(n9917), .B2(n9969), .A(n9916), .ZN(P1_U3272) );
  XOR2_X1 U11122 ( .A(n9918), .B(n9931), .Z(n9921) );
  AOI222_X1 U11123 ( .A1(n10152), .A2(n9921), .B1(n9920), .B2(n10149), .C1(
        n9919), .C2(n10147), .ZN(n10028) );
  INV_X1 U11124 ( .A(n9938), .ZN(n9924) );
  INV_X1 U11125 ( .A(n9922), .ZN(n9923) );
  AOI21_X1 U11126 ( .B1(n10025), .B2(n9924), .A(n9923), .ZN(n10026) );
  NOR2_X1 U11127 ( .A1(n9925), .A2(n10159), .ZN(n9930) );
  INV_X1 U11128 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9928) );
  OAI22_X1 U11129 ( .A1(n10161), .A2(n9928), .B1(n9927), .B2(n9926), .ZN(n9929) );
  AOI211_X1 U11130 ( .C1(n10026), .C2(n10143), .A(n9930), .B(n9929), .ZN(n9935) );
  NAND2_X1 U11131 ( .A1(n9932), .A2(n9931), .ZN(n10023) );
  NAND3_X1 U11132 ( .A1(n10024), .A2(n10023), .A3(n9933), .ZN(n9934) );
  OAI211_X1 U11133 ( .C1(n10028), .C2(n10157), .A(n9935), .B(n9934), .ZN(
        P1_U3273) );
  XNOR2_X1 U11134 ( .A(n9937), .B(n9936), .ZN(n10037) );
  AOI21_X1 U11135 ( .B1(n10030), .B2(n4731), .A(n9938), .ZN(n10033) );
  AOI22_X1 U11136 ( .A1(n10157), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9939), 
        .B2(n10155), .ZN(n9940) );
  OAI21_X1 U11137 ( .B1(n9941), .B2(n10159), .A(n9940), .ZN(n9948) );
  XNOR2_X1 U11138 ( .A(n9943), .B(n9942), .ZN(n9946) );
  AOI222_X1 U11139 ( .A1(n10152), .A2(n9946), .B1(n9945), .B2(n10149), .C1(
        n9944), .C2(n10147), .ZN(n10035) );
  NOR2_X1 U11140 ( .A1(n10035), .A2(n10157), .ZN(n9947) );
  AOI211_X1 U11141 ( .C1(n10033), .C2(n10143), .A(n9948), .B(n9947), .ZN(n9949) );
  OAI21_X1 U11142 ( .B1(n9969), .B2(n10037), .A(n9949), .ZN(P1_U3274) );
  XOR2_X1 U11143 ( .A(n9950), .B(n9954), .Z(n10040) );
  INV_X1 U11144 ( .A(n10040), .ZN(n9970) );
  NAND2_X1 U11145 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  XOR2_X1 U11146 ( .A(n9954), .B(n9953), .Z(n9955) );
  OAI222_X1 U11147 ( .A1(n9959), .A2(n9958), .B1(n9957), .B2(n9956), .C1(
        n10128), .C2(n9955), .ZN(n10038) );
  AOI211_X1 U11148 ( .C1(n9962), .C2(n9961), .A(n10313), .B(n9960), .ZN(n10039) );
  NAND2_X1 U11149 ( .A1(n10039), .A2(n9963), .ZN(n9966) );
  AOI22_X1 U11150 ( .A1(n10157), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9964), 
        .B2(n10155), .ZN(n9965) );
  OAI211_X1 U11151 ( .C1(n4729), .C2(n10159), .A(n9966), .B(n9965), .ZN(n9967)
         );
  AOI21_X1 U11152 ( .B1(n10038), .B2(n10161), .A(n9967), .ZN(n9968) );
  OAI21_X1 U11153 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(P1_U3275) );
  INV_X1 U11154 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9972) );
  AOI21_X1 U11155 ( .B1(n9971), .B2(n10032), .A(n9974), .ZN(n10043) );
  MUX2_X1 U11156 ( .A(n9972), .B(n10043), .S(n10344), .Z(n9973) );
  OAI21_X1 U11157 ( .B1(n10046), .B2(n10042), .A(n9973), .ZN(P1_U3554) );
  INV_X1 U11158 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9976) );
  AOI21_X1 U11159 ( .B1(n9975), .B2(n10032), .A(n9974), .ZN(n10047) );
  MUX2_X1 U11160 ( .A(n9976), .B(n10047), .S(n10344), .Z(n9977) );
  OAI21_X1 U11161 ( .B1(n4860), .B2(n10042), .A(n9977), .ZN(P1_U3553) );
  AOI21_X1 U11162 ( .B1(n10031), .B2(n9979), .A(n9978), .ZN(n9980) );
  OAI211_X1 U11163 ( .C1(n9982), .C2(n10036), .A(n9981), .B(n9980), .ZN(n10050) );
  MUX2_X1 U11164 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10050), .S(n10344), .Z(
        P1_U3550) );
  INV_X1 U11165 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9986) );
  AOI211_X1 U11166 ( .C1(n9985), .C2(n10332), .A(n9984), .B(n9983), .ZN(n10051) );
  MUX2_X1 U11167 ( .A(n9986), .B(n10051), .S(n10344), .Z(n9987) );
  OAI21_X1 U11168 ( .B1(n10054), .B2(n10042), .A(n9987), .ZN(P1_U3549) );
  AOI211_X1 U11169 ( .C1(n10031), .C2(n9990), .A(n9989), .B(n9988), .ZN(n9991)
         );
  OAI21_X1 U11170 ( .B1(n9992), .B2(n10036), .A(n9991), .ZN(n10055) );
  MUX2_X1 U11171 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10055), .S(n10344), .Z(
        P1_U3548) );
  INV_X1 U11172 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9996) );
  AOI211_X1 U11173 ( .C1(n9995), .C2(n10332), .A(n9994), .B(n9993), .ZN(n10056) );
  MUX2_X1 U11174 ( .A(n9996), .B(n10056), .S(n10344), .Z(n9997) );
  OAI21_X1 U11175 ( .B1(n10059), .B2(n10042), .A(n9997), .ZN(P1_U3547) );
  AOI22_X1 U11176 ( .A1(n9999), .A2(n10032), .B1(n10031), .B2(n9998), .ZN(
        n10000) );
  OAI211_X1 U11177 ( .C1(n10002), .C2(n10036), .A(n10001), .B(n10000), .ZN(
        n10060) );
  MUX2_X1 U11178 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10060), .S(n10344), .Z(
        P1_U3546) );
  AOI22_X1 U11179 ( .A1(n10004), .A2(n10032), .B1(n10031), .B2(n10003), .ZN(
        n10005) );
  OAI211_X1 U11180 ( .C1(n10007), .C2(n10036), .A(n10006), .B(n10005), .ZN(
        n10061) );
  MUX2_X1 U11181 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10061), .S(n10344), .Z(
        P1_U3545) );
  AOI21_X1 U11182 ( .B1(n10031), .B2(n10009), .A(n10008), .ZN(n10010) );
  OAI211_X1 U11183 ( .C1(n10012), .C2(n10036), .A(n10011), .B(n10010), .ZN(
        n10062) );
  MUX2_X1 U11184 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10062), .S(n10344), .Z(
        P1_U3544) );
  INV_X1 U11185 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10016) );
  AOI211_X1 U11186 ( .C1(n10015), .C2(n10332), .A(n10014), .B(n10013), .ZN(
        n10063) );
  MUX2_X1 U11187 ( .A(n10016), .B(n10063), .S(n10344), .Z(n10017) );
  OAI21_X1 U11188 ( .B1(n10066), .B2(n10042), .A(n10017), .ZN(P1_U3543) );
  AOI211_X1 U11189 ( .C1(n10020), .C2(n10332), .A(n10019), .B(n10018), .ZN(
        n10067) );
  MUX2_X1 U11190 ( .A(n10021), .B(n10067), .S(n10344), .Z(n10022) );
  OAI21_X1 U11191 ( .B1(n10070), .B2(n10042), .A(n10022), .ZN(P1_U3542) );
  NAND3_X1 U11192 ( .A1(n10024), .A2(n10332), .A3(n10023), .ZN(n10029) );
  AOI22_X1 U11193 ( .A1(n10026), .A2(n10032), .B1(n10031), .B2(n10025), .ZN(
        n10027) );
  NAND3_X1 U11194 ( .A1(n10029), .A2(n10028), .A3(n10027), .ZN(n10071) );
  MUX2_X1 U11195 ( .A(n10071), .B(P1_REG1_REG_18__SCAN_IN), .S(n10341), .Z(
        P1_U3541) );
  AOI22_X1 U11196 ( .A1(n10033), .A2(n10032), .B1(n10031), .B2(n10030), .ZN(
        n10034) );
  OAI211_X1 U11197 ( .C1(n10037), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10072) );
  MUX2_X1 U11198 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10072), .S(n10344), .Z(
        P1_U3540) );
  AOI211_X1 U11199 ( .C1(n10040), .C2(n10332), .A(n10039), .B(n10038), .ZN(
        n10073) );
  MUX2_X1 U11200 ( .A(n9696), .B(n10073), .S(n10344), .Z(n10041) );
  OAI21_X1 U11201 ( .B1(n4729), .B2(n10042), .A(n10041), .ZN(P1_U3539) );
  INV_X1 U11202 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10044) );
  MUX2_X1 U11203 ( .A(n10044), .B(n10043), .S(n10336), .Z(n10045) );
  OAI21_X1 U11204 ( .B1(n10046), .B2(n10076), .A(n10045), .ZN(P1_U3522) );
  INV_X1 U11205 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U11206 ( .A(n10048), .B(n10047), .S(n10336), .Z(n10049) );
  OAI21_X1 U11207 ( .B1(n4860), .B2(n10076), .A(n10049), .ZN(P1_U3521) );
  MUX2_X1 U11208 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10050), .S(n10336), .Z(
        P1_U3518) );
  MUX2_X1 U11209 ( .A(n10052), .B(n10051), .S(n10336), .Z(n10053) );
  OAI21_X1 U11210 ( .B1(n10054), .B2(n10076), .A(n10053), .ZN(P1_U3517) );
  MUX2_X1 U11211 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10055), .S(n10336), .Z(
        P1_U3516) );
  MUX2_X1 U11212 ( .A(n10057), .B(n10056), .S(n10336), .Z(n10058) );
  OAI21_X1 U11213 ( .B1(n10059), .B2(n10076), .A(n10058), .ZN(P1_U3515) );
  MUX2_X1 U11214 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10060), .S(n10336), .Z(
        P1_U3514) );
  MUX2_X1 U11215 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10061), .S(n10336), .Z(
        P1_U3513) );
  MUX2_X1 U11216 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10062), .S(n10336), .Z(
        P1_U3512) );
  MUX2_X1 U11217 ( .A(n10064), .B(n10063), .S(n10336), .Z(n10065) );
  OAI21_X1 U11218 ( .B1(n10066), .B2(n10076), .A(n10065), .ZN(P1_U3511) );
  INV_X1 U11219 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10068) );
  MUX2_X1 U11220 ( .A(n10068), .B(n10067), .S(n10336), .Z(n10069) );
  OAI21_X1 U11221 ( .B1(n10070), .B2(n10076), .A(n10069), .ZN(P1_U3510) );
  MUX2_X1 U11222 ( .A(n10071), .B(P1_REG0_REG_18__SCAN_IN), .S(n10334), .Z(
        P1_U3508) );
  MUX2_X1 U11223 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10072), .S(n10336), .Z(
        P1_U3505) );
  INV_X1 U11224 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10074) );
  MUX2_X1 U11225 ( .A(n10074), .B(n10073), .S(n10336), .Z(n10075) );
  OAI21_X1 U11226 ( .B1(n4729), .B2(n10076), .A(n10075), .ZN(P1_U3502) );
  NOR4_X1 U11227 ( .A1(n10077), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n5508), .ZN(n10078) );
  AOI21_X1 U11228 ( .B1(n10079), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10078), 
        .ZN(n10080) );
  OAI21_X1 U11229 ( .B1(n10082), .B2(n10081), .A(n10080), .ZN(P1_U3322) );
  INV_X1 U11230 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10085) );
  OAI222_X1 U11231 ( .A1(n10086), .A2(n10085), .B1(n10090), .B2(n10084), .C1(
        P1_U3084), .C2(n10083), .ZN(P1_U3323) );
  OAI222_X1 U11232 ( .A1(n10090), .A2(n10089), .B1(n5221), .B2(P1_U3084), .C1(
        n10087), .C2(n10100), .ZN(P1_U3324) );
  NAND2_X1 U11233 ( .A1(n10091), .A2(n10095), .ZN(n10093) );
  OAI211_X1 U11234 ( .C1(n10100), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        P1_U3325) );
  NAND2_X1 U11235 ( .A1(n10096), .A2(n10095), .ZN(n10098) );
  OAI211_X1 U11236 ( .C1(n10100), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        P1_U3326) );
  MUX2_X1 U11237 ( .A(n10101), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11238 ( .A(n10102), .ZN(n10318) );
  INV_X1 U11239 ( .A(n10106), .ZN(n10109) );
  OAI211_X1 U11240 ( .C1(n10105), .C2(n10329), .A(n10104), .B(n10103), .ZN(
        n10108) );
  NOR2_X1 U11241 ( .A1(n10106), .A2(n10153), .ZN(n10107) );
  AOI211_X1 U11242 ( .C1(n10318), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10112) );
  INV_X1 U11243 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11244 ( .A1(n10336), .A2(n10112), .B1(n10110), .B2(n10334), .ZN(
        P1_U3484) );
  AOI22_X1 U11245 ( .A1(n10344), .A2(n10112), .B1(n10111), .B2(n10341), .ZN(
        P1_U3533) );
  OAI21_X1 U11246 ( .B1(n4979), .B2(n10434), .A(n10113), .ZN(n10114) );
  AOI21_X1 U11247 ( .B1(n10115), .B2(n10411), .A(n10114), .ZN(n10118) );
  INV_X1 U11248 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11249 ( .A1(n10455), .A2(n10118), .B1(n10116), .B2(n10453), .ZN(
        P2_U3550) );
  INV_X1 U11250 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U11251 ( .A1(n10444), .A2(n10118), .B1(n10117), .B2(n10442), .ZN(
        P2_U3518) );
  XNOR2_X1 U11252 ( .A(n10119), .B(n10124), .ZN(n10174) );
  NOR2_X1 U11253 ( .A1(n10120), .A2(n10171), .ZN(n10121) );
  OR2_X1 U11254 ( .A1(n10122), .A2(n10121), .ZN(n10172) );
  INV_X1 U11255 ( .A(n10172), .ZN(n10123) );
  AOI22_X1 U11256 ( .A1(n10174), .A2(n10144), .B1(n10143), .B2(n10123), .ZN(
        n10137) );
  XNOR2_X1 U11257 ( .A(n10125), .B(n4606), .ZN(n10129) );
  AOI22_X1 U11258 ( .A1(n10147), .A2(n10150), .B1(n10126), .B2(n10149), .ZN(
        n10127) );
  OAI21_X1 U11259 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(n10130) );
  AOI21_X1 U11260 ( .B1(n10174), .B2(n10131), .A(n10130), .ZN(n10176) );
  INV_X1 U11261 ( .A(n10176), .ZN(n10135) );
  AOI22_X1 U11262 ( .A1(n10157), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10132), 
        .B2(n10155), .ZN(n10133) );
  OAI21_X1 U11263 ( .B1(n10171), .B2(n10159), .A(n10133), .ZN(n10134) );
  AOI21_X1 U11264 ( .B1(n10135), .B2(n10161), .A(n10134), .ZN(n10136) );
  NAND2_X1 U11265 ( .A1(n10137), .A2(n10136), .ZN(P1_U3278) );
  XNOR2_X1 U11266 ( .A(n10138), .B(n10145), .ZN(n10154) );
  INV_X1 U11267 ( .A(n10154), .ZN(n10182) );
  OAI21_X1 U11268 ( .B1(n4725), .B2(n4724), .A(n10141), .ZN(n10178) );
  INV_X1 U11269 ( .A(n10178), .ZN(n10142) );
  AOI22_X1 U11270 ( .A1(n10182), .A2(n10144), .B1(n10143), .B2(n10142), .ZN(
        n10164) );
  XNOR2_X1 U11271 ( .A(n10146), .B(n10145), .ZN(n10151) );
  AOI222_X1 U11272 ( .A1(n10152), .A2(n10151), .B1(n10150), .B2(n10149), .C1(
        n10148), .C2(n10147), .ZN(n10179) );
  OAI21_X1 U11273 ( .B1(n10154), .B2(n10153), .A(n10179), .ZN(n10162) );
  AOI22_X1 U11274 ( .A1(n10157), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10156), 
        .B2(n10155), .ZN(n10158) );
  OAI21_X1 U11275 ( .B1(n4724), .B2(n10159), .A(n10158), .ZN(n10160) );
  AOI21_X1 U11276 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(n10163) );
  NAND2_X1 U11277 ( .A1(n10164), .A2(n10163), .ZN(P1_U3280) );
  OAI22_X1 U11278 ( .A1(n10166), .A2(n10313), .B1(n10165), .B2(n10329), .ZN(
        n10168) );
  AOI211_X1 U11279 ( .C1(n10332), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10185) );
  AOI22_X1 U11280 ( .A1(n10344), .A2(n10185), .B1(n10170), .B2(n10341), .ZN(
        P1_U3538) );
  OAI22_X1 U11281 ( .A1(n10172), .A2(n10313), .B1(n10171), .B2(n10329), .ZN(
        n10173) );
  AOI21_X1 U11282 ( .B1(n10174), .B2(n10318), .A(n10173), .ZN(n10175) );
  AND2_X1 U11283 ( .A1(n10176), .A2(n10175), .ZN(n10187) );
  AOI22_X1 U11284 ( .A1(n10344), .A2(n10187), .B1(n10177), .B2(n10341), .ZN(
        P1_U3536) );
  OAI22_X1 U11285 ( .A1(n10178), .A2(n10313), .B1(n4724), .B2(n10329), .ZN(
        n10181) );
  INV_X1 U11286 ( .A(n10179), .ZN(n10180) );
  AOI211_X1 U11287 ( .C1(n10182), .C2(n10332), .A(n10181), .B(n10180), .ZN(
        n10189) );
  AOI22_X1 U11288 ( .A1(n10344), .A2(n10189), .B1(n10183), .B2(n10341), .ZN(
        P1_U3534) );
  INV_X1 U11289 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11290 ( .A1(n10336), .A2(n10185), .B1(n10184), .B2(n10334), .ZN(
        P1_U3499) );
  INV_X1 U11291 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U11292 ( .A1(n10336), .A2(n10187), .B1(n10186), .B2(n10334), .ZN(
        P1_U3493) );
  INV_X1 U11293 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U11294 ( .A1(n10336), .A2(n10189), .B1(n10188), .B2(n10334), .ZN(
        P1_U3487) );
  XOR2_X1 U11295 ( .A(n10190), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11296 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11297 ( .B1(n10192), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10191), .ZN(
        n10197) );
  OAI21_X1 U11298 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n10207), .A(n10208), .ZN(
        n10193) );
  XOR2_X1 U11299 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10193), .Z(n10212) );
  AOI22_X1 U11300 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10306), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10196) );
  NAND3_X1 U11301 ( .A1(n10302), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10194), .ZN(
        n10195) );
  OAI211_X1 U11302 ( .C1(n10197), .C2(n10212), .A(n10196), .B(n10195), .ZN(
        P1_U3241) );
  AOI211_X1 U11303 ( .C1(n10200), .C2(n10199), .A(n10198), .B(n10288), .ZN(
        n10201) );
  AOI21_X1 U11304 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n10201), 
        .ZN(n10217) );
  INV_X1 U11305 ( .A(n10202), .ZN(n10204) );
  NAND2_X1 U11306 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  AND3_X1 U11307 ( .A1(n10206), .A2(n10284), .A3(n10205), .ZN(n10214) );
  NAND2_X1 U11308 ( .A1(n10208), .A2(n10207), .ZN(n10213) );
  NOR2_X1 U11309 ( .A1(n10209), .A2(n10213), .ZN(n10210) );
  AOI211_X1 U11310 ( .C1(n10213), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10225) );
  AOI211_X1 U11311 ( .C1(n10305), .C2(n10215), .A(n10214), .B(n10225), .ZN(
        n10216) );
  OAI211_X1 U11312 ( .C1(n10231), .C2(n10218), .A(n10217), .B(n10216), .ZN(
        P1_U3243) );
  XNOR2_X1 U11313 ( .A(n10220), .B(n10219), .ZN(n10221) );
  AOI22_X1 U11314 ( .A1(n10305), .A2(n10222), .B1(n10284), .B2(n10221), .ZN(
        n10229) );
  XOR2_X1 U11315 ( .A(n10224), .B(n10223), .Z(n10227) );
  AOI211_X1 U11316 ( .C1(n10302), .C2(n10227), .A(n10226), .B(n10225), .ZN(
        n10228) );
  OAI211_X1 U11317 ( .C1(n10231), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        P1_U3245) );
  AND2_X1 U11318 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  OR3_X1 U11319 ( .A1(n10288), .A2(n10235), .A3(n10234), .ZN(n10238) );
  INV_X1 U11320 ( .A(n10236), .ZN(n10237) );
  OAI211_X1 U11321 ( .C1(n10254), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10240) );
  INV_X1 U11322 ( .A(n10240), .ZN(n10246) );
  OAI21_X1 U11323 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10244) );
  AOI22_X1 U11324 ( .A1(n10306), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10284), 
        .B2(n10244), .ZN(n10245) );
  NAND2_X1 U11325 ( .A1(n10246), .A2(n10245), .ZN(P1_U3246) );
  INV_X1 U11326 ( .A(n10247), .ZN(n10248) );
  OAI211_X1 U11327 ( .C1(n10250), .C2(n10249), .A(n10284), .B(n10248), .ZN(
        n10252) );
  OAI211_X1 U11328 ( .C1(n10254), .C2(n10253), .A(n10252), .B(n10251), .ZN(
        n10255) );
  INV_X1 U11329 ( .A(n10255), .ZN(n10260) );
  XNOR2_X1 U11330 ( .A(n10257), .B(n10256), .ZN(n10258) );
  AOI22_X1 U11331 ( .A1(n10306), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n10302), 
        .B2(n10258), .ZN(n10259) );
  NAND2_X1 U11332 ( .A1(n10260), .A2(n10259), .ZN(P1_U3247) );
  OAI21_X1 U11333 ( .B1(n10263), .B2(n10262), .A(n10261), .ZN(n10270) );
  OAI21_X1 U11334 ( .B1(n10266), .B2(n10265), .A(n10264), .ZN(n10267) );
  NAND2_X1 U11335 ( .A1(n10284), .A2(n10267), .ZN(n10269) );
  OAI211_X1 U11336 ( .C1(n10288), .C2(n10270), .A(n10269), .B(n10268), .ZN(
        n10271) );
  INV_X1 U11337 ( .A(n10271), .ZN(n10274) );
  AOI22_X1 U11338 ( .A1(n10306), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n10305), 
        .B2(n10272), .ZN(n10273) );
  NAND2_X1 U11339 ( .A1(n10274), .A2(n10273), .ZN(P1_U3249) );
  OAI21_X1 U11340 ( .B1(n10277), .B2(n10276), .A(n10275), .ZN(n10278) );
  INV_X1 U11341 ( .A(n10278), .ZN(n10287) );
  INV_X1 U11342 ( .A(n10279), .ZN(n10283) );
  NAND2_X1 U11343 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NAND3_X1 U11344 ( .A1(n10284), .A2(n10283), .A3(n10282), .ZN(n10286) );
  OAI211_X1 U11345 ( .C1(n10288), .C2(n10287), .A(n10286), .B(n10285), .ZN(
        n10289) );
  INV_X1 U11346 ( .A(n10289), .ZN(n10292) );
  AOI22_X1 U11347 ( .A1(n10306), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n10305), 
        .B2(n10290), .ZN(n10291) );
  NAND2_X1 U11348 ( .A1(n10292), .A2(n10291), .ZN(P1_U3250) );
  OAI21_X1 U11349 ( .B1(n10295), .B2(n10294), .A(n10293), .ZN(n10303) );
  AOI211_X1 U11350 ( .C1(n10299), .C2(n10298), .A(n10297), .B(n10296), .ZN(
        n10300) );
  AOI211_X1 U11351 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10308) );
  AOI22_X1 U11352 ( .A1(n10306), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n10305), 
        .B2(n10304), .ZN(n10307) );
  NAND2_X1 U11353 ( .A1(n10308), .A2(n10307), .ZN(P1_U3251) );
  AND2_X1 U11354 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10309), .ZN(P1_U3292) );
  AND2_X1 U11355 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10309), .ZN(P1_U3293) );
  AND2_X1 U11356 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10309), .ZN(P1_U3294) );
  AND2_X1 U11357 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10309), .ZN(P1_U3295) );
  AND2_X1 U11358 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10309), .ZN(P1_U3296) );
  AND2_X1 U11359 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10309), .ZN(P1_U3297) );
  AND2_X1 U11360 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10309), .ZN(P1_U3298) );
  AND2_X1 U11361 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10309), .ZN(P1_U3299) );
  AND2_X1 U11362 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10309), .ZN(P1_U3300) );
  AND2_X1 U11363 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10309), .ZN(P1_U3301) );
  AND2_X1 U11364 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10309), .ZN(P1_U3302) );
  AND2_X1 U11365 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10309), .ZN(P1_U3303) );
  AND2_X1 U11366 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10309), .ZN(P1_U3304) );
  AND2_X1 U11367 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10309), .ZN(P1_U3305) );
  AND2_X1 U11368 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10309), .ZN(P1_U3306) );
  AND2_X1 U11369 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10309), .ZN(P1_U3307) );
  AND2_X1 U11370 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10309), .ZN(P1_U3308) );
  AND2_X1 U11371 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10309), .ZN(P1_U3309) );
  AND2_X1 U11372 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10309), .ZN(P1_U3310) );
  AND2_X1 U11373 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10309), .ZN(P1_U3311) );
  AND2_X1 U11374 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10309), .ZN(P1_U3312) );
  AND2_X1 U11375 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10309), .ZN(P1_U3313) );
  AND2_X1 U11376 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10309), .ZN(P1_U3314) );
  AND2_X1 U11377 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10309), .ZN(P1_U3315) );
  AND2_X1 U11378 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10309), .ZN(P1_U3316) );
  AND2_X1 U11379 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10309), .ZN(P1_U3317) );
  AND2_X1 U11380 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10309), .ZN(P1_U3318) );
  AND2_X1 U11381 ( .A1(n10309), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U11382 ( .A1(n10309), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3320) );
  NOR2_X1 U11383 ( .A1(n10311), .A2(n10310), .ZN(P1_U3321) );
  OAI22_X1 U11384 ( .A1(n10314), .A2(n10313), .B1(n10312), .B2(n10329), .ZN(
        n10316) );
  AOI211_X1 U11385 ( .C1(n10318), .C2(n10317), .A(n10316), .B(n10315), .ZN(
        n10338) );
  INV_X1 U11386 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U11387 ( .A1(n10336), .A2(n10338), .B1(n10319), .B2(n10334), .ZN(
        P1_U3463) );
  OAI21_X1 U11388 ( .B1(n10321), .B2(n10329), .A(n10320), .ZN(n10322) );
  AOI21_X1 U11389 ( .B1(n10323), .B2(n10332), .A(n10322), .ZN(n10324) );
  AND2_X1 U11390 ( .A1(n10325), .A2(n10324), .ZN(n10340) );
  INV_X1 U11391 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U11392 ( .A1(n10336), .A2(n10340), .B1(n10326), .B2(n10334), .ZN(
        P1_U3469) );
  OAI211_X1 U11393 ( .C1(n10330), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10331) );
  AOI21_X1 U11394 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(n10343) );
  INV_X1 U11395 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U11396 ( .A1(n10336), .A2(n10343), .B1(n10335), .B2(n10334), .ZN(
        P1_U3481) );
  INV_X1 U11397 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U11398 ( .A1(n10344), .A2(n10338), .B1(n10337), .B2(n10341), .ZN(
        P1_U3526) );
  INV_X1 U11399 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U11400 ( .A1(n10344), .A2(n10340), .B1(n10339), .B2(n10341), .ZN(
        P1_U3528) );
  INV_X1 U11401 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U11402 ( .A1(n10344), .A2(n10343), .B1(n10342), .B2(n10341), .ZN(
        P1_U3532) );
  NAND2_X1 U11403 ( .A1(n10349), .A2(n10345), .ZN(n10346) );
  NAND2_X1 U11404 ( .A1(n10346), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10348) );
  AOI211_X1 U11405 ( .C1(n10350), .C2(n6158), .A(n10348), .B(n10347), .ZN(
        n10354) );
  AOI22_X1 U11406 ( .A1(n10350), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10349), .ZN(n10353) );
  AOI22_X1 U11407 ( .A1(n10351), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10352) );
  OAI221_X1 U11408 ( .B1(n10354), .B2(n10353), .C1(n10354), .C2(n5034), .A(
        n10352), .ZN(P2_U3245) );
  XNOR2_X1 U11409 ( .A(n10356), .B(n10355), .ZN(n10408) );
  AOI22_X1 U11410 ( .A1(n10408), .A2(n10358), .B1(P2_REG2_REG_5__SCAN_IN), 
        .B2(n10357), .ZN(n10374) );
  OAI21_X1 U11411 ( .B1(n10359), .B2(n4557), .A(n7117), .ZN(n10364) );
  AOI222_X1 U11412 ( .A1(n10365), .A2(n10364), .B1(n10363), .B2(n10362), .C1(
        n10361), .C2(n10360), .ZN(n10405) );
  INV_X1 U11413 ( .A(n10405), .ZN(n10372) );
  OAI211_X1 U11414 ( .C1(n10367), .C2(n10406), .A(n10366), .B(n10411), .ZN(
        n10404) );
  OAI22_X1 U11415 ( .A1(n10404), .A2(n10369), .B1(n10406), .B2(n10368), .ZN(
        n10371) );
  OAI21_X1 U11416 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(n10373) );
  OAI211_X1 U11417 ( .C1(n10376), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        P2_U3291) );
  INV_X1 U11418 ( .A(n10377), .ZN(n10379) );
  AND2_X1 U11419 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10383), .ZN(P2_U3297) );
  AND2_X1 U11420 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10383), .ZN(P2_U3298) );
  AND2_X1 U11421 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10383), .ZN(P2_U3299) );
  AND2_X1 U11422 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10383), .ZN(P2_U3300) );
  AND2_X1 U11423 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10383), .ZN(P2_U3301) );
  AND2_X1 U11424 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10383), .ZN(P2_U3302) );
  AND2_X1 U11425 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10383), .ZN(P2_U3303) );
  AND2_X1 U11426 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10383), .ZN(P2_U3304) );
  AND2_X1 U11427 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10383), .ZN(P2_U3305) );
  AND2_X1 U11428 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10383), .ZN(P2_U3306) );
  AND2_X1 U11429 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10383), .ZN(P2_U3307) );
  AND2_X1 U11430 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10383), .ZN(P2_U3308) );
  AND2_X1 U11431 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10383), .ZN(P2_U3309) );
  AND2_X1 U11432 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10383), .ZN(P2_U3310) );
  AND2_X1 U11433 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10383), .ZN(P2_U3311) );
  AND2_X1 U11434 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10383), .ZN(P2_U3312) );
  AND2_X1 U11435 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10383), .ZN(P2_U3313) );
  AND2_X1 U11436 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10383), .ZN(P2_U3314) );
  AND2_X1 U11437 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10383), .ZN(P2_U3315) );
  AND2_X1 U11438 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10383), .ZN(P2_U3316) );
  AND2_X1 U11439 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10383), .ZN(P2_U3317) );
  AND2_X1 U11440 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10383), .ZN(P2_U3318) );
  AND2_X1 U11441 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10383), .ZN(P2_U3319) );
  AND2_X1 U11442 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10383), .ZN(P2_U3320) );
  AND2_X1 U11443 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10383), .ZN(P2_U3321) );
  AND2_X1 U11444 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10383), .ZN(P2_U3322) );
  AND2_X1 U11445 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10383), .ZN(P2_U3323) );
  AND2_X1 U11446 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10383), .ZN(P2_U3324) );
  AND2_X1 U11447 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10383), .ZN(P2_U3325) );
  AND2_X1 U11448 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10383), .ZN(P2_U3326) );
  INV_X1 U11449 ( .A(n10380), .ZN(n10385) );
  AOI22_X1 U11450 ( .A1(n10382), .A2(n10383), .B1(n10381), .B2(n10385), .ZN(
        P2_U3437) );
  AOI22_X1 U11451 ( .A1(n10386), .A2(n10385), .B1(n10384), .B2(n10383), .ZN(
        P2_U3438) );
  AOI22_X1 U11452 ( .A1(n10388), .A2(n10440), .B1(n6119), .B2(n10387), .ZN(
        n10389) );
  AND2_X1 U11453 ( .A1(n10390), .A2(n10389), .ZN(n10445) );
  INV_X1 U11454 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U11455 ( .A1(n10444), .A2(n10445), .B1(n10391), .B2(n10442), .ZN(
        P2_U3451) );
  OAI21_X1 U11456 ( .B1(n10393), .B2(n10434), .A(n10392), .ZN(n10395) );
  AOI211_X1 U11457 ( .C1(n10396), .C2(n10440), .A(n10395), .B(n10394), .ZN(
        n10447) );
  INV_X1 U11458 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U11459 ( .A1(n10444), .A2(n10447), .B1(n10397), .B2(n10442), .ZN(
        P2_U3457) );
  OAI22_X1 U11460 ( .A1(n10399), .A2(n10436), .B1(n10398), .B2(n10434), .ZN(
        n10401) );
  AOI211_X1 U11461 ( .C1(n10440), .C2(n10402), .A(n10401), .B(n10400), .ZN(
        n10448) );
  INV_X1 U11462 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U11463 ( .A1(n10444), .A2(n10448), .B1(n10403), .B2(n10442), .ZN(
        P2_U3463) );
  OAI211_X1 U11464 ( .C1(n10406), .C2(n10434), .A(n10405), .B(n10404), .ZN(
        n10407) );
  AOI21_X1 U11465 ( .B1(n10440), .B2(n10408), .A(n10407), .ZN(n10449) );
  INV_X1 U11466 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U11467 ( .A1(n10444), .A2(n10449), .B1(n10409), .B2(n10442), .ZN(
        P2_U3466) );
  AOI22_X1 U11468 ( .A1(n10412), .A2(n10411), .B1(n9437), .B2(n10410), .ZN(
        n10413) );
  OAI211_X1 U11469 ( .C1(n10415), .C2(n10426), .A(n10414), .B(n10413), .ZN(
        n10416) );
  INV_X1 U11470 ( .A(n10416), .ZN(n10450) );
  INV_X1 U11471 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U11472 ( .A1(n10444), .A2(n10450), .B1(n10417), .B2(n10442), .ZN(
        P2_U3469) );
  INV_X1 U11473 ( .A(n10418), .ZN(n10424) );
  OAI22_X1 U11474 ( .A1(n10420), .A2(n10436), .B1(n10419), .B2(n10434), .ZN(
        n10422) );
  AOI211_X1 U11475 ( .C1(n10424), .C2(n10423), .A(n10422), .B(n10421), .ZN(
        n10451) );
  INV_X1 U11476 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U11477 ( .A1(n10444), .A2(n10451), .B1(n10425), .B2(n10442), .ZN(
        P2_U3475) );
  OR2_X1 U11478 ( .A1(n10427), .A2(n10426), .ZN(n10432) );
  OAI22_X1 U11479 ( .A1(n10428), .A2(n10436), .B1(n4989), .B2(n10434), .ZN(
        n10429) );
  NOR2_X1 U11480 ( .A1(n10430), .A2(n10429), .ZN(n10431) );
  INV_X1 U11481 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U11482 ( .A1(n10444), .A2(n10452), .B1(n10433), .B2(n10442), .ZN(
        P2_U3481) );
  OAI22_X1 U11483 ( .A1(n10437), .A2(n10436), .B1(n10435), .B2(n10434), .ZN(
        n10439) );
  AOI211_X1 U11484 ( .C1(n10441), .C2(n10440), .A(n10439), .B(n10438), .ZN(
        n10454) );
  INV_X1 U11485 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U11486 ( .A1(n10444), .A2(n10454), .B1(n10443), .B2(n10442), .ZN(
        P2_U3487) );
  AOI22_X1 U11487 ( .A1(n10455), .A2(n10445), .B1(n10345), .B2(n10453), .ZN(
        P2_U3520) );
  INV_X1 U11488 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U11489 ( .A1(n10455), .A2(n10447), .B1(n10446), .B2(n10453), .ZN(
        P2_U3522) );
  AOI22_X1 U11490 ( .A1(n10455), .A2(n10448), .B1(n6209), .B2(n10453), .ZN(
        P2_U3524) );
  AOI22_X1 U11491 ( .A1(n10455), .A2(n10449), .B1(n6221), .B2(n10453), .ZN(
        P2_U3525) );
  AOI22_X1 U11492 ( .A1(n10455), .A2(n10450), .B1(n6249), .B2(n10453), .ZN(
        P2_U3526) );
  AOI22_X1 U11493 ( .A1(n10455), .A2(n10451), .B1(n6659), .B2(n10453), .ZN(
        P2_U3528) );
  AOI22_X1 U11494 ( .A1(n10455), .A2(n10452), .B1(n6855), .B2(n10453), .ZN(
        P2_U3530) );
  AOI22_X1 U11495 ( .A1(n10455), .A2(n10454), .B1(n7277), .B2(n10453), .ZN(
        P2_U3532) );
  INV_X1 U11496 ( .A(n10456), .ZN(n10457) );
  NAND2_X1 U11497 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  XOR2_X1 U11498 ( .A(n10460), .B(n10459), .Z(ADD_1071_U5) );
  XOR2_X1 U11499 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11500 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(ADD_1071_U56) );
  OAI21_X1 U11501 ( .B1(n10466), .B2(n10465), .A(n10464), .ZN(ADD_1071_U57) );
  OAI21_X1 U11502 ( .B1(n10469), .B2(n10468), .A(n10467), .ZN(ADD_1071_U58) );
  OAI21_X1 U11503 ( .B1(n10472), .B2(n10471), .A(n10470), .ZN(ADD_1071_U59) );
  OAI21_X1 U11504 ( .B1(n10475), .B2(n10474), .A(n10473), .ZN(ADD_1071_U60) );
  OAI21_X1 U11505 ( .B1(n10478), .B2(n10477), .A(n10476), .ZN(ADD_1071_U61) );
  AOI21_X1 U11506 ( .B1(n10481), .B2(n10480), .A(n10479), .ZN(ADD_1071_U62) );
  AOI21_X1 U11507 ( .B1(n10484), .B2(n10483), .A(n10482), .ZN(ADD_1071_U63) );
  AOI21_X1 U11508 ( .B1(n10487), .B2(n10486), .A(n10485), .ZN(ADD_1071_U47) );
  XOR2_X1 U11509 ( .A(n10488), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11510 ( .A(n10490), .B(n10489), .Z(ADD_1071_U54) );
  NOR2_X1 U11511 ( .A1(n10492), .A2(n10491), .ZN(n10493) );
  XOR2_X1 U11512 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10493), .Z(ADD_1071_U51) );
  OAI21_X1 U11513 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(n10497) );
  XNOR2_X1 U11514 ( .A(n10497), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11515 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10498), .Z(ADD_1071_U48) );
  XOR2_X1 U11516 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10499), .Z(ADD_1071_U50) );
  XOR2_X1 U11517 ( .A(n10501), .B(n10500), .Z(ADD_1071_U53) );
  XNOR2_X1 U11518 ( .A(n10503), .B(n10502), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U5022 ( .A(n6461), .Z(n4903) );
  CLKBUF_X1 U5643 ( .A(n6304), .Z(n8626) );
  CLKBUF_X1 U6150 ( .A(n7442), .Z(n8141) );
endmodule

