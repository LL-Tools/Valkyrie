

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606;

  INV_X1 U2246 ( .A(n2319), .ZN(n2651) );
  CLKBUF_X1 U2247 ( .A(n4606), .Z(U4043) );
  NOR2_X1 U2248 ( .A1(n2306), .A2(n4388), .ZN(n4606) );
  CLKBUF_X1 U2249 ( .A(n3611), .Z(n2005) );
  NOR2_X1 U2250 ( .A1(n2766), .A2(n4381), .ZN(n3611) );
  INV_X1 U2251 ( .A(n2698), .ZN(n2584) );
  NAND2_X2 U2252 ( .A1(n2755), .A2(n2829), .ZN(n2701) );
  INV_X1 U2253 ( .A(n2300), .ZN(n2353) );
  NAND2_X1 U2254 ( .A1(n4091), .A2(n2814), .ZN(n4068) );
  MUX2_X1 U2255 ( .A(REG1_REG_28__SCAN_IN), .B(n2878), .S(n4453), .Z(n2870) );
  MUX2_X1 U2256 ( .A(REG0_REG_28__SCAN_IN), .B(n2878), .S(n4443), .Z(n2879) );
  AND2_X1 U2257 ( .A1(n2995), .A2(n3779), .ZN(n4440) );
  CLKBUF_X3 U2258 ( .A(n2353), .Z(n2007) );
  OAI21_X2 U2259 ( .B1(n3974), .B2(n2823), .A(n2822), .ZN(n3954) );
  AOI21_X2 U2260 ( .B1(n3507), .B2(n2600), .A(n2599), .ZN(n3524) );
  OAI21_X4 U2261 ( .B1(n2553), .B2(n2156), .A(n2154), .ZN(n3507) );
  AND2_X1 U2262 ( .A1(n2097), .A2(n2047), .ZN(n2553) );
  NAND4_X1 U2263 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .ZN(n3149)
         );
  INV_X4 U2264 ( .A(n2701), .ZN(n2716) );
  INV_X2 U2265 ( .A(n4265), .ZN(n2264) );
  INV_X1 U2266 ( .A(IR_REG_31__SCAN_IN), .ZN(n2759) );
  AND2_X1 U2267 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2254)
         );
  AOI21_X1 U2268 ( .B1(n3938), .B2(n3773), .A(n3701), .ZN(n3922) );
  NAND2_X1 U2269 ( .A1(n2455), .A2(n2165), .ZN(n3370) );
  NAND2_X1 U2270 ( .A1(n2060), .A2(n3749), .ZN(n3645) );
  NAND2_X1 U2271 ( .A1(n3278), .A2(n2206), .ZN(n2204) );
  AND2_X1 U2272 ( .A1(n3041), .A2(n2785), .ZN(n3054) );
  AND2_X1 U2273 ( .A1(n3725), .A2(n3722), .ZN(n3697) );
  NAND2_X1 U2274 ( .A1(n3720), .A2(n3723), .ZN(n2832) );
  NAND2_X1 U2275 ( .A1(n2323), .A2(n2020), .ZN(n3158) );
  INV_X1 U2276 ( .A(n2348), .ZN(n2635) );
  AND2_X2 U2277 ( .A1(n2891), .A2(n4129), .ZN(n4063) );
  NAND2_X1 U2278 ( .A1(n2357), .A2(n2240), .ZN(n3804) );
  AND4_X1 U2279 ( .A1(n2407), .A2(n2406), .A3(n2405), .A4(n2404), .ZN(n3256)
         );
  NOR2_X2 U2280 ( .A1(n2945), .A2(n2944), .ZN(n4345) );
  INV_X1 U2281 ( .A(n4440), .ZN(n4430) );
  AND2_X1 U2282 ( .A1(n3047), .A2(n3109), .ZN(n3064) );
  INV_X2 U2283 ( .A(n2262), .ZN(n2006) );
  INV_X1 U2284 ( .A(n2892), .ZN(n2829) );
  AND2_X1 U2285 ( .A1(n3779), .A2(n4268), .ZN(n2892) );
  INV_X1 U2286 ( .A(n3670), .ZN(n4268) );
  XNOR2_X1 U2287 ( .A(n2280), .B(n2279), .ZN(n3779) );
  AOI21_X1 U2288 ( .B1(n2932), .B2(IR_REG_28__SCAN_IN), .A(n2038), .ZN(n2130)
         );
  OR2_X1 U2289 ( .A1(n2932), .A2(IR_REG_27__SCAN_IN), .ZN(n2131) );
  AND2_X1 U2290 ( .A1(n2292), .A2(n2291), .ZN(n4267) );
  CLKBUF_X2 U2291 ( .A(n2281), .Z(n2932) );
  NOR2_X2 U2292 ( .A1(n2270), .A2(n2258), .ZN(n2761) );
  AND2_X1 U2293 ( .A1(n2560), .A2(n2249), .ZN(n2563) );
  AND2_X1 U2294 ( .A1(n2252), .A2(n2231), .ZN(n2230) );
  NOR2_X1 U2295 ( .A1(n2250), .A2(IR_REG_18__SCAN_IN), .ZN(n2183) );
  NAND2_X1 U2296 ( .A1(n2324), .A2(n2244), .ZN(n2326) );
  AND4_X1 U2297 ( .A1(n2241), .A2(n2243), .A3(n2242), .A4(n2378), .ZN(n2061)
         );
  NOR2_X1 U2298 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2241)
         );
  NOR2_X1 U2299 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2243)
         );
  NOR2_X1 U2300 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2242)
         );
  NOR3_X1 U2301 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .A3(
        IR_REG_24__SCAN_IN), .ZN(n2252) );
  INV_X1 U2302 ( .A(IR_REG_5__SCAN_IN), .ZN(n2378) );
  NOR2_X2 U2303 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2324)
         );
  INV_X1 U2304 ( .A(IR_REG_2__SCAN_IN), .ZN(n2244) );
  INV_X1 U2305 ( .A(IR_REG_22__SCAN_IN), .ZN(n4507) );
  INV_X1 U2306 ( .A(IR_REG_19__SCAN_IN), .ZN(n2293) );
  INV_X1 U2307 ( .A(IR_REG_17__SCAN_IN), .ZN(n2249) );
  INV_X1 U2308 ( .A(IR_REG_20__SCAN_IN), .ZN(n2279) );
  OAI22_X2 U2309 ( .A1(n3178), .A2(n2794), .B1(n3179), .B2(n3802), .ZN(n3232)
         );
  NOR2_X2 U2310 ( .A1(n3280), .A2(n3279), .ZN(n2137) );
  NOR2_X2 U2311 ( .A1(n3081), .A2(n3082), .ZN(n3199) );
  OR2_X2 U2312 ( .A1(n3467), .A2(n2264), .ZN(n2319) );
  NOR3_X2 U2313 ( .A1(n3450), .A2(n3551), .A3(n2127), .ZN(n2129) );
  OR2_X2 U2314 ( .A1(n3408), .A2(n3403), .ZN(n3450) );
  INV_X1 U2315 ( .A(n2262), .ZN(n2008) );
  AND2_X4 U2316 ( .A1(n3467), .A2(n2264), .ZN(n2340) );
  XNOR2_X2 U2317 ( .A(n2255), .B(IR_REG_29__SCAN_IN), .ZN(n3467) );
  NAND2_X1 U2318 ( .A1(n3294), .A2(n3295), .ZN(n2455) );
  AND2_X1 U2319 ( .A1(n2028), .A2(n2801), .ZN(n2206) );
  OR2_X1 U2320 ( .A1(n4079), .A2(n4059), .ZN(n3675) );
  NAND2_X1 U2321 ( .A1(n2204), .A2(n2202), .ZN(n3332) );
  AND2_X1 U2322 ( .A1(n2205), .A2(n2203), .ZN(n2202) );
  INV_X1 U2323 ( .A(n3683), .ZN(n2203) );
  NAND2_X1 U2324 ( .A1(n2229), .A2(IR_REG_31__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2325 ( .A1(n3521), .A2(n2179), .ZN(n2178) );
  XNOR2_X1 U2326 ( .A(n2347), .B(n2701), .ZN(n2349) );
  NAND2_X1 U2327 ( .A1(n3805), .A2(n2698), .ZN(n2310) );
  NAND2_X1 U2328 ( .A1(n3486), .A2(n3487), .ZN(n2097) );
  AOI22_X1 U2329 ( .A1(n3804), .A2(n2698), .B1(n2713), .B2(n2790), .ZN(n2361)
         );
  NAND2_X1 U2330 ( .A1(n2151), .A2(n3204), .ZN(n2150) );
  INV_X1 U2331 ( .A(n3522), .ZN(n2180) );
  XNOR2_X1 U2332 ( .A(n2331), .B(n2716), .ZN(n2336) );
  AND2_X1 U2333 ( .A1(n2698), .A2(n2756), .ZN(n3786) );
  XNOR2_X1 U2334 ( .A(n4275), .B(REG1_REG_2__SCAN_IN), .ZN(n3825) );
  OAI21_X1 U2335 ( .B1(n3006), .B2(n3005), .A(n3008), .ZN(n3009) );
  AOI21_X1 U2336 ( .B1(n3095), .B2(REG1_REG_9__SCAN_IN), .A(n3094), .ZN(n3096)
         );
  OR2_X1 U2337 ( .A1(n3102), .A2(n3101), .ZN(n2139) );
  NAND2_X1 U2338 ( .A1(n2139), .A2(n2105), .ZN(n2104) );
  NOR2_X1 U2339 ( .A1(n2106), .A2(n3873), .ZN(n2105) );
  INV_X1 U2340 ( .A(n2138), .ZN(n2106) );
  AOI21_X1 U2341 ( .B1(n2139), .B2(n2138), .A(n4398), .ZN(n2108) );
  NAND2_X1 U2342 ( .A1(n2043), .A2(n4341), .ZN(n2111) );
  NAND2_X1 U2343 ( .A1(n4366), .A2(n2055), .ZN(n3868) );
  OR2_X1 U2344 ( .A1(n3881), .A2(REG2_REG_17__SCAN_IN), .ZN(n2055) );
  AND2_X1 U2345 ( .A1(n2215), .A2(n2014), .ZN(n2214) );
  NAND2_X1 U2346 ( .A1(n2021), .A2(n2216), .ZN(n2215) );
  NOR2_X1 U2347 ( .A1(n2828), .A2(n2224), .ZN(n2223) );
  NOR2_X1 U2348 ( .A1(n3793), .A2(n3941), .ZN(n2224) );
  AND2_X1 U2349 ( .A1(n3794), .A2(n2871), .ZN(n2811) );
  NAND2_X1 U2350 ( .A1(n3491), .A2(n3423), .ZN(n2806) );
  INV_X1 U2351 ( .A(n3397), .ZN(n2201) );
  NAND2_X1 U2352 ( .A1(n2306), .A2(n2740), .ZN(n2928) );
  INV_X1 U2353 ( .A(n4388), .ZN(n2740) );
  NOR2_X2 U2354 ( .A1(n2010), .A2(n3918), .ZN(n4146) );
  NOR2_X1 U2355 ( .A1(n3984), .A2(n2125), .ZN(n3946) );
  NOR2_X1 U2356 ( .A1(n3984), .A2(n3961), .ZN(n3965) );
  OR2_X1 U2357 ( .A1(n4289), .A2(n4266), .ZN(n4375) );
  INV_X1 U2358 ( .A(n3621), .ZN(n2164) );
  INV_X1 U2359 ( .A(n2552), .ZN(n2163) );
  NAND2_X1 U2360 ( .A1(n3872), .A2(REG1_REG_11__SCAN_IN), .ZN(n2138) );
  INV_X1 U2361 ( .A(n3860), .ZN(n2052) );
  OR2_X1 U2362 ( .A1(n4346), .A2(n2058), .ZN(n2057) );
  AND2_X1 U2363 ( .A1(n4394), .A2(REG2_REG_15__SCAN_IN), .ZN(n2058) );
  NOR2_X1 U2364 ( .A1(n2826), .A2(n2227), .ZN(n2226) );
  INV_X1 U2365 ( .A(n2824), .ZN(n2227) );
  NOR2_X1 U2366 ( .A1(n3652), .A2(n2073), .ZN(n2072) );
  INV_X1 U2367 ( .A(n4126), .ZN(n2871) );
  INV_X1 U2368 ( .A(n2806), .ZN(n2199) );
  NAND2_X1 U2369 ( .A1(n3333), .A2(n3747), .ZN(n2060) );
  AOI21_X1 U2370 ( .B1(n2206), .B2(n2802), .A(n2022), .ZN(n2205) );
  OAI21_X1 U2371 ( .B1(n2795), .B2(n2187), .A(n2798), .ZN(n2186) );
  AND2_X1 U2372 ( .A1(n4267), .A2(n4268), .ZN(n2930) );
  OR2_X1 U2373 ( .A1(n3158), .A2(n3116), .ZN(n3720) );
  OR2_X1 U2374 ( .A1(n2845), .A2(n3489), .ZN(n2128) );
  INV_X1 U2375 ( .A(n3423), .ZN(n3403) );
  INV_X1 U2376 ( .A(n3733), .ZN(n2795) );
  INV_X1 U2377 ( .A(n4267), .ZN(n2764) );
  OR2_X2 U2378 ( .A1(n2290), .A2(n2759), .ZN(n2739) );
  NAND2_X1 U2379 ( .A1(n2279), .A2(n2293), .ZN(n2250) );
  INV_X1 U2380 ( .A(IR_REG_14__SCAN_IN), .ZN(n2245) );
  NOR2_X1 U2381 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2248)
         );
  NOR2_X1 U2382 ( .A1(n3372), .A2(n2166), .ZN(n2165) );
  INV_X1 U2383 ( .A(n2454), .ZN(n2166) );
  OR2_X1 U2384 ( .A1(n2549), .A2(n2548), .ZN(n2554) );
  INV_X1 U2385 ( .A(n2413), .ZN(n2090) );
  NOR2_X1 U2386 ( .A1(n2586), .A2(n3515), .ZN(n2601) );
  OR2_X1 U2387 ( .A1(n2487), .A2(n2486), .ZN(n2501) );
  OR2_X1 U2388 ( .A1(n3582), .A2(n2178), .ZN(n2177) );
  NAND2_X1 U2389 ( .A1(n2698), .A2(n2286), .ZN(n2298) );
  AOI21_X1 U2390 ( .B1(n2015), .B2(n2155), .A(n2044), .ZN(n2154) );
  NAND2_X1 U2391 ( .A1(n2158), .A2(n2157), .ZN(n2156) );
  INV_X1 U2392 ( .A(n3560), .ZN(n2155) );
  NAND2_X1 U2393 ( .A1(n2935), .A2(n2102), .ZN(n2951) );
  NAND2_X1 U2394 ( .A1(n3825), .A2(n3824), .ZN(n2102) );
  NOR2_X1 U2395 ( .A1(n2445), .A2(IR_REG_10__SCAN_IN), .ZN(n2506) );
  NOR2_X1 U2396 ( .A1(n2103), .A2(n2108), .ZN(n4304) );
  NAND2_X1 U2397 ( .A1(n2140), .A2(n4393), .ZN(n2113) );
  OR2_X1 U2398 ( .A1(n4341), .A2(n2546), .ZN(n2112) );
  INV_X1 U2399 ( .A(n2140), .ZN(n2114) );
  XNOR2_X1 U2400 ( .A(n2057), .B(n4393), .ZN(n4357) );
  NAND2_X1 U2401 ( .A1(n2228), .A2(n2226), .ZN(n2225) );
  NAND2_X1 U2402 ( .A1(n3924), .A2(n4101), .ZN(n2082) );
  OR2_X1 U2403 ( .A1(n2630), .A2(n3593), .ZN(n2638) );
  OAI21_X1 U2404 ( .B1(n2848), .B2(n2071), .A(n2069), .ZN(n4031) );
  AOI21_X1 U2405 ( .B1(n3758), .B2(n2070), .A(n2036), .ZN(n2069) );
  INV_X1 U2406 ( .A(n3758), .ZN(n2071) );
  INV_X1 U2407 ( .A(n2072), .ZN(n2070) );
  INV_X1 U2408 ( .A(n2192), .ZN(n2191) );
  OAI21_X1 U2409 ( .B1(n2816), .B2(n2193), .A(n3675), .ZN(n2192) );
  NAND2_X1 U2410 ( .A1(n4068), .A2(n2815), .ZN(n2194) );
  NAND2_X1 U2411 ( .A1(n2807), .A2(n2845), .ZN(n2808) );
  NAND2_X1 U2412 ( .A1(n3422), .A2(n3324), .ZN(n2804) );
  AND2_X1 U2413 ( .A1(n3805), .A2(n3040), .ZN(n3042) );
  NAND2_X1 U2414 ( .A1(n3946), .A2(n3928), .ZN(n3927) );
  OR2_X1 U2415 ( .A1(n4004), .A2(n2872), .ZN(n3984) );
  NAND2_X1 U2416 ( .A1(n4014), .A2(n4005), .ZN(n4004) );
  INV_X1 U2417 ( .A(n4422), .ZN(n4428) );
  AND2_X1 U2418 ( .A1(n2723), .A2(n2918), .ZN(n2916) );
  INV_X1 U2419 ( .A(n2928), .ZN(n3030) );
  NAND2_X1 U2420 ( .A1(n2260), .A2(IR_REG_31__SCAN_IN), .ZN(n2068) );
  NOR2_X1 U2421 ( .A1(n2259), .A2(n2759), .ZN(n2065) );
  NAND2_X1 U2422 ( .A1(IR_REG_30__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2064) );
  INV_X1 U2423 ( .A(IR_REG_28__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U2424 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2253) );
  NAND2_X1 U2425 ( .A1(n2563), .A2(n4463), .ZN(n2278) );
  NOR2_X1 U2426 ( .A1(n2720), .A2(n2182), .ZN(n2181) );
  AND2_X1 U2427 ( .A1(n2504), .A2(n2503), .ZN(n3491) );
  INV_X1 U2428 ( .A(n2167), .ZN(n2098) );
  NAND2_X1 U2429 ( .A1(n3386), .A2(n2170), .ZN(n2099) );
  OAI21_X1 U2430 ( .B1(n2011), .B2(n2169), .A(n2168), .ZN(n2167) );
  AND2_X1 U2431 ( .A1(n2648), .A2(n2174), .ZN(n2173) );
  INV_X1 U2432 ( .A(n3582), .ZN(n2092) );
  NAND2_X1 U2433 ( .A1(n2175), .A2(n2178), .ZN(n2174) );
  NOR2_X1 U2434 ( .A1(n2016), .A2(n3606), .ZN(n2093) );
  AND4_X1 U2435 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), .ZN(n3389)
         );
  NAND2_X1 U2436 ( .A1(n3146), .A2(n2365), .ZN(n3131) );
  OR2_X1 U2437 ( .A1(n2774), .A2(n2763), .ZN(n3625) );
  OAI21_X1 U2438 ( .B1(n3930), .B2(n2300), .A(n2697), .ZN(n3942) );
  NAND2_X1 U2439 ( .A1(n2685), .A2(n2684), .ZN(n3793) );
  INV_X1 U2440 ( .A(n3491), .ZN(n3796) );
  MUX2_X1 U2441 ( .A(n2939), .B(REG2_REG_2__SCAN_IN), .S(n4275), .Z(n3830) );
  AND2_X1 U2442 ( .A1(n2122), .A2(n2120), .ZN(n3094) );
  NAND2_X1 U2443 ( .A1(n2121), .A2(n4544), .ZN(n2122) );
  NAND2_X1 U2444 ( .A1(n3011), .A2(n2119), .ZN(n2118) );
  OAI21_X1 U2445 ( .B1(n4375), .B2(n3885), .A(n2145), .ZN(n2144) );
  AOI21_X1 U2446 ( .B1(n4345), .B2(ADDR_REG_18__SCAN_IN), .A(n3884), .ZN(n2145) );
  XNOR2_X1 U2447 ( .A(n2053), .B(n3891), .ZN(n3896) );
  NOR2_X1 U2448 ( .A1(n3890), .A2(n2054), .ZN(n2053) );
  AND2_X1 U2449 ( .A1(n4270), .A2(REG2_REG_18__SCAN_IN), .ZN(n2054) );
  INV_X1 U2450 ( .A(n2213), .ZN(n3916) );
  NAND2_X1 U2451 ( .A1(n2021), .A2(n2218), .ZN(n2217) );
  INV_X1 U2452 ( .A(IR_REG_29__SCAN_IN), .ZN(n2259) );
  AND2_X1 U2453 ( .A1(n3668), .A2(n3975), .ZN(n3762) );
  INV_X1 U2454 ( .A(IR_REG_21__SCAN_IN), .ZN(n2251) );
  NOR2_X1 U2455 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2246)
         );
  NOR2_X1 U2456 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2247)
         );
  INV_X1 U2457 ( .A(n3205), .ZN(n2152) );
  NOR2_X1 U2458 ( .A1(n3548), .A2(n3560), .ZN(n2157) );
  INV_X1 U2459 ( .A(n2162), .ZN(n2158) );
  OR2_X1 U2460 ( .A1(n4314), .A2(n3875), .ZN(n3877) );
  NAND2_X1 U2461 ( .A1(n3913), .A2(n2221), .ZN(n2220) );
  INV_X1 U2462 ( .A(n2827), .ZN(n2221) );
  AND2_X1 U2463 ( .A1(n3793), .A2(n3948), .ZN(n3701) );
  AND2_X1 U2464 ( .A1(n4047), .A2(n2853), .ZN(n3758) );
  AND2_X1 U2465 ( .A1(n2815), .A2(n3674), .ZN(n2190) );
  NAND2_X1 U2466 ( .A1(n4102), .A2(n4078), .ZN(n2815) );
  NAND2_X1 U2467 ( .A1(n4053), .A2(n4083), .ZN(n2816) );
  NAND2_X1 U2468 ( .A1(n4105), .A2(n4126), .ZN(n2812) );
  INV_X1 U2469 ( .A(n2237), .ZN(n2195) );
  NAND2_X1 U2470 ( .A1(n3645), .A2(n3706), .ZN(n3444) );
  AND2_X1 U2471 ( .A1(n3734), .A2(n2079), .ZN(n2078) );
  NAND2_X1 U2472 ( .A1(n2834), .A2(n3730), .ZN(n2079) );
  INV_X1 U2473 ( .A(n3728), .ZN(n2075) );
  INV_X1 U2474 ( .A(n2791), .ZN(n2212) );
  INV_X1 U2475 ( .A(n2786), .ZN(n2209) );
  NAND2_X1 U2476 ( .A1(n3967), .A2(n3948), .ZN(n2125) );
  AND2_X1 U2477 ( .A1(n2183), .A2(n2249), .ZN(n2135) );
  INV_X1 U2478 ( .A(n2326), .ZN(n2062) );
  NAND2_X1 U2479 ( .A1(n2171), .A2(n3419), .ZN(n2168) );
  NAND2_X1 U2480 ( .A1(n2172), .A2(n3418), .ZN(n2171) );
  NAND2_X1 U2481 ( .A1(n3383), .A2(n3382), .ZN(n2172) );
  INV_X1 U2482 ( .A(n3383), .ZN(n2169) );
  NAND2_X1 U2483 ( .A1(n2041), .A2(n2011), .ZN(n2170) );
  AND2_X1 U2484 ( .A1(n3498), .A2(n3499), .ZN(n2648) );
  INV_X1 U2485 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3515) );
  INV_X1 U2486 ( .A(n2873), .ZN(n3912) );
  NOR2_X1 U2487 ( .A1(n2164), .A2(n2163), .ZN(n2162) );
  NOR2_X1 U2488 ( .A1(n3548), .A2(n2161), .ZN(n2160) );
  NAND2_X1 U2489 ( .A1(n2164), .A2(n2163), .ZN(n2161) );
  AOI21_X1 U2490 ( .B1(n3496), .B2(n2662), .A(n2661), .ZN(n3571) );
  INV_X1 U2491 ( .A(n2713), .ZN(n2659) );
  NOR2_X1 U2492 ( .A1(n2649), .A2(n3574), .ZN(n2663) );
  OR2_X1 U2493 ( .A1(n2435), .A2(n2432), .ZN(n2456) );
  AND2_X1 U2494 ( .A1(n3642), .A2(DATAI_22_), .ZN(n4015) );
  INV_X1 U2495 ( .A(n2553), .ZN(n2159) );
  XNOR2_X1 U2496 ( .A(n2965), .B(n2948), .ZN(n2964) );
  NOR2_X1 U2497 ( .A1(n3013), .A2(n3021), .ZN(n2119) );
  NAND2_X1 U2498 ( .A1(n3011), .A2(n3010), .ZN(n2121) );
  NOR2_X1 U2499 ( .A1(n3003), .A2(n3002), .ZN(n3086) );
  INV_X1 U2500 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4495) );
  OR2_X1 U2501 ( .A1(n3086), .A2(n2056), .ZN(n3088) );
  NOR2_X1 U2502 ( .A1(n3087), .A2(n3283), .ZN(n2056) );
  NOR2_X1 U2503 ( .A1(n4304), .A2(n3874), .ZN(n4316) );
  NAND2_X1 U2504 ( .A1(n2049), .A2(n3861), .ZN(n3863) );
  AOI21_X1 U2505 ( .B1(n3860), .B2(n2051), .A(n2046), .ZN(n2050) );
  AND2_X1 U2506 ( .A1(n3863), .A2(n4334), .ZN(n3864) );
  AND2_X1 U2507 ( .A1(n3642), .A2(n2931), .ZN(n2944) );
  AND2_X1 U2508 ( .A1(n4394), .A2(REG1_REG_15__SCAN_IN), .ZN(n2140) );
  INV_X1 U2509 ( .A(n2057), .ZN(n3866) );
  NOR2_X1 U2510 ( .A1(n3868), .A2(n3869), .ZN(n3890) );
  INV_X1 U2511 ( .A(n2825), .ZN(n2218) );
  NOR2_X1 U2512 ( .A1(n2692), .A2(n4496), .ZN(n2704) );
  OR2_X1 U2513 ( .A1(n2678), .A2(n3612), .ZN(n2692) );
  AND2_X1 U2514 ( .A1(n3955), .A2(n3668), .ZN(n3978) );
  OR2_X1 U2515 ( .A1(n2638), .A2(n3500), .ZN(n2649) );
  AND2_X1 U2516 ( .A1(n3996), .A2(n3995), .ZN(n4021) );
  AND3_X1 U2517 ( .A1(n2634), .A2(n2633), .A3(n2632), .ZN(n4030) );
  NAND2_X1 U2518 ( .A1(n2848), .A2(n2072), .ZN(n4048) );
  NAND2_X1 U2519 ( .A1(n4118), .A2(n2813), .ZN(n2814) );
  OR2_X1 U2520 ( .A1(n2128), .A2(n2871), .ZN(n2127) );
  OR2_X1 U2521 ( .A1(n2574), .A2(n2573), .ZN(n2586) );
  NAND2_X1 U2522 ( .A1(n2848), .A2(n3751), .ZN(n4116) );
  NAND2_X1 U2523 ( .A1(n2810), .A2(n2012), .ZN(n2882) );
  NAND2_X1 U2524 ( .A1(n3555), .A2(n3627), .ZN(n2809) );
  AND2_X1 U2525 ( .A1(n2526), .A2(n2525), .ZN(n2535) );
  AOI21_X1 U2526 ( .B1(n2009), .B2(n2199), .A(n2039), .ZN(n2198) );
  AND4_X1 U2527 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n3563)
         );
  NAND2_X1 U2528 ( .A1(n2473), .A2(REG3_REG_11__SCAN_IN), .ZN(n2487) );
  NOR2_X1 U2529 ( .A1(n2456), .A2(n4495), .ZN(n2473) );
  NAND2_X1 U2530 ( .A1(n2838), .A2(n3743), .ZN(n3333) );
  NAND2_X1 U2531 ( .A1(n2204), .A2(n2205), .ZN(n3330) );
  OAI21_X1 U2532 ( .B1(n3273), .B2(n3744), .A(n3741), .ZN(n3303) );
  INV_X1 U2533 ( .A(n2186), .ZN(n2185) );
  NAND2_X1 U2534 ( .A1(n2084), .A2(n3736), .ZN(n3273) );
  NAND2_X1 U2535 ( .A1(n3238), .A2(n3740), .ZN(n2084) );
  INV_X1 U2536 ( .A(n4101), .ZN(n4117) );
  INV_X1 U2537 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2401) );
  AND2_X1 U2538 ( .A1(n2836), .A2(n3737), .ZN(n3733) );
  OAI21_X1 U2539 ( .B1(n3191), .B2(n2077), .A(n2074), .ZN(n3173) );
  AOI21_X1 U2540 ( .B1(n2078), .B2(n2076), .A(n2075), .ZN(n2074) );
  INV_X1 U2541 ( .A(n2078), .ZN(n2077) );
  INV_X1 U2542 ( .A(n3730), .ZN(n2076) );
  INV_X1 U2543 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2366) );
  NOR2_X1 U2544 ( .A1(n2367), .A2(n2366), .ZN(n2388) );
  INV_X1 U2545 ( .A(n4147), .ZN(n4099) );
  INV_X1 U2546 ( .A(n3804), .ZN(n3164) );
  INV_X1 U2547 ( .A(n3132), .ZN(n3169) );
  INV_X1 U2548 ( .A(n2790), .ZN(n3198) );
  INV_X1 U2549 ( .A(n4121), .ZN(n4104) );
  NOR2_X1 U2550 ( .A1(n4038), .A2(n4015), .ZN(n4014) );
  NAND2_X1 U2551 ( .A1(n3642), .A2(DATAI_23_), .ZN(n4005) );
  NAND2_X1 U2552 ( .A1(n2134), .A2(n4039), .ZN(n4038) );
  AND2_X1 U2553 ( .A1(n3642), .A2(DATAI_20_), .ZN(n4059) );
  NOR2_X1 U2554 ( .A1(n4125), .A2(n4100), .ZN(n4094) );
  NAND2_X1 U2555 ( .A1(n4094), .A2(n4083), .ZN(n4082) );
  NOR2_X1 U2556 ( .A1(n3450), .A2(n2128), .ZN(n3436) );
  NOR2_X1 U2557 ( .A1(n3450), .A2(n3489), .ZN(n3451) );
  NOR2_X1 U2558 ( .A1(n3342), .A2(n3343), .ZN(n3341) );
  NAND2_X1 U2559 ( .A1(n3341), .A2(n3324), .ZN(n3408) );
  NAND2_X1 U2560 ( .A1(n2137), .A2(n2136), .ZN(n3342) );
  AND2_X1 U2561 ( .A1(n3229), .A2(n3265), .ZN(n3244) );
  NAND2_X1 U2562 ( .A1(n3244), .A2(n3243), .ZN(n3280) );
  OR2_X1 U2563 ( .A1(n3197), .A2(n3169), .ZN(n3180) );
  NOR2_X1 U2564 ( .A1(n3180), .A2(n3179), .ZN(n3229) );
  AND2_X1 U2565 ( .A1(n4057), .A2(n4435), .ZN(n4422) );
  AND2_X1 U2566 ( .A1(n2565), .A2(n2564), .ZN(n3881) );
  OR2_X1 U2567 ( .A1(n2508), .A2(IR_REG_13__SCAN_IN), .ZN(n2532) );
  INV_X1 U2568 ( .A(IR_REG_3__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U2569 ( .A1(n2326), .A2(IR_REG_31__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U2570 ( .A1(n2282), .A2(n2141), .ZN(n2936) );
  AOI22_X1 U2571 ( .A1(n2027), .A2(n4401), .B1(n2142), .B2(n2759), .ZN(n2141)
         );
  INV_X1 U2572 ( .A(IR_REG_1__SCAN_IN), .ZN(n2142) );
  NAND2_X1 U2573 ( .A1(n2091), .A2(n2413), .ZN(n3252) );
  NAND2_X1 U2574 ( .A1(n3262), .A2(n3261), .ZN(n2091) );
  NAND2_X1 U2575 ( .A1(n2485), .A2(n2484), .ZN(n3386) );
  INV_X1 U2576 ( .A(n4001), .ZN(n3541) );
  NOR2_X1 U2577 ( .A1(n2153), .A2(n2015), .ZN(n3562) );
  NOR3_X1 U2578 ( .A1(n2553), .A2(n2162), .A3(n3548), .ZN(n2153) );
  NAND2_X1 U2579 ( .A1(n3642), .A2(DATAI_24_), .ZN(n3985) );
  NOR2_X1 U2580 ( .A1(n3145), .A2(n2101), .ZN(n2100) );
  INV_X1 U2581 ( .A(n2352), .ZN(n2101) );
  AOI21_X1 U2582 ( .B1(n2088), .B2(n2087), .A(n2045), .ZN(n2086) );
  INV_X1 U2583 ( .A(n3261), .ZN(n2087) );
  INV_X1 U2584 ( .A(DATAI_0_), .ZN(n2132) );
  INV_X1 U2585 ( .A(n3511), .ZN(n2598) );
  AND2_X1 U2586 ( .A1(n2177), .A2(n2180), .ZN(n3589) );
  INV_X1 U2587 ( .A(n3343), .ZN(n3358) );
  OR2_X1 U2588 ( .A1(n2774), .A2(n2773), .ZN(n3613) );
  OAI21_X1 U2589 ( .B1(n3536), .B2(n3537), .A(n3538), .ZN(n3609) );
  INV_X1 U2590 ( .A(n3613), .ZN(n3629) );
  INV_X1 U2591 ( .A(n3618), .ZN(n3623) );
  OR2_X1 U2592 ( .A1(n3473), .A2(n2300), .ZN(n2712) );
  NAND2_X1 U2593 ( .A1(n2670), .A2(n2669), .ZN(n3981) );
  INV_X1 U2594 ( .A(n4030), .ZN(n3529) );
  NAND4_X1 U2595 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(n4079)
         );
  INV_X1 U2596 ( .A(n3563), .ZN(n4120) );
  INV_X1 U2597 ( .A(n3256), .ZN(n3801) );
  OR2_X1 U2598 ( .A1(n2319), .A2(n2339), .ZN(n2343) );
  NAND2_X1 U2599 ( .A1(n2353), .A2(REG3_REG_2__SCAN_IN), .ZN(n2323) );
  NAND2_X1 U2600 ( .A1(n2006), .A2(REG0_REG_1__SCAN_IN), .ZN(n2268) );
  OR2_X1 U2601 ( .A1(n2319), .A2(n2301), .ZN(n2302) );
  INV_X1 U2602 ( .A(U4043), .ZN(n3819) );
  XNOR2_X1 U2603 ( .A(n2936), .B(REG1_REG_1__SCAN_IN), .ZN(n3810) );
  XNOR2_X1 U2604 ( .A(n2951), .B(n2948), .ZN(n2950) );
  NAND2_X1 U2605 ( .A1(n2960), .A2(n2959), .ZN(n3006) );
  XNOR2_X1 U2606 ( .A(n3009), .B(n3021), .ZN(n3023) );
  NOR2_X1 U2607 ( .A1(n3023), .A2(n4544), .ZN(n3022) );
  NOR2_X1 U2608 ( .A1(n3022), .A2(n2123), .ZN(n3014) );
  INV_X1 U2609 ( .A(n2121), .ZN(n2123) );
  XNOR2_X1 U2610 ( .A(n3088), .B(n4303), .ZN(n4300) );
  NOR2_X1 U2611 ( .A1(n4294), .A2(n3097), .ZN(n3102) );
  INV_X1 U2612 ( .A(n2139), .ZN(n3871) );
  NAND2_X1 U2613 ( .A1(n4311), .A2(REG2_REG_12__SCAN_IN), .ZN(n4310) );
  NAND2_X1 U2614 ( .A1(n2107), .A2(n2104), .ZN(n4305) );
  INV_X1 U2615 ( .A(n2108), .ZN(n2107) );
  NAND2_X1 U2616 ( .A1(n4310), .A2(n3860), .ZN(n4320) );
  INV_X1 U2617 ( .A(n4394), .ZN(n4352) );
  NAND2_X1 U2618 ( .A1(n2024), .A2(n2109), .ZN(n4355) );
  NAND2_X1 U2619 ( .A1(n2111), .A2(n2113), .ZN(n2110) );
  NAND2_X1 U2620 ( .A1(n4355), .A2(n4547), .ZN(n4354) );
  NAND2_X1 U2621 ( .A1(n4363), .A2(n2117), .ZN(n3882) );
  OR2_X1 U2622 ( .A1(n3881), .A2(REG1_REG_17__SCAN_IN), .ZN(n2117) );
  NAND2_X1 U2623 ( .A1(n2116), .A2(n2115), .ZN(n2147) );
  INV_X1 U2624 ( .A(n3883), .ZN(n2115) );
  INV_X1 U2625 ( .A(n3882), .ZN(n2116) );
  INV_X1 U2626 ( .A(n4325), .ZN(n4370) );
  AND2_X1 U2627 ( .A1(n2147), .A2(n3886), .ZN(n3889) );
  NAND2_X1 U2628 ( .A1(n2219), .A2(n2827), .ZN(n3914) );
  NAND2_X1 U2629 ( .A1(n2225), .A2(n2223), .ZN(n2219) );
  NAND2_X1 U2630 ( .A1(n2225), .A2(n2222), .ZN(n3925) );
  INV_X1 U2631 ( .A(n2224), .ZN(n2222) );
  AOI21_X1 U2632 ( .B1(n2083), .B2(n4107), .A(n2080), .ZN(n4159) );
  NAND2_X1 U2633 ( .A1(n2082), .A2(n2081), .ZN(n2080) );
  XNOR2_X1 U2634 ( .A(n3922), .B(n3926), .ZN(n2083) );
  INV_X1 U2635 ( .A(n3923), .ZN(n2081) );
  AND2_X1 U2636 ( .A1(n2200), .A2(n2034), .ZN(n3443) );
  NAND2_X1 U2637 ( .A1(n2200), .A2(n2009), .ZN(n3441) );
  NAND2_X1 U2638 ( .A1(n2201), .A2(n2806), .ZN(n2200) );
  AND2_X1 U2639 ( .A1(n4278), .A2(n2893), .ZN(n4037) );
  INV_X1 U2640 ( .A(n4037), .ZN(n4135) );
  INV_X1 U2641 ( .A(n4282), .ZN(n4127) );
  NAND2_X1 U2642 ( .A1(n3030), .A2(n2765), .ZN(n4129) );
  AND2_X1 U2643 ( .A1(n4278), .A2(n3073), .ZN(n4383) );
  INV_X1 U2644 ( .A(n4129), .ZN(n4381) );
  INV_X2 U2645 ( .A(n4451), .ZN(n4453) );
  AOI21_X1 U2646 ( .B1(n4440), .B2(n4155), .A(n4154), .ZN(n4156) );
  OAI21_X1 U2647 ( .B1(n2874), .B2(n2873), .A(n2010), .ZN(n3471) );
  OAI21_X1 U2648 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n4229) );
  NAND2_X1 U2649 ( .A1(n4443), .A2(n4440), .ZN(n4263) );
  INV_X2 U2650 ( .A(n4441), .ZN(n4443) );
  OAI21_X1 U2651 ( .B1(n2065), .B2(IR_REG_30__SCAN_IN), .A(n2064), .ZN(n2063)
         );
  NAND2_X1 U2652 ( .A1(n2761), .A2(n2025), .ZN(n2066) );
  NOR2_X1 U2653 ( .A1(n2762), .A2(n2761), .ZN(n4266) );
  NAND2_X1 U2654 ( .A1(n2737), .A2(IR_REG_31__SCAN_IN), .ZN(n2269) );
  NAND2_X1 U2655 ( .A1(n2296), .A2(n2295), .ZN(n3894) );
  NOR2_X1 U2656 ( .A1(n2582), .A2(n2581), .ZN(n4270) );
  AND2_X1 U2657 ( .A1(n2482), .A2(n2493), .ZN(n3872) );
  NAND2_X1 U2658 ( .A1(n2327), .A2(n2326), .ZN(n4275) );
  OAI22_X1 U2659 ( .A1(n2324), .A2(n2124), .B1(IR_REG_31__SCAN_IN), .B2(
        IR_REG_2__SCAN_IN), .ZN(n2325) );
  NAND2_X1 U2660 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2124)
         );
  CLKBUF_X1 U2661 ( .A(IR_REG_0__SCAN_IN), .Z(n4401) );
  NAND2_X1 U2662 ( .A1(n2096), .A2(n2782), .ZN(n2095) );
  NAND2_X1 U2663 ( .A1(n2146), .A2(n2143), .ZN(U3258) );
  NAND2_X1 U2664 ( .A1(n2148), .A2(n2147), .ZN(n2146) );
  NOR2_X1 U2665 ( .A1(n2023), .A2(n2144), .ZN(n2143) );
  AOI21_X1 U2666 ( .B1(n3882), .B2(n3883), .A(n4339), .ZN(n2148) );
  AOI22_X1 U2667 ( .A1(n4283), .A2(n4282), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4063), .ZN(n4284) );
  NAND2_X1 U2668 ( .A1(n2761), .A2(n2259), .ZN(n2913) );
  AND2_X1 U2669 ( .A1(n2034), .A2(n3442), .ZN(n2009) );
  OR3_X1 U2670 ( .A1(n3984), .A2(n2125), .A3(n2048), .ZN(n2010) );
  NOR2_X1 U2671 ( .A1(n2159), .A2(n2163), .ZN(n3547) );
  NAND2_X1 U2672 ( .A1(n3382), .A2(n2514), .ZN(n2011) );
  AND2_X1 U2673 ( .A1(n2196), .A2(n2809), .ZN(n2012) );
  AND2_X1 U2674 ( .A1(n2012), .A2(n2812), .ZN(n2013) );
  AND2_X1 U2675 ( .A1(n2220), .A2(n2037), .ZN(n2014) );
  INV_X1 U2676 ( .A(n2089), .ZN(n2088) );
  OR2_X1 U2677 ( .A1(n3250), .A2(n2090), .ZN(n2089) );
  OR2_X1 U2678 ( .A1(n2160), .A2(n2555), .ZN(n2015) );
  INV_X1 U2679 ( .A(n3365), .ZN(n2136) );
  XOR2_X1 U2680 ( .A(n2746), .B(n2744), .Z(n2016) );
  OR2_X1 U2681 ( .A1(n2748), .A2(n3618), .ZN(n2017) );
  XNOR2_X1 U2682 ( .A(n2545), .B(n2544), .ZN(n4393) );
  INV_X1 U2683 ( .A(n3967), .ZN(n3961) );
  OR2_X1 U2684 ( .A1(n2553), .A2(n2552), .ZN(n2018) );
  NAND2_X1 U2685 ( .A1(n2274), .A2(n2251), .ZN(n2019) );
  AND3_X1 U2686 ( .A1(n2322), .A2(n2321), .A3(n2320), .ZN(n2020) );
  AND2_X1 U2687 ( .A1(n3315), .A2(n3317), .ZN(n3683) );
  AND2_X1 U2688 ( .A1(n3913), .A2(n2223), .ZN(n2021) );
  AOI21_X1 U2689 ( .B1(n3569), .B2(n3572), .A(n3571), .ZN(n3536) );
  OAI21_X1 U2690 ( .B1(n2583), .B2(n2285), .A(n2284), .ZN(n3047) );
  AND2_X1 U2691 ( .A1(n3798), .A2(n3365), .ZN(n2022) );
  AND2_X1 U2692 ( .A1(n4370), .A2(n3870), .ZN(n2023) );
  OR2_X1 U2693 ( .A1(n4342), .A2(n2112), .ZN(n2024) );
  INV_X1 U2694 ( .A(n2796), .ZN(n2187) );
  AND2_X1 U2695 ( .A1(IR_REG_30__SCAN_IN), .A2(n2259), .ZN(n2025) );
  AND2_X1 U2696 ( .A1(n2251), .A2(n4507), .ZN(n2231) );
  AND4_X1 U2697 ( .A1(n2248), .A2(n2247), .A3(n2246), .A4(n2245), .ZN(n2026)
         );
  INV_X1 U2698 ( .A(n2059), .ZN(n2377) );
  NOR2_X1 U2699 ( .A1(n2326), .A2(n2375), .ZN(n2059) );
  AND2_X1 U2700 ( .A1(n2560), .A2(n2135), .ZN(n2274) );
  INV_X1 U2701 ( .A(IR_REG_18__SCAN_IN), .ZN(n4463) );
  AND2_X1 U2702 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2027)
         );
  NAND2_X1 U2703 ( .A1(n2177), .A2(n2175), .ZN(n3497) );
  OR2_X1 U2704 ( .A1(n3798), .A2(n3365), .ZN(n2028) );
  INV_X1 U2705 ( .A(IR_REG_30__SCAN_IN), .ZN(n2260) );
  NOR2_X1 U2706 ( .A1(n3582), .A2(n3525), .ZN(n2029) );
  AND2_X1 U2707 ( .A1(n2139), .A2(n2138), .ZN(n2030) );
  AND2_X1 U2708 ( .A1(n2387), .A2(n2152), .ZN(n2031) );
  AND2_X1 U2709 ( .A1(n2230), .A2(n2256), .ZN(n2032) );
  AND2_X1 U2710 ( .A1(n2183), .A2(n2231), .ZN(n2033) );
  NAND2_X1 U2711 ( .A1(n2062), .A2(n2061), .ZN(n2445) );
  INV_X1 U2712 ( .A(n3551), .ZN(n2898) );
  XNOR2_X1 U2713 ( .A(n2269), .B(IR_REG_24__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U2714 ( .A1(n2189), .A2(n2191), .ZN(n4035) );
  OAI21_X1 U2715 ( .B1(n3386), .B2(n3383), .A(n3382), .ZN(n3417) );
  AND2_X1 U2716 ( .A1(n2099), .A2(n2098), .ZN(n3486) );
  NAND2_X1 U2717 ( .A1(n2194), .A2(n2816), .ZN(n4046) );
  NAND2_X1 U2718 ( .A1(n3796), .A2(n3403), .ZN(n2034) );
  INV_X1 U2719 ( .A(n3751), .ZN(n2073) );
  AND2_X1 U2720 ( .A1(n2882), .A2(n2237), .ZN(n2035) );
  NAND2_X1 U2721 ( .A1(n2455), .A2(n2454), .ZN(n3369) );
  AND2_X1 U2722 ( .A1(n4079), .A2(n3584), .ZN(n2036) );
  NAND2_X1 U2723 ( .A1(n2810), .A2(n2809), .ZN(n2881) );
  INV_X1 U2724 ( .A(n2134), .ZN(n4061) );
  NOR2_X1 U2725 ( .A1(n4082), .A2(n4059), .ZN(n2134) );
  NAND2_X1 U2726 ( .A1(n3924), .A2(n3912), .ZN(n2037) );
  INV_X1 U2727 ( .A(n3626), .ZN(n3795) );
  AND4_X1 U2728 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n3626)
         );
  INV_X1 U2729 ( .A(n3555), .ZN(n2807) );
  AND4_X1 U2730 ( .A1(n2531), .A2(n2530), .A3(n2529), .A4(n2528), .ZN(n3555)
         );
  INV_X1 U2731 ( .A(n2176), .ZN(n2175) );
  NAND2_X1 U2732 ( .A1(n3590), .A2(n2180), .ZN(n2176) );
  AND2_X1 U2733 ( .A1(n2758), .A2(IR_REG_27__SCAN_IN), .ZN(n2038) );
  AND2_X1 U2734 ( .A1(n3626), .A2(n3453), .ZN(n2039) );
  AND2_X1 U2735 ( .A1(n2812), .A2(n2195), .ZN(n2040) );
  NAND2_X1 U2736 ( .A1(n3419), .A2(n3382), .ZN(n2041) );
  INV_X1 U2737 ( .A(n3674), .ZN(n2193) );
  AND2_X1 U2738 ( .A1(n2235), .A2(n2778), .ZN(n2042) );
  INV_X1 U2739 ( .A(n3525), .ZN(n2179) );
  XNOR2_X1 U2740 ( .A(n2271), .B(IR_REG_26__SCAN_IN), .ZN(n2918) );
  INV_X1 U2741 ( .A(n2918), .ZN(n2182) );
  INV_X1 U2742 ( .A(n3873), .ZN(n4398) );
  NAND2_X1 U2743 ( .A1(n2188), .A2(n2795), .ZN(n3231) );
  OAI21_X1 U2744 ( .B1(n3278), .B2(n2802), .A(n2801), .ZN(n3307) );
  NAND2_X1 U2745 ( .A1(n3053), .A2(n2786), .ZN(n3071) );
  NAND2_X1 U2746 ( .A1(n3187), .A2(n2791), .ZN(n3161) );
  NAND2_X1 U2747 ( .A1(n3231), .A2(n2796), .ZN(n3242) );
  AND2_X1 U2748 ( .A1(n3644), .A2(n3751), .ZN(n3693) );
  INV_X1 U2749 ( .A(n3693), .ZN(n2196) );
  AND2_X1 U2750 ( .A1(n2114), .A2(n2546), .ZN(n2043) );
  INV_X1 U2751 ( .A(n4303), .ZN(n4399) );
  AND2_X1 U2752 ( .A1(n2570), .A2(n2569), .ZN(n2044) );
  AND3_X1 U2753 ( .A1(n2062), .A2(n2061), .A3(n2026), .ZN(n2560) );
  NAND2_X1 U2754 ( .A1(n3054), .A2(n2832), .ZN(n3053) );
  AND2_X1 U2755 ( .A1(n2431), .A2(n2430), .ZN(n2045) );
  NAND2_X1 U2756 ( .A1(n2149), .A2(n2352), .ZN(n3144) );
  INV_X1 U2757 ( .A(n2126), .ZN(n4202) );
  NOR3_X1 U2758 ( .A1(n3450), .A2(n3551), .A3(n2128), .ZN(n2126) );
  NAND2_X1 U2759 ( .A1(n2789), .A2(n3189), .ZN(n3187) );
  INV_X1 U2760 ( .A(n2137), .ZN(n3308) );
  AND2_X1 U2761 ( .A1(n3411), .A2(n4324), .ZN(n2046) );
  INV_X1 U2762 ( .A(n4107), .ZN(n4123) );
  NAND2_X1 U2763 ( .A1(n2859), .A2(n3634), .ZN(n4107) );
  NAND2_X1 U2764 ( .A1(n3642), .A2(DATAI_27_), .ZN(n3928) );
  INV_X1 U2765 ( .A(n3928), .ZN(n3767) );
  NAND3_X1 U2766 ( .A1(n2302), .A2(n2303), .A3(n2085), .ZN(n3805) );
  NAND2_X1 U2767 ( .A1(n3642), .A2(DATAI_26_), .ZN(n3948) );
  NAND2_X1 U2768 ( .A1(n2524), .A2(n2523), .ZN(n2047) );
  OR2_X1 U2769 ( .A1(n3912), .A2(n3767), .ZN(n2048) );
  INV_X1 U2770 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2051) );
  INV_X1 U2771 ( .A(n2720), .ZN(n2921) );
  XNOR2_X1 U2772 ( .A(n2273), .B(IR_REG_25__SCAN_IN), .ZN(n2720) );
  INV_X1 U2773 ( .A(n4401), .ZN(n2133) );
  OAI21_X1 U2774 ( .B1(n2052), .B2(n4311), .A(n2050), .ZN(n2049) );
  NOR2_X1 U2775 ( .A1(n4347), .A2(n4348), .ZN(n4346) );
  NOR2_X1 U2776 ( .A1(n4326), .A2(n3864), .ZN(n4347) );
  OR2_X1 U2777 ( .A1(n2761), .A2(n2068), .ZN(n2067) );
  NAND3_X1 U2778 ( .A1(n2067), .A2(n2066), .A3(n2063), .ZN(n4265) );
  OAI21_X1 U2779 ( .B1(n3191), .B2(n2834), .A(n3730), .ZN(n3162) );
  AND2_X1 U2780 ( .A1(n2305), .A2(n2304), .ZN(n2085) );
  NAND2_X1 U2781 ( .A1(n2348), .A2(n3805), .ZN(n2308) );
  OAI21_X1 U2782 ( .B1(n3262), .B2(n2089), .A(n2086), .ZN(n3294) );
  OAI21_X2 U2783 ( .B1(n2092), .B2(n2176), .A(n2173), .ZN(n3496) );
  NAND2_X1 U2784 ( .A1(n2094), .A2(n3605), .ZN(n3479) );
  OR2_X2 U2785 ( .A1(n3609), .A2(n3607), .ZN(n2094) );
  NAND2_X1 U2786 ( .A1(n2094), .A2(n2093), .ZN(n2096) );
  OAI211_X1 U2787 ( .C1(n2096), .C2(n2017), .A(n2095), .B(n2042), .ZN(U3217)
         );
  NAND2_X1 U2788 ( .A1(n2149), .A2(n2100), .ZN(n3146) );
  NAND2_X2 U2789 ( .A1(n2306), .A2(n2892), .ZN(n2636) );
  NAND2_X1 U2790 ( .A1(n2104), .A2(REG1_REG_12__SCAN_IN), .ZN(n2103) );
  NOR2_X1 U2791 ( .A1(n4342), .A2(n4341), .ZN(n4340) );
  AOI21_X1 U2792 ( .B1(n4342), .B2(n2043), .A(n2110), .ZN(n2109) );
  NOR2_X1 U2793 ( .A1(n4340), .A2(n2140), .ZN(n3879) );
  OAI21_X1 U2794 ( .B1(n3023), .B2(n3013), .A(n2118), .ZN(n2120) );
  INV_X1 U2795 ( .A(n2129), .ZN(n4125) );
  NAND2_X4 U2796 ( .A1(n2131), .A2(n2130), .ZN(n2583) );
  INV_X1 U2797 ( .A(n3109), .ZN(n3040) );
  MUX2_X1 U2798 ( .A(n2133), .B(n2132), .S(n2583), .Z(n3109) );
  AND2_X1 U2799 ( .A1(n2563), .A2(n2033), .ZN(n2290) );
  BUF_X4 U2800 ( .A(n2583), .Z(n3642) );
  NAND2_X1 U2801 ( .A1(n2950), .A2(REG1_REG_3__SCAN_IN), .ZN(n2953) );
  NAND2_X1 U2802 ( .A1(n3152), .A2(n3153), .ZN(n2149) );
  NAND2_X1 U2803 ( .A1(n2400), .A2(n2150), .ZN(n3262) );
  NAND2_X1 U2804 ( .A1(n3129), .A2(n2031), .ZN(n2151) );
  NAND2_X1 U2805 ( .A1(n3129), .A2(n2387), .ZN(n3207) );
  NAND2_X1 U2806 ( .A1(n3370), .A2(n2472), .ZN(n3353) );
  NAND2_X2 U2807 ( .A1(n2181), .A2(n2721), .ZN(n2306) );
  INV_X1 U2808 ( .A(n3232), .ZN(n2188) );
  NAND2_X1 U2809 ( .A1(n2184), .A2(n2185), .ZN(n2800) );
  NAND2_X1 U2810 ( .A1(n3232), .A2(n2796), .ZN(n2184) );
  NAND2_X1 U2811 ( .A1(n4068), .A2(n2190), .ZN(n2189) );
  AOI211_X2 U2812 ( .C1(n2810), .C2(n2013), .A(n2040), .B(n2811), .ZN(n4090)
         );
  NAND2_X1 U2813 ( .A1(n3397), .A2(n2009), .ZN(n2197) );
  NAND2_X1 U2814 ( .A1(n2197), .A2(n2198), .ZN(n3429) );
  NAND3_X1 U2815 ( .A1(n3054), .A2(n2832), .A3(n2787), .ZN(n2207) );
  NAND3_X1 U2816 ( .A1(n2208), .A2(n2788), .A3(n2207), .ZN(n3188) );
  NAND2_X1 U2817 ( .A1(n2787), .A2(n2209), .ZN(n2208) );
  NAND3_X1 U2818 ( .A1(n2211), .A2(n2793), .A3(n2210), .ZN(n3178) );
  NAND2_X1 U2819 ( .A1(n2792), .A2(n2212), .ZN(n2210) );
  NAND3_X1 U2820 ( .A1(n2789), .A2(n2792), .A3(n3189), .ZN(n2211) );
  OR2_X1 U2821 ( .A1(n3954), .A2(n2825), .ZN(n2228) );
  OAI21_X1 U2822 ( .B1(n3954), .B2(n2217), .A(n2214), .ZN(n2213) );
  INV_X1 U2823 ( .A(n2226), .ZN(n2216) );
  NAND2_X1 U2824 ( .A1(n2228), .A2(n2824), .ZN(n3935) );
  NAND2_X1 U2825 ( .A1(n2274), .A2(n2230), .ZN(n2270) );
  NAND2_X1 U2826 ( .A1(n2274), .A2(n2032), .ZN(n2229) );
  NOR2_X2 U2827 ( .A1(n2760), .A2(n2254), .ZN(n2255) );
  NAND2_X1 U2828 ( .A1(n2281), .A2(n2253), .ZN(n2760) );
  XNOR2_X1 U2829 ( .A(n3914), .B(n3913), .ZN(n3470) );
  NAND2_X1 U2830 ( .A1(n2315), .A2(n2317), .ZN(n2318) );
  NAND2_X1 U2831 ( .A1(n3467), .A2(n4265), .ZN(n2300) );
  OR3_X1 U2832 ( .A1(n3512), .A2(n3508), .A3(n3599), .ZN(n2232) );
  INV_X1 U2833 ( .A(n4053), .ZN(n4102) );
  INV_X1 U2834 ( .A(n4118), .ZN(n3565) );
  OR2_X1 U2835 ( .A1(n2306), .A2(n2311), .ZN(n2233) );
  NAND2_X1 U2836 ( .A1(n2739), .A2(n2738), .ZN(n2737) );
  INV_X1 U2837 ( .A(n2936), .ZN(n2285) );
  OR2_X1 U2838 ( .A1(n4022), .A2(n3680), .ZN(n2234) );
  OR3_X1 U2839 ( .A1(n2748), .A2(n3618), .A3(n2747), .ZN(n2235) );
  INV_X1 U2840 ( .A(n3798), .ZN(n3335) );
  INV_X1 U2841 ( .A(n4100), .ZN(n2813) );
  INV_X1 U2842 ( .A(n3422), .ZN(n3797) );
  AND4_X1 U2843 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .ZN(n3422)
         );
  OR2_X1 U2844 ( .A1(n3422), .A2(n3324), .ZN(n2236) );
  NAND2_X1 U2845 ( .A1(n4120), .A2(n3551), .ZN(n2237) );
  XNOR2_X1 U2846 ( .A(n2297), .B(n2701), .ZN(n2315) );
  XNOR2_X1 U2847 ( .A(n2315), .B(n2316), .ZN(n3034) );
  OR2_X1 U2848 ( .A1(n3471), .A2(n4263), .ZN(n2238) );
  OR2_X1 U2849 ( .A1(n3471), .A2(n4214), .ZN(n2239) );
  AND3_X1 U2850 ( .A1(n2356), .A2(n2355), .A3(n2354), .ZN(n2240) );
  INV_X1 U2851 ( .A(n3418), .ZN(n2514) );
  NAND2_X1 U2852 ( .A1(n2330), .A2(n2329), .ZN(n2331) );
  NAND2_X1 U2853 ( .A1(n2784), .A2(n2348), .ZN(n2299) );
  INV_X1 U2854 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U2855 ( .A1(n4079), .A2(n4059), .ZN(n3674) );
  OR2_X1 U2856 ( .A1(n2408), .A2(IR_REG_6__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U2857 ( .A1(n2583), .A2(n2283), .ZN(n2284) );
  NAND2_X1 U2858 ( .A1(n2232), .A2(n2598), .ZN(n2599) );
  INV_X1 U2859 ( .A(n2316), .ZN(n2317) );
  INV_X1 U2860 ( .A(n4005), .ZN(n3680) );
  INV_X1 U2861 ( .A(n4083), .ZN(n4078) );
  OR2_X1 U2862 ( .A1(n4435), .A2(n4268), .ZN(n2865) );
  INV_X1 U2863 ( .A(n3226), .ZN(n3265) );
  OR2_X1 U2864 ( .A1(n2779), .A2(n3618), .ZN(n2781) );
  AND2_X1 U2865 ( .A1(n2601), .A2(REG3_REG_20__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U2866 ( .A1(n2613), .A2(REG3_REG_21__SCAN_IN), .ZN(n2630) );
  INV_X1 U2867 ( .A(n3794), .ZN(n4105) );
  NOR2_X1 U2868 ( .A1(n2501), .A2(n3421), .ZN(n2526) );
  INV_X1 U2869 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3421) );
  OR2_X1 U2870 ( .A1(n4289), .A2(n3818), .ZN(n4325) );
  INV_X1 U2871 ( .A(n3793), .ZN(n3964) );
  AND4_X1 U2872 ( .A1(n2579), .A2(n2578), .A3(n2577), .A4(n2576), .ZN(n4118)
         );
  NAND2_X1 U2873 ( .A1(n2535), .A2(REG3_REG_16__SCAN_IN), .ZN(n2574) );
  INV_X1 U2874 ( .A(n2865), .ZN(n2765) );
  INV_X1 U2875 ( .A(n3894), .ZN(n3887) );
  OR2_X1 U2876 ( .A1(n2749), .A2(n3779), .ZN(n4147) );
  AND2_X1 U2877 ( .A1(n3642), .A2(DATAI_21_), .ZN(n3531) );
  XNOR2_X1 U2878 ( .A(n2419), .B(IR_REG_7__SCAN_IN), .ZN(n3007) );
  OR2_X1 U2879 ( .A1(n2402), .A2(n2401), .ZN(n2435) );
  AND2_X1 U2880 ( .A1(n2692), .A2(n2679), .ZN(n3949) );
  OAI21_X1 U2881 ( .B1(n2739), .B2(n2738), .A(n2737), .ZN(n2929) );
  OR2_X1 U2882 ( .A1(n2693), .A2(n2704), .ZN(n3930) );
  AND2_X1 U2883 ( .A1(n2589), .A2(n2588), .ZN(n4053) );
  INV_X1 U2884 ( .A(n4339), .ZN(n4372) );
  AND2_X1 U2885 ( .A1(n4266), .A2(n2930), .ZN(n4121) );
  AND2_X1 U2886 ( .A1(n4278), .A2(n3894), .ZN(n4111) );
  AND2_X1 U2887 ( .A1(n4111), .A2(n4440), .ZN(n4282) );
  NAND2_X1 U2888 ( .A1(n2726), .A2(n2725), .ZN(n2888) );
  NAND2_X1 U2889 ( .A1(n3642), .A2(DATAI_25_), .ZN(n3967) );
  INV_X1 U2890 ( .A(n2888), .ZN(n2876) );
  AND2_X1 U2891 ( .A1(n2509), .A2(n2532), .ZN(n4396) );
  NAND2_X1 U2892 ( .A1(n2929), .A2(STATE_REG_SCAN_IN), .ZN(n4388) );
  XNOR2_X1 U2893 ( .A(n3479), .B(n2016), .ZN(n3485) );
  OR2_X1 U2894 ( .A1(n2774), .A2(n2743), .ZN(n3618) );
  NAND2_X1 U2895 ( .A1(n2712), .A2(n2711), .ZN(n3924) );
  OAI211_X1 U2896 ( .C1(n4006), .C2(n2300), .A(n2641), .B(n2640), .ZN(n4022)
         );
  NAND4_X1 U2897 ( .A1(n2559), .A2(n2558), .A3(n2557), .A4(n2556), .ZN(n3794)
         );
  OR2_X1 U2898 ( .A1(n2447), .A2(n2446), .ZN(n3087) );
  INV_X1 U2899 ( .A(n4396), .ZN(n4324) );
  OR2_X1 U2900 ( .A1(n4289), .A2(n4287), .ZN(n4339) );
  NAND2_X1 U2901 ( .A1(n4453), .A2(n4440), .ZN(n4214) );
  OR2_X1 U2902 ( .A1(n2877), .A2(n2888), .ZN(n4451) );
  AND3_X1 U2903 ( .A1(n4434), .A2(n4433), .A3(n4432), .ZN(n4450) );
  OR2_X1 U2904 ( .A1(n2877), .A2(n2876), .ZN(n4441) );
  NAND2_X1 U2905 ( .A1(n2917), .A2(n3030), .ZN(n4387) );
  INV_X1 U2906 ( .A(n3881), .ZN(n4391) );
  OR4_X1 U2907 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(U3274) );
  INV_X2 U2908 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2909 ( .A(n3467), .ZN(n2261) );
  INV_X1 U2910 ( .A(IR_REG_27__SCAN_IN), .ZN(n2257) );
  INV_X1 U2911 ( .A(IR_REG_26__SCAN_IN), .ZN(n2256) );
  NAND3_X1 U2912 ( .A1(n2257), .A2(n2758), .A3(n2256), .ZN(n2258) );
  NAND2_X1 U2913 ( .A1(n2261), .A2(n2264), .ZN(n2262) );
  INV_X1 U2914 ( .A(n2319), .ZN(n2263) );
  NAND2_X1 U2915 ( .A1(n2263), .A2(REG2_REG_1__SCAN_IN), .ZN(n2267) );
  NAND2_X1 U2916 ( .A1(n2353), .A2(REG3_REG_1__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2917 ( .A1(n2340), .A2(REG1_REG_1__SCAN_IN), .ZN(n2265) );
  NAND4_X2 U2918 ( .A1(n2268), .A2(n2267), .A3(n2266), .A4(n2265), .ZN(n2784)
         );
  INV_X1 U2919 ( .A(IR_REG_23__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U2920 ( .A1(n2270), .A2(IR_REG_31__SCAN_IN), .ZN(n2271) );
  OAI21_X1 U2921 ( .B1(IR_REG_23__SCAN_IN), .B2(IR_REG_24__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2272) );
  NAND2_X1 U2922 ( .A1(n2739), .A2(n2272), .ZN(n2273) );
  INV_X1 U2923 ( .A(n2274), .ZN(n2275) );
  NAND2_X1 U2924 ( .A1(n2275), .A2(IR_REG_31__SCAN_IN), .ZN(n2276) );
  MUX2_X1 U2925 ( .A(IR_REG_31__SCAN_IN), .B(n2276), .S(IR_REG_21__SCAN_IN), 
        .Z(n2277) );
  NAND2_X1 U2926 ( .A1(n2277), .A2(n2019), .ZN(n3670) );
  NAND2_X1 U2927 ( .A1(n2278), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2928 ( .A1(n2294), .A2(n2293), .ZN(n2296) );
  NAND2_X1 U2929 ( .A1(n2296), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  NAND2_X1 U2930 ( .A1(n2784), .A2(n2698), .ZN(n2288) );
  INV_X1 U2931 ( .A(n2324), .ZN(n2282) );
  INV_X1 U2932 ( .A(DATAI_1_), .ZN(n2283) );
  INV_X1 U2933 ( .A(n3047), .ZN(n2286) );
  AND2_X4 U2934 ( .A1(n2306), .A2(n2829), .ZN(n2713) );
  NAND2_X1 U2935 ( .A1(n2286), .A2(n2713), .ZN(n2287) );
  NAND2_X1 U2936 ( .A1(n2288), .A2(n2287), .ZN(n2297) );
  NAND2_X1 U2937 ( .A1(n2019), .A2(IR_REG_31__SCAN_IN), .ZN(n2289) );
  MUX2_X1 U2938 ( .A(IR_REG_31__SCAN_IN), .B(n2289), .S(IR_REG_22__SCAN_IN), 
        .Z(n2292) );
  INV_X1 U2939 ( .A(n2290), .ZN(n2291) );
  OR2_X1 U2940 ( .A1(n2294), .A2(n2293), .ZN(n2295) );
  NAND2_X1 U2941 ( .A1(n4267), .A2(n3894), .ZN(n2755) );
  NAND2_X1 U2942 ( .A1(n2764), .A2(n3670), .ZN(n2749) );
  INV_X1 U2943 ( .A(n2749), .ZN(n2995) );
  AND2_X4 U2944 ( .A1(n2713), .A2(n4430), .ZN(n2348) );
  AND2_X1 U2945 ( .A1(n2299), .A2(n2298), .ZN(n2316) );
  NAND2_X1 U2946 ( .A1(n2008), .A2(REG0_REG_0__SCAN_IN), .ZN(n2305) );
  NAND2_X1 U2947 ( .A1(n2340), .A2(REG1_REG_0__SCAN_IN), .ZN(n2304) );
  NAND2_X1 U2948 ( .A1(n2353), .A2(REG3_REG_0__SCAN_IN), .ZN(n2303) );
  INV_X1 U2949 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2301) );
  INV_X4 U2950 ( .A(n2636), .ZN(n2698) );
  INV_X1 U2951 ( .A(n2306), .ZN(n2753) );
  AOI22_X1 U2952 ( .A1(n3040), .A2(n2698), .B1(n4401), .B2(n2753), .ZN(n2307)
         );
  NAND2_X1 U2953 ( .A1(n2308), .A2(n2307), .ZN(n3108) );
  NAND2_X1 U2954 ( .A1(n3040), .A2(n2713), .ZN(n2309) );
  AND2_X1 U2955 ( .A1(n2310), .A2(n2309), .ZN(n2312) );
  INV_X1 U2956 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2311) );
  NAND2_X1 U2957 ( .A1(n2312), .A2(n2233), .ZN(n3107) );
  NAND2_X1 U2958 ( .A1(n3108), .A2(n3107), .ZN(n2314) );
  NAND2_X1 U2959 ( .A1(n2312), .A2(n2716), .ZN(n2313) );
  NAND2_X1 U2960 ( .A1(n2314), .A2(n2313), .ZN(n3036) );
  NAND2_X1 U2961 ( .A1(n3034), .A2(n3036), .ZN(n3035) );
  NAND2_X1 U2962 ( .A1(n3035), .A2(n2318), .ZN(n3115) );
  INV_X1 U2963 ( .A(n3115), .ZN(n2334) );
  INV_X1 U2964 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2939) );
  OR2_X1 U2965 ( .A1(n2319), .A2(n2939), .ZN(n2322) );
  NAND2_X1 U2966 ( .A1(n2340), .A2(REG1_REG_2__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2967 ( .A1(n2006), .A2(REG0_REG_2__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2968 ( .A1(n3158), .A2(n2698), .ZN(n2330) );
  INV_X1 U2969 ( .A(n2325), .ZN(n2327) );
  INV_X1 U2970 ( .A(DATAI_2_), .ZN(n2328) );
  MUX2_X1 U2971 ( .A(n4275), .B(n2328), .S(n2583), .Z(n3116) );
  INV_X1 U2972 ( .A(n3116), .ZN(n2332) );
  NAND2_X1 U2973 ( .A1(n2332), .A2(n2713), .ZN(n2329) );
  AOI22_X1 U2974 ( .A1(n3158), .A2(n2348), .B1(n2332), .B2(n2698), .ZN(n2335)
         );
  XNOR2_X1 U2975 ( .A(n2336), .B(n2335), .ZN(n3112) );
  INV_X1 U2976 ( .A(n3112), .ZN(n2333) );
  NAND2_X1 U2977 ( .A1(n2334), .A2(n2333), .ZN(n3113) );
  NAND2_X1 U2978 ( .A1(n2336), .A2(n2335), .ZN(n2337) );
  NAND2_X1 U2979 ( .A1(n3113), .A2(n2337), .ZN(n3152) );
  INV_X1 U2980 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2338) );
  NAND2_X1 U2981 ( .A1(n2007), .A2(n2338), .ZN(n2344) );
  INV_X1 U2982 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U2983 ( .A1(n2008), .A2(REG0_REG_3__SCAN_IN), .ZN(n2342) );
  INV_X1 U2984 ( .A(n2340), .ZN(n2654) );
  NAND2_X1 U2985 ( .A1(n2340), .A2(REG1_REG_3__SCAN_IN), .ZN(n2341) );
  NAND2_X1 U2986 ( .A1(n3149), .A2(n2698), .ZN(n2346) );
  XNOR2_X1 U2987 ( .A(n2358), .B(IR_REG_3__SCAN_IN), .ZN(n4274) );
  MUX2_X1 U2988 ( .A(n4274), .B(DATAI_3_), .S(n3642), .Z(n3082) );
  NAND2_X1 U2989 ( .A1(n3082), .A2(n2713), .ZN(n2345) );
  NAND2_X1 U2990 ( .A1(n2346), .A2(n2345), .ZN(n2347) );
  AOI22_X1 U2991 ( .A1(n3149), .A2(n2348), .B1(n2698), .B2(n3082), .ZN(n2350)
         );
  XNOR2_X1 U2992 ( .A(n2349), .B(n2350), .ZN(n3153) );
  INV_X1 U2993 ( .A(n2349), .ZN(n2351) );
  NAND2_X1 U2994 ( .A1(n2351), .A2(n2350), .ZN(n2352) );
  NAND2_X1 U2995 ( .A1(n2651), .A2(REG2_REG_4__SCAN_IN), .ZN(n2357) );
  NAND2_X1 U2996 ( .A1(n2340), .A2(REG1_REG_4__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U2997 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2367) );
  OAI21_X1 U2998 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2367), .ZN(n3200) );
  OR2_X1 U2999 ( .A1(n2300), .A2(n3200), .ZN(n2355) );
  NAND2_X1 U3000 ( .A1(n2006), .A2(REG0_REG_4__SCAN_IN), .ZN(n2354) );
  NAND2_X1 U3001 ( .A1(n2358), .A2(n2373), .ZN(n2359) );
  NAND2_X1 U3002 ( .A1(n2359), .A2(IR_REG_31__SCAN_IN), .ZN(n2360) );
  XNOR2_X1 U3003 ( .A(n2360), .B(IR_REG_4__SCAN_IN), .ZN(n4273) );
  MUX2_X1 U3004 ( .A(n4273), .B(DATAI_4_), .S(n2583), .Z(n2790) );
  INV_X1 U3005 ( .A(n2361), .ZN(n2362) );
  XNOR2_X1 U3006 ( .A(n2362), .B(n2701), .ZN(n2364) );
  OAI22_X1 U3007 ( .A1(n3164), .A2(n2635), .B1(n2584), .B2(n3198), .ZN(n2363)
         );
  XNOR2_X1 U3008 ( .A(n2364), .B(n2363), .ZN(n3145) );
  NAND2_X1 U3009 ( .A1(n2364), .A2(n2363), .ZN(n2365) );
  AND2_X1 U3010 ( .A1(n2367), .A2(n2366), .ZN(n2368) );
  NOR2_X1 U3011 ( .A1(n2388), .A2(n2368), .ZN(n3170) );
  NAND2_X1 U3012 ( .A1(n2007), .A2(n3170), .ZN(n2372) );
  NAND2_X1 U3013 ( .A1(n2651), .A2(REG2_REG_5__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3014 ( .A1(n2006), .A2(REG0_REG_5__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3015 ( .A1(n2340), .A2(REG1_REG_5__SCAN_IN), .ZN(n2369) );
  NAND4_X1 U3016 ( .A1(n2372), .A2(n2371), .A3(n2370), .A4(n2369), .ZN(n3803)
         );
  NAND2_X1 U3017 ( .A1(n3803), .A2(n2698), .ZN(n2382) );
  INV_X1 U3018 ( .A(IR_REG_4__SCAN_IN), .ZN(n2374) );
  NAND2_X1 U3019 ( .A1(n2374), .A2(n2373), .ZN(n2375) );
  NAND2_X1 U3020 ( .A1(n2377), .A2(IR_REG_31__SCAN_IN), .ZN(n2376) );
  MUX2_X1 U3021 ( .A(n2376), .B(IR_REG_31__SCAN_IN), .S(n2378), .Z(n2379) );
  NAND2_X1 U3022 ( .A1(n2059), .A2(n2378), .ZN(n2408) );
  NAND2_X1 U3023 ( .A1(n2379), .A2(n2408), .ZN(n3844) );
  INV_X1 U3024 ( .A(DATAI_5_), .ZN(n2380) );
  MUX2_X1 U3025 ( .A(n3844), .B(n2380), .S(n2583), .Z(n3132) );
  NAND2_X1 U3026 ( .A1(n3169), .A2(n2713), .ZN(n2381) );
  NAND2_X1 U3027 ( .A1(n2382), .A2(n2381), .ZN(n2383) );
  XNOR2_X1 U3028 ( .A(n2383), .B(n2701), .ZN(n2386) );
  AOI22_X1 U3029 ( .A1(n3803), .A2(n2348), .B1(n3169), .B2(n2698), .ZN(n2384)
         );
  XNOR2_X1 U3030 ( .A(n2386), .B(n2384), .ZN(n3130) );
  NAND2_X1 U3031 ( .A1(n3131), .A2(n3130), .ZN(n3129) );
  INV_X1 U3032 ( .A(n2384), .ZN(n2385) );
  NAND2_X1 U3033 ( .A1(n2386), .A2(n2385), .ZN(n2387) );
  NAND2_X1 U3034 ( .A1(n2651), .A2(REG2_REG_6__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3035 ( .A1(n2388), .A2(REG3_REG_6__SCAN_IN), .ZN(n2402) );
  OR2_X1 U3036 ( .A1(n2388), .A2(REG3_REG_6__SCAN_IN), .ZN(n2389) );
  AND2_X1 U3037 ( .A1(n2402), .A2(n2389), .ZN(n3211) );
  NAND2_X1 U3038 ( .A1(n2007), .A2(n3211), .ZN(n2392) );
  NAND2_X1 U3039 ( .A1(n2006), .A2(REG0_REG_6__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U3040 ( .A1(n2340), .A2(REG1_REG_6__SCAN_IN), .ZN(n2390) );
  NAND4_X1 U3041 ( .A1(n2393), .A2(n2392), .A3(n2391), .A4(n2390), .ZN(n3802)
         );
  NAND2_X1 U3042 ( .A1(n3802), .A2(n2348), .ZN(n2396) );
  NAND2_X1 U3043 ( .A1(n2408), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  XNOR2_X1 U3044 ( .A(n2394), .B(IR_REG_6__SCAN_IN), .ZN(n4271) );
  MUX2_X1 U3045 ( .A(n4271), .B(DATAI_6_), .S(n2583), .Z(n3179) );
  NAND2_X1 U3046 ( .A1(n3179), .A2(n2698), .ZN(n2395) );
  NAND2_X1 U3047 ( .A1(n2396), .A2(n2395), .ZN(n3205) );
  NAND2_X1 U3048 ( .A1(n3802), .A2(n2698), .ZN(n2398) );
  NAND2_X1 U3049 ( .A1(n3179), .A2(n2713), .ZN(n2397) );
  NAND2_X1 U3050 ( .A1(n2398), .A2(n2397), .ZN(n2399) );
  XNOR2_X1 U3051 ( .A(n2399), .B(n2701), .ZN(n3204) );
  NAND2_X1 U3052 ( .A1(n3207), .A2(n3205), .ZN(n2400) );
  NAND2_X1 U3053 ( .A1(n2651), .A2(REG2_REG_7__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3054 ( .A1(n2006), .A2(REG0_REG_7__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3055 ( .A1(n2402), .A2(n2401), .ZN(n2403) );
  NAND2_X1 U3056 ( .A1(n2435), .A2(n2403), .ZN(n3270) );
  OR2_X1 U3057 ( .A1(n2300), .A2(n3270), .ZN(n2405) );
  NAND2_X1 U3058 ( .A1(n2340), .A2(REG1_REG_7__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3059 ( .A1(n2441), .A2(IR_REG_31__SCAN_IN), .ZN(n2419) );
  MUX2_X1 U3060 ( .A(n3007), .B(DATAI_7_), .S(n2583), .Z(n3226) );
  OAI22_X1 U3061 ( .A1(n3256), .A2(n2584), .B1(n2659), .B2(n3265), .ZN(n2409)
         );
  XNOR2_X1 U3062 ( .A(n2409), .B(n2716), .ZN(n2410) );
  OAI22_X1 U3063 ( .A1(n3256), .A2(n2635), .B1(n2584), .B2(n3265), .ZN(n2411)
         );
  XNOR2_X1 U3064 ( .A(n2410), .B(n2411), .ZN(n3261) );
  INV_X1 U3065 ( .A(n2410), .ZN(n2412) );
  NAND2_X1 U3066 ( .A1(n2412), .A2(n2411), .ZN(n2413) );
  XNOR2_X1 U3067 ( .A(n2435), .B(REG3_REG_8__SCAN_IN), .ZN(n3258) );
  NAND2_X1 U3068 ( .A1(n2007), .A2(n3258), .ZN(n2417) );
  NAND2_X1 U3069 ( .A1(n2651), .A2(REG2_REG_8__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3070 ( .A1(n2008), .A2(REG0_REG_8__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3071 ( .A1(n2340), .A2(REG1_REG_8__SCAN_IN), .ZN(n2414) );
  NAND4_X1 U3072 ( .A1(n2417), .A2(n2416), .A3(n2415), .A4(n2414), .ZN(n3800)
         );
  NAND2_X1 U3073 ( .A1(n3800), .A2(n2698), .ZN(n2424) );
  INV_X1 U3074 ( .A(IR_REG_7__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3075 ( .A1(n2419), .A2(n2418), .ZN(n2420) );
  NAND2_X1 U3076 ( .A1(n2420), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  INV_X1 U3077 ( .A(IR_REG_8__SCAN_IN), .ZN(n2421) );
  XNOR2_X1 U3078 ( .A(n2422), .B(n2421), .ZN(n3021) );
  INV_X1 U3079 ( .A(DATAI_8_), .ZN(n2905) );
  MUX2_X1 U3080 ( .A(n3021), .B(n2905), .S(n2583), .Z(n3243) );
  INV_X1 U3081 ( .A(n3243), .ZN(n3253) );
  NAND2_X1 U3082 ( .A1(n3253), .A2(n2713), .ZN(n2423) );
  NAND2_X1 U3083 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  XNOR2_X1 U3084 ( .A(n2425), .B(n2701), .ZN(n2428) );
  NAND2_X1 U3085 ( .A1(n3800), .A2(n2348), .ZN(n2427) );
  NAND2_X1 U3086 ( .A1(n3253), .A2(n2698), .ZN(n2426) );
  NAND2_X1 U3087 ( .A1(n2427), .A2(n2426), .ZN(n2429) );
  AND2_X1 U3088 ( .A1(n2428), .A2(n2429), .ZN(n3250) );
  INV_X1 U3089 ( .A(n2428), .ZN(n2431) );
  INV_X1 U3090 ( .A(n2429), .ZN(n2430) );
  NAND2_X1 U3091 ( .A1(n2651), .A2(REG2_REG_9__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U3092 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2432) );
  INV_X1 U3093 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2434) );
  INV_X1 U3094 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2433) );
  OAI21_X1 U3095 ( .B1(n2435), .B2(n2434), .A(n2433), .ZN(n2436) );
  AND2_X1 U3096 ( .A1(n2456), .A2(n2436), .ZN(n3299) );
  NAND2_X1 U3097 ( .A1(n2007), .A2(n3299), .ZN(n2439) );
  NAND2_X1 U3098 ( .A1(n2006), .A2(REG0_REG_9__SCAN_IN), .ZN(n2438) );
  NAND2_X1 U3099 ( .A1(n2340), .A2(REG1_REG_9__SCAN_IN), .ZN(n2437) );
  NAND4_X1 U3100 ( .A1(n2440), .A2(n2439), .A3(n2438), .A4(n2437), .ZN(n3799)
         );
  NAND2_X1 U3101 ( .A1(n3799), .A2(n2698), .ZN(n2449) );
  INV_X1 U3102 ( .A(n2441), .ZN(n2443) );
  NOR2_X1 U3103 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2442)
         );
  AOI21_X1 U3104 ( .B1(n2443), .B2(n2442), .A(n2759), .ZN(n2444) );
  MUX2_X1 U3105 ( .A(n2759), .B(n2444), .S(IR_REG_9__SCAN_IN), .Z(n2447) );
  INV_X1 U3106 ( .A(n2445), .ZN(n2446) );
  INV_X1 U3107 ( .A(n3087), .ZN(n3095) );
  MUX2_X1 U3108 ( .A(n3095), .B(DATAI_9_), .S(n3642), .Z(n3279) );
  NAND2_X1 U3109 ( .A1(n3279), .A2(n2713), .ZN(n2448) );
  NAND2_X1 U3110 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  XNOR2_X1 U3111 ( .A(n2450), .B(n2701), .ZN(n2451) );
  AOI22_X1 U3112 ( .A1(n3799), .A2(n2348), .B1(n2698), .B2(n3279), .ZN(n2452)
         );
  XNOR2_X1 U3113 ( .A(n2451), .B(n2452), .ZN(n3295) );
  INV_X1 U3114 ( .A(n2451), .ZN(n2453) );
  NAND2_X1 U3115 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  AND2_X1 U3116 ( .A1(n2456), .A2(n4495), .ZN(n2457) );
  NOR2_X1 U3117 ( .A1(n2473), .A2(n2457), .ZN(n3375) );
  NAND2_X1 U3118 ( .A1(n2007), .A2(n3375), .ZN(n2461) );
  NAND2_X1 U3119 ( .A1(n2651), .A2(REG2_REG_10__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3120 ( .A1(n2008), .A2(REG0_REG_10__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3121 ( .A1(n2340), .A2(REG1_REG_10__SCAN_IN), .ZN(n2458) );
  NAND4_X1 U3122 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3798)
         );
  NAND2_X1 U3123 ( .A1(n3798), .A2(n2698), .ZN(n2466) );
  NAND2_X1 U3124 ( .A1(n2445), .A2(IR_REG_31__SCAN_IN), .ZN(n2462) );
  MUX2_X1 U3125 ( .A(IR_REG_31__SCAN_IN), .B(n2462), .S(IR_REG_10__SCAN_IN), 
        .Z(n2464) );
  INV_X1 U3126 ( .A(n2506), .ZN(n2463) );
  NAND2_X1 U3127 ( .A1(n2464), .A2(n2463), .ZN(n4303) );
  MUX2_X1 U3128 ( .A(n4399), .B(DATAI_10_), .S(n2583), .Z(n3365) );
  NAND2_X1 U3129 ( .A1(n3365), .A2(n2713), .ZN(n2465) );
  NAND2_X1 U3130 ( .A1(n2466), .A2(n2465), .ZN(n2467) );
  XNOR2_X1 U3131 ( .A(n2467), .B(n2716), .ZN(n2468) );
  AOI22_X1 U3132 ( .A1(n3798), .A2(n2348), .B1(n2698), .B2(n3365), .ZN(n2469)
         );
  XNOR2_X1 U3133 ( .A(n2468), .B(n2469), .ZN(n3372) );
  INV_X1 U3134 ( .A(n2468), .ZN(n2471) );
  INV_X1 U3135 ( .A(n2469), .ZN(n2470) );
  NAND2_X1 U3136 ( .A1(n2471), .A2(n2470), .ZN(n2472) );
  NAND2_X1 U3137 ( .A1(n2651), .A2(REG2_REG_11__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U3138 ( .A1(n2006), .A2(REG0_REG_11__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3139 ( .A1(n2340), .A2(REG1_REG_11__SCAN_IN), .ZN(n2476) );
  OR2_X1 U3140 ( .A1(n2473), .A2(REG3_REG_11__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3141 ( .A1(n2487), .A2(n2474), .ZN(n3363) );
  OR2_X1 U3142 ( .A1(n2300), .A2(n3363), .ZN(n2475) );
  OR2_X1 U3143 ( .A1(n2506), .A2(n2759), .ZN(n2481) );
  INV_X1 U3144 ( .A(n2481), .ZN(n2479) );
  NAND2_X1 U3145 ( .A1(n2479), .A2(IR_REG_11__SCAN_IN), .ZN(n2482) );
  INV_X1 U3146 ( .A(IR_REG_11__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3147 ( .A1(n2481), .A2(n2480), .ZN(n2493) );
  MUX2_X1 U31480 ( .A(n3872), .B(DATAI_11_), .S(n2583), .Z(n3343) );
  OAI22_X1 U31490 ( .A1(n3389), .A2(n2635), .B1(n2584), .B2(n3358), .ZN(n3354)
         );
  OAI22_X1 U3150 ( .A1(n3389), .A2(n2584), .B1(n2659), .B2(n3358), .ZN(n2483)
         );
  XNOR2_X1 U3151 ( .A(n2483), .B(n2701), .ZN(n3355) );
  OAI21_X1 U3152 ( .B1(n3353), .B2(n3354), .A(n3355), .ZN(n2485) );
  NAND2_X1 U3153 ( .A1(n3353), .A2(n3354), .ZN(n2484) );
  NAND2_X1 U3154 ( .A1(n2651), .A2(REG2_REG_12__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3155 ( .A1(n2006), .A2(REG0_REG_12__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U3156 ( .A1(n2487), .A2(n2486), .ZN(n2488) );
  NAND2_X1 U3157 ( .A1(n2501), .A2(n2488), .ZN(n3326) );
  OR2_X1 U3158 ( .A1(n2300), .A2(n3326), .ZN(n2490) );
  NAND2_X1 U3159 ( .A1(n2340), .A2(REG1_REG_12__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3160 ( .A1(n2493), .A2(IR_REG_31__SCAN_IN), .ZN(n2494) );
  XNOR2_X1 U3161 ( .A(n2494), .B(IR_REG_12__SCAN_IN), .ZN(n3873) );
  INV_X1 U3162 ( .A(DATAI_12_), .ZN(n2495) );
  MUX2_X1 U3163 ( .A(n4398), .B(n2495), .S(n2583), .Z(n3324) );
  OAI22_X1 U3164 ( .A1(n3422), .A2(n2584), .B1(n2659), .B2(n3324), .ZN(n2496)
         );
  XNOR2_X1 U3165 ( .A(n2496), .B(n2701), .ZN(n2497) );
  OAI22_X1 U3166 ( .A1(n3422), .A2(n2635), .B1(n2584), .B2(n3324), .ZN(n2498)
         );
  AND2_X1 U3167 ( .A1(n2497), .A2(n2498), .ZN(n3383) );
  INV_X1 U3168 ( .A(n2497), .ZN(n2500) );
  INV_X1 U3169 ( .A(n2498), .ZN(n2499) );
  NAND2_X1 U3170 ( .A1(n2500), .A2(n2499), .ZN(n3382) );
  AOI22_X1 U3171 ( .A1(n2651), .A2(REG2_REG_13__SCAN_IN), .B1(n2008), .B2(
        REG0_REG_13__SCAN_IN), .ZN(n2504) );
  AND2_X1 U3172 ( .A1(n2501), .A2(n3421), .ZN(n2502) );
  NOR2_X1 U3173 ( .A1(n2526), .A2(n2502), .ZN(n3425) );
  AOI22_X1 U3174 ( .A1(n2007), .A2(n3425), .B1(n2340), .B2(
        REG1_REG_13__SCAN_IN), .ZN(n2503) );
  NOR2_X1 U3175 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2505)
         );
  NAND2_X1 U3176 ( .A1(n2506), .A2(n2505), .ZN(n2508) );
  NAND2_X1 U3177 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2507) );
  MUX2_X1 U3178 ( .A(IR_REG_31__SCAN_IN), .B(n2507), .S(IR_REG_13__SCAN_IN), 
        .Z(n2509) );
  INV_X1 U3179 ( .A(DATAI_13_), .ZN(n2510) );
  MUX2_X1 U3180 ( .A(n4324), .B(n2510), .S(n3642), .Z(n3423) );
  OAI22_X1 U3181 ( .A1(n3491), .A2(n2584), .B1(n2659), .B2(n3423), .ZN(n2511)
         );
  XNOR2_X1 U3182 ( .A(n2511), .B(n2716), .ZN(n3418) );
  OR2_X1 U3183 ( .A1(n3491), .A2(n2635), .ZN(n2513) );
  NAND2_X1 U3184 ( .A1(n3403), .A2(n2698), .ZN(n2512) );
  NAND2_X1 U3185 ( .A1(n2513), .A2(n2512), .ZN(n3419) );
  NAND2_X1 U3186 ( .A1(n2651), .A2(REG2_REG_14__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3187 ( .A1(n2008), .A2(REG0_REG_14__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3188 ( .A1(n2340), .A2(REG1_REG_14__SCAN_IN), .ZN(n2516) );
  XNOR2_X1 U3189 ( .A(n2526), .B(REG3_REG_14__SCAN_IN), .ZN(n3455) );
  OR2_X1 U3190 ( .A1(n2300), .A2(n3455), .ZN(n2515) );
  NAND2_X1 U3191 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2519) );
  XNOR2_X1 U3192 ( .A(n2519), .B(IR_REG_14__SCAN_IN), .ZN(n4334) );
  MUX2_X1 U3193 ( .A(n4334), .B(DATAI_14_), .S(n2583), .Z(n3489) );
  INV_X1 U3194 ( .A(n3489), .ZN(n3453) );
  OAI22_X1 U3195 ( .A1(n3626), .A2(n2584), .B1(n3453), .B2(n2659), .ZN(n2520)
         );
  XNOR2_X1 U3196 ( .A(n2520), .B(n2716), .ZN(n2524) );
  INV_X1 U3197 ( .A(n2524), .ZN(n2521) );
  OAI22_X1 U3198 ( .A1(n3626), .A2(n2635), .B1(n3453), .B2(n2584), .ZN(n2522)
         );
  NAND2_X1 U3199 ( .A1(n2521), .A2(n2522), .ZN(n3487) );
  INV_X1 U3200 ( .A(n2522), .ZN(n2523) );
  NAND2_X1 U3201 ( .A1(n2651), .A2(REG2_REG_15__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U3202 ( .A1(n2006), .A2(REG0_REG_15__SCAN_IN), .ZN(n2530) );
  AND2_X1 U3203 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2525) );
  AOI21_X1 U3204 ( .B1(n2526), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2527) );
  OR2_X1 U3205 ( .A1(n2535), .A2(n2527), .ZN(n3632) );
  OR2_X1 U3206 ( .A1(n2300), .A2(n3632), .ZN(n2529) );
  NAND2_X1 U3207 ( .A1(n2340), .A2(REG1_REG_15__SCAN_IN), .ZN(n2528) );
  OAI21_X1 U3208 ( .B1(n2532), .B2(IR_REG_14__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2542) );
  XNOR2_X1 U3209 ( .A(n2542), .B(IR_REG_15__SCAN_IN), .ZN(n4394) );
  INV_X1 U32100 ( .A(DATAI_15_), .ZN(n2533) );
  MUX2_X1 U32110 ( .A(n4352), .B(n2533), .S(n2583), .Z(n3627) );
  OAI22_X1 U32120 ( .A1(n3555), .A2(n2584), .B1(n2659), .B2(n3627), .ZN(n2534)
         );
  XNOR2_X1 U32130 ( .A(n2534), .B(n2701), .ZN(n2552) );
  NAND2_X1 U32140 ( .A1(n2651), .A2(REG2_REG_16__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32150 ( .A1(n2006), .A2(REG0_REG_16__SCAN_IN), .ZN(n2539) );
  OR2_X1 U32160 ( .A1(n2535), .A2(REG3_REG_16__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32170 ( .A1(n2574), .A2(n2536), .ZN(n3550) );
  OR2_X1 U32180 ( .A1(n2300), .A2(n3550), .ZN(n2538) );
  NAND2_X1 U32190 ( .A1(n2340), .A2(REG1_REG_16__SCAN_IN), .ZN(n2537) );
  INV_X1 U32200 ( .A(IR_REG_15__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32210 ( .A1(n2542), .A2(n2541), .ZN(n2543) );
  NAND2_X1 U32220 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2545) );
  INV_X1 U32230 ( .A(IR_REG_16__SCAN_IN), .ZN(n2544) );
  INV_X1 U32240 ( .A(n4393), .ZN(n2546) );
  MUX2_X1 U32250 ( .A(n2546), .B(DATAI_16_), .S(n2583), .Z(n3551) );
  OAI22_X1 U32260 ( .A1(n3563), .A2(n2584), .B1(n2898), .B2(n2659), .ZN(n2547)
         );
  XNOR2_X1 U32270 ( .A(n2547), .B(n2701), .ZN(n2549) );
  INV_X1 U32280 ( .A(n2549), .ZN(n2551) );
  OAI22_X1 U32290 ( .A1(n3563), .A2(n2635), .B1(n2898), .B2(n2584), .ZN(n2548)
         );
  INV_X1 U32300 ( .A(n2548), .ZN(n2550) );
  OAI21_X1 U32310 ( .B1(n2551), .B2(n2550), .A(n2554), .ZN(n3548) );
  OAI22_X1 U32320 ( .A1(n3555), .A2(n2635), .B1(n2584), .B2(n3627), .ZN(n3621)
         );
  INV_X1 U32330 ( .A(n2554), .ZN(n2555) );
  XNOR2_X1 U32340 ( .A(n2574), .B(REG3_REG_17__SCAN_IN), .ZN(n4128) );
  NAND2_X1 U32350 ( .A1(n2007), .A2(n4128), .ZN(n2559) );
  NAND2_X1 U32360 ( .A1(n2651), .A2(REG2_REG_17__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U32370 ( .A1(n2008), .A2(REG0_REG_17__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U32380 ( .A1(n2340), .A2(REG1_REG_17__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U32390 ( .A1(n3794), .A2(n2698), .ZN(n2567) );
  NOR2_X1 U32400 ( .A1(n2560), .A2(n2759), .ZN(n2561) );
  MUX2_X1 U32410 ( .A(n2759), .B(n2561), .S(IR_REG_17__SCAN_IN), .Z(n2562) );
  INV_X1 U32420 ( .A(n2562), .ZN(n2565) );
  INV_X1 U32430 ( .A(n2563), .ZN(n2564) );
  INV_X1 U32440 ( .A(DATAI_17_), .ZN(n4390) );
  MUX2_X1 U32450 ( .A(n4391), .B(n4390), .S(n2583), .Z(n4126) );
  NAND2_X1 U32460 ( .A1(n2871), .A2(n2713), .ZN(n2566) );
  NAND2_X1 U32470 ( .A1(n2567), .A2(n2566), .ZN(n2568) );
  XNOR2_X1 U32480 ( .A(n2568), .B(n2716), .ZN(n2570) );
  AOI22_X1 U32490 ( .A1(n3794), .A2(n2348), .B1(n2871), .B2(n2698), .ZN(n2569)
         );
  NOR2_X1 U32500 ( .A1(n2570), .A2(n2569), .ZN(n3560) );
  NAND2_X1 U32510 ( .A1(n2651), .A2(REG2_REG_18__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32520 ( .A1(n2006), .A2(REG0_REG_18__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32530 ( .A1(n2340), .A2(REG1_REG_18__SCAN_IN), .ZN(n2577) );
  INV_X1 U32540 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2572) );
  INV_X1 U32550 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2571) );
  OAI21_X1 U32560 ( .B1(n2574), .B2(n2572), .A(n2571), .ZN(n2575) );
  NAND2_X1 U32570 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2573) );
  NAND2_X1 U32580 ( .A1(n2575), .A2(n2586), .ZN(n4096) );
  OR2_X1 U32590 ( .A1(n2300), .A2(n4096), .ZN(n2576) );
  NOR2_X1 U32600 ( .A1(n2563), .A2(n2759), .ZN(n2580) );
  MUX2_X1 U32610 ( .A(n2759), .B(n2580), .S(IR_REG_18__SCAN_IN), .Z(n2582) );
  INV_X1 U32620 ( .A(n2278), .ZN(n2581) );
  MUX2_X1 U32630 ( .A(n4270), .B(DATAI_18_), .S(n2583), .Z(n4100) );
  OAI22_X1 U32640 ( .A1(n4118), .A2(n2635), .B1(n2584), .B2(n2813), .ZN(n3508)
         );
  OAI22_X1 U32650 ( .A1(n4118), .A2(n2584), .B1(n2659), .B2(n2813), .ZN(n2585)
         );
  XNOR2_X1 U32660 ( .A(n2585), .B(n2701), .ZN(n3599) );
  AOI22_X1 U32670 ( .A1(n2651), .A2(REG2_REG_19__SCAN_IN), .B1(n2008), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2589) );
  AND2_X1 U32680 ( .A1(n2586), .A2(n3515), .ZN(n2587) );
  NOR2_X1 U32690 ( .A1(n2601), .A2(n2587), .ZN(n4084) );
  AOI22_X1 U32700 ( .A1(n2007), .A2(n4084), .B1(n2340), .B2(
        REG1_REG_19__SCAN_IN), .ZN(n2588) );
  INV_X1 U32710 ( .A(DATAI_19_), .ZN(n2590) );
  MUX2_X1 U32720 ( .A(n3894), .B(n2590), .S(n3642), .Z(n4083) );
  OAI22_X1 U32730 ( .A1(n4053), .A2(n2636), .B1(n2659), .B2(n4083), .ZN(n2591)
         );
  XNOR2_X1 U32740 ( .A(n2591), .B(n2716), .ZN(n2594) );
  OR2_X1 U32750 ( .A1(n4053), .A2(n2635), .ZN(n2593) );
  NAND2_X1 U32760 ( .A1(n4078), .A2(n2698), .ZN(n2592) );
  AND2_X1 U32770 ( .A1(n2593), .A2(n2592), .ZN(n2595) );
  NOR2_X1 U32780 ( .A1(n2594), .A2(n2595), .ZN(n3512) );
  AOI21_X1 U32790 ( .B1(n3508), .B2(n3599), .A(n3512), .ZN(n2600) );
  INV_X1 U32800 ( .A(n2594), .ZN(n2597) );
  INV_X1 U32810 ( .A(n2595), .ZN(n2596) );
  NOR2_X1 U32820 ( .A1(n2597), .A2(n2596), .ZN(n3511) );
  NAND2_X1 U32830 ( .A1(n2651), .A2(REG2_REG_20__SCAN_IN), .ZN(n2606) );
  NOR2_X1 U32840 ( .A1(n2601), .A2(REG3_REG_20__SCAN_IN), .ZN(n2602) );
  NOR2_X1 U32850 ( .A1(n2613), .A2(n2602), .ZN(n4062) );
  NAND2_X1 U32860 ( .A1(n2007), .A2(n4062), .ZN(n2605) );
  NAND2_X1 U32870 ( .A1(n2008), .A2(REG0_REG_20__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U32880 ( .A1(n2340), .A2(REG1_REG_20__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U32890 ( .A1(n4079), .A2(n2698), .ZN(n2608) );
  NAND2_X1 U32900 ( .A1(n4059), .A2(n2713), .ZN(n2607) );
  NAND2_X1 U32910 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  XNOR2_X1 U32920 ( .A(n2609), .B(n2716), .ZN(n2612) );
  AND2_X1 U32930 ( .A1(n2698), .A2(n4059), .ZN(n2610) );
  AOI21_X1 U32940 ( .B1(n4079), .B2(n2348), .A(n2610), .ZN(n2611) );
  NOR2_X1 U32950 ( .A1(n2612), .A2(n2611), .ZN(n3579) );
  NOR2_X2 U32960 ( .A1(n3524), .A2(n3579), .ZN(n3582) );
  AND2_X1 U32970 ( .A1(n2612), .A2(n2611), .ZN(n3525) );
  NAND2_X1 U32980 ( .A1(n2651), .A2(REG2_REG_21__SCAN_IN), .ZN(n2618) );
  OR2_X1 U32990 ( .A1(n2613), .A2(REG3_REG_21__SCAN_IN), .ZN(n2614) );
  AND2_X1 U33000 ( .A1(n2630), .A2(n2614), .ZN(n3528) );
  NAND2_X1 U33010 ( .A1(n2007), .A2(n3528), .ZN(n2617) );
  NAND2_X1 U33020 ( .A1(n2006), .A2(REG0_REG_21__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U33030 ( .A1(n2340), .A2(REG1_REG_21__SCAN_IN), .ZN(n2615) );
  NAND4_X1 U33040 ( .A1(n2618), .A2(n2617), .A3(n2616), .A4(n2615), .ZN(n4051)
         );
  NAND2_X1 U33050 ( .A1(n4051), .A2(n2698), .ZN(n2620) );
  NAND2_X1 U33060 ( .A1(n3531), .A2(n2713), .ZN(n2619) );
  NAND2_X1 U33070 ( .A1(n2620), .A2(n2619), .ZN(n2621) );
  XNOR2_X1 U33080 ( .A(n2621), .B(n2701), .ZN(n2627) );
  INV_X1 U33090 ( .A(n2627), .ZN(n2625) );
  NAND2_X1 U33100 ( .A1(n4051), .A2(n2348), .ZN(n2623) );
  NAND2_X1 U33110 ( .A1(n3531), .A2(n2698), .ZN(n2622) );
  NAND2_X1 U33120 ( .A1(n2623), .A2(n2622), .ZN(n2626) );
  INV_X1 U33130 ( .A(n2626), .ZN(n2624) );
  NAND2_X1 U33140 ( .A1(n2625), .A2(n2624), .ZN(n3521) );
  AND2_X1 U33150 ( .A1(n2627), .A2(n2626), .ZN(n3522) );
  NAND2_X1 U33160 ( .A1(n2006), .A2(REG0_REG_22__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U33170 ( .A1(n2340), .A2(REG1_REG_22__SCAN_IN), .ZN(n2628) );
  AND2_X1 U33180 ( .A1(n2629), .A2(n2628), .ZN(n2634) );
  INV_X1 U33190 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U33200 ( .A1(n2630), .A2(n3593), .ZN(n2631) );
  NAND2_X1 U33210 ( .A1(n2638), .A2(n2631), .ZN(n4016) );
  OR2_X1 U33220 ( .A1(n4016), .A2(n2300), .ZN(n2633) );
  NAND2_X1 U33230 ( .A1(n2651), .A2(REG2_REG_22__SCAN_IN), .ZN(n2632) );
  INV_X1 U33240 ( .A(n4015), .ZN(n4025) );
  OAI22_X1 U33250 ( .A1(n4030), .A2(n2635), .B1(n4025), .B2(n2584), .ZN(n2646)
         );
  OAI22_X1 U33260 ( .A1(n4030), .A2(n2636), .B1(n4025), .B2(n2659), .ZN(n2637)
         );
  XNOR2_X1 U33270 ( .A(n2637), .B(n2701), .ZN(n2647) );
  XOR2_X1 U33280 ( .A(n2646), .B(n2647), .Z(n3590) );
  INV_X1 U33290 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U33300 ( .A1(n2638), .A2(n3500), .ZN(n2639) );
  NAND2_X1 U33310 ( .A1(n2649), .A2(n2639), .ZN(n4006) );
  AOI22_X1 U33320 ( .A1(n2651), .A2(REG2_REG_23__SCAN_IN), .B1(n2006), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33330 ( .A1(n2340), .A2(REG1_REG_23__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U33340 ( .A1(n4022), .A2(n2698), .ZN(n2643) );
  NAND2_X1 U33350 ( .A1(n3680), .A2(n2713), .ZN(n2642) );
  NAND2_X1 U33360 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
  XNOR2_X1 U33370 ( .A(n2644), .B(n2701), .ZN(n2658) );
  NOR2_X1 U33380 ( .A1(n4005), .A2(n2584), .ZN(n2645) );
  AOI21_X1 U33390 ( .B1(n4022), .B2(n2348), .A(n2645), .ZN(n2656) );
  XNOR2_X1 U33400 ( .A(n2658), .B(n2656), .ZN(n3498) );
  OR2_X1 U33410 ( .A1(n2647), .A2(n2646), .ZN(n3499) );
  INV_X1 U33420 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4172) );
  INV_X1 U33430 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3574) );
  AND2_X1 U33440 ( .A1(n2649), .A2(n3574), .ZN(n2650) );
  NOR2_X1 U33450 ( .A1(n2663), .A2(n2650), .ZN(n3987) );
  NAND2_X1 U33460 ( .A1(n3987), .A2(n2007), .ZN(n2653) );
  AOI22_X1 U33470 ( .A1(n2651), .A2(REG2_REG_24__SCAN_IN), .B1(n2006), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2652) );
  OAI211_X1 U33480 ( .C1(n2654), .C2(n4172), .A(n2653), .B(n2652), .ZN(n4001)
         );
  NOR2_X1 U33490 ( .A1(n3985), .A2(n2584), .ZN(n2655) );
  AOI21_X1 U33500 ( .B1(n4001), .B2(n2348), .A(n2655), .ZN(n2661) );
  INV_X1 U33510 ( .A(n2656), .ZN(n2657) );
  NAND2_X1 U33520 ( .A1(n2658), .A2(n2657), .ZN(n2662) );
  NAND3_X1 U3353 ( .A1(n3496), .A2(n2661), .A3(n2662), .ZN(n3569) );
  OAI22_X1 U33540 ( .A1(n3541), .A2(n2584), .B1(n2659), .B2(n3985), .ZN(n2660)
         );
  XNOR2_X1 U3355 ( .A(n2660), .B(n2701), .ZN(n3572) );
  OR2_X1 U3356 ( .A1(n2663), .A2(REG3_REG_25__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3357 ( .A1(n2663), .A2(REG3_REG_25__SCAN_IN), .ZN(n2678) );
  AND2_X1 U3358 ( .A1(n2664), .A2(n2678), .ZN(n3969) );
  NAND2_X1 U3359 ( .A1(n3969), .A2(n2007), .ZN(n2670) );
  INV_X1 U3360 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3361 ( .A1(n2340), .A2(REG1_REG_25__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3362 ( .A1(n2008), .A2(REG0_REG_25__SCAN_IN), .ZN(n2665) );
  OAI211_X1 U3363 ( .C1(n2319), .C2(n2667), .A(n2666), .B(n2665), .ZN(n2668)
         );
  INV_X1 U3364 ( .A(n2668), .ZN(n2669) );
  NAND2_X1 U3365 ( .A1(n3981), .A2(n2698), .ZN(n2672) );
  NAND2_X1 U3366 ( .A1(n3961), .A2(n2713), .ZN(n2671) );
  NAND2_X1 U3367 ( .A1(n2672), .A2(n2671), .ZN(n2673) );
  XNOR2_X1 U3368 ( .A(n2673), .B(n2701), .ZN(n2677) );
  NAND2_X1 U3369 ( .A1(n3981), .A2(n2348), .ZN(n2675) );
  NAND2_X1 U3370 ( .A1(n3961), .A2(n2698), .ZN(n2674) );
  NAND2_X1 U3371 ( .A1(n2675), .A2(n2674), .ZN(n2676) );
  NOR2_X1 U3372 ( .A1(n2677), .A2(n2676), .ZN(n3537) );
  NAND2_X1 U3373 ( .A1(n2677), .A2(n2676), .ZN(n3538) );
  INV_X1 U3374 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3612) );
  NAND2_X1 U3375 ( .A1(n2678), .A2(n3612), .ZN(n2679) );
  NAND2_X1 U3376 ( .A1(n3949), .A2(n2007), .ZN(n2685) );
  INV_X1 U3377 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3378 ( .A1(n2340), .A2(REG1_REG_26__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3379 ( .A1(n2008), .A2(REG0_REG_26__SCAN_IN), .ZN(n2680) );
  OAI211_X1 U3380 ( .C1(n2319), .C2(n2682), .A(n2681), .B(n2680), .ZN(n2683)
         );
  INV_X1 U3381 ( .A(n2683), .ZN(n2684) );
  NAND2_X1 U3382 ( .A1(n3793), .A2(n2698), .ZN(n2687) );
  INV_X1 U3383 ( .A(n3948), .ZN(n3941) );
  NAND2_X1 U3384 ( .A1(n3941), .A2(n2713), .ZN(n2686) );
  NAND2_X1 U3385 ( .A1(n2687), .A2(n2686), .ZN(n2688) );
  XNOR2_X1 U3386 ( .A(n2688), .B(n2716), .ZN(n2691) );
  NOR2_X1 U3387 ( .A1(n3948), .A2(n2584), .ZN(n2689) );
  AOI21_X1 U3388 ( .B1(n3793), .B2(n2348), .A(n2689), .ZN(n2690) );
  NOR2_X1 U3389 ( .A1(n2691), .A2(n2690), .ZN(n3607) );
  NAND2_X1 U3390 ( .A1(n2691), .A2(n2690), .ZN(n3605) );
  INV_X1 U3391 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4496) );
  AND2_X1 U3392 ( .A1(n2692), .A2(n4496), .ZN(n2693) );
  INV_X1 U3393 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U3394 ( .A1(n2340), .A2(REG1_REG_27__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U3395 ( .A1(n2006), .A2(REG0_REG_27__SCAN_IN), .ZN(n2694) );
  OAI211_X1 U3396 ( .C1(n2319), .C2(n3929), .A(n2695), .B(n2694), .ZN(n2696)
         );
  INV_X1 U3397 ( .A(n2696), .ZN(n2697) );
  NAND2_X1 U3398 ( .A1(n3942), .A2(n2698), .ZN(n2700) );
  NAND2_X1 U3399 ( .A1(n3767), .A2(n2713), .ZN(n2699) );
  NAND2_X1 U3400 ( .A1(n2700), .A2(n2699), .ZN(n2702) );
  XNOR2_X1 U3401 ( .A(n2702), .B(n2701), .ZN(n2746) );
  NOR2_X1 U3402 ( .A1(n3928), .A2(n2584), .ZN(n2703) );
  AOI21_X1 U3403 ( .B1(n3942), .B2(n2348), .A(n2703), .ZN(n2744) );
  NAND2_X1 U3404 ( .A1(n2704), .A2(REG3_REG_28__SCAN_IN), .ZN(n3899) );
  INV_X1 U3405 ( .A(n2704), .ZN(n2706) );
  INV_X1 U3406 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3407 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  NAND2_X1 U3408 ( .A1(n3899), .A2(n2707), .ZN(n3473) );
  INV_X1 U3409 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U3410 ( .A1(n2340), .A2(REG1_REG_28__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U3411 ( .A1(n2008), .A2(REG0_REG_28__SCAN_IN), .ZN(n2708) );
  OAI211_X1 U3412 ( .C1(n2319), .C2(n3472), .A(n2709), .B(n2708), .ZN(n2710)
         );
  INV_X1 U3413 ( .A(n2710), .ZN(n2711) );
  NAND2_X1 U3414 ( .A1(n3924), .A2(n2698), .ZN(n2715) );
  NAND2_X1 U3415 ( .A1(n3642), .A2(DATAI_28_), .ZN(n2873) );
  NAND2_X1 U3416 ( .A1(n3912), .A2(n2713), .ZN(n2714) );
  NAND2_X1 U3417 ( .A1(n2715), .A2(n2714), .ZN(n2717) );
  XNOR2_X1 U3418 ( .A(n2717), .B(n2716), .ZN(n2719) );
  AOI22_X1 U3419 ( .A1(n3924), .A2(n2348), .B1(n3912), .B2(n2698), .ZN(n2718)
         );
  XNOR2_X1 U3420 ( .A(n2719), .B(n2718), .ZN(n2780) );
  INV_X1 U3421 ( .A(n2780), .ZN(n2748) );
  NAND2_X1 U3422 ( .A1(n2720), .A2(B_REG_SCAN_IN), .ZN(n2722) );
  MUX2_X1 U3423 ( .A(n2722), .B(B_REG_SCAN_IN), .S(n2721), .Z(n2723) );
  INV_X1 U3424 ( .A(D_REG_0__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3425 ( .A1(n2916), .A2(n2920), .ZN(n2726) );
  INV_X1 U3426 ( .A(n2721), .ZN(n2724) );
  NAND2_X1 U3427 ( .A1(n2724), .A2(n2182), .ZN(n2725) );
  NOR4_X1 U3428 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2730) );
  NOR4_X1 U3429 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2729) );
  NOR4_X1 U3430 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2728) );
  NOR4_X1 U3431 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2727) );
  NAND4_X1 U3432 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(n2736)
         );
  NOR2_X1 U3433 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_25__SCAN_IN), .ZN(n2734)
         );
  NOR4_X1 U3434 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2733) );
  NOR4_X1 U3435 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2732) );
  NOR4_X1 U3436 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2731) );
  NAND4_X1 U3437 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .ZN(n2735)
         );
  OAI21_X1 U3438 ( .B1(n2736), .B2(n2735), .A(n2916), .ZN(n2867) );
  NAND2_X1 U3439 ( .A1(n2720), .A2(n2182), .ZN(n2864) );
  AND2_X1 U3440 ( .A1(n2867), .A2(n2864), .ZN(n2890) );
  INV_X1 U3441 ( .A(D_REG_1__SCAN_IN), .ZN(n2923) );
  NAND2_X1 U3442 ( .A1(n2916), .A2(n2923), .ZN(n2887) );
  NAND3_X1 U3443 ( .A1(n2876), .A2(n2890), .A3(n2887), .ZN(n2774) );
  NAND2_X1 U3444 ( .A1(n3779), .A2(n3894), .ZN(n2751) );
  INV_X1 U3445 ( .A(n2751), .ZN(n2741) );
  NOR2_X1 U3446 ( .A1(n2749), .A2(n2741), .ZN(n2742) );
  NOR2_X1 U3447 ( .A1(n2742), .A2(n2930), .ZN(n2750) );
  NAND2_X1 U3448 ( .A1(n3030), .A2(n2750), .ZN(n2743) );
  INV_X1 U3449 ( .A(n2744), .ZN(n2745) );
  AND2_X1 U3450 ( .A1(n2746), .A2(n2745), .ZN(n2779) );
  INV_X1 U3451 ( .A(n2779), .ZN(n2747) );
  OAI21_X1 U3452 ( .B1(n4099), .B2(n2750), .A(n2774), .ZN(n2752) );
  NAND2_X1 U3453 ( .A1(n2930), .A2(n2751), .ZN(n2885) );
  NAND2_X1 U3454 ( .A1(n2752), .A2(n2885), .ZN(n3028) );
  INV_X1 U3455 ( .A(n2929), .ZN(n2754) );
  NOR3_X1 U3456 ( .A1(n3028), .A2(n2754), .A3(n2753), .ZN(n2757) );
  NOR2_X1 U3457 ( .A1(n4388), .A2(n2755), .ZN(n2756) );
  NAND2_X1 U34580 ( .A1(n2774), .A2(n3786), .ZN(n3029) );
  OAI21_X2 U34590 ( .B1(n2757), .B2(U3149), .A(n3029), .ZN(n3616) );
  INV_X1 U3460 ( .A(n3616), .ZN(n3633) );
  MUX2_X1 U3461 ( .A(n2760), .B(n2759), .S(n2758), .Z(n2762) );
  NAND2_X1 U3462 ( .A1(n3786), .A2(n4266), .ZN(n2763) );
  INV_X1 U3463 ( .A(n3625), .ZN(n3530) );
  AOI22_X1 U3464 ( .A1(n3942), .A2(n3530), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2776) );
  NOR3_X1 U3465 ( .A1(n2774), .A2(n4147), .A3(n2928), .ZN(n2766) );
  AND2_X1 U3466 ( .A1(n3779), .A2(n3887), .ZN(n4376) );
  NAND2_X1 U34670 ( .A1(n4376), .A2(n2764), .ZN(n4435) );
  INV_X1 U3468 ( .A(n2005), .ZN(n3552) );
  OR2_X1 U34690 ( .A1(n3899), .A2(n2300), .ZN(n2772) );
  INV_X1 U3470 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U34710 ( .A1(n2340), .A2(REG1_REG_29__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U3472 ( .A1(n2006), .A2(REG0_REG_29__SCAN_IN), .ZN(n2767) );
  OAI211_X1 U34730 ( .C1(n2319), .C2(n2769), .A(n2768), .B(n2767), .ZN(n2770)
         );
  INV_X1 U3474 ( .A(n2770), .ZN(n2771) );
  NAND2_X1 U34750 ( .A1(n2772), .A2(n2771), .ZN(n3792) );
  INV_X1 U3476 ( .A(n4266), .ZN(n3815) );
  NAND2_X1 U34770 ( .A1(n3786), .A2(n3815), .ZN(n2773) );
  AOI22_X1 U3478 ( .A1(n3912), .A2(n3552), .B1(n3792), .B2(n3629), .ZN(n2775)
         );
  OAI211_X1 U34790 ( .C1(n3633), .C2(n3473), .A(n2776), .B(n2775), .ZN(n2777)
         );
  INV_X1 U3480 ( .A(n2777), .ZN(n2778) );
  NOR2_X1 U34810 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  INV_X1 U3482 ( .A(n2784), .ZN(n2783) );
  NAND2_X1 U34830 ( .A1(n2783), .A2(n2286), .ZN(n2831) );
  NAND2_X1 U3484 ( .A1(n2784), .A2(n3047), .ZN(n3717) );
  NAND2_X1 U34850 ( .A1(n2831), .A2(n3717), .ZN(n3043) );
  NAND2_X1 U3486 ( .A1(n3042), .A2(n3043), .ZN(n3041) );
  NAND2_X1 U34870 ( .A1(n2784), .A2(n2286), .ZN(n2785) );
  NAND2_X1 U3488 ( .A1(n3158), .A2(n3116), .ZN(n3723) );
  INV_X1 U34890 ( .A(n3158), .ZN(n3077) );
  NAND2_X1 U3490 ( .A1(n3077), .A2(n3116), .ZN(n2786) );
  NAND2_X1 U34910 ( .A1(n3149), .A2(n3082), .ZN(n2787) );
  INV_X1 U3492 ( .A(n3149), .ZN(n3192) );
  INV_X1 U34930 ( .A(n3082), .ZN(n3155) );
  NAND2_X1 U3494 ( .A1(n3192), .A2(n3155), .ZN(n2788) );
  INV_X1 U34950 ( .A(n3188), .ZN(n2789) );
  NAND2_X1 U3496 ( .A1(n3804), .A2(n3198), .ZN(n3730) );
  NAND2_X1 U34970 ( .A1(n3164), .A2(n2790), .ZN(n3726) );
  NAND2_X1 U3498 ( .A1(n3730), .A2(n3726), .ZN(n3189) );
  NAND2_X1 U34990 ( .A1(n3804), .A2(n2790), .ZN(n2791) );
  INV_X1 U3500 ( .A(n3803), .ZN(n3175) );
  NAND2_X1 U35010 ( .A1(n3175), .A2(n3132), .ZN(n2792) );
  NAND2_X1 U3502 ( .A1(n3803), .A2(n3169), .ZN(n2793) );
  AND2_X1 U35030 ( .A1(n3802), .A2(n3179), .ZN(n2794) );
  NAND2_X1 U3504 ( .A1(n3256), .A2(n3226), .ZN(n2836) );
  NAND2_X1 U35050 ( .A1(n3801), .A2(n3265), .ZN(n3737) );
  NAND2_X1 U35060 ( .A1(n3801), .A2(n3226), .ZN(n2796) );
  INV_X1 U35070 ( .A(n3800), .ZN(n2797) );
  NAND2_X1 U35080 ( .A1(n2797), .A2(n3243), .ZN(n2798) );
  NAND2_X1 U35090 ( .A1(n3800), .A2(n3253), .ZN(n2799) );
  NAND2_X1 U35100 ( .A1(n2800), .A2(n2799), .ZN(n3278) );
  AND2_X1 U35110 ( .A1(n3799), .A2(n3279), .ZN(n2802) );
  INV_X1 U35120 ( .A(n3799), .ZN(n3368) );
  INV_X1 U35130 ( .A(n3279), .ZN(n3296) );
  NAND2_X1 U35140 ( .A1(n3368), .A2(n3296), .ZN(n2801) );
  NAND2_X1 U35150 ( .A1(n3389), .A2(n3343), .ZN(n3315) );
  INV_X1 U35160 ( .A(n3389), .ZN(n3364) );
  NAND2_X1 U35170 ( .A1(n3364), .A2(n3358), .ZN(n3317) );
  NAND2_X1 U35180 ( .A1(n3389), .A2(n3358), .ZN(n2803) );
  NAND2_X1 U35190 ( .A1(n3332), .A2(n2803), .ZN(n3322) );
  NAND2_X1 U35200 ( .A1(n3322), .A2(n2236), .ZN(n2805) );
  INV_X1 U35210 ( .A(n3324), .ZN(n3387) );
  NAND2_X1 U35220 ( .A1(n2805), .A2(n2804), .ZN(n3397) );
  NAND2_X1 U35230 ( .A1(n3626), .A2(n3489), .ZN(n3430) );
  NAND2_X1 U35240 ( .A1(n3795), .A2(n3453), .ZN(n3650) );
  NAND2_X1 U35250 ( .A1(n3430), .A2(n3650), .ZN(n3442) );
  NAND2_X1 U35260 ( .A1(n3429), .A2(n2808), .ZN(n2810) );
  INV_X1 U35270 ( .A(n3627), .ZN(n2845) );
  NAND2_X1 U35280 ( .A1(n3563), .A2(n3551), .ZN(n3644) );
  NAND2_X1 U35290 ( .A1(n4120), .A2(n2898), .ZN(n3751) );
  NAND2_X1 U35300 ( .A1(n4118), .A2(n4100), .ZN(n4072) );
  NAND2_X1 U35310 ( .A1(n3565), .A2(n2813), .ZN(n4073) );
  NAND2_X1 U35320 ( .A1(n4072), .A2(n4073), .ZN(n4092) );
  NAND2_X1 U35330 ( .A1(n4090), .A2(n4092), .ZN(n4091) );
  NAND2_X1 U35340 ( .A1(n4051), .A2(n3531), .ZN(n2818) );
  NOR2_X1 U35350 ( .A1(n4051), .A2(n3531), .ZN(n2817) );
  AOI21_X1 U35360 ( .B1(n4035), .B2(n2818), .A(n2817), .ZN(n4013) );
  NAND2_X1 U35370 ( .A1(n4030), .A2(n4015), .ZN(n3997) );
  NAND2_X1 U35380 ( .A1(n3529), .A2(n4025), .ZN(n2855) );
  NAND2_X1 U35390 ( .A1(n3997), .A2(n2855), .ZN(n4020) );
  NAND2_X1 U35400 ( .A1(n4013), .A2(n4020), .ZN(n4012) );
  NAND2_X1 U35410 ( .A1(n3529), .A2(n4015), .ZN(n2819) );
  NAND2_X1 U35420 ( .A1(n4012), .A2(n2819), .ZN(n3992) );
  NAND2_X1 U35430 ( .A1(n3992), .A2(n2234), .ZN(n2821) );
  NAND2_X1 U35440 ( .A1(n4022), .A2(n3680), .ZN(n2820) );
  NAND2_X1 U35450 ( .A1(n2821), .A2(n2820), .ZN(n3974) );
  NOR2_X1 U35460 ( .A1(n3541), .A2(n3985), .ZN(n2823) );
  NAND2_X1 U35470 ( .A1(n3541), .A2(n3985), .ZN(n2822) );
  NOR2_X1 U35480 ( .A1(n3981), .A2(n3961), .ZN(n2825) );
  NAND2_X1 U35490 ( .A1(n3981), .A2(n3961), .ZN(n2824) );
  NOR2_X1 U35500 ( .A1(n3964), .A2(n3948), .ZN(n2826) );
  NOR2_X1 U35510 ( .A1(n3942), .A2(n3767), .ZN(n2828) );
  NAND2_X1 U35520 ( .A1(n3942), .A2(n3767), .ZN(n2827) );
  NOR2_X1 U35530 ( .A1(n3924), .A2(n2873), .ZN(n3900) );
  NAND2_X1 U35540 ( .A1(n3924), .A2(n2873), .ZN(n3635) );
  INV_X1 U35550 ( .A(n3635), .ZN(n3902) );
  OR2_X1 U35560 ( .A1(n3900), .A2(n3902), .ZN(n3913) );
  XNOR2_X1 U35570 ( .A(n4267), .B(n2829), .ZN(n2830) );
  NAND2_X1 U35580 ( .A1(n2830), .A2(n3894), .ZN(n4057) );
  INV_X1 U35590 ( .A(n3043), .ZN(n3705) );
  NOR2_X1 U35600 ( .A1(n3805), .A2(n3109), .ZN(n3719) );
  NAND2_X1 U35610 ( .A1(n3705), .A2(n3719), .ZN(n3055) );
  NAND2_X1 U35620 ( .A1(n3055), .A2(n2831), .ZN(n2833) );
  INV_X1 U35630 ( .A(n2832), .ZN(n3696) );
  NAND2_X1 U35640 ( .A1(n2833), .A2(n3696), .ZN(n3057) );
  NAND2_X1 U35650 ( .A1(n3057), .A2(n3720), .ZN(n3075) );
  NAND2_X1 U35660 ( .A1(n3192), .A2(n3082), .ZN(n3725) );
  NAND2_X1 U35670 ( .A1(n3149), .A2(n3155), .ZN(n3722) );
  NAND2_X1 U35680 ( .A1(n3075), .A2(n3697), .ZN(n3074) );
  NAND2_X1 U35690 ( .A1(n3074), .A2(n3725), .ZN(n3191) );
  INV_X1 U35700 ( .A(n3726), .ZN(n2834) );
  OR2_X1 U35710 ( .A1(n3803), .A2(n3132), .ZN(n3734) );
  NAND2_X1 U35720 ( .A1(n3803), .A2(n3132), .ZN(n3728) );
  INV_X1 U35730 ( .A(n3179), .ZN(n3208) );
  AND2_X1 U35740 ( .A1(n3802), .A2(n3208), .ZN(n3735) );
  OR2_X1 U35750 ( .A1(n3173), .A2(n3735), .ZN(n2835) );
  INV_X1 U35760 ( .A(n3802), .ZN(n3264) );
  NAND2_X1 U35770 ( .A1(n3264), .A2(n3179), .ZN(n3732) );
  NAND2_X1 U35780 ( .A1(n2835), .A2(n3732), .ZN(n3224) );
  INV_X1 U35790 ( .A(n2836), .ZN(n2837) );
  OAI21_X1 U35800 ( .B1(n3224), .B2(n2837), .A(n3737), .ZN(n3238) );
  OR2_X1 U35810 ( .A1(n3800), .A2(n3243), .ZN(n3740) );
  NAND2_X1 U3582 ( .A1(n3800), .A2(n3243), .ZN(n3736) );
  AND2_X1 U3583 ( .A1(n3799), .A2(n3296), .ZN(n3744) );
  NAND2_X1 U3584 ( .A1(n3368), .A2(n3279), .ZN(n3741) );
  NAND2_X1 U3585 ( .A1(n3798), .A2(n2136), .ZN(n3746) );
  NAND2_X1 U3586 ( .A1(n3303), .A2(n3746), .ZN(n2838) );
  NAND2_X1 U3587 ( .A1(n3335), .A2(n3365), .ZN(n3743) );
  NAND2_X1 U3588 ( .A1(n3797), .A2(n3324), .ZN(n3398) );
  NAND2_X1 U3589 ( .A1(n3796), .A2(n3423), .ZN(n2839) );
  NAND2_X1 U3590 ( .A1(n3398), .A2(n2839), .ZN(n2841) );
  INV_X1 U3591 ( .A(n3317), .ZN(n2840) );
  NOR2_X1 U3592 ( .A1(n2841), .A2(n2840), .ZN(n3747) );
  NAND2_X1 U3593 ( .A1(n3422), .A2(n3387), .ZN(n3400) );
  NAND2_X1 U3594 ( .A1(n3315), .A2(n3400), .ZN(n2844) );
  INV_X1 U3595 ( .A(n2841), .ZN(n2843) );
  NOR2_X1 U3596 ( .A1(n3796), .A2(n3423), .ZN(n2842) );
  AOI21_X1 U3597 ( .B1(n2844), .B2(n2843), .A(n2842), .ZN(n3749) );
  INV_X1 U3598 ( .A(n3442), .ZN(n3706) );
  NAND2_X1 U3599 ( .A1(n3555), .A2(n2845), .ZN(n3646) );
  NAND2_X1 U3600 ( .A1(n2807), .A2(n3627), .ZN(n3649) );
  NAND2_X1 U3601 ( .A1(n3646), .A2(n3649), .ZN(n3703) );
  INV_X1 U3602 ( .A(n3430), .ZN(n3647) );
  NOR2_X1 U3603 ( .A1(n3703), .A2(n3647), .ZN(n2846) );
  NAND2_X1 U3604 ( .A1(n3444), .A2(n2846), .ZN(n2847) );
  NAND2_X1 U3605 ( .A1(n2847), .A2(n3649), .ZN(n2894) );
  NAND2_X1 U3606 ( .A1(n2894), .A2(n3693), .ZN(n2848) );
  NAND2_X1 U3607 ( .A1(n4102), .A2(n4083), .ZN(n2849) );
  AND2_X1 U3608 ( .A1(n4073), .A2(n2849), .ZN(n2851) );
  NAND2_X1 U3609 ( .A1(n3794), .A2(n4126), .ZN(n4069) );
  NAND2_X1 U3610 ( .A1(n2851), .A2(n4069), .ZN(n3652) );
  OR2_X1 U3611 ( .A1(n3794), .A2(n4126), .ZN(n4070) );
  NAND2_X1 U3612 ( .A1(n4072), .A2(n4070), .ZN(n2852) );
  NOR2_X1 U3613 ( .A1(n4102), .A2(n4083), .ZN(n2850) );
  AOI21_X1 U3614 ( .B1(n2852), .B2(n2851), .A(n2850), .ZN(n4047) );
  INV_X1 U3615 ( .A(n4079), .ZN(n3516) );
  NAND2_X1 U3616 ( .A1(n3516), .A2(n4059), .ZN(n2853) );
  INV_X1 U3617 ( .A(n4059), .ZN(n3584) );
  INV_X1 U3618 ( .A(n4051), .ZN(n3592) );
  NAND2_X1 U3619 ( .A1(n3592), .A2(n3531), .ZN(n3995) );
  NAND2_X1 U3620 ( .A1(n3997), .A2(n3995), .ZN(n3760) );
  INV_X1 U3621 ( .A(n3760), .ZN(n2854) );
  NAND2_X1 U3622 ( .A1(n4031), .A2(n2854), .ZN(n2858) );
  NAND2_X1 U3623 ( .A1(n4022), .A2(n4005), .ZN(n2856) );
  NAND2_X1 U3624 ( .A1(n2856), .A2(n2855), .ZN(n3763) );
  INV_X1 U3625 ( .A(n3531), .ZN(n4039) );
  AND2_X1 U3626 ( .A1(n4051), .A2(n4039), .ZN(n3994) );
  AND2_X1 U3627 ( .A1(n3997), .A2(n3994), .ZN(n2857) );
  NOR2_X1 U3628 ( .A1(n3763), .A2(n2857), .ZN(n3655) );
  NAND2_X1 U3629 ( .A1(n2858), .A2(n3655), .ZN(n3976) );
  OR2_X1 U3630 ( .A1(n4001), .A2(n3985), .ZN(n3668) );
  OR2_X1 U3631 ( .A1(n4022), .A2(n4005), .ZN(n3975) );
  NAND2_X1 U3632 ( .A1(n3976), .A2(n3762), .ZN(n3956) );
  AND2_X1 U3633 ( .A1(n3981), .A2(n3967), .ZN(n3671) );
  AND2_X1 U3634 ( .A1(n4001), .A2(n3985), .ZN(n3667) );
  NOR2_X1 U3635 ( .A1(n3671), .A2(n3667), .ZN(n3766) );
  NAND2_X1 U3636 ( .A1(n3956), .A2(n3766), .ZN(n3938) );
  NOR2_X1 U3637 ( .A1(n3793), .A2(n3948), .ZN(n3702) );
  NOR2_X1 U3638 ( .A1(n3981), .A2(n3967), .ZN(n3936) );
  NOR2_X1 U3639 ( .A1(n3702), .A2(n3936), .ZN(n3773) );
  XNOR2_X1 U3640 ( .A(n3942), .B(n3767), .ZN(n3926) );
  NOR2_X1 U3641 ( .A1(n3942), .A2(n3928), .ZN(n3636) );
  AOI21_X1 U3642 ( .B1(n3922), .B2(n3926), .A(n3636), .ZN(n3903) );
  XNOR2_X1 U3643 ( .A(n3903), .B(n3913), .ZN(n2863) );
  NAND2_X1 U3644 ( .A1(n4267), .A2(n3887), .ZN(n2859) );
  INV_X1 U3645 ( .A(n3779), .ZN(n4269) );
  NAND2_X1 U3646 ( .A1(n4268), .A2(n4269), .ZN(n3634) );
  NAND2_X1 U3647 ( .A1(n3942), .A2(n4121), .ZN(n2861) );
  AND2_X2 U3648 ( .A1(n3815), .A2(n2930), .ZN(n4101) );
  NAND2_X1 U3649 ( .A1(n3792), .A2(n4101), .ZN(n2860) );
  OAI211_X1 U3650 ( .C1(n4147), .C2(n2873), .A(n2861), .B(n2860), .ZN(n2862)
         );
  AOI21_X1 U3651 ( .B1(n2863), .B2(n4107), .A(n2862), .ZN(n3474) );
  OAI21_X1 U3652 ( .B1(n3470), .B2(n4422), .A(n3474), .ZN(n2878) );
  NAND2_X1 U3653 ( .A1(n2887), .A2(n2864), .ZN(n2869) );
  NAND2_X1 U3654 ( .A1(n2885), .A2(n2865), .ZN(n2866) );
  NOR2_X1 U3655 ( .A1(n2928), .A2(n2866), .ZN(n2868) );
  NAND3_X1 U3656 ( .A1(n2869), .A2(n2868), .A3(n2867), .ZN(n2877) );
  INV_X1 U3657 ( .A(n2870), .ZN(n2875) );
  NAND2_X1 U3658 ( .A1(n3064), .A2(n3116), .ZN(n3081) );
  NAND2_X1 U3659 ( .A1(n3199), .A2(n3198), .ZN(n3197) );
  INV_X1 U3660 ( .A(n3985), .ZN(n2872) );
  INV_X1 U3661 ( .A(n3927), .ZN(n2874) );
  NAND2_X1 U3662 ( .A1(n2875), .A2(n2239), .ZN(U3546) );
  INV_X1 U3663 ( .A(n2879), .ZN(n2880) );
  NAND2_X1 U3664 ( .A1(n2880), .A2(n2238), .ZN(U3514) );
  INV_X1 U3665 ( .A(n2882), .ZN(n2883) );
  AOI21_X1 U3666 ( .B1(n3693), .B2(n2881), .A(n2883), .ZN(n2884) );
  INV_X1 U3667 ( .A(n2884), .ZN(n4206) );
  INV_X1 U3668 ( .A(n2885), .ZN(n2886) );
  NOR2_X1 U3669 ( .A1(n2928), .A2(n2886), .ZN(n2889) );
  NAND4_X1 U3670 ( .A1(n2890), .A2(n2889), .A3(n2888), .A4(n2887), .ZN(n2891)
         );
  INV_X2 U3671 ( .A(n4063), .ZN(n4278) );
  NAND2_X1 U3672 ( .A1(n2892), .A2(n3887), .ZN(n3072) );
  NAND2_X1 U3673 ( .A1(n4057), .A2(n3072), .ZN(n2893) );
  NOR2_X1 U3674 ( .A1(n4206), .A2(n4135), .ZN(n2903) );
  XNOR2_X1 U3675 ( .A(n2894), .B(n2196), .ZN(n2897) );
  AOI22_X1 U3676 ( .A1(n3794), .A2(n4101), .B1(n3551), .B2(n4099), .ZN(n2895)
         );
  OAI21_X1 U3677 ( .B1(n3555), .B2(n4104), .A(n2895), .ZN(n2896) );
  AOI21_X1 U3678 ( .B1(n2897), .B2(n4107), .A(n2896), .ZN(n4205) );
  NOR2_X1 U3679 ( .A1(n4205), .A2(n4063), .ZN(n2902) );
  OR2_X1 U3680 ( .A1(n3436), .A2(n2898), .ZN(n4203) );
  AND3_X1 U3681 ( .A1(n4203), .A2(n4202), .A3(n4282), .ZN(n2901) );
  INV_X1 U3682 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2899) );
  OAI22_X1 U3683 ( .A1(n4278), .A2(n2899), .B1(n3550), .B2(n4129), .ZN(n2900)
         );
  INV_X1 U3684 ( .A(DATAI_11_), .ZN(n4481) );
  NAND2_X1 U3685 ( .A1(n3872), .A2(STATE_REG_SCAN_IN), .ZN(n2904) );
  OAI21_X1 U3686 ( .B1(STATE_REG_SCAN_IN), .B2(n4481), .A(n2904), .ZN(U3341)
         );
  MUX2_X1 U3687 ( .A(n2905), .B(n3021), .S(STATE_REG_SCAN_IN), .Z(n2906) );
  INV_X1 U3688 ( .A(n2906), .ZN(U3344) );
  MUX2_X1 U3689 ( .A(n3894), .B(n2590), .S(U3149), .Z(n2907) );
  INV_X1 U3690 ( .A(n2907), .ZN(U3333) );
  INV_X1 U3691 ( .A(DATAI_7_), .ZN(n2908) );
  INV_X1 U3692 ( .A(n3007), .ZN(n2962) );
  MUX2_X1 U3693 ( .A(n2908), .B(n2962), .S(STATE_REG_SCAN_IN), .Z(n2909) );
  INV_X1 U3694 ( .A(n2909), .ZN(U3345) );
  INV_X1 U3695 ( .A(DATAI_9_), .ZN(n2910) );
  MUX2_X1 U3696 ( .A(n3087), .B(n2910), .S(U3149), .Z(n2911) );
  INV_X1 U3697 ( .A(n2911), .ZN(U3343) );
  INV_X1 U3698 ( .A(DATAI_26_), .ZN(n4485) );
  NAND2_X1 U3699 ( .A1(n2918), .A2(STATE_REG_SCAN_IN), .ZN(n2912) );
  OAI21_X1 U3700 ( .B1(STATE_REG_SCAN_IN), .B2(n4485), .A(n2912), .ZN(U3326)
         );
  INV_X1 U3701 ( .A(DATAI_31_), .ZN(n2915) );
  OR4_X1 U3702 ( .A1(n2913), .A2(IR_REG_30__SCAN_IN), .A3(n2759), .A4(U3149), 
        .ZN(n2914) );
  OAI21_X1 U3703 ( .B1(STATE_REG_SCAN_IN), .B2(n2915), .A(n2914), .ZN(U3321)
         );
  INV_X1 U3704 ( .A(n2916), .ZN(n2917) );
  NOR3_X1 U3705 ( .A1(n2721), .A2(n4388), .A3(n2918), .ZN(n2919) );
  AOI21_X1 U3706 ( .B1(n4387), .B2(n2920), .A(n2919), .ZN(U3458) );
  NOR2_X1 U3707 ( .A1(n2921), .A2(n4388), .ZN(n2922) );
  AOI22_X1 U3708 ( .A1(n4387), .A2(n2923), .B1(n2922), .B2(n2182), .ZN(U3459)
         );
  INV_X1 U3709 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4581) );
  NAND2_X1 U3710 ( .A1(n3158), .A2(U4043), .ZN(n2924) );
  OAI21_X1 U3711 ( .B1(U4043), .B2(n4581), .A(n2924), .ZN(U3552) );
  INV_X1 U3712 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U3713 ( .A1(n3149), .A2(U4043), .ZN(n2925) );
  OAI21_X1 U3714 ( .B1(U4043), .B2(n4585), .A(n2925), .ZN(U3553) );
  INV_X1 U3715 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U3716 ( .A1(n3565), .A2(U4043), .ZN(n2926) );
  OAI21_X1 U3717 ( .B1(U4043), .B2(n4588), .A(n2926), .ZN(U3568) );
  INV_X1 U3718 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U3719 ( .A1(n3529), .A2(U4043), .ZN(n2927) );
  OAI21_X1 U3720 ( .B1(U4043), .B2(n4587), .A(n2927), .ZN(U3572) );
  INV_X1 U3721 ( .A(n4274), .ZN(n2948) );
  OR2_X1 U3722 ( .A1(n2929), .A2(U3149), .ZN(n3790) );
  NAND2_X1 U3723 ( .A1(n2928), .A2(n3790), .ZN(n2943) );
  NAND2_X1 U3724 ( .A1(n2930), .A2(n2929), .ZN(n2931) );
  NAND2_X1 U3725 ( .A1(n2943), .A2(n2944), .ZN(n4289) );
  XNOR2_X1 U3726 ( .A(n2932), .B(IR_REG_27__SCAN_IN), .ZN(n4287) );
  AND2_X1 U3727 ( .A1(n4401), .A2(REG1_REG_0__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U3728 ( .A1(n3810), .A2(n3809), .ZN(n3808) );
  NAND2_X1 U3729 ( .A1(n2285), .A2(REG1_REG_1__SCAN_IN), .ZN(n2933) );
  NAND2_X1 U3730 ( .A1(n3808), .A2(n2933), .ZN(n3824) );
  INV_X1 U3731 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2934) );
  OR2_X1 U3732 ( .A1(n4275), .A2(n2934), .ZN(n2935) );
  XOR2_X1 U3733 ( .A(REG1_REG_3__SCAN_IN), .B(n2950), .Z(n2942) );
  NAND2_X1 U3734 ( .A1(n4266), .A2(n4287), .ZN(n3818) );
  INV_X1 U3735 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2937) );
  MUX2_X1 U3736 ( .A(n2937), .B(REG2_REG_1__SCAN_IN), .S(n2936), .Z(n3807) );
  AND2_X1 U3737 ( .A1(n4401), .A2(REG2_REG_0__SCAN_IN), .ZN(n3820) );
  NAND2_X1 U3738 ( .A1(n3807), .A2(n3820), .ZN(n3806) );
  NAND2_X1 U3739 ( .A1(n2285), .A2(REG2_REG_1__SCAN_IN), .ZN(n2938) );
  NAND2_X1 U3740 ( .A1(n3806), .A2(n2938), .ZN(n3829) );
  NAND2_X1 U3741 ( .A1(n3830), .A2(n3829), .ZN(n3828) );
  OR2_X1 U3742 ( .A1(n4275), .A2(n2939), .ZN(n2940) );
  NAND2_X1 U3743 ( .A1(n3828), .A2(n2940), .ZN(n2965) );
  XNOR2_X1 U3744 ( .A(n2964), .B(n2339), .ZN(n2941) );
  AOI22_X1 U3745 ( .A1(n4372), .A2(n2942), .B1(n4370), .B2(n2941), .ZN(n2947)
         );
  INV_X1 U3746 ( .A(n2943), .ZN(n2945) );
  NOR2_X1 U3747 ( .A1(STATE_REG_SCAN_IN), .A2(n2338), .ZN(n3157) );
  AOI21_X1 U3748 ( .B1(n4345), .B2(ADDR_REG_3__SCAN_IN), .A(n3157), .ZN(n2946)
         );
  OAI211_X1 U3749 ( .C1(n2948), .C2(n4375), .A(n2947), .B(n2946), .ZN(U3243)
         );
  INV_X1 U3750 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U3751 ( .A1(n3364), .A2(U4043), .ZN(n2949) );
  OAI21_X1 U3752 ( .B1(U4043), .B2(n4584), .A(n2949), .ZN(U3561) );
  INV_X1 U3753 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4545) );
  MUX2_X1 U3754 ( .A(n4545), .B(REG1_REG_7__SCAN_IN), .S(n3007), .Z(n2961) );
  NAND2_X1 U3755 ( .A1(n2951), .A2(n4274), .ZN(n2952) );
  NAND2_X1 U3756 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  INV_X1 U3757 ( .A(n4273), .ZN(n2968) );
  XNOR2_X1 U3758 ( .A(n2954), .B(n2968), .ZN(n3834) );
  NAND2_X1 U3759 ( .A1(n3834), .A2(REG1_REG_4__SCAN_IN), .ZN(n2956) );
  NAND2_X1 U3760 ( .A1(n2954), .A2(n4273), .ZN(n2955) );
  NAND2_X1 U3761 ( .A1(n2956), .A2(n2955), .ZN(n3848) );
  MUX2_X1 U3762 ( .A(n4541), .B(REG1_REG_5__SCAN_IN), .S(n3844), .Z(n3849) );
  NAND2_X1 U3763 ( .A1(n3848), .A2(n3849), .ZN(n3847) );
  INV_X1 U3764 ( .A(n3844), .ZN(n4272) );
  NAND2_X1 U3765 ( .A1(n4272), .A2(REG1_REG_5__SCAN_IN), .ZN(n2957) );
  NAND2_X1 U3766 ( .A1(n3847), .A2(n2957), .ZN(n2958) );
  INV_X1 U3767 ( .A(n4271), .ZN(n2987) );
  XNOR2_X1 U3768 ( .A(n2958), .B(n2987), .ZN(n2984) );
  NAND2_X1 U3769 ( .A1(n2984), .A2(REG1_REG_6__SCAN_IN), .ZN(n2960) );
  NAND2_X1 U3770 ( .A1(n2958), .A2(n4271), .ZN(n2959) );
  XOR2_X1 U3771 ( .A(n2961), .B(n3006), .Z(n2983) );
  AND2_X1 U3772 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3267) );
  NOR2_X1 U3773 ( .A1(n4375), .A2(n2962), .ZN(n2963) );
  AOI211_X1 U3774 ( .C1(n4345), .C2(ADDR_REG_7__SCAN_IN), .A(n3267), .B(n2963), 
        .ZN(n2982) );
  NAND2_X1 U3775 ( .A1(n2964), .A2(REG2_REG_3__SCAN_IN), .ZN(n2967) );
  NAND2_X1 U3776 ( .A1(n2965), .A2(n4274), .ZN(n2966) );
  NAND2_X1 U3777 ( .A1(n2967), .A2(n2966), .ZN(n2969) );
  XNOR2_X1 U3778 ( .A(n2969), .B(n2968), .ZN(n3835) );
  NAND2_X1 U3779 ( .A1(n3835), .A2(REG2_REG_4__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3780 ( .A1(n2969), .A2(n4273), .ZN(n2970) );
  NAND2_X1 U3781 ( .A1(n2971), .A2(n2970), .ZN(n3851) );
  INV_X1 U3782 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3167) );
  MUX2_X1 U3783 ( .A(n3167), .B(REG2_REG_5__SCAN_IN), .S(n3844), .Z(n3852) );
  NAND2_X1 U3784 ( .A1(n3851), .A2(n3852), .ZN(n3850) );
  NAND2_X1 U3785 ( .A1(n4272), .A2(REG2_REG_5__SCAN_IN), .ZN(n2972) );
  NAND2_X1 U3786 ( .A1(n3850), .A2(n2972), .ZN(n2973) );
  XNOR2_X1 U3787 ( .A(n2973), .B(n2987), .ZN(n2985) );
  NAND2_X1 U3788 ( .A1(n2985), .A2(REG2_REG_6__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3789 ( .A1(n2973), .A2(n4271), .ZN(n2974) );
  NAND2_X1 U3790 ( .A1(n2975), .A2(n2974), .ZN(n2980) );
  MUX2_X1 U3791 ( .A(n2977), .B(REG2_REG_7__SCAN_IN), .S(n3007), .Z(n2976) );
  INV_X1 U3792 ( .A(n2976), .ZN(n2979) );
  INV_X1 U3793 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2977) );
  MUX2_X1 U3794 ( .A(REG2_REG_7__SCAN_IN), .B(n2977), .S(n3007), .Z(n2978) );
  NAND2_X1 U3795 ( .A1(n2980), .A2(n2978), .ZN(n2999) );
  OAI211_X1 U3796 ( .C1(n2980), .C2(n2979), .A(n2999), .B(n4370), .ZN(n2981)
         );
  OAI211_X1 U3797 ( .C1(n2983), .C2(n4339), .A(n2982), .B(n2981), .ZN(U3247)
         );
  XNOR2_X1 U3798 ( .A(n2984), .B(REG1_REG_6__SCAN_IN), .ZN(n2991) );
  XOR2_X1 U3799 ( .A(REG2_REG_6__SCAN_IN), .B(n2985), .Z(n2989) );
  AND2_X1 U3800 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3210) );
  AOI21_X1 U3801 ( .B1(n4345), .B2(ADDR_REG_6__SCAN_IN), .A(n3210), .ZN(n2986)
         );
  OAI21_X1 U3802 ( .B1(n2987), .B2(n4375), .A(n2986), .ZN(n2988) );
  AOI21_X1 U3803 ( .B1(n4370), .B2(n2989), .A(n2988), .ZN(n2990) );
  OAI21_X1 U3804 ( .B1(n2991), .B2(n4339), .A(n2990), .ZN(U3246) );
  INV_X1 U3805 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U3806 ( .A1(n4001), .A2(U4043), .ZN(n2992) );
  OAI21_X1 U3807 ( .B1(U4043), .B2(n4590), .A(n2992), .ZN(U3574) );
  NOR2_X1 U3808 ( .A1(n4345), .A2(U4043), .ZN(U3148) );
  AND2_X1 U3809 ( .A1(n3805), .A2(n3109), .ZN(n3716) );
  OR2_X1 U3810 ( .A1(n3716), .A2(n3719), .ZN(n4382) );
  NAND2_X1 U3811 ( .A1(n4057), .A2(n4123), .ZN(n2994) );
  AND2_X1 U3812 ( .A1(n2784), .A2(n4101), .ZN(n2993) );
  AOI21_X1 U3813 ( .B1(n4382), .B2(n2994), .A(n2993), .ZN(n4377) );
  INV_X1 U3814 ( .A(n4435), .ZN(n4414) );
  AND2_X1 U3815 ( .A1(n3040), .A2(n2995), .ZN(n4380) );
  AOI21_X1 U3816 ( .B1(n4382), .B2(n4414), .A(n4380), .ZN(n2996) );
  AND2_X1 U3817 ( .A1(n4377), .A2(n2996), .ZN(n4403) );
  NAND2_X1 U3818 ( .A1(n4451), .A2(REG1_REG_0__SCAN_IN), .ZN(n2997) );
  OAI21_X1 U3819 ( .B1(n4403), .B2(n4451), .A(n2997), .ZN(U3518) );
  NAND2_X1 U3820 ( .A1(n3007), .A2(REG2_REG_7__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3821 ( .A1(n2999), .A2(n2998), .ZN(n3000) );
  XNOR2_X1 U3822 ( .A(n3000), .B(n3021), .ZN(n3018) );
  INV_X1 U3823 ( .A(n3021), .ZN(n3010) );
  AND2_X1 U3824 ( .A1(n3000), .A2(n3010), .ZN(n3001) );
  AOI21_X1 U3825 ( .B1(n3018), .B2(REG2_REG_8__SCAN_IN), .A(n3001), .ZN(n3003)
         );
  INV_X1 U3826 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3283) );
  MUX2_X1 U3827 ( .A(REG2_REG_9__SCAN_IN), .B(n3283), .S(n3087), .Z(n3002) );
  AOI211_X1 U3828 ( .C1(n3003), .C2(n3002), .A(n4325), .B(n3086), .ZN(n3004)
         );
  INV_X1 U3829 ( .A(n3004), .ZN(n3017) );
  AND2_X1 U3830 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3298) );
  AND2_X1 U3831 ( .A1(n3007), .A2(REG1_REG_7__SCAN_IN), .ZN(n3005) );
  OR2_X1 U3832 ( .A1(n3007), .A2(REG1_REG_7__SCAN_IN), .ZN(n3008) );
  INV_X1 U3833 ( .A(n3009), .ZN(n3011) );
  INV_X1 U3834 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4544) );
  INV_X1 U3835 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3012) );
  MUX2_X1 U3836 ( .A(REG1_REG_9__SCAN_IN), .B(n3012), .S(n3087), .Z(n3013) );
  AOI211_X1 U3837 ( .C1(n3014), .C2(n3013), .A(n3094), .B(n4339), .ZN(n3015)
         );
  AOI211_X1 U3838 ( .C1(n4345), .C2(ADDR_REG_9__SCAN_IN), .A(n3298), .B(n3015), 
        .ZN(n3016) );
  OAI211_X1 U3839 ( .C1(n4375), .C2(n3087), .A(n3017), .B(n3016), .ZN(U3249)
         );
  XOR2_X1 U3840 ( .A(REG2_REG_8__SCAN_IN), .B(n3018), .Z(n3026) );
  NAND2_X1 U3841 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3254) );
  INV_X1 U3842 ( .A(n3254), .ZN(n3019) );
  AOI21_X1 U3843 ( .B1(n4345), .B2(ADDR_REG_8__SCAN_IN), .A(n3019), .ZN(n3020)
         );
  OAI21_X1 U3844 ( .B1(n3021), .B2(n4375), .A(n3020), .ZN(n3025) );
  AOI211_X1 U3845 ( .C1(n4544), .C2(n3023), .A(n4339), .B(n3022), .ZN(n3024)
         );
  AOI211_X1 U3846 ( .C1(n4370), .C2(n3026), .A(n3025), .B(n3024), .ZN(n3027)
         );
  INV_X1 U3847 ( .A(n3027), .ZN(U3248) );
  INV_X1 U3848 ( .A(n3028), .ZN(n3031) );
  NAND3_X1 U3849 ( .A1(n3031), .A2(n3030), .A3(n3029), .ZN(n3119) );
  INV_X1 U3850 ( .A(n3119), .ZN(n3039) );
  INV_X1 U3851 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3122) );
  INV_X1 U3852 ( .A(n3805), .ZN(n3032) );
  OAI22_X1 U3853 ( .A1(n3032), .A2(n3625), .B1(n3613), .B2(n3077), .ZN(n3033)
         );
  AOI21_X1 U3854 ( .B1(n3552), .B2(n2286), .A(n3033), .ZN(n3038) );
  OAI211_X1 U3855 ( .C1(n3034), .C2(n3036), .A(n3035), .B(n3623), .ZN(n3037)
         );
  OAI211_X1 U3856 ( .C1(n3039), .C2(n3122), .A(n3038), .B(n3037), .ZN(U3219)
         );
  AOI21_X1 U3857 ( .B1(n3040), .B2(n2286), .A(n3064), .ZN(n3127) );
  OAI21_X1 U3858 ( .B1(n3043), .B2(n3042), .A(n3041), .ZN(n3123) );
  NOR2_X1 U3859 ( .A1(n3123), .A2(n4435), .ZN(n3051) );
  OAI21_X1 U3860 ( .B1(n3705), .B2(n3719), .A(n3055), .ZN(n3044) );
  NAND2_X1 U3861 ( .A1(n3044), .A2(n4107), .ZN(n3050) );
  NAND2_X1 U3862 ( .A1(n3805), .A2(n4121), .ZN(n3046) );
  NAND2_X1 U3863 ( .A1(n3158), .A2(n4101), .ZN(n3045) );
  OAI211_X1 U3864 ( .C1(n4147), .C2(n3047), .A(n3046), .B(n3045), .ZN(n3048)
         );
  INV_X1 U3865 ( .A(n3048), .ZN(n3049) );
  OAI211_X1 U3866 ( .C1(n3123), .C2(n4057), .A(n3050), .B(n3049), .ZN(n3124)
         );
  AOI211_X1 U3867 ( .C1(n4440), .C2(n3127), .A(n3051), .B(n3124), .ZN(n4404)
         );
  NAND2_X1 U3868 ( .A1(n4451), .A2(REG1_REG_1__SCAN_IN), .ZN(n3052) );
  OAI21_X1 U3869 ( .B1(n4404), .B2(n4451), .A(n3052), .ZN(U3519) );
  OAI21_X1 U3870 ( .B1(n3054), .B2(n2832), .A(n3053), .ZN(n3142) );
  NAND3_X1 U3871 ( .A1(n3055), .A2(n2832), .A3(n2831), .ZN(n3056) );
  NAND2_X1 U3872 ( .A1(n3057), .A2(n3056), .ZN(n3061) );
  NAND2_X1 U3873 ( .A1(n2784), .A2(n4121), .ZN(n3059) );
  NAND2_X1 U3874 ( .A1(n3149), .A2(n4101), .ZN(n3058) );
  OAI211_X1 U3875 ( .C1(n4147), .C2(n3116), .A(n3059), .B(n3058), .ZN(n3060)
         );
  AOI21_X1 U3876 ( .B1(n3061), .B2(n4107), .A(n3060), .ZN(n3063) );
  INV_X1 U3877 ( .A(n4057), .ZN(n3337) );
  NAND2_X1 U3878 ( .A1(n3142), .A2(n3337), .ZN(n3062) );
  NAND2_X1 U3879 ( .A1(n3063), .A2(n3062), .ZN(n3139) );
  AOI21_X1 U3880 ( .B1(n4414), .B2(n3142), .A(n3139), .ZN(n3070) );
  OAI21_X1 U3881 ( .B1(n3064), .B2(n3116), .A(n3081), .ZN(n3138) );
  INV_X1 U3882 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3065) );
  OAI22_X1 U3883 ( .A1(n4263), .A2(n3138), .B1(n4443), .B2(n3065), .ZN(n3066)
         );
  INV_X1 U3884 ( .A(n3066), .ZN(n3067) );
  OAI21_X1 U3885 ( .B1(n3070), .B2(n4441), .A(n3067), .ZN(U3471) );
  INV_X1 U3886 ( .A(n4214), .ZN(n4137) );
  INV_X1 U3887 ( .A(n3138), .ZN(n3068) );
  AOI22_X1 U3888 ( .A1(n4137), .A2(n3068), .B1(REG1_REG_2__SCAN_IN), .B2(n4451), .ZN(n3069) );
  OAI21_X1 U3889 ( .B1(n3070), .B2(n4451), .A(n3069), .ZN(U3520) );
  XNOR2_X1 U3890 ( .A(n3071), .B(n3697), .ZN(n4405) );
  INV_X1 U3891 ( .A(n3072), .ZN(n3073) );
  INV_X1 U3892 ( .A(n4383), .ZN(n3416) );
  OAI21_X1 U3893 ( .B1(n3697), .B2(n3075), .A(n3074), .ZN(n3079) );
  AOI22_X1 U3894 ( .A1(n3804), .A2(n4101), .B1(n4099), .B2(n3082), .ZN(n3076)
         );
  OAI21_X1 U3895 ( .B1(n3077), .B2(n4104), .A(n3076), .ZN(n3078) );
  AOI21_X1 U3896 ( .B1(n3079), .B2(n4107), .A(n3078), .ZN(n3080) );
  OAI21_X1 U3897 ( .B1(n4405), .B2(n4057), .A(n3080), .ZN(n4406) );
  NAND2_X1 U3898 ( .A1(n4406), .A2(n4278), .ZN(n3085) );
  AOI21_X1 U3899 ( .B1(n3082), .B2(n3081), .A(n3199), .ZN(n4408) );
  OAI22_X1 U3900 ( .A1(n4278), .A2(n2339), .B1(n4129), .B2(REG3_REG_3__SCAN_IN), .ZN(n3083) );
  AOI21_X1 U3901 ( .B1(n4408), .B2(n4282), .A(n3083), .ZN(n3084) );
  OAI211_X1 U3902 ( .C1(n4405), .C2(n3416), .A(n3085), .B(n3084), .ZN(U3287)
         );
  INV_X1 U3903 ( .A(n3872), .ZN(n3106) );
  NAND2_X1 U3904 ( .A1(n4399), .A2(n3088), .ZN(n3089) );
  NAND2_X1 U3905 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4300), .ZN(n4299) );
  NAND2_X1 U3906 ( .A1(n3089), .A2(n4299), .ZN(n3093) );
  INV_X1 U3907 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3908 ( .A1(n3872), .A2(REG2_REG_11__SCAN_IN), .ZN(n3858) );
  INV_X1 U3909 ( .A(n3858), .ZN(n3090) );
  AOI21_X1 U3910 ( .B1(n3091), .B2(n3106), .A(n3090), .ZN(n3092) );
  NAND2_X1 U3911 ( .A1(n3092), .A2(n3093), .ZN(n3857) );
  OAI211_X1 U3912 ( .C1(n3093), .C2(n3092), .A(n4370), .B(n3857), .ZN(n3105)
         );
  INV_X1 U3913 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4591) );
  NOR2_X1 U3914 ( .A1(STATE_REG_SCAN_IN), .A2(n4591), .ZN(n3360) );
  NOR2_X1 U3915 ( .A1(n3096), .A2(n4303), .ZN(n3097) );
  INV_X1 U3916 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4296) );
  XNOR2_X1 U3917 ( .A(n4303), .B(n3096), .ZN(n4295) );
  NOR2_X1 U3918 ( .A1(n4296), .A2(n4295), .ZN(n4294) );
  INV_X1 U3919 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3098) );
  OR2_X1 U3920 ( .A1(n3872), .A2(n3098), .ZN(n3100) );
  NAND2_X1 U3921 ( .A1(n3872), .A2(n3098), .ZN(n3099) );
  AND2_X1 U3922 ( .A1(n3100), .A2(n3099), .ZN(n3101) );
  AOI211_X1 U3923 ( .C1(n3102), .C2(n3101), .A(n3871), .B(n4339), .ZN(n3103)
         );
  AOI211_X1 U3924 ( .C1(n4345), .C2(ADDR_REG_11__SCAN_IN), .A(n3360), .B(n3103), .ZN(n3104) );
  OAI211_X1 U3925 ( .C1(n4375), .C2(n3106), .A(n3105), .B(n3104), .ZN(U3251)
         );
  XNOR2_X1 U3926 ( .A(n3108), .B(n3107), .ZN(n3817) );
  OAI22_X1 U3927 ( .A1(n2005), .A2(n3109), .B1(n2783), .B2(n3613), .ZN(n3110)
         );
  AOI21_X1 U3928 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3119), .A(n3110), .ZN(n3111)
         );
  OAI21_X1 U3929 ( .B1(n3618), .B2(n3817), .A(n3111), .ZN(U3229) );
  INV_X1 U3930 ( .A(n3113), .ZN(n3114) );
  AOI21_X1 U3931 ( .B1(n3112), .B2(n3115), .A(n3114), .ZN(n3121) );
  OAI22_X1 U3932 ( .A1(n3192), .A2(n3613), .B1(n3625), .B2(n2783), .ZN(n3118)
         );
  NOR2_X1 U3933 ( .A1(n2005), .A2(n3116), .ZN(n3117) );
  AOI211_X1 U3934 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3119), .A(n3118), .B(n3117), 
        .ZN(n3120) );
  OAI21_X1 U3935 ( .B1(n3121), .B2(n3618), .A(n3120), .ZN(U3234) );
  OAI22_X1 U3936 ( .A1(n3416), .A2(n3123), .B1(n3122), .B2(n4129), .ZN(n3126)
         );
  MUX2_X1 U3937 ( .A(n3124), .B(REG2_REG_1__SCAN_IN), .S(n4063), .Z(n3125) );
  AOI211_X1 U3938 ( .C1(n4282), .C2(n3127), .A(n3126), .B(n3125), .ZN(n3128)
         );
  INV_X1 U3939 ( .A(n3128), .ZN(U3289) );
  INV_X1 U3940 ( .A(n3170), .ZN(n3136) );
  OAI211_X1 U3941 ( .C1(n3131), .C2(n3130), .A(n3129), .B(n3623), .ZN(n3135)
         );
  AND2_X1 U3942 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3846) );
  OAI22_X1 U3943 ( .A1(n2005), .A2(n3132), .B1(n3164), .B2(n3625), .ZN(n3133)
         );
  AOI211_X1 U3944 ( .C1(n3629), .C2(n3802), .A(n3846), .B(n3133), .ZN(n3134)
         );
  OAI211_X1 U3945 ( .C1(n3633), .C2(n3136), .A(n3135), .B(n3134), .ZN(U3224)
         );
  INV_X1 U3946 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3137) );
  OAI22_X1 U3947 ( .A1(n4127), .A2(n3138), .B1(n3137), .B2(n4129), .ZN(n3141)
         );
  MUX2_X1 U3948 ( .A(n3139), .B(REG2_REG_2__SCAN_IN), .S(n4063), .Z(n3140) );
  AOI211_X1 U3949 ( .C1(n4383), .C2(n3142), .A(n3141), .B(n3140), .ZN(n3143)
         );
  INV_X1 U3950 ( .A(n3143), .ZN(U3288) );
  AOI21_X1 U3951 ( .B1(n3144), .B2(n3145), .A(n3618), .ZN(n3147) );
  NAND2_X1 U3952 ( .A1(n3147), .A2(n3146), .ZN(n3151) );
  AND2_X1 U3953 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3836) );
  OAI22_X1 U3954 ( .A1(n2005), .A2(n3198), .B1(n3175), .B2(n3613), .ZN(n3148)
         );
  AOI211_X1 U3955 ( .C1(n3530), .C2(n3149), .A(n3836), .B(n3148), .ZN(n3150)
         );
  OAI211_X1 U3956 ( .C1(n3633), .C2(n3200), .A(n3151), .B(n3150), .ZN(U3227)
         );
  XNOR2_X1 U3957 ( .A(n3153), .B(n3152), .ZN(n3154) );
  NAND2_X1 U3958 ( .A1(n3154), .A2(n3623), .ZN(n3160) );
  OAI22_X1 U3959 ( .A1(n2005), .A2(n3155), .B1(n3164), .B2(n3613), .ZN(n3156)
         );
  AOI211_X1 U3960 ( .C1(n3530), .C2(n3158), .A(n3157), .B(n3156), .ZN(n3159)
         );
  OAI211_X1 U3961 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3633), .A(n3160), .B(n3159), 
        .ZN(U3215) );
  NAND2_X1 U3962 ( .A1(n3734), .A2(n3728), .ZN(n3685) );
  XNOR2_X1 U3963 ( .A(n3161), .B(n3685), .ZN(n4417) );
  XNOR2_X1 U3964 ( .A(n3162), .B(n3685), .ZN(n3166) );
  AOI22_X1 U3965 ( .A1(n3802), .A2(n4101), .B1(n3169), .B2(n4099), .ZN(n3163)
         );
  OAI21_X1 U3966 ( .B1(n3164), .B2(n4104), .A(n3163), .ZN(n3165) );
  AOI21_X1 U3967 ( .B1(n3166), .B2(n4107), .A(n3165), .ZN(n4418) );
  MUX2_X1 U3968 ( .A(n4418), .B(n3167), .S(n4063), .Z(n3172) );
  INV_X1 U3969 ( .A(n3180), .ZN(n3168) );
  AOI21_X1 U3970 ( .B1(n3169), .B2(n3197), .A(n3168), .ZN(n4421) );
  AOI22_X1 U3971 ( .A1(n4421), .A2(n4282), .B1(n3170), .B2(n4381), .ZN(n3171)
         );
  OAI211_X1 U3972 ( .C1(n4135), .C2(n4417), .A(n3172), .B(n3171), .ZN(U3285)
         );
  INV_X1 U3973 ( .A(n3735), .ZN(n3729) );
  AND2_X1 U3974 ( .A1(n3729), .A2(n3732), .ZN(n3692) );
  XOR2_X1 U3975 ( .A(n3692), .B(n3173), .Z(n3177) );
  AOI22_X1 U3976 ( .A1(n3801), .A2(n4101), .B1(n4099), .B2(n3179), .ZN(n3174)
         );
  OAI21_X1 U3977 ( .B1(n3175), .B2(n4104), .A(n3174), .ZN(n3176) );
  AOI21_X1 U3978 ( .B1(n3177), .B2(n4107), .A(n3176), .ZN(n3215) );
  XOR2_X1 U3979 ( .A(n3178), .B(n3692), .Z(n3216) );
  INV_X1 U3980 ( .A(n3216), .ZN(n3185) );
  AND2_X1 U3981 ( .A1(n3180), .A2(n3179), .ZN(n3181) );
  NOR2_X1 U3982 ( .A1(n3229), .A2(n3181), .ZN(n3220) );
  INV_X1 U3983 ( .A(n3220), .ZN(n3183) );
  AOI22_X1 U3984 ( .A1(n4063), .A2(REG2_REG_6__SCAN_IN), .B1(n3211), .B2(n4381), .ZN(n3182) );
  OAI21_X1 U3985 ( .B1(n3183), .B2(n4127), .A(n3182), .ZN(n3184) );
  AOI21_X1 U3986 ( .B1(n3185), .B2(n4037), .A(n3184), .ZN(n3186) );
  OAI21_X1 U3987 ( .B1(n4063), .B2(n3215), .A(n3186), .ZN(U3284) );
  INV_X1 U3988 ( .A(n3189), .ZN(n3698) );
  NAND2_X1 U3989 ( .A1(n3188), .A2(n3698), .ZN(n3190) );
  NAND2_X1 U3990 ( .A1(n3187), .A2(n3190), .ZN(n4410) );
  XOR2_X1 U3991 ( .A(n3698), .B(n3191), .Z(n3196) );
  OAI22_X1 U3992 ( .A1(n3192), .A2(n4104), .B1(n3198), .B2(n4147), .ZN(n3194)
         );
  NOR2_X1 U3993 ( .A1(n4410), .A2(n4057), .ZN(n3193) );
  AOI211_X1 U3994 ( .C1(n4101), .C2(n3803), .A(n3194), .B(n3193), .ZN(n3195)
         );
  OAI21_X1 U3995 ( .B1(n4123), .B2(n3196), .A(n3195), .ZN(n4412) );
  OAI211_X1 U3996 ( .C1(n3199), .C2(n3198), .A(n3197), .B(n4440), .ZN(n4411)
         );
  OAI22_X1 U3997 ( .A1(n4411), .A2(n3887), .B1(n4129), .B2(n3200), .ZN(n3201)
         );
  OAI21_X1 U3998 ( .B1(n4412), .B2(n3201), .A(n4278), .ZN(n3203) );
  NAND2_X1 U3999 ( .A1(n4063), .A2(REG2_REG_4__SCAN_IN), .ZN(n3202) );
  OAI211_X1 U4000 ( .C1(n4410), .C2(n3416), .A(n3203), .B(n3202), .ZN(U3286)
         );
  XOR2_X1 U4001 ( .A(n3205), .B(n3204), .Z(n3206) );
  XNOR2_X1 U4002 ( .A(n3207), .B(n3206), .ZN(n3214) );
  OAI22_X1 U4003 ( .A1(n2005), .A2(n3208), .B1(n3256), .B2(n3613), .ZN(n3209)
         );
  AOI211_X1 U4004 ( .C1(n3530), .C2(n3803), .A(n3210), .B(n3209), .ZN(n3213)
         );
  NAND2_X1 U4005 ( .A1(n3616), .A2(n3211), .ZN(n3212) );
  OAI211_X1 U4006 ( .C1(n3214), .C2(n3618), .A(n3213), .B(n3212), .ZN(U3236)
         );
  INV_X1 U4007 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4542) );
  OAI21_X1 U4008 ( .B1(n3216), .B2(n4422), .A(n3215), .ZN(n3219) );
  NAND2_X1 U4009 ( .A1(n3219), .A2(n4453), .ZN(n3218) );
  NAND2_X1 U4010 ( .A1(n3220), .A2(n4137), .ZN(n3217) );
  OAI211_X1 U4011 ( .C1(n4453), .C2(n4542), .A(n3218), .B(n3217), .ZN(U3524)
         );
  INV_X1 U4012 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4013 ( .A1(n3219), .A2(n4443), .ZN(n3222) );
  INV_X1 U4014 ( .A(n4263), .ZN(n4215) );
  NAND2_X1 U4015 ( .A1(n3220), .A2(n4215), .ZN(n3221) );
  OAI211_X1 U4016 ( .C1(n4443), .C2(n3223), .A(n3222), .B(n3221), .ZN(U3479)
         );
  XNOR2_X1 U4017 ( .A(n3224), .B(n3733), .ZN(n3225) );
  NAND2_X1 U4018 ( .A1(n3225), .A2(n4107), .ZN(n3228) );
  AOI22_X1 U4019 ( .A1(n3800), .A2(n4101), .B1(n3226), .B2(n4099), .ZN(n3227)
         );
  OAI211_X1 U4020 ( .C1(n3264), .C2(n4104), .A(n3228), .B(n3227), .ZN(n4424)
         );
  INV_X1 U4021 ( .A(n4424), .ZN(n3237) );
  OAI21_X1 U4022 ( .B1(n3229), .B2(n3265), .A(n4440), .ZN(n3230) );
  NOR2_X1 U4023 ( .A1(n3230), .A2(n3244), .ZN(n4425) );
  OAI22_X1 U4024 ( .A1(n4278), .A2(n2977), .B1(n3270), .B2(n4129), .ZN(n3235)
         );
  INV_X1 U4025 ( .A(n3231), .ZN(n3233) );
  AND2_X1 U4026 ( .A1(n3232), .A2(n3733), .ZN(n4423) );
  NOR3_X1 U4027 ( .A1(n3233), .A2(n4423), .A3(n4135), .ZN(n3234) );
  AOI211_X1 U4028 ( .C1(n4111), .C2(n4425), .A(n3235), .B(n3234), .ZN(n3236)
         );
  OAI21_X1 U4029 ( .B1(n4063), .B2(n3237), .A(n3236), .ZN(U3283) );
  AND2_X1 U4030 ( .A1(n3740), .A2(n3736), .ZN(n3682) );
  XNOR2_X1 U4031 ( .A(n3238), .B(n3682), .ZN(n3241) );
  OAI22_X1 U4032 ( .A1(n3368), .A2(n4117), .B1(n4147), .B2(n3243), .ZN(n3239)
         );
  AOI21_X1 U4033 ( .B1(n4121), .B2(n3801), .A(n3239), .ZN(n3240) );
  OAI21_X1 U4034 ( .B1(n3241), .B2(n4123), .A(n3240), .ZN(n3287) );
  INV_X1 U4035 ( .A(n3287), .ZN(n3249) );
  XNOR2_X1 U4036 ( .A(n3242), .B(n3682), .ZN(n3288) );
  OR2_X1 U4037 ( .A1(n3244), .A2(n3243), .ZN(n3245) );
  NAND2_X1 U4038 ( .A1(n3280), .A2(n3245), .ZN(n3293) );
  AOI22_X1 U4039 ( .A1(n4063), .A2(REG2_REG_8__SCAN_IN), .B1(n3258), .B2(n4381), .ZN(n3246) );
  OAI21_X1 U4040 ( .B1(n3293), .B2(n4127), .A(n3246), .ZN(n3247) );
  AOI21_X1 U4041 ( .B1(n3288), .B2(n4037), .A(n3247), .ZN(n3248) );
  OAI21_X1 U4042 ( .B1(n3249), .B2(n4063), .A(n3248), .ZN(U3282) );
  NOR2_X1 U40430 ( .A1(n2045), .A2(n3250), .ZN(n3251) );
  XNOR2_X1 U4044 ( .A(n3252), .B(n3251), .ZN(n3260) );
  AOI22_X1 U4045 ( .A1(n3552), .A2(n3253), .B1(n3629), .B2(n3799), .ZN(n3255)
         );
  OAI211_X1 U4046 ( .C1(n3256), .C2(n3625), .A(n3255), .B(n3254), .ZN(n3257)
         );
  AOI21_X1 U4047 ( .B1(n3258), .B2(n3616), .A(n3257), .ZN(n3259) );
  OAI21_X1 U4048 ( .B1(n3260), .B2(n3618), .A(n3259), .ZN(U3218) );
  XOR2_X1 U4049 ( .A(n3262), .B(n3261), .Z(n3263) );
  NAND2_X1 U4050 ( .A1(n3263), .A2(n3623), .ZN(n3269) );
  OAI22_X1 U4051 ( .A1(n2005), .A2(n3265), .B1(n3264), .B2(n3625), .ZN(n3266)
         );
  AOI211_X1 U4052 ( .C1(n3629), .C2(n3800), .A(n3267), .B(n3266), .ZN(n3268)
         );
  OAI211_X1 U4053 ( .C1(n3633), .C2(n3270), .A(n3269), .B(n3268), .ZN(U3210)
         );
  INV_X1 U4054 ( .A(n3744), .ZN(n3271) );
  AND2_X1 U4055 ( .A1(n3271), .A2(n3741), .ZN(n3684) );
  INV_X1 U4056 ( .A(n3684), .ZN(n3272) );
  XNOR2_X1 U4057 ( .A(n3273), .B(n3272), .ZN(n3277) );
  NAND2_X1 U4058 ( .A1(n3800), .A2(n4121), .ZN(n3275) );
  NAND2_X1 U4059 ( .A1(n3798), .A2(n4101), .ZN(n3274) );
  OAI211_X1 U4060 ( .C1(n4147), .C2(n3296), .A(n3275), .B(n3274), .ZN(n3276)
         );
  AOI21_X1 U4061 ( .B1(n3277), .B2(n4107), .A(n3276), .ZN(n4434) );
  XNOR2_X1 U4062 ( .A(n3278), .B(n3684), .ZN(n4429) );
  NAND2_X1 U4063 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  NAND2_X1 U4064 ( .A1(n3308), .A2(n3281), .ZN(n4431) );
  NOR2_X1 U4065 ( .A1(n4431), .A2(n4127), .ZN(n3285) );
  INV_X1 U4066 ( .A(n3299), .ZN(n3282) );
  OAI22_X1 U4067 ( .A1(n4278), .A2(n3283), .B1(n3282), .B2(n4129), .ZN(n3284)
         );
  AOI211_X1 U4068 ( .C1(n4429), .C2(n4037), .A(n3285), .B(n3284), .ZN(n3286)
         );
  OAI21_X1 U4069 ( .B1(n4434), .B2(n4063), .A(n3286), .ZN(U3281) );
  AOI21_X1 U4070 ( .B1(n3288), .B2(n4428), .A(n3287), .ZN(n3290) );
  MUX2_X1 U4071 ( .A(n4544), .B(n3290), .S(n4453), .Z(n3289) );
  OAI21_X1 U4072 ( .B1(n3293), .B2(n4214), .A(n3289), .ZN(U3526) );
  INV_X1 U4073 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3291) );
  MUX2_X1 U4074 ( .A(n3291), .B(n3290), .S(n4443), .Z(n3292) );
  OAI21_X1 U4075 ( .B1(n3293), .B2(n4263), .A(n3292), .ZN(U3483) );
  XOR2_X1 U4076 ( .A(n3294), .B(n3295), .Z(n3302) );
  OAI22_X1 U4077 ( .A1(n2005), .A2(n3296), .B1(n3335), .B2(n3613), .ZN(n3297)
         );
  AOI211_X1 U4078 ( .C1(n3530), .C2(n3800), .A(n3298), .B(n3297), .ZN(n3301)
         );
  NAND2_X1 U4079 ( .A1(n3616), .A2(n3299), .ZN(n3300) );
  OAI211_X1 U4080 ( .C1(n3302), .C2(n3618), .A(n3301), .B(n3300), .ZN(U3228)
         );
  AND2_X1 U4081 ( .A1(n3743), .A2(n3746), .ZN(n3687) );
  XOR2_X1 U4082 ( .A(n3687), .B(n3303), .Z(n3306) );
  OAI22_X1 U4083 ( .A1(n3389), .A2(n4117), .B1(n4147), .B2(n2136), .ZN(n3304)
         );
  AOI21_X1 U4084 ( .B1(n4121), .B2(n3799), .A(n3304), .ZN(n3305) );
  OAI21_X1 U4085 ( .B1(n3306), .B2(n4123), .A(n3305), .ZN(n3347) );
  INV_X1 U4086 ( .A(n3347), .ZN(n3314) );
  XOR2_X1 U4087 ( .A(n3307), .B(n3687), .Z(n3348) );
  OAI21_X1 U4088 ( .B1(n2137), .B2(n2136), .A(n3342), .ZN(n3352) );
  NOR2_X1 U4089 ( .A1(n3352), .A2(n4127), .ZN(n3312) );
  INV_X1 U4090 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3310) );
  INV_X1 U4091 ( .A(n3375), .ZN(n3309) );
  OAI22_X1 U4092 ( .A1(n4278), .A2(n3310), .B1(n3309), .B2(n4129), .ZN(n3311)
         );
  AOI211_X1 U4093 ( .C1(n3348), .C2(n4037), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OAI21_X1 U4094 ( .B1(n3314), .B2(n4063), .A(n3313), .ZN(U3280) );
  INV_X1 U4095 ( .A(n3315), .ZN(n3316) );
  AOI21_X1 U4096 ( .B1(n3333), .B2(n3317), .A(n3316), .ZN(n3401) );
  AND2_X1 U4097 ( .A1(n3400), .A2(n3398), .ZN(n3688) );
  INV_X1 U4098 ( .A(n3688), .ZN(n3323) );
  XNOR2_X1 U4099 ( .A(n3401), .B(n3323), .ZN(n3321) );
  OR2_X1 U4100 ( .A1(n3491), .A2(n4117), .ZN(n3319) );
  NAND2_X1 U4101 ( .A1(n3387), .A2(n4099), .ZN(n3318) );
  OAI211_X1 U4102 ( .C1(n3389), .C2(n4104), .A(n3319), .B(n3318), .ZN(n3320)
         );
  AOI21_X1 U4103 ( .B1(n3321), .B2(n4107), .A(n3320), .ZN(n3379) );
  XNOR2_X1 U4104 ( .A(n3322), .B(n3323), .ZN(n3377) );
  OR2_X1 U4105 ( .A1(n3341), .A2(n3324), .ZN(n3325) );
  NAND2_X1 U4106 ( .A1(n3408), .A2(n3325), .ZN(n3396) );
  INV_X1 U4107 ( .A(n3326), .ZN(n3391) );
  AOI22_X1 U4108 ( .A1(n4063), .A2(REG2_REG_12__SCAN_IN), .B1(n3391), .B2(
        n4381), .ZN(n3327) );
  OAI21_X1 U4109 ( .B1(n3396), .B2(n4127), .A(n3327), .ZN(n3328) );
  AOI21_X1 U4110 ( .B1(n3377), .B2(n4037), .A(n3328), .ZN(n3329) );
  OAI21_X1 U4111 ( .B1(n3379), .B2(n4063), .A(n3329), .ZN(U3278) );
  NAND2_X1 U4112 ( .A1(n3330), .A2(n3683), .ZN(n3331) );
  NAND2_X1 U4113 ( .A1(n3332), .A2(n3331), .ZN(n3338) );
  INV_X1 U4114 ( .A(n3338), .ZN(n4436) );
  XOR2_X1 U4115 ( .A(n3683), .B(n3333), .Z(n3340) );
  AOI22_X1 U4116 ( .A1(n3797), .A2(n4101), .B1(n3343), .B2(n4099), .ZN(n3334)
         );
  OAI21_X1 U4117 ( .B1(n3335), .B2(n4104), .A(n3334), .ZN(n3336) );
  AOI21_X1 U4118 ( .B1(n3338), .B2(n3337), .A(n3336), .ZN(n3339) );
  OAI21_X1 U4119 ( .B1(n3340), .B2(n4123), .A(n3339), .ZN(n4437) );
  NAND2_X1 U4120 ( .A1(n4437), .A2(n4278), .ZN(n3346) );
  AOI21_X1 U4121 ( .B1(n3343), .B2(n3342), .A(n3341), .ZN(n4439) );
  OAI22_X1 U4122 ( .A1(n4278), .A2(n3091), .B1(n3363), .B2(n4129), .ZN(n3344)
         );
  AOI21_X1 U4123 ( .B1(n4439), .B2(n4282), .A(n3344), .ZN(n3345) );
  OAI211_X1 U4124 ( .C1(n4436), .C2(n3416), .A(n3346), .B(n3345), .ZN(U3279)
         );
  INV_X1 U4125 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4528) );
  AOI21_X1 U4126 ( .B1(n4428), .B2(n3348), .A(n3347), .ZN(n3350) );
  MUX2_X1 U4127 ( .A(n4528), .B(n3350), .S(n4443), .Z(n3349) );
  OAI21_X1 U4128 ( .B1(n3352), .B2(n4263), .A(n3349), .ZN(U3487) );
  MUX2_X1 U4129 ( .A(n4296), .B(n3350), .S(n4453), .Z(n3351) );
  OAI21_X1 U4130 ( .B1(n3352), .B2(n4214), .A(n3351), .ZN(U3528) );
  XNOR2_X1 U4131 ( .A(n3355), .B(n3354), .ZN(n3356) );
  XNOR2_X1 U4132 ( .A(n3353), .B(n3356), .ZN(n3357) );
  NAND2_X1 U4133 ( .A1(n3357), .A2(n3623), .ZN(n3362) );
  OAI22_X1 U4134 ( .A1(n2005), .A2(n3358), .B1(n3422), .B2(n3613), .ZN(n3359)
         );
  AOI211_X1 U4135 ( .C1(n3530), .C2(n3798), .A(n3360), .B(n3359), .ZN(n3361)
         );
  OAI211_X1 U4136 ( .C1(n3633), .C2(n3363), .A(n3362), .B(n3361), .ZN(U3233)
         );
  AOI22_X1 U4137 ( .A1(n3552), .A2(n3365), .B1(n3629), .B2(n3364), .ZN(n3367)
         );
  NOR2_X1 U4138 ( .A1(n4495), .A2(STATE_REG_SCAN_IN), .ZN(n4297) );
  INV_X1 U4139 ( .A(n4297), .ZN(n3366) );
  OAI211_X1 U4140 ( .C1(n3368), .C2(n3625), .A(n3367), .B(n3366), .ZN(n3374)
         );
  INV_X1 U4141 ( .A(n3370), .ZN(n3371) );
  AOI211_X1 U4142 ( .C1(n3372), .C2(n3369), .A(n3618), .B(n3371), .ZN(n3373)
         );
  AOI211_X1 U4143 ( .C1(n3375), .C2(n3616), .A(n3374), .B(n3373), .ZN(n3376)
         );
  INV_X1 U4144 ( .A(n3376), .ZN(U3214) );
  NAND2_X1 U4145 ( .A1(n3377), .A2(n4428), .ZN(n3378) );
  AND2_X1 U4146 ( .A1(n3379), .A2(n3378), .ZN(n3394) );
  INV_X1 U4147 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3380) );
  MUX2_X1 U4148 ( .A(n3394), .B(n3380), .S(n4441), .Z(n3381) );
  OAI21_X1 U4149 ( .B1(n3396), .B2(n4263), .A(n3381), .ZN(U3491) );
  INV_X1 U4150 ( .A(n3382), .ZN(n3384) );
  NOR2_X1 U4151 ( .A1(n3384), .A2(n3383), .ZN(n3385) );
  XNOR2_X1 U4152 ( .A(n3386), .B(n3385), .ZN(n3393) );
  AOI22_X1 U4153 ( .A1(n3552), .A2(n3387), .B1(n3629), .B2(n3796), .ZN(n3388)
         );
  NAND2_X1 U4154 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4307) );
  OAI211_X1 U4155 ( .C1(n3389), .C2(n3625), .A(n3388), .B(n4307), .ZN(n3390)
         );
  AOI21_X1 U4156 ( .B1(n3391), .B2(n3616), .A(n3390), .ZN(n3392) );
  OAI21_X1 U4157 ( .B1(n3393), .B2(n3618), .A(n3392), .ZN(U3221) );
  INV_X1 U4158 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4306) );
  MUX2_X1 U4159 ( .A(n4306), .B(n3394), .S(n4453), .Z(n3395) );
  OAI21_X1 U4160 ( .B1(n3396), .B2(n4214), .A(n3395), .ZN(U3530) );
  XNOR2_X1 U4161 ( .A(n3491), .B(n3403), .ZN(n3677) );
  XOR2_X1 U4162 ( .A(n3677), .B(n3397), .Z(n3460) );
  INV_X1 U4163 ( .A(n3398), .ZN(n3399) );
  AOI21_X1 U4164 ( .B1(n3401), .B2(n3400), .A(n3399), .ZN(n3402) );
  XOR2_X1 U4165 ( .A(n3677), .B(n3402), .Z(n3406) );
  AOI22_X1 U4166 ( .A1(n3795), .A2(n4101), .B1(n4099), .B2(n3403), .ZN(n3404)
         );
  OAI21_X1 U4167 ( .B1(n3422), .B2(n4104), .A(n3404), .ZN(n3405) );
  AOI21_X1 U4168 ( .B1(n3406), .B2(n4107), .A(n3405), .ZN(n3407) );
  OAI21_X1 U4169 ( .B1(n3460), .B2(n4057), .A(n3407), .ZN(n3461) );
  NAND2_X1 U4170 ( .A1(n3461), .A2(n4278), .ZN(n3415) );
  INV_X1 U4171 ( .A(n3408), .ZN(n3409) );
  OAI21_X1 U4172 ( .B1(n3409), .B2(n3423), .A(n3450), .ZN(n3466) );
  INV_X1 U4173 ( .A(n3466), .ZN(n3413) );
  INV_X1 U4174 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3411) );
  INV_X1 U4175 ( .A(n3425), .ZN(n3410) );
  OAI22_X1 U4176 ( .A1(n4278), .A2(n3411), .B1(n3410), .B2(n4129), .ZN(n3412)
         );
  AOI21_X1 U4177 ( .B1(n3413), .B2(n4282), .A(n3412), .ZN(n3414) );
  OAI211_X1 U4178 ( .C1(n3460), .C2(n3416), .A(n3415), .B(n3414), .ZN(U3277)
         );
  XOR2_X1 U4179 ( .A(n3419), .B(n3418), .Z(n3420) );
  XNOR2_X1 U4180 ( .A(n3417), .B(n3420), .ZN(n3428) );
  NOR2_X1 U4181 ( .A1(STATE_REG_SCAN_IN), .A2(n3421), .ZN(n4317) );
  OAI22_X1 U4182 ( .A1(n2005), .A2(n3423), .B1(n3422), .B2(n3625), .ZN(n3424)
         );
  AOI211_X1 U4183 ( .C1(n3629), .C2(n3795), .A(n4317), .B(n3424), .ZN(n3427)
         );
  NAND2_X1 U4184 ( .A1(n3616), .A2(n3425), .ZN(n3426) );
  OAI211_X1 U4185 ( .C1(n3428), .C2(n3618), .A(n3427), .B(n3426), .ZN(U3231)
         );
  XNOR2_X1 U4186 ( .A(n3429), .B(n3703), .ZN(n4208) );
  INV_X1 U4187 ( .A(n4208), .ZN(n3440) );
  NAND2_X1 U4188 ( .A1(n3444), .A2(n3430), .ZN(n3431) );
  XNOR2_X1 U4189 ( .A(n3431), .B(n3703), .ZN(n3434) );
  OAI22_X1 U4190 ( .A1(n3563), .A2(n4117), .B1(n4147), .B2(n3627), .ZN(n3432)
         );
  AOI21_X1 U4191 ( .B1(n4121), .B2(n3795), .A(n3432), .ZN(n3433) );
  OAI21_X1 U4192 ( .B1(n3434), .B2(n4123), .A(n3433), .ZN(n4207) );
  NOR2_X1 U4193 ( .A1(n3451), .A2(n3627), .ZN(n3435) );
  OR2_X1 U4194 ( .A1(n3436), .A2(n3435), .ZN(n4259) );
  NOR2_X1 U4195 ( .A1(n4259), .A2(n4127), .ZN(n3438) );
  INV_X1 U4196 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3865) );
  OAI22_X1 U4197 ( .A1(n4278), .A2(n3865), .B1(n3632), .B2(n4129), .ZN(n3437)
         );
  AOI211_X1 U4198 ( .C1(n4207), .C2(n4278), .A(n3438), .B(n3437), .ZN(n3439)
         );
  OAI21_X1 U4199 ( .B1(n3440), .B2(n4135), .A(n3439), .ZN(U3275) );
  OAI21_X1 U4200 ( .B1(n3443), .B2(n3442), .A(n3441), .ZN(n4212) );
  INV_X1 U4201 ( .A(n4212), .ZN(n3449) );
  OAI21_X1 U4202 ( .B1(n3706), .B2(n3645), .A(n3444), .ZN(n3447) );
  AOI22_X1 U4203 ( .A1(n2807), .A2(n4101), .B1(n3489), .B2(n4099), .ZN(n3445)
         );
  OAI21_X1 U4204 ( .B1(n3491), .B2(n4104), .A(n3445), .ZN(n3446) );
  AOI21_X1 U4205 ( .B1(n3447), .B2(n4107), .A(n3446), .ZN(n3448) );
  OAI21_X1 U4206 ( .B1(n3449), .B2(n4057), .A(n3448), .ZN(n4211) );
  INV_X1 U4207 ( .A(n4211), .ZN(n3459) );
  INV_X1 U4208 ( .A(n3450), .ZN(n3454) );
  INV_X1 U4209 ( .A(n3451), .ZN(n3452) );
  OAI21_X1 U4210 ( .B1(n3454), .B2(n3453), .A(n3452), .ZN(n4264) );
  INV_X1 U4211 ( .A(n3455), .ZN(n3493) );
  AOI22_X1 U4212 ( .A1(n4063), .A2(REG2_REG_14__SCAN_IN), .B1(n3493), .B2(
        n4381), .ZN(n3456) );
  OAI21_X1 U4213 ( .B1(n4264), .B2(n4127), .A(n3456), .ZN(n3457) );
  AOI21_X1 U4214 ( .B1(n4212), .B2(n4383), .A(n3457), .ZN(n3458) );
  OAI21_X1 U4215 ( .B1(n3459), .B2(n4063), .A(n3458), .ZN(U3276) );
  INV_X1 U4216 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4548) );
  INV_X1 U4217 ( .A(n3460), .ZN(n3462) );
  AOI21_X1 U4218 ( .B1(n4414), .B2(n3462), .A(n3461), .ZN(n3464) );
  MUX2_X1 U4219 ( .A(n4548), .B(n3464), .S(n4453), .Z(n3463) );
  OAI21_X1 U4220 ( .B1(n4214), .B2(n3466), .A(n3463), .ZN(U3531) );
  INV_X1 U4221 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4527) );
  MUX2_X1 U4222 ( .A(n4527), .B(n3464), .S(n4443), .Z(n3465) );
  OAI21_X1 U4223 ( .B1(n3466), .B2(n4263), .A(n3465), .ZN(U3493) );
  INV_X1 U4224 ( .A(DATAI_29_), .ZN(n3469) );
  NAND2_X1 U4225 ( .A1(n3467), .A2(STATE_REG_SCAN_IN), .ZN(n3468) );
  OAI21_X1 U4226 ( .B1(STATE_REG_SCAN_IN), .B2(n3469), .A(n3468), .ZN(U3323)
         );
  INV_X1 U4227 ( .A(n3471), .ZN(n3477) );
  OAI22_X1 U4228 ( .A1(n3473), .A2(n4129), .B1(n3472), .B2(n4278), .ZN(n3476)
         );
  NOR2_X1 U4229 ( .A1(n3474), .A2(n4063), .ZN(n3475) );
  AOI211_X1 U4230 ( .C1(n4282), .C2(n3477), .A(n3476), .B(n3475), .ZN(n3478)
         );
  OAI21_X1 U4231 ( .B1(n3470), .B2(n4135), .A(n3478), .ZN(U3262) );
  INV_X1 U4232 ( .A(n3930), .ZN(n3483) );
  OAI22_X1 U4233 ( .A1(n3964), .A2(n3625), .B1(n2005), .B2(n3928), .ZN(n3482)
         );
  INV_X1 U4234 ( .A(n3924), .ZN(n3480) );
  OAI22_X1 U4235 ( .A1(n3480), .A2(n3613), .B1(STATE_REG_SCAN_IN), .B2(n4496), 
        .ZN(n3481) );
  AOI211_X1 U4236 ( .C1(n3483), .C2(n3616), .A(n3482), .B(n3481), .ZN(n3484)
         );
  OAI21_X1 U4237 ( .B1(n3485), .B2(n3618), .A(n3484), .ZN(U3211) );
  NAND2_X1 U4238 ( .A1(n2047), .A2(n3487), .ZN(n3488) );
  XNOR2_X1 U4239 ( .A(n3486), .B(n3488), .ZN(n3495) );
  AOI22_X1 U4240 ( .A1(n3552), .A2(n3489), .B1(n3629), .B2(n2807), .ZN(n3490)
         );
  NAND2_X1 U4241 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4336) );
  OAI211_X1 U4242 ( .C1(n3491), .C2(n3625), .A(n3490), .B(n4336), .ZN(n3492)
         );
  AOI21_X1 U4243 ( .B1(n3493), .B2(n3616), .A(n3492), .ZN(n3494) );
  OAI21_X1 U4244 ( .B1(n3495), .B2(n3618), .A(n3494), .ZN(U3212) );
  NAND2_X1 U4245 ( .A1(n3496), .A2(n3623), .ZN(n3506) );
  AOI21_X1 U4246 ( .B1(n3497), .B2(n3499), .A(n3498), .ZN(n3505) );
  INV_X1 U4247 ( .A(n4006), .ZN(n3503) );
  OAI22_X1 U4248 ( .A1(n3541), .A2(n3613), .B1(STATE_REG_SCAN_IN), .B2(n3500), 
        .ZN(n3502) );
  OAI22_X1 U4249 ( .A1(n2005), .A2(n4005), .B1(n4030), .B2(n3625), .ZN(n3501)
         );
  AOI211_X1 U4250 ( .C1(n3503), .C2(n3616), .A(n3502), .B(n3501), .ZN(n3504)
         );
  OAI21_X1 U4251 ( .B1(n3506), .B2(n3505), .A(n3504), .ZN(U3213) );
  INV_X1 U4252 ( .A(n3508), .ZN(n3598) );
  INV_X1 U4253 ( .A(n3507), .ZN(n3509) );
  OAI21_X1 U4254 ( .B1(n3509), .B2(n3508), .A(n3599), .ZN(n3510) );
  OAI21_X1 U4255 ( .B1(n3598), .B2(n3507), .A(n3510), .ZN(n3514) );
  NOR2_X1 U4256 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  XNOR2_X1 U4257 ( .A(n3514), .B(n3513), .ZN(n3520) );
  NOR2_X1 U4258 ( .A1(STATE_REG_SCAN_IN), .A2(n3515), .ZN(n3892) );
  OAI22_X1 U4259 ( .A1(n2005), .A2(n4083), .B1(n3516), .B2(n3613), .ZN(n3517)
         );
  AOI211_X1 U4260 ( .C1(n3530), .C2(n3565), .A(n3892), .B(n3517), .ZN(n3519)
         );
  NAND2_X1 U4261 ( .A1(n3616), .A2(n4084), .ZN(n3518) );
  OAI211_X1 U4262 ( .C1(n3520), .C2(n3618), .A(n3519), .B(n3518), .ZN(U3216)
         );
  INV_X1 U4263 ( .A(n3521), .ZN(n3523) );
  NOR2_X1 U4264 ( .A1(n3523), .A2(n3522), .ZN(n3527) );
  AOI211_X1 U4265 ( .C1(n3524), .C2(n2179), .A(n3579), .B(n3527), .ZN(n3526)
         );
  AOI211_X1 U4266 ( .C1(n2029), .C2(n3527), .A(n3618), .B(n3526), .ZN(n3535)
         );
  INV_X1 U4267 ( .A(n3528), .ZN(n4040) );
  AOI22_X1 U4268 ( .A1(n3629), .A2(n3529), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3533) );
  AOI22_X1 U4269 ( .A1(n3552), .A2(n3531), .B1(n3530), .B2(n4079), .ZN(n3532)
         );
  OAI211_X1 U4270 ( .C1(n3633), .C2(n4040), .A(n3533), .B(n3532), .ZN(n3534)
         );
  OR2_X1 U4271 ( .A1(n3535), .A2(n3534), .ZN(U3220) );
  INV_X1 U4272 ( .A(n3537), .ZN(n3539) );
  NAND2_X1 U4273 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  XNOR2_X1 U4274 ( .A(n3536), .B(n3540), .ZN(n3546) );
  OAI22_X1 U4275 ( .A1(n2005), .A2(n3967), .B1(n3541), .B2(n3625), .ZN(n3544)
         );
  INV_X1 U4276 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3542) );
  OAI22_X1 U4277 ( .A1(n3964), .A2(n3613), .B1(STATE_REG_SCAN_IN), .B2(n3542), 
        .ZN(n3543) );
  AOI211_X1 U4278 ( .C1(n3969), .C2(n3616), .A(n3544), .B(n3543), .ZN(n3545)
         );
  OAI21_X1 U4279 ( .B1(n3546), .B2(n3618), .A(n3545), .ZN(U3222) );
  OAI21_X1 U4280 ( .B1(n3547), .B2(n3621), .A(n2018), .ZN(n3549) );
  XNOR2_X1 U4281 ( .A(n3549), .B(n3548), .ZN(n3559) );
  INV_X1 U4282 ( .A(n3550), .ZN(n3557) );
  AOI22_X1 U4283 ( .A1(n3552), .A2(n3551), .B1(n3629), .B2(n3794), .ZN(n3554)
         );
  INV_X1 U4284 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4493) );
  NOR2_X1 U4285 ( .A1(n4493), .A2(STATE_REG_SCAN_IN), .ZN(n4353) );
  INV_X1 U4286 ( .A(n4353), .ZN(n3553) );
  OAI211_X1 U4287 ( .C1(n3555), .C2(n3625), .A(n3554), .B(n3553), .ZN(n3556)
         );
  AOI21_X1 U4288 ( .B1(n3557), .B2(n3616), .A(n3556), .ZN(n3558) );
  OAI21_X1 U4289 ( .B1(n3559), .B2(n3618), .A(n3558), .ZN(U3223) );
  NOR2_X1 U4290 ( .A1(n3560), .A2(n2044), .ZN(n3561) );
  XNOR2_X1 U4291 ( .A(n3562), .B(n3561), .ZN(n3568) );
  NOR2_X1 U4292 ( .A1(STATE_REG_SCAN_IN), .A2(n2572), .ZN(n4362) );
  OAI22_X1 U4293 ( .A1(n2005), .A2(n4126), .B1(n3563), .B2(n3625), .ZN(n3564)
         );
  AOI211_X1 U4294 ( .C1(n3629), .C2(n3565), .A(n4362), .B(n3564), .ZN(n3567)
         );
  NAND2_X1 U4295 ( .A1(n3616), .A2(n4128), .ZN(n3566) );
  OAI211_X1 U4296 ( .C1(n3568), .C2(n3618), .A(n3567), .B(n3566), .ZN(U3225)
         );
  INV_X1 U4297 ( .A(n3569), .ZN(n3570) );
  NOR2_X1 U4298 ( .A1(n3571), .A2(n3570), .ZN(n3573) );
  XNOR2_X1 U4299 ( .A(n3573), .B(n3572), .ZN(n3578) );
  INV_X1 U4300 ( .A(n3981), .ZN(n3610) );
  OAI22_X1 U4301 ( .A1(n3610), .A2(n3613), .B1(STATE_REG_SCAN_IN), .B2(n3574), 
        .ZN(n3576) );
  INV_X1 U4302 ( .A(n4022), .ZN(n3979) );
  OAI22_X1 U4303 ( .A1(n2005), .A2(n3985), .B1(n3979), .B2(n3625), .ZN(n3575)
         );
  AOI211_X1 U4304 ( .C1(n3987), .C2(n3616), .A(n3576), .B(n3575), .ZN(n3577)
         );
  OAI21_X1 U4305 ( .B1(n3578), .B2(n3618), .A(n3577), .ZN(U3226) );
  INV_X1 U4306 ( .A(n3579), .ZN(n3580) );
  NAND2_X1 U4307 ( .A1(n3580), .A2(n2179), .ZN(n3581) );
  AOI22_X1 U4308 ( .A1(n3582), .A2(n2179), .B1(n3524), .B2(n3581), .ZN(n3588)
         );
  INV_X1 U4309 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3583) );
  OAI22_X1 U4310 ( .A1(n3613), .A2(n3592), .B1(STATE_REG_SCAN_IN), .B2(n3583), 
        .ZN(n3586) );
  OAI22_X1 U4311 ( .A1(n2005), .A2(n3584), .B1(n4053), .B2(n3625), .ZN(n3585)
         );
  AOI211_X1 U4312 ( .C1(n4062), .C2(n3616), .A(n3586), .B(n3585), .ZN(n3587)
         );
  OAI21_X1 U4313 ( .B1(n3588), .B2(n3618), .A(n3587), .ZN(U3230) );
  OAI21_X1 U4314 ( .B1(n3590), .B2(n3589), .A(n3497), .ZN(n3591) );
  NAND2_X1 U4315 ( .A1(n3591), .A2(n3623), .ZN(n3597) );
  OAI22_X1 U4316 ( .A1(n2005), .A2(n4025), .B1(n3592), .B2(n3625), .ZN(n3595)
         );
  OAI22_X1 U4317 ( .A1(n3613), .A2(n3979), .B1(STATE_REG_SCAN_IN), .B2(n3593), 
        .ZN(n3594) );
  NOR2_X1 U4318 ( .A1(n3595), .A2(n3594), .ZN(n3596) );
  OAI211_X1 U4319 ( .C1(n3633), .C2(n4016), .A(n3597), .B(n3596), .ZN(U3232)
         );
  XNOR2_X1 U4320 ( .A(n3599), .B(n3598), .ZN(n3600) );
  XNOR2_X1 U4321 ( .A(n3507), .B(n3600), .ZN(n3601) );
  NAND2_X1 U4322 ( .A1(n3601), .A2(n3623), .ZN(n3604) );
  AND2_X1 U4323 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3884) );
  OAI22_X1 U4324 ( .A1(n2005), .A2(n2813), .B1(n4105), .B2(n3625), .ZN(n3602)
         );
  AOI211_X1 U4325 ( .C1(n3629), .C2(n4102), .A(n3884), .B(n3602), .ZN(n3603)
         );
  OAI211_X1 U4326 ( .C1(n3633), .C2(n4096), .A(n3604), .B(n3603), .ZN(U3235)
         );
  INV_X1 U4327 ( .A(n3605), .ZN(n3606) );
  NOR2_X1 U4328 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  XNOR2_X1 U4329 ( .A(n3609), .B(n3608), .ZN(n3619) );
  OAI22_X1 U4330 ( .A1(n2005), .A2(n3948), .B1(n3610), .B2(n3625), .ZN(n3615)
         );
  INV_X1 U4331 ( .A(n3942), .ZN(n3768) );
  OAI22_X1 U4332 ( .A1(n3768), .A2(n3613), .B1(STATE_REG_SCAN_IN), .B2(n3612), 
        .ZN(n3614) );
  AOI211_X1 U4333 ( .C1(n3949), .C2(n3616), .A(n3615), .B(n3614), .ZN(n3617)
         );
  OAI21_X1 U4334 ( .B1(n3619), .B2(n3618), .A(n3617), .ZN(U3237) );
  INV_X1 U4335 ( .A(n3547), .ZN(n3620) );
  NAND2_X1 U4336 ( .A1(n3620), .A2(n2018), .ZN(n3622) );
  XNOR2_X1 U4337 ( .A(n3622), .B(n3621), .ZN(n3624) );
  NAND2_X1 U4338 ( .A1(n3624), .A2(n3623), .ZN(n3631) );
  AND2_X1 U4339 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4344) );
  OAI22_X1 U4340 ( .A1(n2005), .A2(n3627), .B1(n3626), .B2(n3625), .ZN(n3628)
         );
  AOI211_X1 U4341 ( .C1(n3629), .C2(n4120), .A(n4344), .B(n3628), .ZN(n3630)
         );
  OAI211_X1 U4342 ( .C1(n3633), .C2(n3632), .A(n3631), .B(n3630), .ZN(U3238)
         );
  INV_X1 U4343 ( .A(n3634), .ZN(n3784) );
  NAND2_X1 U4344 ( .A1(n3642), .A2(DATAI_29_), .ZN(n3917) );
  NAND2_X1 U4345 ( .A1(n3792), .A2(n3917), .ZN(n3707) );
  NAND2_X1 U4346 ( .A1(n3707), .A2(n3635), .ZN(n3643) );
  NOR2_X1 U4347 ( .A1(n3701), .A2(n3643), .ZN(n3769) );
  NOR2_X1 U4348 ( .A1(n3900), .A2(n3636), .ZN(n3660) );
  INV_X1 U4349 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4350 ( .A1(n2340), .A2(REG1_REG_30__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4351 ( .A1(n2006), .A2(REG0_REG_30__SCAN_IN), .ZN(n3637) );
  OAI211_X1 U4352 ( .C1(n2319), .C2(n3639), .A(n3638), .B(n3637), .ZN(n3905)
         );
  NAND2_X1 U4353 ( .A1(n3642), .A2(DATAI_30_), .ZN(n4148) );
  OR2_X1 U4354 ( .A1(n3905), .A2(n4148), .ZN(n3669) );
  NAND2_X1 U4355 ( .A1(n2340), .A2(REG1_REG_31__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U4356 ( .A1(n2006), .A2(REG0_REG_31__SCAN_IN), .ZN(n3640) );
  OAI211_X1 U4357 ( .C1(n2319), .C2(n4566), .A(n3641), .B(n3640), .ZN(n4140)
         );
  NAND2_X1 U4358 ( .A1(n3642), .A2(DATAI_31_), .ZN(n4141) );
  NAND2_X1 U4359 ( .A1(n4140), .A2(n4141), .ZN(n3778) );
  AND2_X1 U4360 ( .A1(n3669), .A2(n3778), .ZN(n3661) );
  OR2_X1 U4361 ( .A1(n3792), .A2(n3917), .ZN(n3708) );
  OAI211_X1 U4362 ( .C1(n3660), .C2(n3643), .A(n3661), .B(n3708), .ZN(n3774)
         );
  AOI21_X1 U4363 ( .B1(n3926), .B2(n3769), .A(n3774), .ZN(n3666) );
  NAND2_X1 U4364 ( .A1(n3905), .A2(n4148), .ZN(n3672) );
  INV_X1 U4365 ( .A(n3644), .ZN(n3756) );
  INV_X1 U4366 ( .A(n3645), .ZN(n3651) );
  INV_X1 U4367 ( .A(n3646), .ZN(n3648) );
  NOR2_X1 U4368 ( .A1(n3647), .A2(n3648), .ZN(n3753) );
  AOI21_X1 U4369 ( .B1(n3650), .B2(n3649), .A(n3648), .ZN(n3752) );
  AOI21_X1 U4370 ( .B1(n3651), .B2(n3753), .A(n3752), .ZN(n3653) );
  INV_X1 U4371 ( .A(n3652), .ZN(n3755) );
  OAI211_X1 U4372 ( .C1(n3756), .C2(n3653), .A(n3755), .B(n3751), .ZN(n3654)
         );
  AOI21_X1 U4373 ( .B1(n3758), .B2(n3654), .A(n2036), .ZN(n3656) );
  OAI21_X1 U4374 ( .B1(n3760), .B2(n3656), .A(n3655), .ZN(n3657) );
  NAND2_X1 U4375 ( .A1(n3762), .A2(n3657), .ZN(n3659) );
  INV_X1 U4376 ( .A(n3708), .ZN(n3658) );
  AOI21_X1 U4377 ( .B1(n3766), .B2(n3659), .A(n3658), .ZN(n3662) );
  NAND4_X1 U4378 ( .A1(n3662), .A2(n3773), .A3(n3661), .A4(n3660), .ZN(n3663)
         );
  OR2_X1 U4379 ( .A1(n4140), .A2(n4141), .ZN(n3673) );
  OAI211_X1 U4380 ( .C1(n4141), .C2(n3672), .A(n3663), .B(n3673), .ZN(n3665)
         );
  INV_X1 U4381 ( .A(n4141), .ZN(n3664) );
  OAI22_X1 U4382 ( .A1(n3666), .A2(n3665), .B1(n3664), .B2(n4148), .ZN(n3783)
         );
  INV_X1 U4383 ( .A(n3667), .ZN(n3955) );
  NAND4_X1 U4384 ( .A1(n3978), .A2(n3670), .A3(n3778), .A4(n3669), .ZN(n3679)
         );
  NOR2_X1 U4385 ( .A1(n3936), .A2(n3671), .ZN(n3957) );
  NAND2_X1 U4386 ( .A1(n3673), .A2(n3672), .ZN(n3777) );
  INV_X1 U4387 ( .A(n3777), .ZN(n3676) );
  NAND2_X1 U4388 ( .A1(n3675), .A2(n3674), .ZN(n4049) );
  NAND3_X1 U4389 ( .A1(n3957), .A2(n3676), .A3(n4049), .ZN(n3678) );
  OR3_X1 U4390 ( .A1(n3679), .A2(n3678), .A3(n3677), .ZN(n3681) );
  XNOR2_X1 U4391 ( .A(n4022), .B(n3680), .ZN(n3993) );
  INV_X1 U4392 ( .A(n3993), .ZN(n3998) );
  XNOR2_X1 U4393 ( .A(n4053), .B(n4078), .ZN(n4075) );
  NOR4_X1 U4394 ( .A1(n3913), .A2(n3681), .A3(n3998), .A4(n4075), .ZN(n3713)
         );
  INV_X1 U4395 ( .A(n4092), .ZN(n4097) );
  NAND4_X1 U4396 ( .A1(n3684), .A2(n4097), .A3(n3683), .A4(n3682), .ZN(n3690)
         );
  INV_X1 U4397 ( .A(n3685), .ZN(n3686) );
  NAND2_X1 U4398 ( .A1(n4070), .A2(n4069), .ZN(n4114) );
  INV_X1 U4399 ( .A(n4114), .ZN(n4115) );
  NAND4_X1 U4400 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n4115), .ZN(n3689)
         );
  NOR2_X1 U4401 ( .A1(n3690), .A2(n3689), .ZN(n3712) );
  INV_X1 U4402 ( .A(n3994), .ZN(n3691) );
  NAND2_X1 U4403 ( .A1(n3691), .A2(n3995), .ZN(n4036) );
  INV_X1 U4404 ( .A(n4036), .ZN(n3695) );
  INV_X1 U4405 ( .A(n4020), .ZN(n3694) );
  NAND4_X1 U4406 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3700)
         );
  NAND4_X1 U4407 ( .A1(n3698), .A2(n3697), .A3(n3733), .A4(n3696), .ZN(n3699)
         );
  NOR2_X1 U4408 ( .A1(n3700), .A2(n3699), .ZN(n3711) );
  NOR2_X1 U4409 ( .A1(n3702), .A2(n3701), .ZN(n3940) );
  NOR2_X1 U4410 ( .A1(n4382), .A2(n3703), .ZN(n3704) );
  NAND4_X1 U4411 ( .A1(n3940), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3709)
         );
  NAND2_X1 U4412 ( .A1(n3708), .A2(n3707), .ZN(n3915) );
  NOR2_X1 U4413 ( .A1(n3709), .A2(n3915), .ZN(n3710) );
  NAND4_X1 U4414 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3715)
         );
  INV_X1 U4415 ( .A(n3926), .ZN(n3714) );
  NOR2_X1 U4416 ( .A1(n3715), .A2(n3714), .ZN(n3781) );
  INV_X1 U4417 ( .A(n3716), .ZN(n3718) );
  OAI211_X1 U4418 ( .C1(n3719), .C2(n4268), .A(n3718), .B(n3717), .ZN(n3721)
         );
  NAND3_X1 U4419 ( .A1(n3721), .A2(n3720), .A3(n2831), .ZN(n3724) );
  NAND3_X1 U4420 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3727) );
  NAND3_X1 U4421 ( .A1(n3727), .A2(n3726), .A3(n3725), .ZN(n3731) );
  AND4_X1 U4422 ( .A1(n3731), .A2(n3730), .A3(n3729), .A4(n3728), .ZN(n3739)
         );
  OAI211_X1 U4423 ( .C1(n3735), .C2(n3734), .A(n3733), .B(n3732), .ZN(n3738)
         );
  OAI211_X1 U4424 ( .C1(n3739), .C2(n3738), .A(n3737), .B(n3736), .ZN(n3742)
         );
  AND3_X1 U4425 ( .A1(n3742), .A2(n3741), .A3(n3740), .ZN(n3745) );
  OAI21_X1 U4426 ( .B1(n3745), .B2(n3744), .A(n3743), .ZN(n3748) );
  NAND3_X1 U4427 ( .A1(n3748), .A2(n3747), .A3(n3746), .ZN(n3750) );
  AND2_X1 U4428 ( .A1(n3750), .A2(n3749), .ZN(n3754) );
  AOI211_X1 U4429 ( .C1(n3754), .C2(n3753), .A(n2073), .B(n3752), .ZN(n3757)
         );
  OAI21_X1 U4430 ( .B1(n3757), .B2(n3756), .A(n3755), .ZN(n3759) );
  AOI211_X1 U4431 ( .C1(n3759), .C2(n3758), .A(n2036), .B(n3994), .ZN(n3761)
         );
  NOR2_X1 U4432 ( .A1(n3761), .A2(n3760), .ZN(n3764) );
  OAI21_X1 U4433 ( .B1(n3764), .B2(n3763), .A(n3762), .ZN(n3765) );
  NAND2_X1 U4434 ( .A1(n3766), .A2(n3765), .ZN(n3772) );
  NOR2_X1 U4435 ( .A1(n3768), .A2(n3767), .ZN(n3771) );
  INV_X1 U4436 ( .A(n3769), .ZN(n3770) );
  AOI211_X1 U4437 ( .C1(n3773), .C2(n3772), .A(n3771), .B(n3770), .ZN(n3775)
         );
  NOR2_X1 U4438 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  AOI21_X1 U4439 ( .B1(n3778), .B2(n3777), .A(n3776), .ZN(n3780) );
  MUX2_X1 U4440 ( .A(n3781), .B(n3780), .S(n3779), .Z(n3782) );
  AOI21_X1 U4441 ( .B1(n3784), .B2(n3783), .A(n3782), .ZN(n3785) );
  XNOR2_X1 U4442 ( .A(n3785), .B(n3894), .ZN(n3791) );
  INV_X1 U4443 ( .A(n3786), .ZN(n3787) );
  NOR2_X1 U4444 ( .A1(n3787), .A2(n3818), .ZN(n3789) );
  OAI21_X1 U4445 ( .B1(n3790), .B2(n4267), .A(B_REG_SCAN_IN), .ZN(n3788) );
  OAI22_X1 U4446 ( .A1(n3791), .A2(n3790), .B1(n3789), .B2(n3788), .ZN(U3239)
         );
  MUX2_X1 U4447 ( .A(n4140), .B(DATAO_REG_31__SCAN_IN), .S(n3819), .Z(U3581)
         );
  MUX2_X1 U4448 ( .A(n3905), .B(DATAO_REG_30__SCAN_IN), .S(n3819), .Z(U3580)
         );
  MUX2_X1 U4449 ( .A(DATAO_REG_29__SCAN_IN), .B(n3792), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4450 ( .A(DATAO_REG_28__SCAN_IN), .B(n3924), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4451 ( .A(DATAO_REG_27__SCAN_IN), .B(n3942), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4452 ( .A(n3793), .B(DATAO_REG_26__SCAN_IN), .S(n3819), .Z(U3576)
         );
  MUX2_X1 U4453 ( .A(n3981), .B(DATAO_REG_25__SCAN_IN), .S(n3819), .Z(U3575)
         );
  MUX2_X1 U4454 ( .A(DATAO_REG_23__SCAN_IN), .B(n4022), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4455 ( .A(n4051), .B(DATAO_REG_21__SCAN_IN), .S(n3819), .Z(U3571)
         );
  MUX2_X1 U4456 ( .A(n4079), .B(DATAO_REG_20__SCAN_IN), .S(n3819), .Z(U3570)
         );
  MUX2_X1 U4457 ( .A(DATAO_REG_19__SCAN_IN), .B(n4102), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4458 ( .A(n3794), .B(DATAO_REG_17__SCAN_IN), .S(n3819), .Z(U3567)
         );
  MUX2_X1 U4459 ( .A(n4120), .B(DATAO_REG_16__SCAN_IN), .S(n3819), .Z(U3566)
         );
  MUX2_X1 U4460 ( .A(n2807), .B(DATAO_REG_15__SCAN_IN), .S(n3819), .Z(U3565)
         );
  MUX2_X1 U4461 ( .A(n3795), .B(DATAO_REG_14__SCAN_IN), .S(n3819), .Z(U3564)
         );
  MUX2_X1 U4462 ( .A(DATAO_REG_13__SCAN_IN), .B(n3796), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4463 ( .A(n3797), .B(DATAO_REG_12__SCAN_IN), .S(n3819), .Z(U3562)
         );
  MUX2_X1 U4464 ( .A(n3798), .B(DATAO_REG_10__SCAN_IN), .S(n3819), .Z(U3560)
         );
  MUX2_X1 U4465 ( .A(n3799), .B(DATAO_REG_9__SCAN_IN), .S(n3819), .Z(U3559) );
  MUX2_X1 U4466 ( .A(n3800), .B(DATAO_REG_8__SCAN_IN), .S(n3819), .Z(U3558) );
  MUX2_X1 U4467 ( .A(n3801), .B(DATAO_REG_7__SCAN_IN), .S(n3819), .Z(U3557) );
  MUX2_X1 U4468 ( .A(n3802), .B(DATAO_REG_6__SCAN_IN), .S(n3819), .Z(U3556) );
  MUX2_X1 U4469 ( .A(n3803), .B(DATAO_REG_5__SCAN_IN), .S(n3819), .Z(U3555) );
  MUX2_X1 U4470 ( .A(n3804), .B(DATAO_REG_4__SCAN_IN), .S(n3819), .Z(U3554) );
  MUX2_X1 U4471 ( .A(n2784), .B(DATAO_REG_1__SCAN_IN), .S(n3819), .Z(U3551) );
  MUX2_X1 U4472 ( .A(n3805), .B(DATAO_REG_0__SCAN_IN), .S(n3819), .Z(U3550) );
  AOI22_X1 U4473 ( .A1(n4345), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3814) );
  INV_X1 U4474 ( .A(n4375), .ZN(n4335) );
  NAND2_X1 U4475 ( .A1(n4335), .A2(n2285), .ZN(n3813) );
  OAI211_X1 U4476 ( .C1(n3820), .C2(n3807), .A(n4370), .B(n3806), .ZN(n3812)
         );
  OAI211_X1 U4477 ( .C1(n3810), .C2(n3809), .A(n4372), .B(n3808), .ZN(n3811)
         );
  NAND4_X1 U4478 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(U3241)
         );
  AOI21_X1 U4479 ( .B1(n4287), .B2(n2301), .A(n3815), .ZN(n4288) );
  INV_X1 U4480 ( .A(n4287), .ZN(n3816) );
  NAND3_X1 U4481 ( .A1(n3817), .A2(n4266), .A3(n3816), .ZN(n3823) );
  INV_X1 U4482 ( .A(n3818), .ZN(n3821) );
  AOI21_X1 U4483 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n3822) );
  OAI211_X1 U4484 ( .C1(n4401), .C2(n4288), .A(n3823), .B(n3822), .ZN(n3843)
         );
  AOI22_X1 U4485 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4345), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3833) );
  XNOR2_X1 U4486 ( .A(n3825), .B(n3824), .ZN(n3826) );
  OAI22_X1 U4487 ( .A1(n3826), .A2(n4339), .B1(n4375), .B2(n4275), .ZN(n3827)
         );
  INV_X1 U4488 ( .A(n3827), .ZN(n3832) );
  OAI211_X1 U4489 ( .C1(n3830), .C2(n3829), .A(n4370), .B(n3828), .ZN(n3831)
         );
  NAND4_X1 U4490 ( .A1(n3843), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(U3242)
         );
  NAND2_X1 U4491 ( .A1(n4345), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3842) );
  XOR2_X1 U4492 ( .A(REG1_REG_4__SCAN_IN), .B(n3834), .Z(n3840) );
  XNOR2_X1 U4493 ( .A(n3835), .B(REG2_REG_4__SCAN_IN), .ZN(n3838) );
  AOI21_X1 U4494 ( .B1(n4335), .B2(n4273), .A(n3836), .ZN(n3837) );
  OAI21_X1 U4495 ( .B1(n3838), .B2(n4325), .A(n3837), .ZN(n3839) );
  AOI21_X1 U4496 ( .B1(n4372), .B2(n3840), .A(n3839), .ZN(n3841) );
  NAND3_X1 U4497 ( .A1(n3843), .A2(n3842), .A3(n3841), .ZN(U3244) );
  NOR2_X1 U4498 ( .A1(n4375), .A2(n3844), .ZN(n3845) );
  AOI211_X1 U4499 ( .C1(n4345), .C2(ADDR_REG_5__SCAN_IN), .A(n3846), .B(n3845), 
        .ZN(n3855) );
  OAI211_X1 U4500 ( .C1(n3849), .C2(n3848), .A(n4372), .B(n3847), .ZN(n3854)
         );
  OAI211_X1 U4501 ( .C1(n3852), .C2(n3851), .A(n4370), .B(n3850), .ZN(n3853)
         );
  NAND3_X1 U4502 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(U3245) );
  INV_X1 U4503 ( .A(n4270), .ZN(n3885) );
  XNOR2_X1 U4504 ( .A(n4270), .B(REG2_REG_18__SCAN_IN), .ZN(n3869) );
  NOR2_X1 U4505 ( .A1(n3881), .A2(REG2_REG_17__SCAN_IN), .ZN(n3856) );
  AOI21_X1 U4506 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3881), .A(n3856), .ZN(n4368) );
  NAND2_X1 U4507 ( .A1(n3858), .A2(n3857), .ZN(n3859) );
  NAND2_X1 U4508 ( .A1(n3873), .A2(n3859), .ZN(n3860) );
  XNOR2_X1 U4509 ( .A(n3859), .B(n4398), .ZN(n4311) );
  NAND2_X1 U4510 ( .A1(n4396), .A2(REG2_REG_13__SCAN_IN), .ZN(n3861) );
  INV_X1 U4511 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4327) );
  INV_X1 U4512 ( .A(n3864), .ZN(n3862) );
  OAI21_X1 U4513 ( .B1(n4334), .B2(n3863), .A(n3862), .ZN(n4328) );
  NOR2_X1 U4514 ( .A1(n4327), .A2(n4328), .ZN(n4326) );
  AOI22_X1 U4515 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4352), .B1(n4394), .B2(
        n3865), .ZN(n4348) );
  NAND2_X1 U4516 ( .A1(n3866), .A2(n4393), .ZN(n3867) );
  NAND2_X1 U4517 ( .A1(n4357), .A2(n2899), .ZN(n4356) );
  NAND2_X1 U4518 ( .A1(n3867), .A2(n4356), .ZN(n4367) );
  NAND2_X1 U4519 ( .A1(n4368), .A2(n4367), .ZN(n4366) );
  AOI21_X1 U4520 ( .B1(n3869), .B2(n3868), .A(n3890), .ZN(n3870) );
  NAND2_X1 U4521 ( .A1(n4270), .A2(REG1_REG_18__SCAN_IN), .ZN(n3886) );
  OAI21_X1 U4522 ( .B1(n4270), .B2(REG1_REG_18__SCAN_IN), .A(n3886), .ZN(n3883) );
  INV_X1 U4523 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U4524 ( .A1(n3881), .A2(REG1_REG_17__SCAN_IN), .B1(n4200), .B2(
        n4391), .ZN(n4365) );
  NOR2_X1 U4525 ( .A1(n2030), .A2(n4398), .ZN(n3874) );
  AOI22_X1 U4526 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4324), .B1(n4396), .B2(
        n4548), .ZN(n4315) );
  NOR2_X1 U4527 ( .A1(n4316), .A2(n4315), .ZN(n4314) );
  AND2_X1 U4528 ( .A1(n4396), .A2(REG1_REG_13__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4529 ( .A1(n3877), .A2(n4334), .ZN(n3876) );
  INV_X1 U4530 ( .A(n3876), .ZN(n3878) );
  INV_X1 U4531 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4330) );
  OAI21_X1 U4532 ( .B1(n3877), .B2(n4334), .A(n3876), .ZN(n4331) );
  NOR2_X1 U4533 ( .A1(n4330), .A2(n4331), .ZN(n4329) );
  NOR2_X1 U4534 ( .A1(n3878), .A2(n4329), .ZN(n4342) );
  INV_X1 U4535 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4536 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4352), .B1(n4394), .B2(
        n4209), .ZN(n4341) );
  NAND2_X1 U4537 ( .A1(n3879), .A2(n4393), .ZN(n3880) );
  INV_X1 U4538 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U4539 ( .A1(n3880), .A2(n4354), .ZN(n4364) );
  NAND2_X1 U4540 ( .A1(n4365), .A2(n4364), .ZN(n4363) );
  XNOR2_X1 U4541 ( .A(n3887), .B(REG1_REG_19__SCAN_IN), .ZN(n3888) );
  XNOR2_X1 U4542 ( .A(n3889), .B(n3888), .ZN(n3898) );
  INV_X1 U4543 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4558) );
  MUX2_X1 U4544 ( .A(n4558), .B(REG2_REG_19__SCAN_IN), .S(n3894), .Z(n3891) );
  AOI21_X1 U4545 ( .B1(n4345), .B2(ADDR_REG_19__SCAN_IN), .A(n3892), .ZN(n3893) );
  OAI21_X1 U4546 ( .B1(n3894), .B2(n4375), .A(n3893), .ZN(n3895) );
  AOI21_X1 U4547 ( .B1(n3896), .B2(n4370), .A(n3895), .ZN(n3897) );
  OAI21_X1 U4548 ( .B1(n3898), .B2(n4339), .A(n3897), .ZN(U3259) );
  INV_X1 U4549 ( .A(n3899), .ZN(n3911) );
  INV_X1 U4550 ( .A(n3900), .ZN(n3901) );
  OAI21_X1 U4551 ( .B1(n3903), .B2(n3902), .A(n3901), .ZN(n3904) );
  XNOR2_X1 U4552 ( .A(n3904), .B(n3915), .ZN(n3910) );
  INV_X1 U4553 ( .A(n3905), .ZN(n3907) );
  NAND2_X1 U4554 ( .A1(n4287), .A2(B_REG_SCAN_IN), .ZN(n3906) );
  NAND2_X1 U4555 ( .A1(n4101), .A2(n3906), .ZN(n4138) );
  OAI22_X1 U4556 ( .A1(n3907), .A2(n4138), .B1(n3917), .B2(n4147), .ZN(n3908)
         );
  AOI21_X1 U4557 ( .B1(n3924), .B2(n4121), .A(n3908), .ZN(n3909) );
  OAI21_X1 U4558 ( .B1(n3910), .B2(n4123), .A(n3909), .ZN(n4154) );
  AOI21_X1 U4559 ( .B1(n3911), .B2(n4381), .A(n4154), .ZN(n3921) );
  XNOR2_X1 U4560 ( .A(n3916), .B(n3915), .ZN(n4153) );
  NAND2_X1 U4561 ( .A1(n4153), .A2(n4037), .ZN(n3920) );
  INV_X1 U4562 ( .A(n3917), .ZN(n3918) );
  AOI21_X1 U4563 ( .B1(n3918), .B2(n2010), .A(n4146), .ZN(n4155) );
  AOI22_X1 U4564 ( .A1(n4155), .A2(n4282), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4063), .ZN(n3919) );
  OAI211_X1 U4565 ( .C1(n4063), .C2(n3921), .A(n3920), .B(n3919), .ZN(U3354)
         );
  OAI22_X1 U4566 ( .A1(n3964), .A2(n4104), .B1(n3928), .B2(n4147), .ZN(n3923)
         );
  XOR2_X1 U4567 ( .A(n3926), .B(n3925), .Z(n4158) );
  NAND2_X1 U4568 ( .A1(n4158), .A2(n4037), .ZN(n3934) );
  OAI21_X1 U4569 ( .B1(n3946), .B2(n3928), .A(n3927), .ZN(n4161) );
  INV_X1 U4570 ( .A(n4161), .ZN(n3932) );
  OAI22_X1 U4571 ( .A1(n3930), .A2(n4129), .B1(n3929), .B2(n4278), .ZN(n3931)
         );
  AOI21_X1 U4572 ( .B1(n3932), .B2(n4282), .A(n3931), .ZN(n3933) );
  OAI211_X1 U4573 ( .C1(n4159), .C2(n4063), .A(n3934), .B(n3933), .ZN(U3263)
         );
  XNOR2_X1 U4574 ( .A(n3935), .B(n3940), .ZN(n4163) );
  INV_X1 U4575 ( .A(n4163), .ZN(n3953) );
  INV_X1 U4576 ( .A(n3936), .ZN(n3937) );
  NAND2_X1 U4577 ( .A1(n3938), .A2(n3937), .ZN(n3939) );
  XOR2_X1 U4578 ( .A(n3940), .B(n3939), .Z(n3945) );
  AOI22_X1 U4579 ( .A1(n3981), .A2(n4121), .B1(n3941), .B2(n4099), .ZN(n3944)
         );
  NAND2_X1 U4580 ( .A1(n3942), .A2(n4101), .ZN(n3943) );
  OAI211_X1 U4581 ( .C1(n3945), .C2(n4123), .A(n3944), .B(n3943), .ZN(n4162)
         );
  INV_X1 U4582 ( .A(n3946), .ZN(n3947) );
  OAI21_X1 U4583 ( .B1(n3965), .B2(n3948), .A(n3947), .ZN(n4225) );
  AOI22_X1 U4584 ( .A1(n3949), .A2(n4381), .B1(n4063), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n3950) );
  OAI21_X1 U4585 ( .B1(n4225), .B2(n4127), .A(n3950), .ZN(n3951) );
  AOI21_X1 U4586 ( .B1(n4162), .B2(n4278), .A(n3951), .ZN(n3952) );
  OAI21_X1 U4587 ( .B1(n3953), .B2(n4135), .A(n3952), .ZN(U3264) );
  XOR2_X1 U4588 ( .A(n3957), .B(n3954), .Z(n4167) );
  INV_X1 U4589 ( .A(n4167), .ZN(n3973) );
  NAND2_X1 U4590 ( .A1(n3956), .A2(n3955), .ZN(n3959) );
  INV_X1 U4591 ( .A(n3957), .ZN(n3958) );
  XNOR2_X1 U4592 ( .A(n3959), .B(n3958), .ZN(n3960) );
  NAND2_X1 U4593 ( .A1(n3960), .A2(n4107), .ZN(n3963) );
  AOI22_X1 U4594 ( .A1(n4001), .A2(n4121), .B1(n3961), .B2(n4099), .ZN(n3962)
         );
  OAI211_X1 U4595 ( .C1(n3964), .C2(n4117), .A(n3963), .B(n3962), .ZN(n4166)
         );
  INV_X1 U4596 ( .A(n3984), .ZN(n3968) );
  INV_X1 U4597 ( .A(n3965), .ZN(n3966) );
  AOI22_X1 U4598 ( .A1(n4063), .A2(REG2_REG_25__SCAN_IN), .B1(n3969), .B2(
        n4381), .ZN(n3970) );
  OAI21_X1 U4599 ( .B1(n4229), .B2(n4127), .A(n3970), .ZN(n3971) );
  AOI21_X1 U4600 ( .B1(n4278), .B2(n4166), .A(n3971), .ZN(n3972) );
  OAI21_X1 U4601 ( .B1(n3973), .B2(n4135), .A(n3972), .ZN(U3265) );
  XNOR2_X1 U4602 ( .A(n3974), .B(n3978), .ZN(n4171) );
  INV_X1 U4603 ( .A(n4171), .ZN(n3991) );
  NAND2_X1 U4604 ( .A1(n3976), .A2(n3975), .ZN(n3977) );
  XOR2_X1 U4605 ( .A(n3978), .B(n3977), .Z(n3983) );
  OAI22_X1 U4606 ( .A1(n3979), .A2(n4104), .B1(n3985), .B2(n4147), .ZN(n3980)
         );
  AOI21_X1 U4607 ( .B1(n4101), .B2(n3981), .A(n3980), .ZN(n3982) );
  OAI21_X1 U4608 ( .B1(n3983), .B2(n4123), .A(n3982), .ZN(n4170) );
  INV_X1 U4609 ( .A(n4004), .ZN(n3986) );
  OAI21_X1 U4610 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n4233) );
  AOI22_X1 U4611 ( .A1(n4063), .A2(REG2_REG_24__SCAN_IN), .B1(n3987), .B2(
        n4381), .ZN(n3988) );
  OAI21_X1 U4612 ( .B1(n4233), .B2(n4127), .A(n3988), .ZN(n3989) );
  AOI21_X1 U4613 ( .B1(n4170), .B2(n4278), .A(n3989), .ZN(n3990) );
  OAI21_X1 U4614 ( .B1(n3991), .B2(n4135), .A(n3990), .ZN(U3266) );
  XNOR2_X1 U4615 ( .A(n3992), .B(n3993), .ZN(n4175) );
  INV_X1 U4616 ( .A(n4175), .ZN(n4011) );
  OR2_X1 U4617 ( .A1(n4031), .A2(n3994), .ZN(n3996) );
  OAI21_X1 U4618 ( .B1(n4021), .B2(n4020), .A(n3997), .ZN(n3999) );
  XNOR2_X1 U4619 ( .A(n3999), .B(n3998), .ZN(n4003) );
  OAI22_X1 U4620 ( .A1(n4030), .A2(n4104), .B1(n4147), .B2(n4005), .ZN(n4000)
         );
  AOI21_X1 U4621 ( .B1(n4001), .B2(n4101), .A(n4000), .ZN(n4002) );
  OAI21_X1 U4622 ( .B1(n4003), .B2(n4123), .A(n4002), .ZN(n4174) );
  OAI21_X1 U4623 ( .B1(n4014), .B2(n4005), .A(n4004), .ZN(n4237) );
  NOR2_X1 U4624 ( .A1(n4237), .A2(n4127), .ZN(n4009) );
  INV_X1 U4625 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4007) );
  OAI22_X1 U4626 ( .A1(n4278), .A2(n4007), .B1(n4006), .B2(n4129), .ZN(n4008)
         );
  AOI211_X1 U4627 ( .C1(n4174), .C2(n4278), .A(n4009), .B(n4008), .ZN(n4010)
         );
  OAI21_X1 U4628 ( .B1(n4011), .B2(n4135), .A(n4010), .ZN(U3267) );
  OAI21_X1 U4629 ( .B1(n4013), .B2(n4020), .A(n4012), .ZN(n4182) );
  INV_X1 U4630 ( .A(n4014), .ZN(n4179) );
  NAND2_X1 U4631 ( .A1(n4038), .A2(n4015), .ZN(n4178) );
  AND2_X1 U4632 ( .A1(n4178), .A2(n4282), .ZN(n4019) );
  INV_X1 U4633 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4017) );
  OAI22_X1 U4634 ( .A1(n4278), .A2(n4017), .B1(n4016), .B2(n4129), .ZN(n4018)
         );
  AOI21_X1 U4635 ( .B1(n4179), .B2(n4019), .A(n4018), .ZN(n4029) );
  XNOR2_X1 U4636 ( .A(n4021), .B(n4020), .ZN(n4027) );
  NAND2_X1 U4637 ( .A1(n4022), .A2(n4101), .ZN(n4024) );
  NAND2_X1 U4638 ( .A1(n4051), .A2(n4121), .ZN(n4023) );
  OAI211_X1 U4639 ( .C1(n4147), .C2(n4025), .A(n4024), .B(n4023), .ZN(n4026)
         );
  AOI21_X1 U4640 ( .B1(n4027), .B2(n4107), .A(n4026), .ZN(n4181) );
  OR2_X1 U4641 ( .A1(n4181), .A2(n4063), .ZN(n4028) );
  OAI211_X1 U4642 ( .C1(n4182), .C2(n4135), .A(n4029), .B(n4028), .ZN(U3268)
         );
  OAI22_X1 U4643 ( .A1(n4030), .A2(n4117), .B1(n4147), .B2(n4039), .ZN(n4034)
         );
  XOR2_X1 U4644 ( .A(n4036), .B(n4031), .Z(n4032) );
  NOR2_X1 U4645 ( .A1(n4032), .A2(n4123), .ZN(n4033) );
  AOI211_X1 U4646 ( .C1(n4121), .C2(n4079), .A(n4034), .B(n4033), .ZN(n4183)
         );
  XNOR2_X1 U4647 ( .A(n4035), .B(n4036), .ZN(n4185) );
  NAND2_X1 U4648 ( .A1(n4185), .A2(n4037), .ZN(n4045) );
  OAI21_X1 U4649 ( .B1(n2134), .B2(n4039), .A(n4038), .ZN(n4242) );
  INV_X1 U4650 ( .A(n4242), .ZN(n4043) );
  INV_X1 U4651 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4041) );
  OAI22_X1 U4652 ( .A1(n4278), .A2(n4041), .B1(n4040), .B2(n4129), .ZN(n4042)
         );
  AOI21_X1 U4653 ( .B1(n4043), .B2(n4282), .A(n4042), .ZN(n4044) );
  OAI211_X1 U4654 ( .C1(n4063), .C2(n4183), .A(n4045), .B(n4044), .ZN(U3269)
         );
  XNOR2_X1 U4655 ( .A(n4046), .B(n4049), .ZN(n4058) );
  NAND2_X1 U4656 ( .A1(n4048), .A2(n4047), .ZN(n4050) );
  XNOR2_X1 U4657 ( .A(n4050), .B(n4049), .ZN(n4055) );
  AOI22_X1 U4658 ( .A1(n4051), .A2(n4101), .B1(n4059), .B2(n4099), .ZN(n4052)
         );
  OAI21_X1 U4659 ( .B1(n4053), .B2(n4104), .A(n4052), .ZN(n4054) );
  AOI21_X1 U4660 ( .B1(n4055), .B2(n4107), .A(n4054), .ZN(n4056) );
  OAI21_X1 U4661 ( .B1(n4058), .B2(n4057), .A(n4056), .ZN(n4188) );
  INV_X1 U4662 ( .A(n4188), .ZN(n4067) );
  INV_X1 U4663 ( .A(n4058), .ZN(n4189) );
  NAND2_X1 U4664 ( .A1(n4082), .A2(n4059), .ZN(n4060) );
  NAND2_X1 U4665 ( .A1(n4061), .A2(n4060), .ZN(n4246) );
  AOI22_X1 U4666 ( .A1(n4063), .A2(REG2_REG_20__SCAN_IN), .B1(n4062), .B2(
        n4381), .ZN(n4064) );
  OAI21_X1 U4667 ( .B1(n4246), .B2(n4127), .A(n4064), .ZN(n4065) );
  AOI21_X1 U4668 ( .B1(n4189), .B2(n4383), .A(n4065), .ZN(n4066) );
  OAI21_X1 U4669 ( .B1(n4067), .B2(n4063), .A(n4066), .ZN(U3270) );
  XNOR2_X1 U4670 ( .A(n4068), .B(n4075), .ZN(n4192) );
  INV_X1 U4671 ( .A(n4192), .ZN(n4089) );
  INV_X1 U4672 ( .A(n4069), .ZN(n4071) );
  OAI21_X1 U4673 ( .B1(n4116), .B2(n4071), .A(n4070), .ZN(n4098) );
  INV_X1 U4674 ( .A(n4072), .ZN(n4074) );
  OAI21_X1 U4675 ( .B1(n4098), .B2(n4074), .A(n4073), .ZN(n4076) );
  XNOR2_X1 U4676 ( .A(n4076), .B(n4075), .ZN(n4077) );
  NAND2_X1 U4677 ( .A1(n4077), .A2(n4107), .ZN(n4081) );
  AOI22_X1 U4678 ( .A1(n4079), .A2(n4101), .B1(n4078), .B2(n4099), .ZN(n4080)
         );
  OAI211_X1 U4679 ( .C1(n4118), .C2(n4104), .A(n4081), .B(n4080), .ZN(n4191)
         );
  OAI21_X1 U4680 ( .B1(n4094), .B2(n4083), .A(n4082), .ZN(n4249) );
  NOR2_X1 U4681 ( .A1(n4249), .A2(n4127), .ZN(n4087) );
  INV_X1 U4682 ( .A(n4084), .ZN(n4085) );
  OAI22_X1 U4683 ( .A1(n4278), .A2(n4558), .B1(n4085), .B2(n4129), .ZN(n4086)
         );
  AOI211_X1 U4684 ( .C1(n4191), .C2(n4278), .A(n4087), .B(n4086), .ZN(n4088)
         );
  OAI21_X1 U4685 ( .B1(n4089), .B2(n4135), .A(n4088), .ZN(U3271) );
  OAI21_X1 U4686 ( .B1(n4090), .B2(n4092), .A(n4091), .ZN(n4093) );
  INV_X1 U4687 ( .A(n4093), .ZN(n4197) );
  INV_X1 U4688 ( .A(n4094), .ZN(n4095) );
  OAI211_X1 U4689 ( .C1(n2129), .C2(n2813), .A(n4095), .B(n4440), .ZN(n4195)
         );
  INV_X1 U4690 ( .A(n4195), .ZN(n4112) );
  OAI22_X1 U4691 ( .A1(n4278), .A2(n4557), .B1(n4096), .B2(n4129), .ZN(n4110)
         );
  XNOR2_X1 U4692 ( .A(n4098), .B(n4097), .ZN(n4108) );
  AOI22_X1 U4693 ( .A1(n4102), .A2(n4101), .B1(n4100), .B2(n4099), .ZN(n4103)
         );
  OAI21_X1 U4694 ( .B1(n4105), .B2(n4104), .A(n4103), .ZN(n4106) );
  AOI21_X1 U4695 ( .B1(n4108), .B2(n4107), .A(n4106), .ZN(n4196) );
  NOR2_X1 U4696 ( .A1(n4196), .A2(n4063), .ZN(n4109) );
  AOI211_X1 U4697 ( .C1(n4112), .C2(n4111), .A(n4110), .B(n4109), .ZN(n4113)
         );
  OAI21_X1 U4698 ( .B1(n4197), .B2(n4135), .A(n4113), .ZN(U3272) );
  XNOR2_X1 U4699 ( .A(n2035), .B(n4114), .ZN(n4199) );
  INV_X1 U4700 ( .A(n4199), .ZN(n4136) );
  XNOR2_X1 U4701 ( .A(n4116), .B(n4115), .ZN(n4124) );
  OAI22_X1 U4702 ( .A1(n4118), .A2(n4117), .B1(n4147), .B2(n4126), .ZN(n4119)
         );
  AOI21_X1 U4703 ( .B1(n4121), .B2(n4120), .A(n4119), .ZN(n4122) );
  OAI21_X1 U4704 ( .B1(n4124), .B2(n4123), .A(n4122), .ZN(n4198) );
  OAI21_X1 U4705 ( .B1(n2126), .B2(n4126), .A(n4125), .ZN(n4254) );
  NOR2_X1 U4706 ( .A1(n4254), .A2(n4127), .ZN(n4133) );
  INV_X1 U4707 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4131) );
  INV_X1 U4708 ( .A(n4128), .ZN(n4130) );
  OAI22_X1 U4709 ( .A1(n4278), .A2(n4131), .B1(n4130), .B2(n4129), .ZN(n4132)
         );
  AOI211_X1 U4710 ( .C1(n4198), .C2(n4278), .A(n4133), .B(n4132), .ZN(n4134)
         );
  OAI21_X1 U4711 ( .B1(n4136), .B2(n4135), .A(n4134), .ZN(U3273) );
  INV_X1 U4712 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4144) );
  NAND2_X1 U4713 ( .A1(n4146), .A2(n4148), .ZN(n4145) );
  XNOR2_X1 U4714 ( .A(n4145), .B(n4141), .ZN(n4279) );
  NAND2_X1 U4715 ( .A1(n4279), .A2(n4137), .ZN(n4143) );
  INV_X1 U4716 ( .A(n4138), .ZN(n4139) );
  NAND2_X1 U4717 ( .A1(n4140), .A2(n4139), .ZN(n4150) );
  OAI21_X1 U4718 ( .B1(n4141), .B2(n4147), .A(n4150), .ZN(n4277) );
  NAND2_X1 U4719 ( .A1(n4453), .A2(n4277), .ZN(n4142) );
  OAI211_X1 U4720 ( .C1(n4453), .C2(n4144), .A(n4143), .B(n4142), .ZN(U3549)
         );
  OAI21_X1 U4721 ( .B1(n4146), .B2(n4148), .A(n4145), .ZN(n4281) );
  OR2_X1 U4722 ( .A1(n4148), .A2(n4147), .ZN(n4149) );
  AND2_X1 U4723 ( .A1(n4150), .A2(n4149), .ZN(n4285) );
  INV_X1 U4724 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4151) );
  MUX2_X1 U4725 ( .A(n4285), .B(n4151), .S(n4451), .Z(n4152) );
  OAI21_X1 U4726 ( .B1(n4281), .B2(n4214), .A(n4152), .ZN(U3548) );
  NAND2_X1 U4727 ( .A1(n4153), .A2(n4428), .ZN(n4157) );
  NAND2_X1 U4728 ( .A1(n4157), .A2(n4156), .ZN(n4220) );
  MUX2_X1 U4729 ( .A(REG1_REG_29__SCAN_IN), .B(n4220), .S(n4453), .Z(U3547) );
  NAND2_X1 U4730 ( .A1(n4158), .A2(n4428), .ZN(n4160) );
  OAI211_X1 U4731 ( .C1(n4430), .C2(n4161), .A(n4160), .B(n4159), .ZN(n4221)
         );
  MUX2_X1 U4732 ( .A(REG1_REG_27__SCAN_IN), .B(n4221), .S(n4453), .Z(U3545) );
  INV_X1 U4733 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4164) );
  AOI21_X1 U4734 ( .B1(n4163), .B2(n4428), .A(n4162), .ZN(n4222) );
  MUX2_X1 U4735 ( .A(n4164), .B(n4222), .S(n4453), .Z(n4165) );
  OAI21_X1 U4736 ( .B1(n4214), .B2(n4225), .A(n4165), .ZN(U3544) );
  INV_X1 U4737 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4168) );
  AOI21_X1 U4738 ( .B1(n4167), .B2(n4428), .A(n4166), .ZN(n4226) );
  MUX2_X1 U4739 ( .A(n4168), .B(n4226), .S(n4453), .Z(n4169) );
  OAI21_X1 U4740 ( .B1(n4214), .B2(n4229), .A(n4169), .ZN(U3543) );
  AOI21_X1 U4741 ( .B1(n4171), .B2(n4428), .A(n4170), .ZN(n4230) );
  MUX2_X1 U4742 ( .A(n4172), .B(n4230), .S(n4453), .Z(n4173) );
  OAI21_X1 U4743 ( .B1(n4214), .B2(n4233), .A(n4173), .ZN(U3542) );
  INV_X1 U4744 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4176) );
  AOI21_X1 U4745 ( .B1(n4175), .B2(n4428), .A(n4174), .ZN(n4234) );
  MUX2_X1 U4746 ( .A(n4176), .B(n4234), .S(n4453), .Z(n4177) );
  OAI21_X1 U4747 ( .B1(n4214), .B2(n4237), .A(n4177), .ZN(U3541) );
  NAND3_X1 U4748 ( .A1(n4179), .A2(n4440), .A3(n4178), .ZN(n4180) );
  OAI211_X1 U4749 ( .C1(n4182), .C2(n4422), .A(n4181), .B(n4180), .ZN(n4238)
         );
  MUX2_X1 U4750 ( .A(REG1_REG_22__SCAN_IN), .B(n4238), .S(n4453), .Z(U3540) );
  INV_X1 U4751 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4186) );
  INV_X1 U4752 ( .A(n4183), .ZN(n4184) );
  AOI21_X1 U4753 ( .B1(n4185), .B2(n4428), .A(n4184), .ZN(n4239) );
  MUX2_X1 U4754 ( .A(n4186), .B(n4239), .S(n4453), .Z(n4187) );
  OAI21_X1 U4755 ( .B1(n4214), .B2(n4242), .A(n4187), .ZN(U3539) );
  INV_X1 U4756 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4554) );
  AOI21_X1 U4757 ( .B1(n4414), .B2(n4189), .A(n4188), .ZN(n4243) );
  MUX2_X1 U4758 ( .A(n4554), .B(n4243), .S(n4453), .Z(n4190) );
  OAI21_X1 U4759 ( .B1(n4214), .B2(n4246), .A(n4190), .ZN(U3538) );
  INV_X1 U4760 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4193) );
  AOI21_X1 U4761 ( .B1(n4192), .B2(n4428), .A(n4191), .ZN(n4247) );
  MUX2_X1 U4762 ( .A(n4193), .B(n4247), .S(n4453), .Z(n4194) );
  OAI21_X1 U4763 ( .B1(n4214), .B2(n4249), .A(n4194), .ZN(U3537) );
  OAI211_X1 U4764 ( .C1(n4197), .C2(n4422), .A(n4196), .B(n4195), .ZN(n4250)
         );
  MUX2_X1 U4765 ( .A(REG1_REG_18__SCAN_IN), .B(n4250), .S(n4453), .Z(U3536) );
  AOI21_X1 U4766 ( .B1(n4199), .B2(n4428), .A(n4198), .ZN(n4251) );
  MUX2_X1 U4767 ( .A(n4200), .B(n4251), .S(n4453), .Z(n4201) );
  OAI21_X1 U4768 ( .B1(n4214), .B2(n4254), .A(n4201), .ZN(U3535) );
  NAND3_X1 U4769 ( .A1(n4203), .A2(n4440), .A3(n4202), .ZN(n4204) );
  OAI211_X1 U4770 ( .C1(n4206), .C2(n4422), .A(n4205), .B(n4204), .ZN(n4255)
         );
  MUX2_X1 U4771 ( .A(REG1_REG_16__SCAN_IN), .B(n4255), .S(n4453), .Z(U3534) );
  AOI21_X1 U4772 ( .B1(n4208), .B2(n4428), .A(n4207), .ZN(n4256) );
  MUX2_X1 U4773 ( .A(n4209), .B(n4256), .S(n4453), .Z(n4210) );
  OAI21_X1 U4774 ( .B1(n4214), .B2(n4259), .A(n4210), .ZN(U3533) );
  AOI21_X1 U4775 ( .B1(n4414), .B2(n4212), .A(n4211), .ZN(n4260) );
  MUX2_X1 U4776 ( .A(n4330), .B(n4260), .S(n4453), .Z(n4213) );
  OAI21_X1 U4777 ( .B1(n4214), .B2(n4264), .A(n4213), .ZN(U3532) );
  INV_X1 U4778 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U4779 ( .A1(n4279), .A2(n4215), .ZN(n4217) );
  NAND2_X1 U4780 ( .A1(n4443), .A2(n4277), .ZN(n4216) );
  OAI211_X1 U4781 ( .C1(n4443), .C2(n4538), .A(n4217), .B(n4216), .ZN(U3517)
         );
  INV_X1 U4782 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4218) );
  MUX2_X1 U4783 ( .A(n4285), .B(n4218), .S(n4441), .Z(n4219) );
  OAI21_X1 U4784 ( .B1(n4281), .B2(n4263), .A(n4219), .ZN(U3516) );
  MUX2_X1 U4785 ( .A(REG0_REG_29__SCAN_IN), .B(n4220), .S(n4443), .Z(U3515) );
  MUX2_X1 U4786 ( .A(REG0_REG_27__SCAN_IN), .B(n4221), .S(n4443), .Z(U3513) );
  INV_X1 U4787 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4223) );
  MUX2_X1 U4788 ( .A(n4223), .B(n4222), .S(n4443), .Z(n4224) );
  OAI21_X1 U4789 ( .B1(n4225), .B2(n4263), .A(n4224), .ZN(U3512) );
  INV_X1 U4790 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4227) );
  MUX2_X1 U4791 ( .A(n4227), .B(n4226), .S(n4443), .Z(n4228) );
  OAI21_X1 U4792 ( .B1(n4229), .B2(n4263), .A(n4228), .ZN(U3511) );
  INV_X1 U4793 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4231) );
  MUX2_X1 U4794 ( .A(n4231), .B(n4230), .S(n4443), .Z(n4232) );
  OAI21_X1 U4795 ( .B1(n4233), .B2(n4263), .A(n4232), .ZN(U3510) );
  INV_X1 U4796 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4235) );
  MUX2_X1 U4797 ( .A(n4235), .B(n4234), .S(n4443), .Z(n4236) );
  OAI21_X1 U4798 ( .B1(n4237), .B2(n4263), .A(n4236), .ZN(U3509) );
  MUX2_X1 U4799 ( .A(REG0_REG_22__SCAN_IN), .B(n4238), .S(n4443), .Z(U3508) );
  INV_X1 U4800 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4240) );
  MUX2_X1 U4801 ( .A(n4240), .B(n4239), .S(n4443), .Z(n4241) );
  OAI21_X1 U4802 ( .B1(n4242), .B2(n4263), .A(n4241), .ZN(U3507) );
  INV_X1 U4803 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4244) );
  MUX2_X1 U4804 ( .A(n4244), .B(n4243), .S(n4443), .Z(n4245) );
  OAI21_X1 U4805 ( .B1(n4246), .B2(n4263), .A(n4245), .ZN(U3506) );
  INV_X1 U4806 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4539) );
  MUX2_X1 U4807 ( .A(n4539), .B(n4247), .S(n4443), .Z(n4248) );
  OAI21_X1 U4808 ( .B1(n4249), .B2(n4263), .A(n4248), .ZN(U3505) );
  MUX2_X1 U4809 ( .A(REG0_REG_18__SCAN_IN), .B(n4250), .S(n4443), .Z(U3503) );
  INV_X1 U4810 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4252) );
  MUX2_X1 U4811 ( .A(n4252), .B(n4251), .S(n4443), .Z(n4253) );
  OAI21_X1 U4812 ( .B1(n4254), .B2(n4263), .A(n4253), .ZN(U3501) );
  MUX2_X1 U4813 ( .A(REG0_REG_16__SCAN_IN), .B(n4255), .S(n4443), .Z(U3499) );
  INV_X1 U4814 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4257) );
  MUX2_X1 U4815 ( .A(n4257), .B(n4256), .S(n4443), .Z(n4258) );
  OAI21_X1 U4816 ( .B1(n4259), .B2(n4263), .A(n4258), .ZN(U3497) );
  INV_X1 U4817 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4261) );
  MUX2_X1 U4818 ( .A(n4261), .B(n4260), .S(n4443), .Z(n4262) );
  OAI21_X1 U4819 ( .B1(n4264), .B2(n4263), .A(n4262), .ZN(U3495) );
  MUX2_X1 U4820 ( .A(n4265), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4821 ( .A(DATAI_28_), .B(n4266), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4822 ( .A(n4287), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4823 ( .A(DATAI_25_), .B(n2921), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4824 ( .A(n2721), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4825 ( .A(n4267), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4826 ( .A(n4268), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4827 ( .A(DATAI_20_), .B(n4269), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4828 ( .A(n4270), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U4829 ( .A(n4334), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U4830 ( .A(DATAI_6_), .B(n4271), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U4831 ( .A(n4272), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4832 ( .A(DATAI_4_), .B(n4273), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4833 ( .A(DATAI_3_), .B(n4274), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  INV_X1 U4834 ( .A(n4275), .ZN(n4276) );
  MUX2_X1 U4835 ( .A(DATAI_2_), .B(n4276), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  INV_X1 U4836 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U4837 ( .A1(n4279), .A2(n4282), .B1(n4278), .B2(n4277), .ZN(n4280)
         );
  OAI21_X1 U4838 ( .B1(n4278), .B2(n4566), .A(n4280), .ZN(U3260) );
  INV_X1 U4839 ( .A(n4281), .ZN(n4283) );
  OAI21_X1 U4840 ( .B1(n4063), .B2(n4285), .A(n4284), .ZN(U3261) );
  INV_X1 U4841 ( .A(n4289), .ZN(n4286) );
  OAI211_X1 U4842 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4287), .A(n4288), .B(n4286), 
        .ZN(n4293) );
  OAI22_X1 U4843 ( .A1(n4289), .A2(n4288), .B1(n4339), .B2(REG1_REG_0__SCAN_IN), .ZN(n4290) );
  INV_X1 U4844 ( .A(n4290), .ZN(n4292) );
  AOI22_X1 U4845 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4345), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4291) );
  OAI221_X1 U4846 ( .B1(n4401), .B2(n4293), .C1(n2133), .C2(n4292), .A(n4291), 
        .ZN(U3240) );
  AOI211_X1 U4847 ( .C1(n4296), .C2(n4295), .A(n4294), .B(n4339), .ZN(n4298)
         );
  AOI211_X1 U4848 ( .C1(n4345), .C2(ADDR_REG_10__SCAN_IN), .A(n4298), .B(n4297), .ZN(n4302) );
  OAI211_X1 U4849 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4300), .A(n4370), .B(n4299), .ZN(n4301) );
  OAI211_X1 U4850 ( .C1(n4375), .C2(n4303), .A(n4302), .B(n4301), .ZN(U3250)
         );
  AOI211_X1 U4851 ( .C1(n4306), .C2(n4305), .A(n4304), .B(n4339), .ZN(n4309)
         );
  INV_X1 U4852 ( .A(n4307), .ZN(n4308) );
  AOI211_X1 U4853 ( .C1(n4345), .C2(ADDR_REG_12__SCAN_IN), .A(n4309), .B(n4308), .ZN(n4313) );
  OAI211_X1 U4854 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4311), .A(n4370), .B(n4310), .ZN(n4312) );
  OAI211_X1 U4855 ( .C1(n4375), .C2(n4398), .A(n4313), .B(n4312), .ZN(U3252)
         );
  AOI211_X1 U4856 ( .C1(n4316), .C2(n4315), .A(n4314), .B(n4339), .ZN(n4318)
         );
  AOI211_X1 U4857 ( .C1(n4345), .C2(ADDR_REG_13__SCAN_IN), .A(n4318), .B(n4317), .ZN(n4323) );
  AOI22_X1 U4858 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4396), .B1(n4324), .B2(
        n3411), .ZN(n4321) );
  AOI21_X1 U4859 ( .B1(n4321), .B2(n4320), .A(n4325), .ZN(n4319) );
  OAI21_X1 U4860 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4322) );
  OAI211_X1 U4861 ( .C1(n4375), .C2(n4324), .A(n4323), .B(n4322), .ZN(U3253)
         );
  NAND2_X1 U4862 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4345), .ZN(n4338) );
  AOI211_X1 U4863 ( .C1(n4328), .C2(n4327), .A(n4326), .B(n4325), .ZN(n4333)
         );
  AOI211_X1 U4864 ( .C1(n4331), .C2(n4330), .A(n4329), .B(n4339), .ZN(n4332)
         );
  AOI211_X1 U4865 ( .C1(n4335), .C2(n4334), .A(n4333), .B(n4332), .ZN(n4337)
         );
  NAND3_X1 U4866 ( .A1(n4338), .A2(n4337), .A3(n4336), .ZN(U3254) );
  AOI211_X1 U4867 ( .C1(n4342), .C2(n4341), .A(n4340), .B(n4339), .ZN(n4343)
         );
  AOI211_X1 U4868 ( .C1(n4345), .C2(ADDR_REG_15__SCAN_IN), .A(n4344), .B(n4343), .ZN(n4351) );
  AOI21_X1 U4869 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4349) );
  NAND2_X1 U4870 ( .A1(n4370), .A2(n4349), .ZN(n4350) );
  OAI211_X1 U4871 ( .C1(n4375), .C2(n4352), .A(n4351), .B(n4350), .ZN(U3255)
         );
  AOI21_X1 U4872 ( .B1(n4345), .B2(ADDR_REG_16__SCAN_IN), .A(n4353), .ZN(n4361) );
  OAI21_X1 U4873 ( .B1(n4355), .B2(n4547), .A(n4354), .ZN(n4359) );
  OAI21_X1 U4874 ( .B1(n4357), .B2(n2899), .A(n4356), .ZN(n4358) );
  AOI22_X1 U4875 ( .A1(n4372), .A2(n4359), .B1(n4370), .B2(n4358), .ZN(n4360)
         );
  OAI211_X1 U4876 ( .C1(n4393), .C2(n4375), .A(n4361), .B(n4360), .ZN(U3256)
         );
  AOI21_X1 U4877 ( .B1(n4345), .B2(ADDR_REG_17__SCAN_IN), .A(n4362), .ZN(n4374) );
  OAI21_X1 U4878 ( .B1(n4365), .B2(n4364), .A(n4363), .ZN(n4371) );
  OAI21_X1 U4879 ( .B1(n4368), .B2(n4367), .A(n4366), .ZN(n4369) );
  AOI22_X1 U4880 ( .A1(n4372), .A2(n4371), .B1(n4370), .B2(n4369), .ZN(n4373)
         );
  OAI211_X1 U4881 ( .C1(n4391), .C2(n4375), .A(n4374), .B(n4373), .ZN(U3257)
         );
  INV_X1 U4882 ( .A(n4376), .ZN(n4379) );
  INV_X1 U4883 ( .A(n4377), .ZN(n4378) );
  AOI21_X1 U4884 ( .B1(n4380), .B2(n4379), .A(n4378), .ZN(n4385) );
  AOI22_X1 U4885 ( .A1(n4383), .A2(n4382), .B1(REG3_REG_0__SCAN_IN), .B2(n4381), .ZN(n4384) );
  OAI221_X1 U4886 ( .B1(n4063), .B2(n4385), .C1(n4278), .C2(n2301), .A(n4384), 
        .ZN(U3290) );
  INV_X1 U4887 ( .A(n4387), .ZN(n4386) );
  INV_X1 U4888 ( .A(D_REG_31__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U4889 ( .A1(n4386), .A2(n4519), .ZN(U3291) );
  AND2_X1 U4890 ( .A1(D_REG_30__SCAN_IN), .A2(n4387), .ZN(U3292) );
  AND2_X1 U4891 ( .A1(D_REG_29__SCAN_IN), .A2(n4387), .ZN(U3293) );
  AND2_X1 U4892 ( .A1(D_REG_28__SCAN_IN), .A2(n4387), .ZN(U3294) );
  AND2_X1 U4893 ( .A1(D_REG_27__SCAN_IN), .A2(n4387), .ZN(U3295) );
  AND2_X1 U4894 ( .A1(D_REG_26__SCAN_IN), .A2(n4387), .ZN(U3296) );
  INV_X1 U4895 ( .A(D_REG_25__SCAN_IN), .ZN(n4518) );
  NOR2_X1 U4896 ( .A1(n4386), .A2(n4518), .ZN(U3297) );
  INV_X1 U4897 ( .A(D_REG_24__SCAN_IN), .ZN(n4506) );
  NOR2_X1 U4898 ( .A1(n4386), .A2(n4506), .ZN(U3298) );
  AND2_X1 U4899 ( .A1(D_REG_23__SCAN_IN), .A2(n4387), .ZN(U3299) );
  AND2_X1 U4900 ( .A1(D_REG_22__SCAN_IN), .A2(n4387), .ZN(U3300) );
  AND2_X1 U4901 ( .A1(D_REG_21__SCAN_IN), .A2(n4387), .ZN(U3301) );
  AND2_X1 U4902 ( .A1(D_REG_20__SCAN_IN), .A2(n4387), .ZN(U3302) );
  AND2_X1 U4903 ( .A1(D_REG_19__SCAN_IN), .A2(n4387), .ZN(U3303) );
  AND2_X1 U4904 ( .A1(D_REG_18__SCAN_IN), .A2(n4387), .ZN(U3304) );
  AND2_X1 U4905 ( .A1(D_REG_17__SCAN_IN), .A2(n4387), .ZN(U3305) );
  AND2_X1 U4906 ( .A1(D_REG_16__SCAN_IN), .A2(n4387), .ZN(U3306) );
  AND2_X1 U4907 ( .A1(D_REG_15__SCAN_IN), .A2(n4387), .ZN(U3307) );
  INV_X1 U4908 ( .A(D_REG_14__SCAN_IN), .ZN(n4505) );
  NOR2_X1 U4909 ( .A1(n4386), .A2(n4505), .ZN(U3308) );
  AND2_X1 U4910 ( .A1(D_REG_13__SCAN_IN), .A2(n4387), .ZN(U3309) );
  AND2_X1 U4911 ( .A1(D_REG_12__SCAN_IN), .A2(n4387), .ZN(U3310) );
  INV_X1 U4912 ( .A(D_REG_11__SCAN_IN), .ZN(n4508) );
  NOR2_X1 U4913 ( .A1(n4386), .A2(n4508), .ZN(U3311) );
  AND2_X1 U4914 ( .A1(D_REG_10__SCAN_IN), .A2(n4387), .ZN(U3312) );
  AND2_X1 U4915 ( .A1(D_REG_9__SCAN_IN), .A2(n4387), .ZN(U3313) );
  AND2_X1 U4916 ( .A1(D_REG_8__SCAN_IN), .A2(n4387), .ZN(U3314) );
  AND2_X1 U4917 ( .A1(D_REG_7__SCAN_IN), .A2(n4387), .ZN(U3315) );
  AND2_X1 U4918 ( .A1(D_REG_6__SCAN_IN), .A2(n4387), .ZN(U3316) );
  AND2_X1 U4919 ( .A1(D_REG_5__SCAN_IN), .A2(n4387), .ZN(U3317) );
  AND2_X1 U4920 ( .A1(D_REG_4__SCAN_IN), .A2(n4387), .ZN(U3318) );
  AND2_X1 U4921 ( .A1(D_REG_3__SCAN_IN), .A2(n4387), .ZN(U3319) );
  AND2_X1 U4922 ( .A1(D_REG_2__SCAN_IN), .A2(n4387), .ZN(U3320) );
  OAI21_X1 U4923 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4388), .ZN(
        n4389) );
  INV_X1 U4924 ( .A(n4389), .ZN(U3329) );
  AOI22_X1 U4925 ( .A1(STATE_REG_SCAN_IN), .A2(n4391), .B1(n4390), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4926 ( .A(DATAI_16_), .ZN(n4392) );
  AOI22_X1 U4927 ( .A1(STATE_REG_SCAN_IN), .A2(n4393), .B1(n4392), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U4928 ( .A1(U3149), .A2(n4394), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4395) );
  INV_X1 U4929 ( .A(n4395), .ZN(U3337) );
  OAI22_X1 U4930 ( .A1(U3149), .A2(n4396), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4397) );
  INV_X1 U4931 ( .A(n4397), .ZN(U3339) );
  AOI22_X1 U4932 ( .A1(STATE_REG_SCAN_IN), .A2(n4398), .B1(n2495), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U4933 ( .A1(U3149), .A2(n4399), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4400) );
  INV_X1 U4934 ( .A(n4400), .ZN(U3342) );
  OAI22_X1 U4935 ( .A1(U3149), .A2(n4401), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4402) );
  INV_X1 U4936 ( .A(n4402), .ZN(U3352) );
  INV_X1 U4937 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U4938 ( .A1(n4443), .A2(n4403), .B1(n4522), .B2(n4441), .ZN(U3467)
         );
  INV_X1 U4939 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U4940 ( .A1(n4443), .A2(n4404), .B1(n4521), .B2(n4441), .ZN(U3469)
         );
  NOR2_X1 U4941 ( .A1(n4405), .A2(n4435), .ZN(n4407) );
  AOI211_X1 U4942 ( .C1(n4440), .C2(n4408), .A(n4407), .B(n4406), .ZN(n4445)
         );
  INV_X1 U4943 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4944 ( .A1(n4443), .A2(n4445), .B1(n4409), .B2(n4441), .ZN(U3473)
         );
  INV_X1 U4945 ( .A(n4410), .ZN(n4415) );
  INV_X1 U4946 ( .A(n4411), .ZN(n4413) );
  AOI211_X1 U4947 ( .C1(n4415), .C2(n4414), .A(n4413), .B(n4412), .ZN(n4447)
         );
  INV_X1 U4948 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U4949 ( .A1(n4443), .A2(n4447), .B1(n4416), .B2(n4441), .ZN(U3475)
         );
  NOR2_X1 U4950 ( .A1(n4417), .A2(n4422), .ZN(n4420) );
  INV_X1 U4951 ( .A(n4418), .ZN(n4419) );
  AOI211_X1 U4952 ( .C1(n4440), .C2(n4421), .A(n4420), .B(n4419), .ZN(n4448)
         );
  INV_X1 U4953 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U4954 ( .A1(n4443), .A2(n4448), .B1(n4525), .B2(n4441), .ZN(U3477)
         );
  NOR2_X1 U4955 ( .A1(n4423), .A2(n4422), .ZN(n4426) );
  AOI211_X1 U4956 ( .C1(n4426), .C2(n3231), .A(n4425), .B(n4424), .ZN(n4449)
         );
  INV_X1 U4957 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4427) );
  AOI22_X1 U4958 ( .A1(n4443), .A2(n4449), .B1(n4427), .B2(n4441), .ZN(U3481)
         );
  NAND2_X1 U4959 ( .A1(n4429), .A2(n4428), .ZN(n4433) );
  OR2_X1 U4960 ( .A1(n4431), .A2(n4430), .ZN(n4432) );
  INV_X1 U4961 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U4962 ( .A1(n4443), .A2(n4450), .B1(n4524), .B2(n4441), .ZN(U3485)
         );
  NOR2_X1 U4963 ( .A1(n4436), .A2(n4435), .ZN(n4438) );
  AOI211_X1 U4964 ( .C1(n4440), .C2(n4439), .A(n4438), .B(n4437), .ZN(n4452)
         );
  INV_X1 U4965 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U4966 ( .A1(n4443), .A2(n4452), .B1(n4442), .B2(n4441), .ZN(U3489)
         );
  INV_X1 U4967 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U4968 ( .A1(n4453), .A2(n4445), .B1(n4444), .B2(n4451), .ZN(U3521)
         );
  INV_X1 U4969 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4446) );
  AOI22_X1 U4970 ( .A1(n4453), .A2(n4447), .B1(n4446), .B2(n4451), .ZN(U3522)
         );
  INV_X1 U4971 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U4972 ( .A1(n4453), .A2(n4448), .B1(n4541), .B2(n4451), .ZN(U3523)
         );
  AOI22_X1 U4973 ( .A1(n4453), .A2(n4449), .B1(n4545), .B2(n4451), .ZN(U3525)
         );
  AOI22_X1 U4974 ( .A1(n4453), .A2(n4450), .B1(n3012), .B2(n4451), .ZN(U3527)
         );
  AOI22_X1 U4975 ( .A1(n4453), .A2(n4452), .B1(n3098), .B2(n4451), .ZN(U3529)
         );
  NAND4_X1 U4976 ( .A1(REG1_REG_6__SCAN_IN), .A2(REG0_REG_31__SCAN_IN), .A3(
        n4539), .A4(n4541), .ZN(n4476) );
  NOR4_X1 U4977 ( .A1(REG2_REG_12__SCAN_IN), .A2(REG2_REG_3__SCAN_IN), .A3(
        n2899), .A4(n4554), .ZN(n4456) );
  NOR3_X1 U4978 ( .A1(REG2_REG_22__SCAN_IN), .A2(REG2_REG_19__SCAN_IN), .A3(
        REG2_REG_18__SCAN_IN), .ZN(n4455) );
  NOR4_X1 U4979 ( .A1(REG1_REG_16__SCAN_IN), .A2(REG1_REG_7__SCAN_IN), .A3(
        n4548), .A4(n4544), .ZN(n4454) );
  NAND4_X1 U4980 ( .A1(REG2_REG_24__SCAN_IN), .A2(n4456), .A3(n4455), .A4(
        n4454), .ZN(n4475) );
  INV_X1 U4981 ( .A(DATAI_25_), .ZN(n4484) );
  NOR4_X1 U4982 ( .A1(DATAI_6_), .A2(n4481), .A3(n4484), .A4(n4485), .ZN(n4459) );
  NOR4_X1 U4983 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .A3(
        IR_REG_9__SCAN_IN), .A4(IR_REG_4__SCAN_IN), .ZN(n4458) );
  NOR4_X1 U4984 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .A3(
        n4496), .A4(n4495), .ZN(n4457) );
  NAND4_X1 U4985 ( .A1(REG3_REG_7__SCAN_IN), .A2(n4459), .A3(n4458), .A4(n4457), .ZN(n4460) );
  OR4_X1 U4986 ( .A1(n4460), .A2(DATAI_4_), .A3(DATAI_2_), .A4(DATAI_3_), .ZN(
        n4474) );
  NOR4_X1 U4987 ( .A1(DATAO_REG_3__SCAN_IN), .A2(ADDR_REG_1__SCAN_IN), .A3(
        n4584), .A4(n4581), .ZN(n4472) );
  NOR4_X1 U4988 ( .A1(REG2_REG_28__SCAN_IN), .A2(REG2_REG_31__SCAN_IN), .A3(
        ADDR_REG_16__SCAN_IN), .A4(ADDR_REG_13__SCAN_IN), .ZN(n4471) );
  NAND4_X1 U4989 ( .A1(DATAO_REG_18__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .A3(
        n4587), .A4(n4590), .ZN(n4462) );
  NAND3_X1 U4990 ( .A1(ADDR_REG_12__SCAN_IN), .A2(ADDR_REG_5__SCAN_IN), .A3(
        ADDR_REG_7__SCAN_IN), .ZN(n4461) );
  NOR3_X1 U4991 ( .A1(ADDR_REG_3__SCAN_IN), .A2(n4462), .A3(n4461), .ZN(n4470)
         );
  AND4_X1 U4992 ( .A1(D_REG_31__SCAN_IN), .A2(n4521), .A3(n4518), .A4(n4522), 
        .ZN(n4468) );
  AND4_X1 U4993 ( .A1(REG0_REG_10__SCAN_IN), .A2(REG0_REG_5__SCAN_IN), .A3(
        n4527), .A4(n4524), .ZN(n4467) );
  NAND4_X1 U4994 ( .A1(n4463), .A2(IR_REG_16__SCAN_IN), .A3(IR_REG_19__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n4465) );
  NAND3_X1 U4995 ( .A1(n4507), .A2(IR_REG_20__SCAN_IN), .A3(D_REG_11__SCAN_IN), 
        .ZN(n4464) );
  NOR2_X1 U4996 ( .A1(n4465), .A2(n4464), .ZN(n4466) );
  AND4_X1 U4997 ( .A1(n4468), .A2(n4467), .A3(n4466), .A4(n4505), .ZN(n4469)
         );
  NAND4_X1 U4998 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(n4473)
         );
  NOR4_X1 U4999 ( .A1(n4476), .A2(n4475), .A3(n4474), .A4(n4473), .ZN(n4605)
         );
  INV_X1 U5000 ( .A(DATAI_4_), .ZN(n4479) );
  INV_X1 U5001 ( .A(DATAI_3_), .ZN(n4478) );
  AOI22_X1 U5002 ( .A1(n4479), .A2(keyinput24), .B1(keyinput45), .B2(n4478), 
        .ZN(n4477) );
  OAI221_X1 U5003 ( .B1(n4479), .B2(keyinput24), .C1(n4478), .C2(keyinput45), 
        .A(n4477), .ZN(n4491) );
  INV_X1 U5004 ( .A(DATAI_6_), .ZN(n4482) );
  AOI22_X1 U5005 ( .A1(n4482), .A2(keyinput4), .B1(n4481), .B2(keyinput9), 
        .ZN(n4480) );
  OAI221_X1 U5006 ( .B1(n4482), .B2(keyinput4), .C1(n4481), .C2(keyinput9), 
        .A(n4480), .ZN(n4490) );
  AOI22_X1 U5007 ( .A1(n4485), .A2(keyinput18), .B1(n4484), .B2(keyinput11), 
        .ZN(n4483) );
  OAI221_X1 U5008 ( .B1(n4485), .B2(keyinput18), .C1(n4484), .C2(keyinput11), 
        .A(n4483), .ZN(n4489) );
  XNOR2_X1 U5009 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput60), .ZN(n4487) );
  XNOR2_X1 U5010 ( .A(DATAI_2_), .B(keyinput51), .ZN(n4486) );
  NAND2_X1 U5011 ( .A1(n4487), .A2(n4486), .ZN(n4488) );
  NOR4_X1 U5012 ( .A1(n4491), .A2(n4490), .A3(n4489), .A4(n4488), .ZN(n4536)
         );
  AOI22_X1 U5013 ( .A1(n2572), .A2(keyinput13), .B1(keyinput61), .B2(n4493), 
        .ZN(n4492) );
  OAI221_X1 U5014 ( .B1(n2572), .B2(keyinput13), .C1(n4493), .C2(keyinput61), 
        .A(n4492), .ZN(n4503) );
  AOI22_X1 U5015 ( .A1(n4496), .A2(keyinput57), .B1(keyinput21), .B2(n4495), 
        .ZN(n4494) );
  OAI221_X1 U5016 ( .B1(n4496), .B2(keyinput57), .C1(n4495), .C2(keyinput21), 
        .A(n4494), .ZN(n4502) );
  XNOR2_X1 U5017 ( .A(IR_REG_4__SCAN_IN), .B(keyinput47), .ZN(n4500) );
  XNOR2_X1 U5018 ( .A(IR_REG_9__SCAN_IN), .B(keyinput3), .ZN(n4499) );
  XNOR2_X1 U5019 ( .A(IR_REG_14__SCAN_IN), .B(keyinput56), .ZN(n4498) );
  XNOR2_X1 U5020 ( .A(IR_REG_11__SCAN_IN), .B(keyinput44), .ZN(n4497) );
  NAND4_X1 U5021 ( .A1(n4500), .A2(n4499), .A3(n4498), .A4(n4497), .ZN(n4501)
         );
  NOR3_X1 U5022 ( .A1(n4503), .A2(n4502), .A3(n4501), .ZN(n4535) );
  AOI22_X1 U5023 ( .A1(n4506), .A2(keyinput46), .B1(keyinput49), .B2(n4505), 
        .ZN(n4504) );
  OAI221_X1 U5024 ( .B1(n4506), .B2(keyinput46), .C1(n4505), .C2(keyinput49), 
        .A(n4504), .ZN(n4516) );
  XNOR2_X1 U5025 ( .A(n4507), .B(keyinput50), .ZN(n4515) );
  XNOR2_X1 U5026 ( .A(keyinput63), .B(n4508), .ZN(n4514) );
  XNOR2_X1 U5027 ( .A(IR_REG_18__SCAN_IN), .B(keyinput26), .ZN(n4512) );
  XNOR2_X1 U5028 ( .A(IR_REG_16__SCAN_IN), .B(keyinput23), .ZN(n4511) );
  XNOR2_X1 U5029 ( .A(IR_REG_20__SCAN_IN), .B(keyinput36), .ZN(n4510) );
  XNOR2_X1 U5030 ( .A(IR_REG_19__SCAN_IN), .B(keyinput25), .ZN(n4509) );
  NAND4_X1 U5031 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n4513)
         );
  NOR4_X1 U5032 ( .A1(n4516), .A2(n4515), .A3(n4514), .A4(n4513), .ZN(n4534)
         );
  AOI22_X1 U5033 ( .A1(n4519), .A2(keyinput37), .B1(keyinput27), .B2(n4518), 
        .ZN(n4517) );
  OAI221_X1 U5034 ( .B1(n4519), .B2(keyinput37), .C1(n4518), .C2(keyinput27), 
        .A(n4517), .ZN(n4532) );
  AOI22_X1 U5035 ( .A1(n4522), .A2(keyinput32), .B1(n4521), .B2(keyinput30), 
        .ZN(n4520) );
  OAI221_X1 U5036 ( .B1(n4522), .B2(keyinput32), .C1(n4521), .C2(keyinput30), 
        .A(n4520), .ZN(n4531) );
  AOI22_X1 U5037 ( .A1(n4525), .A2(keyinput15), .B1(n4524), .B2(keyinput34), 
        .ZN(n4523) );
  OAI221_X1 U5038 ( .B1(n4525), .B2(keyinput15), .C1(n4524), .C2(keyinput34), 
        .A(n4523), .ZN(n4530) );
  AOI22_X1 U5039 ( .A1(n4528), .A2(keyinput31), .B1(n4527), .B2(keyinput22), 
        .ZN(n4526) );
  OAI221_X1 U5040 ( .B1(n4528), .B2(keyinput31), .C1(n4527), .C2(keyinput22), 
        .A(n4526), .ZN(n4529) );
  NOR4_X1 U5041 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(n4533)
         );
  NAND4_X1 U5042 ( .A1(n4536), .A2(n4535), .A3(n4534), .A4(n4533), .ZN(n4601)
         );
  AOI22_X1 U5043 ( .A1(n4539), .A2(keyinput28), .B1(keyinput41), .B2(n4538), 
        .ZN(n4537) );
  OAI221_X1 U5044 ( .B1(n4539), .B2(keyinput28), .C1(n4538), .C2(keyinput41), 
        .A(n4537), .ZN(n4552) );
  AOI22_X1 U5045 ( .A1(n4542), .A2(keyinput12), .B1(keyinput48), .B2(n4541), 
        .ZN(n4540) );
  OAI221_X1 U5046 ( .B1(n4542), .B2(keyinput12), .C1(n4541), .C2(keyinput48), 
        .A(n4540), .ZN(n4551) );
  AOI22_X1 U5047 ( .A1(n4545), .A2(keyinput0), .B1(n4544), .B2(keyinput62), 
        .ZN(n4543) );
  OAI221_X1 U5048 ( .B1(n4545), .B2(keyinput0), .C1(n4544), .C2(keyinput62), 
        .A(n4543), .ZN(n4550) );
  AOI22_X1 U5049 ( .A1(n4548), .A2(keyinput53), .B1(n4547), .B2(keyinput52), 
        .ZN(n4546) );
  OAI221_X1 U5050 ( .B1(n4548), .B2(keyinput53), .C1(n4547), .C2(keyinput52), 
        .A(n4546), .ZN(n4549) );
  NOR4_X1 U5051 ( .A1(n4552), .A2(n4551), .A3(n4550), .A4(n4549), .ZN(n4599)
         );
  AOI22_X1 U5052 ( .A1(n2339), .A2(keyinput29), .B1(n4554), .B2(keyinput19), 
        .ZN(n4553) );
  OAI221_X1 U5053 ( .B1(n2339), .B2(keyinput29), .C1(n4554), .C2(keyinput19), 
        .A(n4553), .ZN(n4564) );
  AOI22_X1 U5054 ( .A1(n2899), .A2(keyinput14), .B1(keyinput38), .B2(n2051), 
        .ZN(n4555) );
  OAI221_X1 U5055 ( .B1(n2899), .B2(keyinput14), .C1(n2051), .C2(keyinput38), 
        .A(n4555), .ZN(n4563) );
  INV_X1 U5056 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5057 ( .A1(n4558), .A2(keyinput33), .B1(keyinput54), .B2(n4557), 
        .ZN(n4556) );
  OAI221_X1 U5058 ( .B1(n4558), .B2(keyinput33), .C1(n4557), .C2(keyinput54), 
        .A(n4556), .ZN(n4562) );
  INV_X1 U5059 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5060 ( .A1(n4017), .A2(keyinput10), .B1(keyinput58), .B2(n4560), 
        .ZN(n4559) );
  OAI221_X1 U5061 ( .B1(n4017), .B2(keyinput10), .C1(n4560), .C2(keyinput58), 
        .A(n4559), .ZN(n4561) );
  NOR4_X1 U5062 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), .ZN(n4598)
         );
  AOI22_X1 U5063 ( .A1(n3472), .A2(keyinput55), .B1(keyinput20), .B2(n4566), 
        .ZN(n4565) );
  OAI221_X1 U5064 ( .B1(n3472), .B2(keyinput55), .C1(n4566), .C2(keyinput20), 
        .A(n4565), .ZN(n4579) );
  INV_X1 U5065 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4569) );
  INV_X1 U5066 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5067 ( .A1(n4569), .A2(keyinput8), .B1(keyinput16), .B2(n4568), 
        .ZN(n4567) );
  OAI221_X1 U5068 ( .B1(n4569), .B2(keyinput8), .C1(n4568), .C2(keyinput16), 
        .A(n4567), .ZN(n4578) );
  INV_X1 U5069 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4572) );
  INV_X1 U5070 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5071 ( .A1(n4572), .A2(keyinput35), .B1(n4571), .B2(keyinput59), 
        .ZN(n4570) );
  OAI221_X1 U5072 ( .B1(n4572), .B2(keyinput35), .C1(n4571), .C2(keyinput59), 
        .A(n4570), .ZN(n4577) );
  INV_X1 U5073 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4575) );
  INV_X1 U5074 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5075 ( .A1(n4575), .A2(keyinput40), .B1(keyinput42), .B2(n4574), 
        .ZN(n4573) );
  OAI221_X1 U5076 ( .B1(n4575), .B2(keyinput40), .C1(n4574), .C2(keyinput42), 
        .A(n4573), .ZN(n4576) );
  NOR4_X1 U5077 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4597)
         );
  INV_X1 U5078 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4582) );
  AOI22_X1 U5079 ( .A1(n4582), .A2(keyinput1), .B1(n4581), .B2(keyinput39), 
        .ZN(n4580) );
  OAI221_X1 U5080 ( .B1(n4582), .B2(keyinput1), .C1(n4581), .C2(keyinput39), 
        .A(n4580), .ZN(n4595) );
  AOI22_X1 U5081 ( .A1(n4585), .A2(keyinput5), .B1(keyinput2), .B2(n4584), 
        .ZN(n4583) );
  OAI221_X1 U5082 ( .B1(n4585), .B2(keyinput5), .C1(n4584), .C2(keyinput2), 
        .A(n4583), .ZN(n4594) );
  AOI22_X1 U5083 ( .A1(n4588), .A2(keyinput17), .B1(keyinput43), .B2(n4587), 
        .ZN(n4586) );
  OAI221_X1 U5084 ( .B1(n4588), .B2(keyinput17), .C1(n4587), .C2(keyinput43), 
        .A(n4586), .ZN(n4593) );
  AOI22_X1 U5085 ( .A1(n4591), .A2(keyinput6), .B1(keyinput7), .B2(n4590), 
        .ZN(n4589) );
  OAI221_X1 U5086 ( .B1(n4591), .B2(keyinput6), .C1(n4590), .C2(keyinput7), 
        .A(n4589), .ZN(n4592) );
  NOR4_X1 U5087 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NAND4_X1 U5088 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4600)
         );
  NOR2_X1 U5089 ( .A1(n4601), .A2(n4600), .ZN(n4603) );
  MUX2_X1 U5090 ( .A(n2285), .B(DATAI_1_), .S(U3149), .Z(n4602) );
  XNOR2_X1 U5091 ( .A(n4603), .B(n4602), .ZN(n4604) );
  XNOR2_X1 U5092 ( .A(n4605), .B(n4604), .ZN(U3351) );
endmodule

