

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5131, n5132, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195;

  OR2_X1 U5195 ( .A1(n6410), .A2(n5593), .ZN(n5590) );
  CLKBUF_X1 U5196 ( .A(n5926), .Z(n8848) );
  INV_X1 U5197 ( .A(n6444), .ZN(n6579) );
  CLKBUF_X2 U5199 ( .A(n5944), .Z(n5960) );
  AND4_X1 U5200 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n6997)
         );
  AND2_X2 U5201 ( .A1(n5870), .A2(n9223), .ZN(n8847) );
  NAND2_X1 U5203 ( .A1(n5869), .A2(n5868), .ZN(n5872) );
  NAND2_X2 U5204 ( .A1(n6429), .A2(n6624), .ZN(n6637) );
  INV_X1 U5205 ( .A(n6637), .ZN(n6455) );
  INV_X1 U5206 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6061) );
  INV_X1 U5207 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U5208 ( .A1(n7158), .A2(n5131), .ZN(n7130) );
  INV_X1 U5210 ( .A(n7156), .ZN(n7548) );
  XNOR2_X1 U5211 ( .A(n8196), .B(n8214), .ZN(n11080) );
  INV_X1 U5212 ( .A(n5134), .ZN(n6258) );
  NAND2_X1 U5213 ( .A1(n10679), .A2(n10685), .ZN(n9019) );
  AND2_X1 U5214 ( .A1(n5940), .A2(n5436), .ZN(n5941) );
  INV_X2 U5215 ( .A(n7130), .ZN(n7534) );
  AND2_X1 U5216 ( .A1(n9016), .A2(n5604), .ZN(n9045) );
  INV_X1 U5217 ( .A(n7153), .ZN(n8787) );
  INV_X1 U5218 ( .A(n7250), .ZN(n8795) );
  XNOR2_X2 U5219 ( .A(n9189), .B(n9188), .ZN(n9204) );
  OAI21_X2 U5220 ( .B1(n9897), .B2(n5331), .A(n5220), .ZN(n5337) );
  AOI21_X2 U5221 ( .B1(n5164), .B2(n5408), .A(n5407), .ZN(n5406) );
  NAND2_X2 U5222 ( .A1(n5922), .A2(n5921), .ZN(n6426) );
  XNOR2_X1 U5223 ( .A(n7112), .B(n7111), .ZN(n5131) );
  OAI21_X2 U5224 ( .B1(n6239), .B2(SI_22_), .A(n5818), .ZN(n6252) );
  NOR2_X2 U5225 ( .A1(n10930), .A2(n10931), .ZN(n10929) );
  NOR2_X2 U5226 ( .A1(n8361), .A2(n9451), .ZN(n9472) );
  XNOR2_X2 U5227 ( .A(n7607), .B(n7747), .ZN(n7210) );
  AOI21_X2 U5228 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n11061), .A(n11068), .ZN(
        n7607) );
  AOI21_X2 U5229 ( .B1(n6794), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6793), .ZN(
        n6929) );
  NOR2_X2 U5230 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  NAND2_X1 U5231 ( .A1(n8410), .A2(n8409), .ZN(n8700) );
  NAND2_X1 U5232 ( .A1(n8931), .A2(n8895), .ZN(n8872) );
  INV_X2 U5233 ( .A(n11160), .ZN(n7821) );
  NAND2_X1 U5234 ( .A1(n6065), .A2(n6064), .ZN(n7744) );
  AOI21_X1 U5235 ( .B1(n7533), .B2(n8854), .A(n5714), .ZN(n11129) );
  NAND2_X1 U5236 ( .A1(n10356), .A2(n7034), .ZN(n9057) );
  NAND2_X1 U5237 ( .A1(n9058), .A2(n8905), .ZN(n6866) );
  INV_X2 U5238 ( .A(n6985), .ZN(n7034) );
  INV_X2 U5239 ( .A(n6258), .ZN(n6289) );
  BUF_X1 U5240 ( .A(n6195), .Z(n5135) );
  INV_X1 U5241 ( .A(n7532), .ZN(n7524) );
  AND2_X1 U5242 ( .A1(n7130), .A2(n8701), .ZN(n7532) );
  INV_X2 U5243 ( .A(n6964), .ZN(n6877) );
  OR2_X1 U5244 ( .A1(n8853), .A2(n6731), .ZN(n5393) );
  CLKBUF_X1 U5245 ( .A(n6325), .Z(n5139) );
  INV_X1 U5246 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10312) );
  AND2_X1 U5247 ( .A1(n5596), .A2(n5158), .ZN(n5591) );
  NAND2_X1 U5248 ( .A1(n8794), .A2(n5349), .ZN(n5348) );
  OR2_X1 U5249 ( .A1(n5351), .A2(n8748), .ZN(n5349) );
  AOI22_X1 U5250 ( .A1(n9501), .A2(n9643), .B1(n7162), .B2(n9716), .ZN(n9710)
         );
  NOR2_X1 U5251 ( .A1(n5272), .A2(n5271), .ZN(n5270) );
  NOR2_X1 U5252 ( .A1(n5315), .A2(n5314), .ZN(n9519) );
  AND2_X1 U5253 ( .A1(n10613), .A2(n8884), .ZN(n10587) );
  INV_X1 U5254 ( .A(n10500), .ZN(n10508) );
  NAND2_X1 U5255 ( .A1(n9262), .A2(n9154), .ZN(n9335) );
  NAND2_X1 U5256 ( .A1(n9852), .A2(n6564), .ZN(n9910) );
  NOR2_X1 U5257 ( .A1(n9527), .A2(n9526), .ZN(n5315) );
  NAND2_X1 U5258 ( .A1(n5640), .A2(n6288), .ZN(n6680) );
  AND2_X1 U5259 ( .A1(n5281), .A2(n5216), .ZN(n9537) );
  NAND2_X1 U5260 ( .A1(n10641), .A2(n10642), .ZN(n10640) );
  OR2_X1 U5261 ( .A1(n9576), .A2(n5282), .ZN(n5281) );
  NOR2_X1 U5262 ( .A1(n8771), .A2(n5733), .ZN(n5728) );
  AND2_X1 U5263 ( .A1(n5414), .A2(n5420), .ZN(n5413) );
  XNOR2_X1 U5264 ( .A(n6267), .B(n6284), .ZN(n8674) );
  NAND2_X1 U5265 ( .A1(n5886), .A2(n5885), .ZN(n10538) );
  NAND2_X1 U5266 ( .A1(n5725), .A2(n5724), .ZN(n9608) );
  AND2_X1 U5267 ( .A1(n8773), .A2(n8772), .ZN(n9553) );
  NAND2_X1 U5268 ( .A1(n9642), .A2(n5306), .ZN(n5303) );
  XNOR2_X1 U5269 ( .A(n8360), .B(n9457), .ZN(n9452) );
  AND2_X1 U5270 ( .A1(n5484), .A2(n5483), .ZN(n8360) );
  NAND2_X1 U5271 ( .A1(n5883), .A2(n5829), .ZN(n6391) );
  AND2_X1 U5272 ( .A1(n8760), .A2(n8759), .ZN(n9638) );
  NAND2_X1 U5273 ( .A1(n5880), .A2(n5828), .ZN(n5883) );
  NAND2_X1 U5274 ( .A1(n6254), .A2(n6253), .ZN(n10579) );
  OR2_X1 U5275 ( .A1(n9423), .A2(n8358), .ZN(n5486) );
  NOR2_X1 U5276 ( .A1(n9415), .A2(n9414), .ZN(n9413) );
  NAND2_X1 U5277 ( .A1(n5266), .A2(n5265), .ZN(n8051) );
  AOI21_X1 U5278 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10948), .A(n10941), .ZN(
        n10901) );
  NAND2_X1 U5279 ( .A1(n6312), .A2(n5587), .ZN(n7664) );
  NAND2_X1 U5280 ( .A1(n7933), .A2(n5277), .ZN(n8023) );
  NOR2_X1 U5281 ( .A1(n8309), .A2(n5225), .ZN(n8351) );
  INV_X1 U5282 ( .A(n6546), .ZN(n10767) );
  NAND2_X1 U5283 ( .A1(n6162), .A2(n6161), .ZN(n10759) );
  AND2_X1 U5284 ( .A1(n9084), .A2(n8942), .ZN(n8943) );
  NOR2_X1 U5285 ( .A1(n8219), .A2(n8218), .ZN(n8309) );
  NAND2_X1 U5286 ( .A1(n6969), .A2(n5994), .ZN(n7027) );
  NAND2_X1 U5287 ( .A1(n6132), .A2(n6131), .ZN(n6540) );
  AND2_X1 U5288 ( .A1(n5673), .A2(n5206), .ZN(n7752) );
  OR2_X1 U5289 ( .A1(n7821), .A2(n10349), .ZN(n8931) );
  NOR2_X1 U5290 ( .A1(n7356), .A2(n8009), .ZN(n5435) );
  AND4_X1 U5291 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .ZN(n9246)
         );
  OAI21_X1 U5292 ( .B1(n7657), .B2(n7656), .A(n7655), .ZN(n7789) );
  NAND4_X2 U5293 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n9593)
         );
  INV_X2 U5294 ( .A(n10659), .ZN(n10632) );
  INV_X1 U5295 ( .A(n11129), .ZN(n7418) );
  OAI211_X1 U5296 ( .C1(n7524), .C2(n7527), .A(n7526), .B(n7525), .ZN(n11117)
         );
  INV_X2 U5297 ( .A(n8232), .ZN(n5132) );
  NAND2_X1 U5298 ( .A1(n6003), .A2(n6002), .ZN(n6005) );
  INV_X1 U5299 ( .A(n6875), .ZN(n7014) );
  NAND2_X1 U5300 ( .A1(n6875), .A2(n5917), .ZN(n9058) );
  NAND2_X1 U5301 ( .A1(n6422), .A2(n5322), .ZN(n6429) );
  AND2_X2 U5302 ( .A1(n6705), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3973) );
  AND4_X2 U5303 ( .A1(n7129), .A2(n7128), .A3(n7127), .A4(n7126), .ZN(n7311)
         );
  OAI211_X1 U5304 ( .C1(n7524), .C2(n7316), .A(n7315), .B(n7314), .ZN(n7562)
         );
  NAND4_X1 U5305 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7305)
         );
  NOR2_X2 U5306 ( .A1(n8464), .A2(n7161), .ZN(n7162) );
  CLKBUF_X2 U5307 ( .A(n6195), .Z(n5134) );
  NOR2_X2 U5308 ( .A1(n8464), .A2(n7336), .ZN(n7160) );
  AOI21_X1 U5309 ( .B1(n11011), .B2(n5474), .A(n5473), .ZN(n11027) );
  NAND2_X1 U5310 ( .A1(n7175), .A2(n7174), .ZN(n7274) );
  AND2_X2 U5311 ( .A1(n7098), .A2(n7097), .ZN(n7539) );
  XNOR2_X1 U5312 ( .A(n7147), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7189) );
  AND2_X2 U5313 ( .A1(n7098), .A2(n7099), .ZN(n7155) );
  XNOR2_X1 U5314 ( .A(n7150), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8746) );
  NAND2_X2 U5315 ( .A1(n6707), .A2(n7113), .ZN(n6396) );
  BUF_X1 U5316 ( .A(n6325), .Z(n5138) );
  XNOR2_X1 U5317 ( .A(n7151), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7153) );
  NAND2_X1 U5318 ( .A1(n5867), .A2(n5866), .ZN(n5869) );
  NAND2_X1 U5319 ( .A1(n7144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U5320 ( .A1(n6334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U5321 ( .A1(n5772), .A2(SI_4_), .ZN(n5774) );
  OR2_X1 U5322 ( .A1(n7946), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U5323 ( .A(n6699), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8828) );
  AND2_X1 U5324 ( .A1(n6773), .A2(n5676), .ZN(n7395) );
  NOR2_X1 U5325 ( .A1(n5678), .A2(n7141), .ZN(n5676) );
  INV_X4 U5326 ( .A(n7113), .ZN(n5823) );
  AND2_X1 U5327 ( .A1(n5386), .A2(n5385), .ZN(n5384) );
  XNOR2_X1 U5328 ( .A(n6742), .B(P2_IR_REG_3__SCAN_IN), .ZN(n11016) );
  INV_X2 U5329 ( .A(n5771), .ZN(n7113) );
  OR2_X1 U5330 ( .A1(n7140), .A2(n7139), .ZN(n7141) );
  AND4_X1 U5331 ( .A1(n6691), .A2(n5748), .A3(n6690), .A4(n6689), .ZN(n6692)
         );
  AND2_X2 U5332 ( .A1(n5637), .A2(n5636), .ZN(n5771) );
  OR2_X1 U5333 ( .A1(n6936), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7140) );
  AND4_X1 U5334 ( .A1(n10284), .A2(n5971), .A3(n6058), .A4(n6061), .ZN(n5832)
         );
  NAND2_X1 U5335 ( .A1(n10325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5866) );
  AND3_X1 U5336 ( .A1(n5839), .A2(n6341), .A3(n5838), .ZN(n5840) );
  NAND3_X1 U5337 ( .A1(n11097), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5636) );
  AND2_X1 U5338 ( .A1(n6688), .A2(n6832), .ZN(n5680) );
  AND2_X1 U5339 ( .A1(n5746), .A2(n6688), .ZN(n5745) );
  CLKBUF_X1 U5340 ( .A(n7132), .Z(n7232) );
  AND2_X1 U5341 ( .A1(n7133), .A2(n5354), .ZN(n5353) );
  INV_X1 U5342 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10311) );
  INV_X1 U5343 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10079) );
  INV_X1 U5344 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6341) );
  NOR3_X1 U5345 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .A3(
        P2_IR_REG_7__SCAN_IN), .ZN(n6687) );
  INV_X1 U5346 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6935) );
  INV_X2 U5347 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5348 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7363) );
  NOR2_X2 U5349 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7132) );
  INV_X1 U5350 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7133) );
  NOR2_X1 U5351 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6686) );
  INV_X1 U5352 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7138) );
  INV_X1 U5353 ( .A(P2_RD_REG_SCAN_IN), .ZN(n11097) );
  NOR2_X1 U5354 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5830) );
  INV_X1 U5355 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10096) );
  INV_X1 U5356 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6949) );
  AND2_X1 U5358 ( .A1(n5871), .A2(n5870), .ZN(n6195) );
  NAND4_X2 U5359 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n9549)
         );
  AND2_X1 U5360 ( .A1(n5870), .A2(n9223), .ZN(n5136) );
  AND2_X1 U5361 ( .A1(n5870), .A2(n9223), .ZN(n5137) );
  NAND3_X2 U5362 ( .A1(n5931), .A2(n5930), .A3(n5929), .ZN(n6434) );
  NOR2_X2 U5363 ( .A1(n10573), .A2(n10579), .ZN(n10574) );
  XNOR2_X2 U5364 ( .A(n7112), .B(n7111), .ZN(n7159) );
  INV_X1 U5365 ( .A(n5871), .ZN(n9223) );
  INV_X4 U5366 ( .A(n9158), .ZN(n7528) );
  XNOR2_X1 U5367 ( .A(n5844), .B(n10321), .ZN(n6325) );
  AND2_X4 U5368 ( .A1(n7130), .A2(n7113), .ZN(n7313) );
  XNOR2_X2 U5369 ( .A(n5949), .B(n10276), .ZN(n6931) );
  AOI211_X2 U5370 ( .C1(n6680), .C2(n6324), .A(n10655), .B(n5159), .ZN(n10495)
         );
  NAND3_X1 U5371 ( .A1(n5731), .A2(n8772), .A3(n5732), .ZN(n5734) );
  AOI21_X1 U5372 ( .B1(n5379), .B2(n8623), .A(n5377), .ZN(n5376) );
  INV_X1 U5373 ( .A(n8638), .ZN(n5377) );
  AND2_X1 U5374 ( .A1(n9565), .A2(n8621), .ZN(n9564) );
  OR2_X1 U5375 ( .A1(n9740), .A2(n9268), .ZN(n8764) );
  NOR2_X1 U5376 ( .A1(n9744), .A2(n9629), .ZN(n9196) );
  NOR2_X1 U5377 ( .A1(n8112), .A2(n8737), .ZN(n5470) );
  INV_X1 U5378 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6832) );
  INV_X1 U5379 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6688) );
  INV_X1 U5380 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5354) );
  AND4_X1 U5381 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n8018), .ZN(n8293)
         );
  NAND2_X1 U5382 ( .A1(n5486), .A2(n5485), .ZN(n5484) );
  INV_X1 U5383 ( .A(n9443), .ZN(n5485) );
  NOR2_X1 U5384 ( .A1(n9536), .A2(n5730), .ZN(n5729) );
  INV_X1 U5385 ( .A(n8773), .ZN(n5730) );
  NAND2_X1 U5386 ( .A1(n10514), .A2(n5182), .ZN(n10479) );
  INV_X1 U5387 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5323) );
  NOR2_X1 U5388 ( .A1(n8494), .A2(n5387), .ZN(n8501) );
  AND2_X1 U5389 ( .A1(n5372), .A2(n5208), .ZN(n5371) );
  NAND2_X1 U5390 ( .A1(n5165), .A2(n5375), .ZN(n5372) );
  INV_X1 U5391 ( .A(n5454), .ZN(n5453) );
  OAI21_X1 U5392 ( .B1(n5455), .B2(n5457), .A(n5181), .ZN(n5454) );
  NAND2_X1 U5393 ( .A1(n5283), .A2(n5290), .ZN(n5282) );
  NOR2_X1 U5394 ( .A1(n9553), .A2(n5287), .ZN(n5284) );
  INV_X1 U5395 ( .A(n9034), .ZN(n5271) );
  OR2_X1 U5396 ( .A1(n9703), .A2(n9505), .ZN(n8779) );
  NAND2_X1 U5397 ( .A1(n5487), .A2(n5488), .ZN(n8357) );
  AOI21_X1 U5398 ( .B1(n8352), .B2(n5489), .A(n5232), .ZN(n5488) );
  OR2_X1 U5399 ( .A1(n9736), .A2(n9337), .ZN(n9565) );
  INV_X1 U5400 ( .A(n5727), .ZN(n5726) );
  OAI21_X1 U5401 ( .B1(n9622), .B2(n8566), .A(n8763), .ZN(n5727) );
  NAND2_X1 U5402 ( .A1(n7829), .A2(n7798), .ZN(n7831) );
  AND2_X1 U5403 ( .A1(n8779), .A2(n8720), .ZN(n9201) );
  INV_X1 U5404 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5746) );
  AND2_X1 U5405 ( .A1(n7005), .A2(n6685), .ZN(n5322) );
  AND2_X1 U5406 ( .A1(n5697), .A2(n5702), .ZN(n5420) );
  OR2_X1 U5407 ( .A1(n10556), .A2(n10710), .ZN(n5702) );
  NAND2_X1 U5408 ( .A1(n5698), .A2(n5700), .ZN(n5697) );
  NAND2_X1 U5409 ( .A1(n6106), .A2(n6105), .ZN(n5411) );
  XNOR2_X1 U5410 ( .A(n5817), .B(n5816), .ZN(n6239) );
  XNOR2_X1 U5411 ( .A(n5805), .B(n10159), .ZN(n6170) );
  AOI21_X1 U5412 ( .B1(n9224), .B2(n5650), .A(n5179), .ZN(n5649) );
  INV_X1 U5413 ( .A(n9166), .ZN(n5650) );
  INV_X1 U5414 ( .A(n9396), .ZN(n5524) );
  NAND2_X1 U5415 ( .A1(n5142), .A2(n8319), .ZN(n5525) );
  INV_X1 U5416 ( .A(n9499), .ZN(n9506) );
  AND2_X1 U5417 ( .A1(n9713), .A2(n9716), .ZN(n5457) );
  INV_X1 U5418 ( .A(n7155), .ZN(n8708) );
  OR2_X1 U5419 ( .A1(n8037), .A2(n9521), .ZN(n8682) );
  NAND2_X1 U5420 ( .A1(n8765), .A2(n5728), .ZN(n5731) );
  INV_X1 U5421 ( .A(n8764), .ZN(n5733) );
  NAND2_X1 U5422 ( .A1(n5463), .A2(n5461), .ZN(n9576) );
  AND2_X1 U5423 ( .A1(n5462), .A2(n5466), .ZN(n5461) );
  AOI21_X1 U5424 ( .B1(n9595), .B2(n9590), .A(n5197), .ZN(n5466) );
  AND2_X1 U5425 ( .A1(n8516), .A2(n9657), .ZN(n9672) );
  NOR2_X1 U5426 ( .A1(n5470), .A2(n5171), .ZN(n5311) );
  AOI21_X1 U5427 ( .B1(n5719), .B2(n8499), .A(n5716), .ZN(n5715) );
  INV_X1 U5428 ( .A(n8491), .ZN(n5716) );
  NAND2_X1 U5429 ( .A1(n8023), .A2(n8735), .ZN(n8026) );
  OR2_X1 U5430 ( .A1(n8785), .A2(n7268), .ZN(n9643) );
  XNOR2_X1 U5431 ( .A(n7149), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8800) );
  INV_X1 U5432 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7143) );
  OR2_X1 U5433 ( .A1(n6222), .A2(n6221), .ZN(n6233) );
  AND2_X1 U5434 ( .A1(n6685), .A2(n8128), .ZN(n6668) );
  INV_X1 U5435 ( .A(n6344), .ZN(n6302) );
  INV_X1 U5436 ( .A(n5584), .ZN(n5581) );
  OR2_X1 U5437 ( .A1(n10556), .A2(n10693), .ZN(n10532) );
  OR2_X1 U5438 ( .A1(n10631), .A2(n10616), .ZN(n5694) );
  OAI22_X1 U5439 ( .A1(n10642), .A2(n5695), .B1(n10742), .B2(n10807), .ZN(
        n5690) );
  NOR2_X1 U5440 ( .A1(n10642), .A2(n5692), .ZN(n5691) );
  INV_X1 U5441 ( .A(n6200), .ZN(n5692) );
  NAND2_X1 U5442 ( .A1(n6317), .A2(n8890), .ZN(n8277) );
  INV_X1 U5443 ( .A(n6105), .ZN(n5408) );
  INV_X1 U5444 ( .A(n5703), .ZN(n5407) );
  AOI21_X1 U5445 ( .B1(n5705), .B2(n5704), .A(n5192), .ZN(n5703) );
  INV_X1 U5446 ( .A(n5164), .ZN(n5409) );
  AND4_X1 U5447 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n7515)
         );
  AOI21_X1 U5448 ( .B1(n8868), .B2(n5396), .A(n5191), .ZN(n5395) );
  INV_X1 U5449 ( .A(n6012), .ZN(n5396) );
  INV_X1 U5450 ( .A(n9913), .ZN(n10745) );
  AND2_X1 U5451 ( .A1(n9011), .A2(n9120), .ZN(n11164) );
  INV_X1 U5452 ( .A(n8853), .ZN(n6206) );
  NAND2_X1 U5453 ( .A1(n5868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U5454 ( .A1(n5607), .A2(n5606), .ZN(n6218) );
  AOI21_X1 U5455 ( .B1(n5608), .B2(n5614), .A(n5223), .ZN(n5606) );
  XNOR2_X1 U5456 ( .A(n5810), .B(n9956), .ZN(n6217) );
  NAND2_X1 U5457 ( .A1(n5610), .A2(n5611), .ZN(n6202) );
  NAND2_X1 U5458 ( .A1(n6159), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6187) );
  NOR2_X1 U5459 ( .A1(n6140), .A2(n5632), .ZN(n5631) );
  AOI21_X1 U5460 ( .B1(n9017), .B2(n10464), .A(n6419), .ZN(n5604) );
  OAI21_X1 U5461 ( .B1(n10509), .B2(n10508), .A(n9019), .ZN(n6322) );
  NAND2_X1 U5462 ( .A1(n10661), .A2(n6421), .ZN(n10576) );
  NAND2_X1 U5463 ( .A1(n8435), .A2(n8854), .ZN(n5640) );
  NAND2_X1 U5464 ( .A1(n5723), .A2(n11104), .ZN(n8462) );
  INV_X1 U5465 ( .A(n8476), .ZN(n5363) );
  NAND2_X1 U5466 ( .A1(n5246), .A2(n5245), .ZN(n5244) );
  NOR2_X1 U5467 ( .A1(n9080), .A2(n9011), .ZN(n5245) );
  NAND2_X1 U5468 ( .A1(n8932), .A2(n8902), .ZN(n5246) );
  NAND2_X1 U5469 ( .A1(n8903), .A2(n9011), .ZN(n5243) );
  OR2_X1 U5470 ( .A1(n8485), .A2(n8727), .ZN(n5392) );
  AND2_X1 U5471 ( .A1(n5585), .A2(n8972), .ZN(n8989) );
  NOR2_X1 U5472 ( .A1(n8977), .A2(n8968), .ZN(n8971) );
  INV_X1 U5473 ( .A(n5165), .ZN(n5369) );
  INV_X1 U5474 ( .A(n5371), .ZN(n5370) );
  INV_X1 U5475 ( .A(n7437), .ZN(n5539) );
  NAND2_X1 U5476 ( .A1(n9155), .A2(n9593), .ZN(n9156) );
  NAND2_X1 U5477 ( .A1(n5291), .A2(n9277), .ZN(n5290) );
  INV_X1 U5478 ( .A(n9725), .ZN(n5291) );
  NOR2_X1 U5479 ( .A1(n5160), .A2(n5289), .ZN(n5283) );
  OR2_X1 U5480 ( .A1(n8104), .A2(n8103), .ZN(n8112) );
  INV_X1 U5481 ( .A(n7438), .ZN(n5538) );
  INV_X1 U5482 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5839) );
  INV_X1 U5483 ( .A(n9156), .ZN(n5656) );
  AND2_X2 U5484 ( .A1(n7303), .A2(n7302), .ZN(n9158) );
  NAND2_X1 U5485 ( .A1(n5255), .A2(n5253), .ZN(n8788) );
  INV_X1 U5486 ( .A(n5254), .ZN(n5253) );
  OAI21_X1 U5487 ( .B1(n9700), .B2(n8786), .A(n8785), .ZN(n5254) );
  NAND2_X1 U5488 ( .A1(n11025), .A2(n7205), .ZN(n5504) );
  NOR2_X1 U5489 ( .A1(n7206), .A2(n7204), .ZN(n5503) );
  NOR2_X1 U5490 ( .A1(n9432), .A2(n8371), .ZN(n8372) );
  NOR2_X1 U5491 ( .A1(n9439), .A2(n8370), .ZN(n8371) );
  OR2_X1 U5492 ( .A1(n9713), .A2(n9531), .ZN(n9185) );
  NOR2_X1 U5493 ( .A1(n9200), .A2(n5456), .ZN(n5455) );
  INV_X1 U5494 ( .A(n5458), .ZN(n5456) );
  AND2_X1 U5495 ( .A1(n9185), .A2(n9184), .ZN(n9200) );
  NOR2_X1 U5496 ( .A1(n9198), .A2(n5468), .ZN(n5467) );
  AND2_X1 U5497 ( .A1(n9667), .A2(n5295), .ZN(n5294) );
  INV_X1 U5498 ( .A(n9194), .ZN(n5295) );
  AND2_X1 U5499 ( .A1(n7940), .A2(n8443), .ZN(n7798) );
  AOI21_X1 U5500 ( .B1(n5453), .B2(n5457), .A(n5202), .ZN(n5451) );
  AOI21_X1 U5501 ( .B1(n9582), .B2(n9199), .A(n5195), .ZN(n5288) );
  OR2_X1 U5502 ( .A1(n9576), .A2(n5279), .ZN(n5285) );
  INV_X1 U5503 ( .A(n5283), .ZN(n5279) );
  INV_X1 U5504 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5679) );
  OR2_X1 U5505 ( .A1(n6680), .A2(n10676), .ZN(n9031) );
  OR2_X1 U5506 ( .A1(n6271), .A2(n6270), .ZN(n6326) );
  NAND2_X1 U5507 ( .A1(n5433), .A2(n10517), .ZN(n5432) );
  NAND2_X1 U5508 ( .A1(n6320), .A2(n10532), .ZN(n8990) );
  NAND2_X1 U5509 ( .A1(n5585), .A2(n8979), .ZN(n5584) );
  OR2_X1 U5510 ( .A1(n10538), .A2(n10684), .ZN(n9027) );
  AND2_X1 U5511 ( .A1(n5684), .A2(n6238), .ZN(n5419) );
  OR2_X1 U5512 ( .A1(n10725), .A2(n10589), .ZN(n6238) );
  NOR2_X1 U5513 ( .A1(n10624), .A2(n5690), .ZN(n5687) );
  AND2_X1 U5514 ( .A1(n8959), .A2(n9094), .ZN(n10642) );
  INV_X1 U5515 ( .A(n5559), .ZN(n5558) );
  OAI21_X1 U5516 ( .B1(n6316), .B2(n5560), .A(n8876), .ZN(n5559) );
  INV_X1 U5517 ( .A(n8948), .ZN(n5560) );
  OR2_X1 U5518 ( .A1(n10759), .A2(n9857), .ZN(n8950) );
  OR2_X1 U5519 ( .A1(n6540), .A2(n10764), .ZN(n9084) );
  INV_X1 U5520 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U5521 ( .A1(n10354), .A2(n11129), .ZN(n9064) );
  NOR2_X1 U5522 ( .A1(n6354), .A2(n8308), .ZN(n6365) );
  NOR2_X1 U5523 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5845) );
  INV_X1 U5524 ( .A(n5625), .ZN(n5620) );
  NOR2_X1 U5525 ( .A1(n6081), .A2(n5626), .ZN(n5625) );
  INV_X1 U5526 ( .A(n5791), .ZN(n5626) );
  INV_X1 U5527 ( .A(n5442), .ZN(n5441) );
  OAI211_X1 U5528 ( .C1(n5974), .C2(n5603), .A(n5602), .B(n5989), .ZN(n5992)
         );
  OAI21_X1 U5529 ( .B1(n9168), .B2(n5183), .A(n5647), .ZN(n5646) );
  INV_X1 U5530 ( .A(n7311), .ZN(n5723) );
  INV_X1 U5531 ( .A(n8297), .ZN(n5664) );
  AND2_X1 U5532 ( .A1(n5144), .A2(n5670), .ZN(n5668) );
  NAND2_X1 U5533 ( .A1(n5205), .A2(n5144), .ZN(n5667) );
  NAND2_X1 U5534 ( .A1(n9282), .A2(n9283), .ZN(n5661) );
  OR2_X1 U5535 ( .A1(n8257), .A2(n9386), .ZN(n5670) );
  AOI22_X1 U5536 ( .A1(n7757), .A2(n5382), .B1(n7156), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n5381) );
  INV_X1 U5537 ( .A(n7241), .ZN(n5474) );
  XNOR2_X1 U5538 ( .A(n7207), .B(n7535), .ZN(n11053) );
  NOR2_X1 U5539 ( .A1(n11053), .A2(n11052), .ZN(n11051) );
  OAI21_X1 U5540 ( .B1(n11043), .B2(n5494), .A(n5493), .ZN(n11059) );
  NAND2_X1 U5541 ( .A1(n5497), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5542 ( .A1(n7245), .A2(n5497), .ZN(n5493) );
  INV_X1 U5543 ( .A(n11060), .ZN(n5497) );
  OR2_X1 U5544 ( .A1(n11043), .A2(n11044), .ZN(n5496) );
  AOI21_X1 U5545 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7771), .A(n7768), .ZN(
        n7974) );
  AOI21_X1 U5546 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8318), .A(n8317), .ZN(
        n8364) );
  AND2_X1 U5547 ( .A1(n9394), .A2(n8367), .ZN(n8368) );
  INV_X1 U5548 ( .A(n8357), .ZN(n8355) );
  NOR2_X1 U5549 ( .A1(n5511), .A2(n5510), .ZN(n9473) );
  NAND2_X1 U5550 ( .A1(n8373), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5511) );
  INV_X1 U5551 ( .A(n5315), .ZN(n5460) );
  NAND2_X1 U5552 ( .A1(n9544), .A2(n8774), .ZN(n9183) );
  OR2_X1 U5553 ( .A1(n9725), .A2(n9277), .ZN(n8773) );
  XNOR2_X1 U5554 ( .A(n9721), .B(n9549), .ZN(n9545) );
  NAND2_X1 U5555 ( .A1(n8770), .A2(n5149), .ZN(n5732) );
  NAND2_X1 U5556 ( .A1(n9576), .A2(n9577), .ZN(n9575) );
  INV_X1 U5557 ( .A(n9564), .ZN(n9595) );
  INV_X1 U5558 ( .A(n5465), .ZN(n5464) );
  OAI21_X1 U5559 ( .B1(n5467), .B2(n9590), .A(n9595), .ZN(n5465) );
  NOR2_X1 U5560 ( .A1(n5300), .A2(n5299), .ZN(n9197) );
  INV_X1 U5561 ( .A(n5302), .ZN(n5299) );
  INV_X1 U5562 ( .A(n5303), .ZN(n5300) );
  NAND2_X1 U5563 ( .A1(n9623), .A2(n9622), .ZN(n9625) );
  NAND2_X1 U5564 ( .A1(n5440), .A2(n9195), .ZN(n9642) );
  NAND2_X1 U5565 ( .A1(n5310), .A2(n5309), .ZN(n9193) );
  AOI21_X1 U5566 ( .B1(n5143), .B2(n5311), .A(n5194), .ZN(n5309) );
  NOR2_X1 U5567 ( .A1(n9685), .A2(n5741), .ZN(n5740) );
  INV_X1 U5568 ( .A(n8754), .ZN(n5741) );
  OR2_X1 U5569 ( .A1(n8110), .A2(n5143), .ZN(n5312) );
  OR2_X1 U5570 ( .A1(n8106), .A2(n7524), .ZN(n8108) );
  XNOR2_X1 U5571 ( .A(n8505), .B(n9384), .ZN(n8737) );
  NAND2_X1 U5572 ( .A1(n8034), .A2(n8498), .ZN(n8122) );
  AOI21_X1 U5573 ( .B1(n5736), .B2(n8496), .A(n8495), .ZN(n5735) );
  AND2_X1 U5574 ( .A1(n8022), .A2(n8123), .ZN(n8739) );
  INV_X1 U5575 ( .A(n5278), .ZN(n5277) );
  OAI21_X1 U5576 ( .B1(n7929), .B2(n7930), .A(n7932), .ZN(n5278) );
  NAND2_X1 U5577 ( .A1(n7942), .A2(n7941), .ZN(n5739) );
  NAND2_X1 U5578 ( .A1(n7429), .A2(n8463), .ZN(n7430) );
  AND2_X1 U5579 ( .A1(n7154), .A2(n7687), .ZN(n9203) );
  XNOR2_X1 U5580 ( .A(n7311), .B(n7428), .ZN(n8469) );
  INV_X1 U5581 ( .A(n7162), .ZN(n9687) );
  NOR2_X1 U5582 ( .A1(n9775), .A2(n7338), .ZN(n7339) );
  OR2_X1 U5583 ( .A1(n8464), .A2(n7192), .ZN(n7677) );
  NAND2_X1 U5584 ( .A1(n8464), .A2(n7171), .ZN(n7679) );
  AND2_X1 U5585 ( .A1(n7270), .A2(n7188), .ZN(n7682) );
  INV_X1 U5586 ( .A(n9201), .ZN(n9188) );
  NAND2_X1 U5587 ( .A1(n8614), .A2(n8613), .ZN(n9732) );
  INV_X1 U5588 ( .A(n9779), .ZN(n9752) );
  AND4_X1 U5589 ( .A1(n7589), .A2(n7588), .A3(n7587), .A4(n7586), .ZN(n7911)
         );
  OR2_X1 U5590 ( .A1(n7189), .A2(n8800), .ZN(n9775) );
  INV_X1 U5591 ( .A(n7160), .ZN(n9773) );
  NAND2_X1 U5592 ( .A1(n5167), .A2(n6764), .ZN(n6765) );
  INV_X1 U5593 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7093) );
  INV_X1 U5594 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5385) );
  AOI21_X1 U5595 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_20__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U5596 ( .A1(n6773), .A2(n5680), .ZN(n6843) );
  AND2_X1 U5597 ( .A1(n6773), .A2(n6688), .ZN(n6833) );
  INV_X1 U5598 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U5599 ( .A1(n6353), .A2(n6347), .ZN(n6685) );
  NOR2_X1 U5600 ( .A1(n8269), .A2(n8245), .ZN(n6347) );
  INV_X1 U5601 ( .A(n6564), .ZN(n5343) );
  OR2_X1 U5602 ( .A1(n9854), .A2(n5343), .ZN(n5342) );
  NAND2_X1 U5603 ( .A1(n5549), .A2(n5548), .ZN(n5547) );
  INV_X1 U5604 ( .A(n9907), .ZN(n5548) );
  INV_X1 U5605 ( .A(n9908), .ZN(n5549) );
  NAND2_X1 U5606 ( .A1(n5542), .A2(n5540), .ZN(n9827) );
  AOI21_X1 U5607 ( .B1(n5543), .B2(n5339), .A(n5541), .ZN(n5540) );
  NAND2_X1 U5608 ( .A1(n9910), .A2(n5543), .ZN(n5542) );
  INV_X1 U5609 ( .A(n6607), .ZN(n5541) );
  AND2_X1 U5610 ( .A1(n6606), .A2(n5544), .ZN(n5543) );
  NAND2_X1 U5611 ( .A1(n5545), .A2(n5546), .ZN(n5544) );
  INV_X1 U5612 ( .A(n5547), .ZN(n5545) );
  NAND2_X1 U5613 ( .A1(n5853), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6099) );
  INV_X1 U5614 ( .A(n5531), .ZN(n5529) );
  NAND2_X1 U5615 ( .A1(n9808), .A2(n5533), .ZN(n5530) );
  NAND2_X1 U5616 ( .A1(n5326), .A2(n5189), .ZN(n9841) );
  OR2_X1 U5617 ( .A1(n6547), .A2(n5329), .ZN(n5328) );
  OR2_X1 U5618 ( .A1(n6035), .A2(n6034), .ZN(n6047) );
  NAND2_X1 U5619 ( .A1(n5325), .A2(n5324), .ZN(n8066) );
  AND2_X1 U5620 ( .A1(n8068), .A2(n7813), .ZN(n5324) );
  NAND2_X1 U5621 ( .A1(n5858), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6243) );
  AND2_X1 U5622 ( .A1(n5528), .A2(n9809), .ZN(n5333) );
  AND2_X1 U5623 ( .A1(n9029), .A2(n9019), .ZN(n10500) );
  NOR2_X1 U5624 ( .A1(n10500), .A2(n5713), .ZN(n5711) );
  NAND2_X1 U5625 ( .A1(n10785), .A2(n10684), .ZN(n5399) );
  NAND2_X1 U5626 ( .A1(n10538), .A2(n10520), .ZN(n5401) );
  INV_X1 U5627 ( .A(n8990), .ZN(n5582) );
  NAND2_X1 U5628 ( .A1(n5200), .A2(n5177), .ZN(n5700) );
  NAND2_X1 U5629 ( .A1(n5200), .A2(n6250), .ZN(n5698) );
  AND2_X1 U5630 ( .A1(n8982), .A2(n8979), .ZN(n10566) );
  NAND2_X1 U5631 ( .A1(n5686), .A2(n5419), .ZN(n10585) );
  NAND2_X1 U5632 ( .A1(n10585), .A2(n10586), .ZN(n10584) );
  NAND2_X1 U5633 ( .A1(n10605), .A2(n5685), .ZN(n5684) );
  INV_X1 U5634 ( .A(n5694), .ZN(n5685) );
  NAND2_X1 U5635 ( .A1(n5687), .A2(n5688), .ZN(n5683) );
  AND2_X1 U5636 ( .A1(n8973), .A2(n8886), .ZN(n10624) );
  AND4_X1 U5637 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n10644)
         );
  AOI21_X1 U5638 ( .B1(n5406), .B2(n5409), .A(n6316), .ZN(n5403) );
  NOR2_X1 U5639 ( .A1(n8943), .A2(n5706), .ZN(n5705) );
  INV_X1 U5640 ( .A(n6124), .ZN(n5706) );
  NAND2_X1 U5641 ( .A1(n5708), .A2(n5161), .ZN(n5707) );
  NAND2_X1 U5642 ( .A1(n6097), .A2(n6096), .ZN(n7671) );
  NAND2_X1 U5643 ( .A1(n7512), .A2(n11160), .ZN(n7669) );
  NOR2_X1 U5644 ( .A1(n8872), .A2(n5588), .ZN(n5587) );
  INV_X1 U5645 ( .A(n8894), .ZN(n5588) );
  NAND2_X1 U5646 ( .A1(n7027), .A2(n8914), .ZN(n7026) );
  AND4_X1 U5647 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n7042)
         );
  NAND2_X1 U5648 ( .A1(n5578), .A2(n9061), .ZN(n5575) );
  NAND2_X1 U5649 ( .A1(n9057), .A2(n9058), .ZN(n5578) );
  XNOR2_X1 U5650 ( .A(n6402), .B(n6401), .ZN(n6410) );
  NAND2_X1 U5651 ( .A1(n5563), .A2(n5561), .ZN(n6402) );
  INV_X1 U5652 ( .A(n5562), .ZN(n5561) );
  NAND2_X1 U5653 ( .A1(n8846), .A2(n8845), .ZN(n10472) );
  INV_X1 U5654 ( .A(n10520), .ZN(n10684) );
  INV_X1 U5655 ( .A(n11156), .ZN(n10763) );
  AND2_X1 U5656 ( .A1(n5139), .A2(n9040), .ZN(n11155) );
  INV_X1 U5657 ( .A(n11155), .ZN(n10741) );
  INV_X1 U5658 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10321) );
  XNOR2_X1 U5659 ( .A(n6287), .B(n6381), .ZN(n8435) );
  AND2_X1 U5660 ( .A1(n6286), .A2(n6380), .ZN(n6287) );
  NAND2_X1 U5661 ( .A1(n5599), .A2(n6386), .ZN(n6286) );
  INV_X1 U5662 ( .A(n5198), .ZN(n5344) );
  AND2_X1 U5663 ( .A1(n5827), .A2(n5879), .ZN(n5828) );
  XNOR2_X1 U5664 ( .A(n6349), .B(n10311), .ZN(n8128) );
  OR2_X1 U5665 ( .A1(n6297), .A2(n10312), .ZN(n6298) );
  NOR2_X1 U5666 ( .A1(n5617), .A2(n6183), .ZN(n5615) );
  NOR2_X1 U5667 ( .A1(n5798), .A2(SI_14_), .ZN(n5632) );
  NAND2_X1 U5668 ( .A1(n6110), .A2(n5634), .ZN(n5633) );
  NOR2_X1 U5669 ( .A1(n6087), .A2(n5623), .ZN(n5622) );
  INV_X1 U5670 ( .A(n5627), .ZN(n5623) );
  NAND2_X1 U5671 ( .A1(n5629), .A2(n5628), .ZN(n5627) );
  INV_X1 U5672 ( .A(SI_11_), .ZN(n5628) );
  INV_X1 U5673 ( .A(n5792), .ZN(n5629) );
  XNOR2_X1 U5674 ( .A(n6082), .B(n6081), .ZN(n8011) );
  XNOR2_X1 U5675 ( .A(n6028), .B(n6027), .ZN(n7825) );
  NAND2_X1 U5676 ( .A1(n5447), .A2(n5448), .ZN(n6028) );
  OR2_X1 U5677 ( .A1(n6005), .A2(n5782), .ZN(n5447) );
  INV_X1 U5678 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U5679 ( .A1(n8579), .A2(n8578), .ZN(n9744) );
  AND4_X1 U5680 ( .A1(n8596), .A2(n8595), .A3(n8594), .A4(n8593), .ZN(n9268)
         );
  INV_X1 U5681 ( .A(n9383), .ZN(n9688) );
  INV_X1 U5682 ( .A(n9392), .ZN(n8474) );
  INV_X1 U5683 ( .A(n9382), .ZN(n9669) );
  INV_X1 U5684 ( .A(n9190), .ZN(n9328) );
  AND2_X1 U5685 ( .A1(n8558), .A2(n8557), .ZN(n9748) );
  AND2_X1 U5686 ( .A1(n8510), .A2(n8509), .ZN(n9768) );
  INV_X1 U5687 ( .A(n8801), .ZN(n5347) );
  AND2_X1 U5688 ( .A1(n8748), .A2(n8792), .ZN(n5350) );
  NOR2_X1 U5689 ( .A1(n8750), .A2(n8749), .ZN(n5252) );
  OR2_X1 U5690 ( .A1(n7769), .A2(n7952), .ZN(n5520) );
  XNOR2_X1 U5691 ( .A(n8368), .B(n9420), .ZN(n9415) );
  AND2_X1 U5692 ( .A1(n11076), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U5693 ( .A1(n5261), .A2(n8380), .ZN(n5250) );
  NAND2_X1 U5694 ( .A1(n11076), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5261) );
  NOR2_X1 U5695 ( .A1(n8401), .A2(n8363), .ZN(n5475) );
  OAI21_X1 U5696 ( .B1(n9472), .B2(n5477), .A(n5476), .ZN(n5248) );
  NAND2_X1 U5697 ( .A1(n5482), .A2(n5235), .ZN(n5476) );
  NAND2_X1 U5698 ( .A1(n5482), .A2(n5236), .ZN(n5477) );
  INV_X1 U5699 ( .A(n8403), .ZN(n5513) );
  NOR2_X1 U5700 ( .A1(n9519), .A2(n5457), .ZN(n9500) );
  AND2_X1 U5701 ( .A1(n8680), .A2(n8679), .ZN(n9521) );
  NAND2_X1 U5702 ( .A1(n8549), .A2(n8548), .ZN(n9755) );
  AND2_X1 U5703 ( .A1(n5878), .A2(n5877), .ZN(n10694) );
  NOR3_X1 U5704 ( .A1(n9921), .A2(n9173), .A3(n9174), .ZN(n9177) );
  NAND2_X1 U5705 ( .A1(n5905), .A2(n5904), .ZN(n10556) );
  AND3_X1 U5706 ( .A1(n6216), .A2(n6215), .A3(n6214), .ZN(n10742) );
  NAND2_X1 U5707 ( .A1(n6220), .A2(n6219), .ZN(n10631) );
  NAND2_X1 U5708 ( .A1(n6241), .A2(n6240), .ZN(n10595) );
  AND4_X1 U5709 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n10740)
         );
  AND2_X1 U5710 ( .A1(n6656), .A2(n6662), .ZN(n9926) );
  INV_X1 U5711 ( .A(n9936), .ZN(n9904) );
  NAND2_X1 U5712 ( .A1(n6302), .A2(n6301), .ZN(n9120) );
  NAND2_X1 U5713 ( .A1(n6295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6300) );
  INV_X1 U5714 ( .A(n9812), .ZN(n10709) );
  AND2_X1 U5715 ( .A1(n6083), .A2(n6063), .ZN(n10963) );
  NAND2_X1 U5716 ( .A1(n9938), .A2(n11156), .ZN(n6409) );
  XNOR2_X1 U5717 ( .A(n6399), .B(n9006), .ZN(n8802) );
  OR2_X1 U5718 ( .A1(n8841), .A2(n6396), .ZN(n6398) );
  AND2_X1 U5719 ( .A1(n6191), .A2(n6190), .ZN(n9913) );
  NAND2_X1 U5720 ( .A1(n6116), .A2(n6115), .ZN(n7907) );
  AND4_X1 U5721 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n9877)
         );
  AND2_X1 U5722 ( .A1(n10601), .A2(n6971), .ZN(n10651) );
  AND2_X1 U5723 ( .A1(n10661), .A2(n6963), .ZN(n10580) );
  INV_X1 U5724 ( .A(n5595), .ZN(n5422) );
  NAND2_X1 U5725 ( .A1(n5201), .A2(n5268), .ZN(n5267) );
  NAND2_X1 U5726 ( .A1(n10485), .A2(n11178), .ZN(n5268) );
  NAND2_X1 U5727 ( .A1(n5437), .A2(n6707), .ZN(n5436) );
  NAND2_X1 U5728 ( .A1(n5438), .A2(n5150), .ZN(n5437) );
  NAND2_X1 U5729 ( .A1(n6203), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U5730 ( .A1(n8479), .A2(n8695), .ZN(n5356) );
  NAND2_X1 U5731 ( .A1(n5362), .A2(n5360), .ZN(n5359) );
  NOR2_X1 U5732 ( .A1(n8478), .A2(n5361), .ZN(n5360) );
  OAI21_X1 U5733 ( .B1(n5364), .B2(n8473), .A(n5363), .ZN(n5362) );
  NAND2_X1 U5734 ( .A1(n5244), .A2(n5243), .ZN(n8935) );
  INV_X1 U5735 ( .A(n5388), .ZN(n5387) );
  AOI21_X1 U5736 ( .B1(n8497), .B2(n8496), .A(n8495), .ZN(n5388) );
  NAND2_X1 U5737 ( .A1(n5361), .A2(n8464), .ZN(n5389) );
  NAND2_X1 U5738 ( .A1(n8487), .A2(n8695), .ZN(n5391) );
  MUX2_X1 U5739 ( .A(n8946), .B(n8945), .S(n9011), .Z(n8954) );
  INV_X1 U5740 ( .A(n5376), .ZN(n5375) );
  INV_X1 U5741 ( .A(n9569), .ZN(n5378) );
  NAND2_X1 U5742 ( .A1(n5376), .A2(n5374), .ZN(n5373) );
  INV_X1 U5743 ( .A(n5379), .ZN(n5374) );
  INV_X1 U5744 ( .A(n9105), .ZN(n5276) );
  AOI21_X1 U5745 ( .B1(n5368), .B2(n5370), .A(n5367), .ZN(n5366) );
  INV_X1 U5746 ( .A(n8661), .ZN(n5367) );
  NAND2_X1 U5747 ( .A1(n9700), .A2(n8716), .ZN(n5256) );
  INV_X1 U5748 ( .A(n9404), .ZN(n5489) );
  INV_X1 U5749 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7137) );
  NOR2_X1 U5750 ( .A1(n5699), .A2(n5418), .ZN(n5417) );
  INV_X1 U5751 ( .A(n5700), .ZN(n5699) );
  INV_X1 U5752 ( .A(SI_17_), .ZN(n10159) );
  NAND2_X1 U5753 ( .A1(n5448), .A2(n5446), .ZN(n5445) );
  INV_X1 U5754 ( .A(n6027), .ZN(n5446) );
  INV_X1 U5755 ( .A(SI_9_), .ZN(n10170) );
  OAI21_X1 U5756 ( .B1(n5771), .B2(n5759), .A(n5758), .ZN(n5760) );
  NAND2_X1 U5757 ( .A1(n9335), .A2(n9156), .ZN(n9244) );
  NOR2_X1 U5758 ( .A1(n11059), .A2(n7247), .ZN(n7612) );
  AOI21_X1 U5759 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7771), .A(n7770), .ZN(
        n7988) );
  NOR2_X1 U5760 ( .A1(n8213), .A2(n8212), .ZN(n8215) );
  OR2_X1 U5761 ( .A1(n9717), .A2(n9162), .ZN(n9182) );
  AND2_X1 U5762 ( .A1(n5168), .A2(n5302), .ZN(n5301) );
  NAND2_X1 U5763 ( .A1(n5168), .A2(n9196), .ZN(n5462) );
  INV_X1 U5764 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U5765 ( .A1(n5305), .A2(n5308), .ZN(n5302) );
  NOR2_X1 U5766 ( .A1(n9748), .A2(n9757), .ZN(n5308) );
  AND2_X1 U5767 ( .A1(n5172), .A2(n5146), .ZN(n5305) );
  AND2_X1 U5768 ( .A1(n5307), .A2(n5172), .ZN(n5306) );
  INV_X1 U5769 ( .A(n9641), .ZN(n5307) );
  NAND2_X1 U5770 ( .A1(n8110), .A2(n5311), .ZN(n5310) );
  INV_X1 U5771 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8321) );
  NOR2_X1 U5772 ( .A1(n8035), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8113) );
  INV_X1 U5773 ( .A(n8735), .ZN(n5738) );
  NAND2_X1 U5774 ( .A1(n8456), .A2(n8458), .ZN(n8725) );
  OR2_X1 U5775 ( .A1(n9708), .A2(n9227), .ZN(n9187) );
  INV_X1 U5776 ( .A(n9545), .ZN(n9536) );
  INV_X1 U5777 ( .A(n5290), .ZN(n5280) );
  NAND2_X1 U5778 ( .A1(n7106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U5779 ( .A1(n8150), .A2(n6535), .ZN(n6541) );
  INV_X1 U5780 ( .A(n8338), .ZN(n5329) );
  AND2_X1 U5781 ( .A1(n6544), .A2(n5173), .ZN(n5327) );
  NAND2_X1 U5782 ( .A1(n5537), .A2(n5187), .ZN(n7857) );
  NOR2_X1 U5783 ( .A1(n6427), .A2(n5752), .ZN(n6433) );
  AND2_X1 U5784 ( .A1(n6637), .A2(n6964), .ZN(n6427) );
  OAI21_X1 U5785 ( .B1(n9037), .B2(n9011), .A(n9118), .ZN(n9008) );
  NOR2_X1 U5786 ( .A1(n10913), .A2(n10914), .ZN(n10912) );
  NAND2_X1 U5787 ( .A1(n10508), .A2(n9019), .ZN(n5570) );
  NOR2_X1 U5788 ( .A1(n6680), .A2(n5432), .ZN(n5431) );
  INV_X1 U5789 ( .A(n10535), .ZN(n5402) );
  INV_X1 U5790 ( .A(n5417), .ZN(n5416) );
  NAND2_X1 U5791 ( .A1(n5417), .A2(n5415), .ZN(n5414) );
  INV_X1 U5792 ( .A(n5419), .ZN(n5415) );
  NAND2_X1 U5793 ( .A1(n10593), .A2(n10797), .ZN(n10573) );
  OAI21_X1 U5794 ( .B1(n8277), .B2(n8957), .A(n8961), .ZN(n10641) );
  NOR2_X1 U5795 ( .A1(n10753), .A2(n5426), .ZN(n5425) );
  INV_X1 U5796 ( .A(n5427), .ZN(n5426) );
  NOR2_X1 U5797 ( .A1(n10759), .A2(n10767), .ZN(n5427) );
  INV_X1 U5798 ( .A(n5161), .ZN(n5704) );
  NOR2_X1 U5799 ( .A1(n6994), .A2(n7418), .ZN(n6972) );
  NAND2_X1 U5800 ( .A1(n5579), .A2(n8905), .ZN(n9060) );
  OAI21_X1 U5801 ( .B1(n5569), .B2(n8992), .A(n5565), .ZN(n5562) );
  AOI21_X1 U5802 ( .B1(n5568), .B2(n5567), .A(n5566), .ZN(n5565) );
  INV_X1 U5803 ( .A(n9019), .ZN(n5567) );
  INV_X1 U5804 ( .A(n9020), .ZN(n5566) );
  NOR2_X1 U5805 ( .A1(n10653), .A2(n10631), .ZN(n5439) );
  OAI21_X1 U5806 ( .B1(n6391), .B2(n6390), .A(n6389), .ZN(n8406) );
  INV_X1 U5807 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10316) );
  INV_X1 U5808 ( .A(n6342), .ZN(n5841) );
  INV_X1 U5809 ( .A(SI_23_), .ZN(n10142) );
  NAND2_X1 U5810 ( .A1(n6296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U5811 ( .A1(n6302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6299) );
  AOI21_X1 U5812 ( .B1(n6218), .B2(n6217), .A(n5811), .ZN(n6227) );
  INV_X1 U5813 ( .A(SI_19_), .ZN(n10154) );
  NOR2_X1 U5814 ( .A1(n5609), .A2(n6201), .ZN(n5608) );
  INV_X1 U5815 ( .A(n5611), .ZN(n5609) );
  AOI21_X1 U5816 ( .B1(n5615), .B2(n5613), .A(n5612), .ZN(n5611) );
  INV_X1 U5817 ( .A(n5807), .ZN(n5612) );
  INV_X1 U5818 ( .A(n6170), .ZN(n5613) );
  INV_X1 U5819 ( .A(n5615), .ZN(n5614) );
  NAND2_X1 U5820 ( .A1(n6142), .A2(n5800), .ZN(n6155) );
  INV_X1 U5821 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10296) );
  AOI21_X1 U5822 ( .B1(n6020), .B2(n5450), .A(n5449), .ZN(n5448) );
  INV_X1 U5823 ( .A(n5783), .ZN(n5449) );
  INV_X1 U5824 ( .A(n5780), .ZN(n5450) );
  OAI21_X1 U5825 ( .B1(n5823), .B2(n5275), .A(n5274), .ZN(n5781) );
  INV_X1 U5826 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U5827 ( .A1(n5823), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5274) );
  OR2_X1 U5828 ( .A1(n6006), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U5829 ( .B1(n5771), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n5761), .ZN(
        n5762) );
  NAND2_X1 U5830 ( .A1(n5771), .A2(n7123), .ZN(n5761) );
  AND2_X1 U5831 ( .A1(n8113), .A2(n8321), .ZN(n8168) );
  NAND2_X1 U5832 ( .A1(n9237), .A2(n8168), .ZN(n8511) );
  INV_X1 U5833 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9237) );
  AOI21_X1 U5834 ( .B1(n9158), .B2(n7686), .A(n7307), .ZN(n7492) );
  AOI21_X1 U5835 ( .B1(n7530), .B2(n7704), .A(n7546), .ZN(n5672) );
  INV_X1 U5836 ( .A(n5655), .ZN(n5654) );
  OAI21_X1 U5837 ( .B1(n9154), .B2(n5656), .A(n9157), .ZN(n5655) );
  NAND2_X1 U5838 ( .A1(n5654), .A2(n5656), .ZN(n5653) );
  INV_X1 U5839 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7835) );
  AND2_X1 U5840 ( .A1(n9149), .A2(n9151), .ZN(n5674) );
  NAND2_X1 U5841 ( .A1(n9255), .A2(n9254), .ZN(n5675) );
  NAND2_X1 U5842 ( .A1(n8414), .A2(n10002), .ZN(n8615) );
  OR2_X1 U5843 ( .A1(n8015), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8035) );
  INV_X1 U5844 ( .A(n9293), .ZN(n9143) );
  AND3_X1 U5845 ( .A1(n7274), .A2(n7678), .A3(n7273), .ZN(n7327) );
  NAND2_X1 U5846 ( .A1(n9234), .A2(n9233), .ZN(n9235) );
  AND4_X1 U5847 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n8751)
         );
  NOR2_X1 U5848 ( .A1(n7092), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n7110) );
  NOR2_X1 U5849 ( .A1(n10977), .A2(n10976), .ZN(n10975) );
  OAI21_X1 U5850 ( .B1(n7237), .B2(P2_REG1_REG_2__SCAN_IN), .A(n7238), .ZN(
        n10998) );
  NOR2_X1 U5851 ( .A1(n11009), .A2(n7697), .ZN(n11008) );
  XNOR2_X1 U5852 ( .A(n7240), .B(n11016), .ZN(n11011) );
  NOR2_X1 U5853 ( .A1(n11011), .A2(n7212), .ZN(n11010) );
  NOR2_X1 U5854 ( .A1(n11008), .A2(n7204), .ZN(n11026) );
  OAI21_X1 U5855 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7243), .A(n7242), .ZN(
        n11028) );
  NAND2_X1 U5856 ( .A1(n11035), .A2(n5259), .ZN(n11048) );
  OR2_X1 U5857 ( .A1(n7222), .A2(n11034), .ZN(n5259) );
  AOI21_X1 U5858 ( .B1(n11048), .B2(n11049), .A(n5257), .ZN(n11066) );
  NOR2_X1 U5859 ( .A1(n5258), .A2(n7535), .ZN(n5257) );
  INV_X1 U5860 ( .A(n7223), .ZN(n5258) );
  NOR2_X1 U5861 ( .A1(n11051), .A2(n7208), .ZN(n11070) );
  XNOR2_X1 U5862 ( .A(n7612), .B(n7747), .ZN(n7248) );
  OAI21_X1 U5863 ( .B1(n7248), .B2(n5499), .A(n5498), .ZN(n7770) );
  NAND2_X1 U5864 ( .A1(n5500), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U5865 ( .A1(n7614), .A2(n5500), .ZN(n5498) );
  INV_X1 U5866 ( .A(n7615), .ZN(n5500) );
  NOR2_X1 U5867 ( .A1(n7248), .A2(n7249), .ZN(n7613) );
  NOR2_X1 U5868 ( .A1(n7980), .A2(n5260), .ZN(n8202) );
  OAI21_X1 U5869 ( .B1(n7772), .B2(n5491), .A(n5490), .ZN(n8213) );
  NAND2_X1 U5870 ( .A1(n5492), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U5871 ( .A1(n7991), .A2(n5492), .ZN(n5490) );
  INV_X1 U5872 ( .A(n7992), .ZN(n5492) );
  NOR2_X1 U5873 ( .A1(n7772), .A2(n7773), .ZN(n7990) );
  AOI21_X1 U5874 ( .B1(n8202), .B2(n8201), .A(n8200), .ZN(n11084) );
  XNOR2_X1 U5875 ( .A(n8357), .B(n8356), .ZN(n9424) );
  NAND2_X1 U5876 ( .A1(n8382), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U5877 ( .A1(n8402), .A2(n5480), .ZN(n5479) );
  NAND2_X1 U5878 ( .A1(n9471), .A2(n8362), .ZN(n5480) );
  INV_X1 U5879 ( .A(n9471), .ZN(n5481) );
  INV_X1 U5880 ( .A(n11090), .ZN(n5482) );
  NAND2_X1 U5881 ( .A1(n8374), .A2(n9486), .ZN(n5509) );
  AND2_X1 U5882 ( .A1(n8373), .A2(n5512), .ZN(n5505) );
  AND2_X1 U5883 ( .A1(n9474), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5512) );
  AND2_X1 U5884 ( .A1(n9213), .A2(n8438), .ZN(n9502) );
  NAND2_X1 U5885 ( .A1(n5459), .A2(n9162), .ZN(n5458) );
  INV_X1 U5886 ( .A(n5455), .ZN(n5314) );
  INV_X1 U5887 ( .A(n9200), .ZN(n9516) );
  OR2_X1 U5888 ( .A1(n9580), .A2(n9577), .ZN(n9581) );
  NAND2_X1 U5889 ( .A1(n8765), .A2(n8764), .ZN(n9563) );
  OR2_X1 U5890 ( .A1(n8591), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8603) );
  AOI21_X1 U5891 ( .B1(n5726), .B2(n8566), .A(n5190), .ZN(n5724) );
  NOR2_X1 U5892 ( .A1(n8550), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8559) );
  NOR2_X1 U5893 ( .A1(n8511), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8534) );
  INV_X1 U5894 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U5895 ( .A1(n9284), .A2(n8534), .ZN(n8550) );
  NOR2_X1 U5896 ( .A1(n5294), .A2(n5162), .ZN(n5293) );
  INV_X1 U5897 ( .A(n9768), .ZN(n9674) );
  OR2_X1 U5898 ( .A1(n9656), .A2(n9667), .ZN(n9671) );
  NAND2_X1 U5899 ( .A1(n8077), .A2(n9389), .ZN(n7940) );
  NAND2_X1 U5900 ( .A1(n7831), .A2(n5747), .ZN(n7929) );
  AND2_X1 U5901 ( .A1(n7827), .A2(n7826), .ZN(n7931) );
  OR2_X1 U5902 ( .A1(n7550), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7584) );
  NOR2_X1 U5903 ( .A1(n7584), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7758) );
  INV_X1 U5904 ( .A(n7798), .ZN(n8727) );
  INV_X1 U5905 ( .A(n8726), .ZN(n7847) );
  INV_X1 U5906 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10210) );
  INV_X1 U5907 ( .A(n8725), .ZN(n7287) );
  OR2_X1 U5908 ( .A1(n8464), .A2(n7191), .ZN(n7687) );
  NAND2_X1 U5909 ( .A1(n7156), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U5910 ( .A1(n5452), .A2(n5451), .ZN(n9202) );
  NAND2_X1 U5911 ( .A1(n8652), .A2(n8651), .ZN(n9721) );
  OR2_X1 U5912 ( .A1(n8830), .A2(n7524), .ZN(n8652) );
  NAND2_X1 U5913 ( .A1(n5285), .A2(n5286), .ZN(n9548) );
  NAND2_X1 U5914 ( .A1(n8628), .A2(n8627), .ZN(n8637) );
  NAND2_X1 U5915 ( .A1(n8601), .A2(n8600), .ZN(n9736) );
  INV_X1 U5916 ( .A(n9694), .ZN(n9774) );
  AND2_X1 U5917 ( .A1(n8163), .A2(n8162), .ZN(n9190) );
  AND2_X1 U5918 ( .A1(n5312), .A2(n5313), .ZN(n8164) );
  NOR2_X1 U5919 ( .A1(n7687), .A2(n7338), .ZN(n8797) );
  NAND2_X1 U5920 ( .A1(n7296), .A2(n6779), .ZN(n7338) );
  INV_X1 U5921 ( .A(n6698), .ZN(n6696) );
  NOR2_X1 U5922 ( .A1(n5743), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U5923 ( .A1(n6695), .A2(n5744), .ZN(n5743) );
  INV_X1 U5924 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5744) );
  INV_X1 U5925 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6694) );
  XNOR2_X1 U5926 ( .A(n6703), .B(P2_IR_REG_23__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U5927 ( .A1(n5659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U5928 ( .A1(n6773), .A2(n5677), .ZN(n7142) );
  NAND2_X1 U5929 ( .A1(n7132), .A2(n7133), .ZN(n6732) );
  NAND2_X1 U5930 ( .A1(n5854), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6147) );
  INV_X1 U5931 ( .A(n6134), .ZN(n5854) );
  NOR2_X1 U5932 ( .A1(n6510), .A2(n5551), .ZN(n5550) );
  INV_X1 U5933 ( .A(n6505), .ZN(n5551) );
  INV_X1 U5934 ( .A(n6212), .ZN(n5857) );
  INV_X1 U5935 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U5936 ( .A1(n5221), .A2(n5532), .ZN(n5531) );
  INV_X1 U5937 ( .A(n9863), .ZN(n5532) );
  NAND2_X1 U5938 ( .A1(n5334), .A2(n5335), .ZN(n9808) );
  INV_X1 U5939 ( .A(n6047), .ZN(n5852) );
  NAND2_X1 U5940 ( .A1(n6839), .A2(n6838), .ZN(n6837) );
  INV_X1 U5941 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U5942 ( .A1(n5321), .A2(n5319), .ZN(n6445) );
  NAND2_X1 U5943 ( .A1(n5320), .A2(n6444), .ZN(n5319) );
  NAND2_X1 U5944 ( .A1(n6637), .A2(n6869), .ZN(n5321) );
  NAND2_X1 U5945 ( .A1(n5330), .A2(n6547), .ZN(n8335) );
  OR2_X1 U5946 ( .A1(n5330), .A2(n6547), .ZN(n8336) );
  AOI21_X1 U5947 ( .B1(n7638), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7637), .ZN(
        n10388) );
  AOI21_X1 U5948 ( .B1(n10891), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10883), .ZN(
        n10415) );
  OR2_X1 U5949 ( .A1(n10944), .A2(n10945), .ZN(n10942) );
  OR2_X1 U5950 ( .A1(n10408), .A2(n10407), .ZN(n10909) );
  AND2_X1 U5951 ( .A1(n10406), .A2(n10917), .ZN(n10408) );
  AND2_X1 U5952 ( .A1(n9031), .A2(n9020), .ZN(n8998) );
  NAND2_X1 U5953 ( .A1(n5398), .A2(n5709), .ZN(n6377) );
  NAND2_X1 U5954 ( .A1(n5710), .A2(n5163), .ZN(n5709) );
  NAND2_X1 U5955 ( .A1(n10513), .A2(n5180), .ZN(n5398) );
  AND2_X1 U5956 ( .A1(n6326), .A2(n6272), .ZN(n10502) );
  INV_X1 U5957 ( .A(n5432), .ZN(n5430) );
  OAI21_X1 U5958 ( .B1(n10587), .B2(n8981), .A(n8978), .ZN(n10563) );
  AND3_X1 U5959 ( .A1(n6237), .A2(n6236), .A3(n6235), .ZN(n10626) );
  AND3_X1 U5960 ( .A1(n6226), .A2(n6225), .A3(n6224), .ZN(n10645) );
  AND2_X1 U5961 ( .A1(n8815), .A2(n5423), .ZN(n10652) );
  NOR2_X1 U5962 ( .A1(n10745), .A2(n5424), .ZN(n5423) );
  INV_X1 U5963 ( .A(n5425), .ZN(n5424) );
  NAND2_X1 U5964 ( .A1(n8815), .A2(n5425), .ZN(n8271) );
  INV_X1 U5965 ( .A(n6177), .ZN(n5856) );
  AOI21_X1 U5966 ( .B1(n5558), .B2(n5560), .A(n5556), .ZN(n5555) );
  INV_X1 U5967 ( .A(n8950), .ZN(n5556) );
  NAND2_X1 U5968 ( .A1(n8815), .A2(n6546), .ZN(n8816) );
  AND2_X1 U5969 ( .A1(n8059), .A2(n8290), .ZN(n8815) );
  INV_X1 U5970 ( .A(n8873), .ZN(n5265) );
  INV_X1 U5971 ( .A(n7898), .ZN(n5266) );
  NOR2_X1 U5972 ( .A1(n7902), .A2(n7907), .ZN(n8059) );
  NAND2_X1 U5973 ( .A1(n5410), .A2(n6105), .ZN(n7899) );
  OR2_X1 U5974 ( .A1(n7662), .A2(n6106), .ZN(n5410) );
  OR2_X1 U5975 ( .A1(n7669), .A2(n7671), .ZN(n7902) );
  AND2_X1 U5976 ( .A1(n8940), .A2(n9078), .ZN(n8870) );
  NAND2_X1 U5977 ( .A1(n5435), .A2(n5434), .ZN(n7386) );
  INV_X1 U5978 ( .A(n5435), .ZN(n7385) );
  AND2_X1 U5979 ( .A1(n6972), .A2(n7064), .ZN(n7048) );
  OR2_X1 U5980 ( .A1(n6993), .A2(n5979), .ZN(n6994) );
  NAND2_X1 U5981 ( .A1(n6867), .A2(n5943), .ZN(n6889) );
  AND2_X1 U5982 ( .A1(n9060), .A2(n9058), .ZN(n6886) );
  NOR2_X1 U5983 ( .A1(n6869), .A2(n6876), .ZN(n6890) );
  NAND2_X1 U5984 ( .A1(n6890), .A2(n7034), .ZN(n6993) );
  NAND2_X1 U5985 ( .A1(n5941), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U5986 ( .A1(n10813), .A2(n6658), .ZN(n10659) );
  NAND2_X1 U5987 ( .A1(n5848), .A2(n5847), .ZN(n10688) );
  AND2_X1 U5988 ( .A1(n6086), .A2(n6085), .ZN(n11160) );
  AND2_X1 U5989 ( .A1(n6655), .A2(n9120), .ZN(n10672) );
  INV_X1 U5990 ( .A(n11178), .ZN(n10770) );
  AND4_X1 U5991 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n7353)
         );
  NAND2_X1 U5992 ( .A1(n5993), .A2(n5170), .ZN(n5714) );
  OR2_X1 U5993 ( .A1(n6739), .A2(n5823), .ZN(n5438) );
  NOR2_X1 U5994 ( .A1(n6958), .A2(n6366), .ZN(n6371) );
  NAND2_X1 U5995 ( .A1(n11166), .A2(n8233), .ZN(n11178) );
  AND2_X1 U5996 ( .A1(n6668), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10813) );
  NAND2_X1 U5997 ( .A1(n5601), .A2(n5600), .ZN(n5599) );
  INV_X1 U5998 ( .A(n6384), .ZN(n5600) );
  AND2_X1 U5999 ( .A1(n6335), .A2(n6334), .ZN(n6353) );
  NOR2_X1 U6000 ( .A1(n6295), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6344) );
  XNOR2_X1 U6001 ( .A(n6299), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8860) );
  INV_X1 U6002 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10303) );
  INV_X1 U6003 ( .A(n5622), .ZN(n5621) );
  AOI21_X1 U6004 ( .B1(n5622), .B2(n5620), .A(n5619), .ZN(n5618) );
  INV_X1 U6005 ( .A(n5794), .ZN(n5619) );
  NAND2_X1 U6006 ( .A1(n6005), .A2(n5780), .ZN(n6021) );
  AND4_X1 U6007 ( .A1(n7555), .A2(n7554), .A3(n7553), .A4(n7552), .ZN(n7793)
         );
  AND4_X1 U6008 ( .A1(n7951), .A2(n7950), .A3(n7949), .A4(n7948), .ZN(n8260)
         );
  XNOR2_X1 U6009 ( .A(n8258), .B(n8257), .ZN(n8259) );
  INV_X1 U6010 ( .A(n5649), .ZN(n5645) );
  NOR2_X1 U6011 ( .A1(n5147), .A2(n9330), .ZN(n5641) );
  NAND2_X1 U6012 ( .A1(n9168), .A2(n9224), .ZN(n5648) );
  OR2_X1 U6013 ( .A1(n7875), .A2(n9389), .ZN(n7876) );
  AND2_X1 U6014 ( .A1(n9359), .A2(n5723), .ZN(n5722) );
  INV_X1 U6015 ( .A(n5667), .ZN(n5666) );
  AOI21_X1 U6016 ( .B1(n5667), .B2(n5665), .A(n5664), .ZN(n5663) );
  INV_X1 U6017 ( .A(n5668), .ZN(n5665) );
  NAND2_X1 U6018 ( .A1(n5662), .A2(n5667), .ZN(n8298) );
  NAND2_X1 U6019 ( .A1(n8258), .A2(n5668), .ZN(n5662) );
  NOR2_X1 U6020 ( .A1(n7703), .A2(n7531), .ZN(n7547) );
  NAND2_X1 U6021 ( .A1(n5661), .A2(n9142), .ZN(n9292) );
  NOR2_X1 U6022 ( .A1(n7705), .A2(n7704), .ZN(n7703) );
  NAND2_X1 U6023 ( .A1(n5675), .A2(n9149), .ZN(n9313) );
  NAND2_X1 U6024 ( .A1(n11105), .A2(n7341), .ZN(n9327) );
  AND2_X1 U6025 ( .A1(n5669), .A2(n5176), .ZN(n8296) );
  NAND2_X1 U6026 ( .A1(n8258), .A2(n5670), .ZN(n5669) );
  NAND2_X1 U6027 ( .A1(n8013), .A2(n8012), .ZN(n8265) );
  INV_X1 U6028 ( .A(n9391), .ZN(n7848) );
  OR2_X1 U6029 ( .A1(n7328), .A2(n7336), .ZN(n9375) );
  INV_X1 U6030 ( .A(n8751), .ZN(n9493) );
  INV_X1 U6031 ( .A(n9246), .ZN(n9578) );
  INV_X1 U6032 ( .A(n9337), .ZN(n9602) );
  AND2_X1 U6033 ( .A1(n5383), .A2(n5381), .ZN(n5380) );
  NAND2_X1 U6034 ( .A1(n7539), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6035 ( .A1(n8711), .A2(n7125), .ZN(n7127) );
  INV_X2 U6036 ( .A(P2_U3893), .ZN(n9483) );
  INV_X1 U6037 ( .A(n5496), .ZN(n11042) );
  INV_X1 U6038 ( .A(n7245), .ZN(n5495) );
  AND2_X1 U6039 ( .A1(n7230), .A2(n7229), .ZN(n7619) );
  NOR2_X1 U6040 ( .A1(n7210), .A2(n7803), .ZN(n7608) );
  NAND2_X1 U6041 ( .A1(n5516), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U6042 ( .A1(n7609), .A2(n5516), .ZN(n5514) );
  INV_X1 U6043 ( .A(n7611), .ZN(n5516) );
  OAI21_X1 U6044 ( .B1(n7769), .B2(n5518), .A(n5517), .ZN(n8195) );
  NAND2_X1 U6045 ( .A1(n7977), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5518) );
  INV_X1 U6046 ( .A(n7975), .ZN(n5519) );
  NOR2_X1 U6047 ( .A1(n11080), .A2(n8017), .ZN(n11079) );
  OAI21_X1 U6048 ( .B1(n11080), .B2(n5522), .A(n5521), .ZN(n8317) );
  NAND2_X1 U6049 ( .A1(n5523), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5522) );
  INV_X1 U6050 ( .A(n8199), .ZN(n5523) );
  OR2_X1 U6051 ( .A1(n8320), .A2(n8319), .ZN(n5527) );
  OR2_X1 U6052 ( .A1(n9405), .A2(n9404), .ZN(n9407) );
  NOR2_X1 U6053 ( .A1(n8353), .A2(n8352), .ZN(n9405) );
  NOR2_X1 U6054 ( .A1(n9413), .A2(n8369), .ZN(n9434) );
  NOR2_X1 U6055 ( .A1(n9434), .A2(n9433), .ZN(n9432) );
  INV_X1 U6056 ( .A(n5486), .ZN(n9444) );
  INV_X1 U6057 ( .A(n5484), .ZN(n9442) );
  NAND2_X1 U6058 ( .A1(n8375), .A2(n8373), .ZN(n9456) );
  AND4_X1 U6059 ( .A1(n8715), .A2(n8433), .A3(n8432), .A4(n8431), .ZN(n9505)
         );
  NAND2_X1 U6060 ( .A1(n8676), .A2(n8675), .ZN(n9713) );
  AND4_X1 U6061 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n9531)
         );
  INV_X1 U6062 ( .A(n9721), .ZN(n9541) );
  NAND2_X1 U6063 ( .A1(n8641), .A2(n8640), .ZN(n9725) );
  NAND2_X1 U6064 ( .A1(n5732), .A2(n5731), .ZN(n9554) );
  NAND2_X1 U6065 ( .A1(n9575), .A2(n9199), .ZN(n9560) );
  OAI21_X1 U6066 ( .B1(n5469), .B2(n9590), .A(n5464), .ZN(n9592) );
  NAND2_X1 U6067 ( .A1(n8589), .A2(n8588), .ZN(n9740) );
  NAND2_X1 U6068 ( .A1(n9625), .A2(n8762), .ZN(n9615) );
  OAI21_X1 U6069 ( .B1(n5292), .B2(n5296), .A(n9194), .ZN(n9668) );
  NAND2_X1 U6070 ( .A1(n8755), .A2(n8754), .ZN(n9684) );
  NAND2_X1 U6071 ( .A1(n5312), .A2(n5311), .ZN(n9191) );
  NAND2_X1 U6072 ( .A1(n5718), .A2(n8123), .ZN(n8160) );
  NAND2_X1 U6073 ( .A1(n8122), .A2(n8739), .ZN(n5718) );
  OAI21_X1 U6074 ( .B1(n8027), .B2(n7524), .A(n8029), .ZN(n8226) );
  AND2_X1 U6075 ( .A1(n7936), .A2(n7935), .ZN(n8024) );
  NAND2_X1 U6076 ( .A1(n5739), .A2(n8446), .ZN(n7944) );
  INV_X1 U6077 ( .A(n7931), .ZN(n7888) );
  INV_X1 U6078 ( .A(n7911), .ZN(n9389) );
  AND3_X1 U6079 ( .A1(n7538), .A2(n7537), .A3(n7536), .ZN(n7723) );
  INV_X1 U6080 ( .A(n7793), .ZN(n9390) );
  INV_X1 U6081 ( .A(n9662), .ZN(n11116) );
  INV_X1 U6082 ( .A(n11105), .ZN(n11118) );
  NAND4_X1 U6083 ( .A1(n7335), .A2(n7334), .A3(n7333), .A4(n7332), .ZN(n9392)
         );
  MUX2_X1 U6084 ( .A(n10974), .B(n9806), .S(n7130), .Z(n7686) );
  NAND2_X1 U6085 ( .A1(n7339), .A2(n7693), .ZN(n11105) );
  OR2_X1 U6086 ( .A1(n7684), .A2(n11103), .ZN(n9662) );
  INV_X1 U6087 ( .A(n9678), .ZN(n9695) );
  NOR2_X1 U6088 ( .A1(n7194), .A2(n7193), .ZN(n8232) );
  OR3_X1 U6089 ( .A1(n9760), .A2(n9759), .A3(n9758), .ZN(n9796) );
  INV_X2 U6090 ( .A(n11192), .ZN(n11195) );
  AND2_X1 U6091 ( .A1(n7295), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6779) );
  NAND2_X1 U6092 ( .A1(n7318), .A2(n6778), .ZN(n6783) );
  NAND2_X1 U6093 ( .A1(n5658), .A2(n5657), .ZN(n7147) );
  AOI21_X1 U6094 ( .B1(n5660), .B2(n7131), .A(n7131), .ZN(n5657) );
  INV_X1 U6095 ( .A(n8556), .ZN(n9486) );
  INV_X1 U6096 ( .A(n7824), .ZN(n7771) );
  INV_X1 U6097 ( .A(n11034), .ZN(n7243) );
  OAI21_X1 U6098 ( .B1(n7399), .B2(n6482), .A(n6481), .ZN(n7440) );
  OAI21_X1 U6099 ( .B1(n9921), .B2(n9173), .A(n9174), .ZN(n9175) );
  NAND2_X1 U6100 ( .A1(n8832), .A2(n6454), .ZN(n6984) );
  NAND2_X1 U6101 ( .A1(n5340), .A2(n5338), .ZN(n9817) );
  AOI21_X1 U6102 ( .B1(n5341), .B2(n5343), .A(n5339), .ZN(n5338) );
  AND2_X1 U6103 ( .A1(n5547), .A2(n5342), .ZN(n5341) );
  NAND2_X1 U6104 ( .A1(n6208), .A2(n6207), .ZN(n10657) );
  AND4_X1 U6105 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(n8002)
         );
  NAND2_X1 U6106 ( .A1(n6033), .A2(n6032), .ZN(n8009) );
  OAI21_X1 U6107 ( .B1(n9910), .B2(n5339), .A(n5543), .ZN(n9826) );
  NAND2_X1 U6108 ( .A1(n6231), .A2(n6230), .ZN(n10725) );
  AND2_X1 U6109 ( .A1(n5325), .A2(n7813), .ZN(n8067) );
  AND2_X1 U6110 ( .A1(n5530), .A2(n5528), .ZN(n9924) );
  NAND2_X1 U6111 ( .A1(n5530), .A2(n5531), .ZN(n9835) );
  OR2_X1 U6112 ( .A1(n8830), .A2(n6396), .ZN(n5886) );
  NAND2_X1 U6113 ( .A1(n5535), .A2(n8336), .ZN(n9843) );
  NAND2_X1 U6114 ( .A1(n8335), .A2(n8338), .ZN(n5535) );
  NAND2_X1 U6115 ( .A1(n9808), .A2(n6614), .ZN(n9865) );
  NAND2_X1 U6116 ( .A1(n5316), .A2(n5317), .ZN(n9876) );
  NAND2_X1 U6117 ( .A1(n5318), .A2(n5157), .ZN(n5317) );
  INV_X1 U6118 ( .A(n6983), .ZN(n5318) );
  NAND2_X1 U6119 ( .A1(n9876), .A2(n9875), .ZN(n9874) );
  AND4_X1 U6120 ( .A1(n6040), .A2(n6039), .A3(n6038), .A4(n6037), .ZN(n7868)
         );
  NAND2_X1 U6121 ( .A1(n8066), .A2(n5552), .ZN(n8150) );
  AND2_X1 U6122 ( .A1(n8151), .A2(n6527), .ZN(n5552) );
  AND2_X1 U6123 ( .A1(n8066), .A2(n6527), .ZN(n8152) );
  NOR2_X1 U6124 ( .A1(n9897), .A2(n9895), .ZN(n9900) );
  AND2_X1 U6125 ( .A1(n6669), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9917) );
  NAND2_X1 U6126 ( .A1(n5332), .A2(n5333), .ZN(n5331) );
  OR2_X1 U6127 ( .A1(n9922), .A2(n9923), .ZN(n6632) );
  INV_X1 U6128 ( .A(n9926), .ZN(n9919) );
  INV_X1 U6129 ( .A(n10685), .ZN(n9933) );
  INV_X1 U6130 ( .A(n10694), .ZN(n10503) );
  OR2_X1 U6131 ( .A1(n10540), .A2(n6258), .ZN(n5894) );
  NAND2_X1 U6132 ( .A1(n5901), .A2(n5900), .ZN(n10710) );
  INV_X1 U6133 ( .A(n10626), .ZN(n10589) );
  AND4_X1 U6134 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n10349)
         );
  INV_X1 U6135 ( .A(n6997), .ZN(n10356) );
  AOI21_X1 U6136 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6800), .A(n6799), .ZN(
        n6803) );
  AOI21_X1 U6137 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6852), .A(n6848), .ZN(
        n6850) );
  AOI21_X1 U6138 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10963), .A(n10953), .ZN(
        n10885) );
  AND2_X1 U6139 ( .A1(n10939), .A2(n10938), .ZN(n10941) );
  OR2_X1 U6140 ( .A1(n6755), .A2(n9124), .ZN(n10952) );
  INV_X1 U6141 ( .A(n10956), .ZN(n10910) );
  NOR2_X1 U6142 ( .A1(n10471), .A2(n10479), .ZN(n10473) );
  AND2_X1 U6143 ( .A1(n6294), .A2(n6293), .ZN(n10676) );
  NAND2_X1 U6144 ( .A1(n10512), .A2(n5712), .ZN(n10499) );
  AND2_X1 U6145 ( .A1(n5583), .A2(n5582), .ZN(n10533) );
  NAND2_X1 U6146 ( .A1(n5696), .A2(n5700), .ZN(n10547) );
  NAND2_X1 U6147 ( .A1(n10584), .A2(n5701), .ZN(n5696) );
  INV_X1 U6148 ( .A(n5698), .ZN(n5701) );
  INV_X1 U6149 ( .A(n10710), .ZN(n10693) );
  NAND2_X1 U6150 ( .A1(n10584), .A2(n6250), .ZN(n10565) );
  NAND2_X1 U6151 ( .A1(n5683), .A2(n5694), .ZN(n10606) );
  AND2_X1 U6152 ( .A1(n5686), .A2(n5684), .ZN(n10604) );
  NAND2_X1 U6153 ( .A1(n5688), .A2(n5689), .ZN(n10621) );
  INV_X1 U6154 ( .A(n5690), .ZN(n5689) );
  AOI21_X1 U6155 ( .B1(n8270), .B2(n6200), .A(n5693), .ZN(n10650) );
  NAND2_X1 U6156 ( .A1(n5557), .A2(n8948), .ZN(n8145) );
  NAND2_X1 U6157 ( .A1(n8822), .A2(n6316), .ZN(n5557) );
  NAND2_X1 U6158 ( .A1(n5405), .A2(n5406), .ZN(n8814) );
  OR2_X1 U6159 ( .A1(n7662), .A2(n5409), .ZN(n5405) );
  NAND2_X1 U6160 ( .A1(n5707), .A2(n5705), .ZN(n8050) );
  NAND2_X1 U6161 ( .A1(n5707), .A2(n6124), .ZN(n8048) );
  NAND2_X1 U6162 ( .A1(n6312), .A2(n8894), .ZN(n7510) );
  NAND2_X1 U6163 ( .A1(n7047), .A2(n8868), .ZN(n7046) );
  NAND2_X1 U6164 ( .A1(n7026), .A2(n6012), .ZN(n7047) );
  NAND2_X1 U6165 ( .A1(n5579), .A2(n5576), .ZN(n5574) );
  INV_X1 U6166 ( .A(n5941), .ZN(n7011) );
  AOI21_X1 U6167 ( .B1(n9219), .B2(n8854), .A(n5226), .ZN(n10779) );
  INV_X1 U6168 ( .A(n10538), .ZN(n10785) );
  INV_X1 U6169 ( .A(n10556), .ZN(n10789) );
  INV_X1 U6170 ( .A(n10657), .ZN(n10807) );
  INV_X1 U6171 ( .A(n6540), .ZN(n8290) );
  INV_X1 U6172 ( .A(n7907), .ZN(n8159) );
  OR2_X1 U6173 ( .A1(n8027), .A2(n6396), .ZN(n6065) );
  INV_X1 U6174 ( .A(n7405), .ZN(n7064) );
  AND2_X1 U6175 ( .A1(n10321), .A2(n10325), .ZN(n5597) );
  XNOR2_X1 U6176 ( .A(n8704), .B(n8703), .ZN(n10821) );
  OAI22_X1 U6177 ( .A1(n8700), .A2(n8699), .B1(SI_30_), .B2(n8698), .ZN(n8704)
         );
  OR2_X1 U6178 ( .A1(n5864), .A2(n5969), .ZN(n5844) );
  INV_X1 U6179 ( .A(n6353), .ZN(n8308) );
  NAND2_X1 U6180 ( .A1(n6340), .A2(n6339), .ZN(n8269) );
  XNOR2_X1 U6181 ( .A(n6346), .B(n5838), .ZN(n8245) );
  NAND2_X1 U6182 ( .A1(n6345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U6183 ( .A1(n6344), .A2(n6343), .ZN(n6345) );
  NOR2_X1 U6184 ( .A1(n6342), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n6343) );
  INV_X1 U6185 ( .A(n6419), .ZN(n8088) );
  INV_X1 U6186 ( .A(n8860), .ZN(n9054) );
  NAND2_X1 U6187 ( .A1(n5616), .A2(n5615), .ZN(n6185) );
  NAND2_X1 U6188 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  AND2_X1 U6189 ( .A1(n6172), .A2(n6160), .ZN(n10441) );
  NAND2_X1 U6190 ( .A1(n5633), .A2(n5630), .ZN(n6141) );
  INV_X1 U6191 ( .A(n5632), .ZN(n5630) );
  AND2_X1 U6192 ( .A1(n6114), .A2(n6128), .ZN(n10948) );
  NAND2_X1 U6193 ( .A1(n5624), .A2(n5622), .ZN(n6089) );
  NAND2_X1 U6194 ( .A1(n6022), .A2(n5297), .ZN(n7750) );
  NAND2_X1 U6195 ( .A1(n6020), .A2(n6021), .ZN(n6022) );
  NAND2_X1 U6196 ( .A1(n5298), .A2(n5782), .ZN(n5297) );
  INV_X1 U6197 ( .A(n6021), .ZN(n5298) );
  NAND2_X1 U6198 ( .A1(n5151), .A2(n5252), .ZN(n5251) );
  OAI21_X1 U6199 ( .B1(n7311), .B2(n9483), .A(n5721), .ZN(P2_U3493) );
  NAND2_X1 U6200 ( .A1(n9483), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5721) );
  INV_X1 U6201 ( .A(n5520), .ZN(n7976) );
  INV_X1 U6202 ( .A(n9489), .ZN(n5264) );
  NAND2_X1 U6203 ( .A1(n5203), .A2(n5247), .ZN(P2_U3201) );
  NOR2_X1 U6204 ( .A1(n5169), .A2(n5248), .ZN(n5247) );
  AOI21_X1 U6205 ( .B1(n5148), .B2(n11086), .A(n5250), .ZN(n5249) );
  OR2_X1 U6206 ( .A1(n9177), .A2(n6653), .ZN(n6683) );
  OR2_X1 U6207 ( .A1(n9128), .A2(n9127), .ZN(n5269) );
  AND2_X1 U6208 ( .A1(n5595), .A2(n5158), .ZN(n8812) );
  NAND2_X1 U6209 ( .A1(n6680), .A2(n7604), .ZN(n6374) );
  NAND2_X1 U6210 ( .A1(n5421), .A2(n6413), .ZN(P1_U3519) );
  NOR2_X1 U6211 ( .A1(n5222), .A2(n6412), .ZN(n6413) );
  OAI21_X1 U6212 ( .B1(n5593), .B2(n5422), .A(n11185), .ZN(n5421) );
  NAND2_X1 U6213 ( .A1(n6680), .A2(n6368), .ZN(n6369) );
  OR2_X1 U6214 ( .A1(n9197), .A2(n9196), .ZN(n5469) );
  NAND2_X1 U6215 ( .A1(n5616), .A2(n5156), .ZN(n5141) );
  OR2_X1 U6216 ( .A1(n8390), .A2(n8364), .ZN(n5142) );
  NAND2_X1 U6217 ( .A1(n8281), .A2(n6544), .ZN(n5330) );
  OR2_X1 U6218 ( .A1(n8111), .A2(n8737), .ZN(n5143) );
  INV_X2 U6219 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5971) );
  INV_X1 U6220 ( .A(n8566), .ZN(n8762) );
  NAND2_X1 U6221 ( .A1(n5570), .A2(n8998), .ZN(n5569) );
  NAND2_X1 U6222 ( .A1(n8294), .A2(n8293), .ZN(n5144) );
  XNOR2_X1 U6223 ( .A(n6701), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6763) );
  OR2_X1 U6224 ( .A1(n5539), .A2(n7438), .ZN(n5145) );
  AND2_X1 U6225 ( .A1(n9755), .A2(n9628), .ZN(n5146) );
  INV_X1 U6226 ( .A(n9199), .ZN(n5289) );
  INV_X1 U6227 ( .A(n8784), .ZN(n9700) );
  AND2_X1 U6228 ( .A1(n5646), .A2(n5648), .ZN(n5147) );
  INV_X1 U6229 ( .A(n9162), .ZN(n9538) );
  AND4_X1 U6230 ( .A1(n8673), .A2(n8672), .A3(n8671), .A4(n8670), .ZN(n9162)
         );
  AND2_X1 U6231 ( .A1(n6146), .A2(n6145), .ZN(n6546) );
  XOR2_X1 U6232 ( .A(n8405), .B(n8404), .Z(n5148) );
  NAND2_X1 U6233 ( .A1(n9564), .A2(n8767), .ZN(n5149) );
  INV_X1 U6234 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7145) );
  NAND2_X1 U6235 ( .A1(n8701), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5150) );
  NOR2_X1 U6236 ( .A1(n5348), .A2(n5352), .ZN(n5151) );
  AND2_X1 U6237 ( .A1(n6186), .A2(n5323), .ZN(n5152) );
  AND2_X1 U6238 ( .A1(n5528), .A2(n5534), .ZN(n5153) );
  INV_X1 U6239 ( .A(n9809), .ZN(n5336) );
  INV_X1 U6240 ( .A(n9517), .ZN(n9227) );
  NAND2_X1 U6241 ( .A1(n9667), .A2(n9685), .ZN(n5154) );
  NAND2_X1 U6242 ( .A1(n5646), .A2(n5188), .ZN(n5155) );
  OR2_X1 U6243 ( .A1(n5805), .A2(SI_17_), .ZN(n5156) );
  XNOR2_X1 U6244 ( .A(n6541), .B(n6542), .ZN(n8280) );
  NAND2_X1 U6245 ( .A1(n6448), .A2(n6449), .ZN(n8832) );
  NAND2_X1 U6246 ( .A1(n6461), .A2(n6460), .ZN(n5157) );
  INV_X1 U6247 ( .A(n9895), .ZN(n5332) );
  AND2_X1 U6248 ( .A1(n6348), .A2(n6298), .ZN(n6419) );
  AND2_X1 U6249 ( .A1(n6409), .A2(n6408), .ZN(n5158) );
  AND2_X1 U6250 ( .A1(n7097), .A2(n8839), .ZN(n7757) );
  AND2_X1 U6251 ( .A1(n10514), .A2(n5431), .ZN(n5159) );
  INV_X1 U6252 ( .A(n8499), .ZN(n8123) );
  AND2_X1 U6253 ( .A1(n8265), .A2(n8293), .ZN(n8499) );
  AND2_X1 U6254 ( .A1(n9572), .A2(n9246), .ZN(n5160) );
  NAND2_X1 U6255 ( .A1(n7907), .A2(n10348), .ZN(n5161) );
  AND2_X1 U6256 ( .A1(n9674), .A2(n9694), .ZN(n5162) );
  OR2_X1 U6257 ( .A1(n10679), .A2(n9933), .ZN(n5163) );
  AND2_X1 U6258 ( .A1(n5705), .A2(n5411), .ZN(n5164) );
  AND2_X1 U6259 ( .A1(n5373), .A2(n5378), .ZN(n5165) );
  AND3_X1 U6260 ( .A1(n7118), .A2(n7117), .A3(n7116), .ZN(n7304) );
  AND2_X1 U6261 ( .A1(n6685), .A2(n6424), .ZN(n5166) );
  XOR2_X1 U6262 ( .A(n6763), .B(P2_B_REG_SCAN_IN), .Z(n5167) );
  INV_X1 U6263 ( .A(n8868), .ZN(n5397) );
  NAND2_X1 U6264 ( .A1(n9908), .A2(n9907), .ZN(n5546) );
  INV_X1 U6265 ( .A(n5546), .ZN(n5339) );
  AND2_X1 U6266 ( .A1(n5467), .A2(n9595), .ZN(n5168) );
  INV_X1 U6267 ( .A(n10586), .ZN(n5418) );
  INV_X1 U6268 ( .A(n7428), .ZN(n11104) );
  OAI211_X1 U6269 ( .C1(n7524), .C2(n8842), .A(n7136), .B(n7135), .ZN(n7428)
         );
  INV_X1 U6270 ( .A(n10550), .ZN(n5585) );
  INV_X1 U6271 ( .A(n9224), .ZN(n5651) );
  AND3_X1 U6272 ( .A1(n9472), .A2(n5475), .A3(n5482), .ZN(n5169) );
  OR2_X1 U6273 ( .A1(n6707), .A2(n6801), .ZN(n5170) );
  XNOR2_X1 U6274 ( .A(n5598), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5871) );
  AND2_X1 U6275 ( .A1(n8505), .A2(n9384), .ZN(n5171) );
  OR2_X1 U6276 ( .A1(n9635), .A2(n9613), .ZN(n5172) );
  OR2_X1 U6277 ( .A1(n6548), .A2(n8338), .ZN(n5173) );
  NOR2_X1 U6278 ( .A1(n5348), .A2(n5350), .ZN(n5174) );
  OR2_X1 U6279 ( .A1(n9617), .A2(n9347), .ZN(n5175) );
  NAND2_X1 U6280 ( .A1(n8257), .A2(n9386), .ZN(n5176) );
  AND2_X1 U6281 ( .A1(n10579), .A2(n10590), .ZN(n5177) );
  INV_X1 U6282 ( .A(n10590), .ZN(n10551) );
  AND2_X1 U6283 ( .A1(n5469), .A2(n5175), .ZN(n5178) );
  INV_X1 U6284 ( .A(n6680), .ZN(n10493) );
  NAND2_X1 U6285 ( .A1(n6398), .A2(n6397), .ZN(n8809) );
  INV_X1 U6286 ( .A(n8809), .ZN(n5429) );
  INV_X1 U6287 ( .A(n9393), .ZN(n7565) );
  NAND2_X1 U6288 ( .A1(n7157), .A2(n5380), .ZN(n9393) );
  AND2_X1 U6289 ( .A1(n9167), .A2(n9716), .ZN(n5179) );
  OR2_X1 U6290 ( .A1(n8372), .A2(n9457), .ZN(n8375) );
  AND2_X1 U6291 ( .A1(n5163), .A2(n10526), .ZN(n5180) );
  OR2_X1 U6292 ( .A1(n9708), .A2(n9517), .ZN(n5181) );
  AND2_X1 U6293 ( .A1(n5431), .A2(n5429), .ZN(n5182) );
  INV_X1 U6294 ( .A(n9277), .ZN(n9561) );
  AND4_X1 U6295 ( .A1(n8649), .A2(n8648), .A3(n8647), .A4(n8646), .ZN(n9277)
         );
  AND2_X1 U6296 ( .A1(n5649), .A2(n5651), .ZN(n5183) );
  INV_X1 U6297 ( .A(n10753), .ZN(n9862) );
  NAND2_X1 U6298 ( .A1(n6175), .A2(n6174), .ZN(n10753) );
  AND2_X1 U6299 ( .A1(n5734), .A2(n8773), .ZN(n5184) );
  AND2_X1 U6300 ( .A1(n5460), .A2(n5458), .ZN(n5185) );
  OR2_X1 U6301 ( .A1(n5538), .A2(n7437), .ZN(n5186) );
  AND2_X1 U6302 ( .A1(n5536), .A2(n5186), .ZN(n5187) );
  INV_X1 U6303 ( .A(n8716), .ZN(n9702) );
  OR2_X1 U6304 ( .A1(n9168), .A2(n5645), .ZN(n5188) );
  AND2_X1 U6305 ( .A1(n6553), .A2(n5328), .ZN(n5189) );
  INV_X1 U6306 ( .A(n5534), .ZN(n5533) );
  NAND2_X1 U6307 ( .A1(n5221), .A2(n6614), .ZN(n5534) );
  NOR2_X1 U6308 ( .A1(n9744), .A2(n9347), .ZN(n5190) );
  NOR2_X1 U6309 ( .A1(n10352), .A2(n7049), .ZN(n5191) );
  NOR2_X1 U6310 ( .A1(n8290), .A2(n10764), .ZN(n5192) );
  AND2_X1 U6311 ( .A1(n6481), .A2(n5145), .ZN(n5193) );
  INV_X1 U6312 ( .A(n5678), .ZN(n5677) );
  NAND2_X1 U6313 ( .A1(n5680), .A2(n5679), .ZN(n5678) );
  INV_X1 U6314 ( .A(n5287), .ZN(n5286) );
  NOR2_X1 U6315 ( .A1(n5288), .A2(n5160), .ZN(n5287) );
  AND2_X1 U6316 ( .A1(n9190), .A2(n9688), .ZN(n5194) );
  AND2_X1 U6317 ( .A1(n8637), .A2(n9578), .ZN(n5195) );
  INV_X1 U6318 ( .A(n5695), .ZN(n5693) );
  NAND2_X1 U6319 ( .A1(n10745), .A2(n10344), .ZN(n5695) );
  NOR2_X1 U6320 ( .A1(n9667), .A2(n8758), .ZN(n5196) );
  NOR2_X1 U6321 ( .A1(n9736), .A2(n9602), .ZN(n5197) );
  INV_X1 U6322 ( .A(n5720), .ZN(n5719) );
  OAI21_X1 U6323 ( .B1(n8739), .B2(n8499), .A(n8737), .ZN(n5720) );
  INV_X1 U6324 ( .A(n5713), .ZN(n5712) );
  NOR2_X1 U6325 ( .A1(n10517), .A2(n10694), .ZN(n5713) );
  AND2_X1 U6326 ( .A1(n5841), .A2(n5840), .ZN(n5198) );
  AND2_X1 U6327 ( .A1(n5469), .A2(n5467), .ZN(n5199) );
  NAND2_X1 U6328 ( .A1(n10538), .A2(n10684), .ZN(n8991) );
  OR2_X1 U6329 ( .A1(n10579), .A2(n10590), .ZN(n5200) );
  INV_X1 U6330 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7111) );
  NOR2_X1 U6331 ( .A1(n10495), .A2(n6331), .ZN(n5201) );
  INV_X1 U6332 ( .A(n5583), .ZN(n10548) );
  OR2_X1 U6333 ( .A1(n5586), .A2(n5584), .ZN(n5583) );
  NAND2_X1 U6334 ( .A1(n8437), .A2(n8436), .ZN(n9708) );
  AND2_X1 U6335 ( .A1(n6636), .A2(n6635), .ZN(n9173) );
  AND2_X1 U6336 ( .A1(n9708), .A2(n9517), .ZN(n5202) );
  AND2_X1 U6337 ( .A1(n8381), .A2(n5249), .ZN(n5203) );
  INV_X1 U6338 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U6339 ( .A1(n8659), .A2(n9545), .ZN(n5204) );
  NAND2_X1 U6340 ( .A1(n5176), .A2(n8295), .ZN(n5205) );
  INV_X1 U6341 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10325) );
  NOR2_X1 U6342 ( .A1(n7579), .A2(n7580), .ZN(n5206) );
  AND2_X1 U6343 ( .A1(n9160), .A2(n5653), .ZN(n5207) );
  AND2_X1 U6344 ( .A1(n9553), .A2(n8650), .ZN(n5208) );
  AND2_X1 U6345 ( .A1(n9083), .A2(n8940), .ZN(n5209) );
  AND2_X1 U6346 ( .A1(n10512), .A2(n5711), .ZN(n5210) );
  INV_X1 U6347 ( .A(n5337), .ZN(n9921) );
  NOR2_X1 U6348 ( .A1(n9490), .A2(n5262), .ZN(n5211) );
  INV_X1 U6349 ( .A(n9685), .ZN(n5296) );
  AND2_X1 U6350 ( .A1(n9194), .A2(n8528), .ZN(n9685) );
  NAND2_X1 U6351 ( .A1(n8265), .A2(n9385), .ZN(n5212) );
  AND2_X1 U6352 ( .A1(n5742), .A2(n7095), .ZN(n5213) );
  AND2_X1 U6353 ( .A1(n5157), .A2(n6454), .ZN(n5214) );
  AND2_X1 U6354 ( .A1(n9143), .A2(n9142), .ZN(n5215) );
  OR2_X1 U6355 ( .A1(n5284), .A2(n5280), .ZN(n5216) );
  AND2_X1 U6356 ( .A1(n5196), .A2(n8756), .ZN(n5217) );
  NAND2_X1 U6357 ( .A1(n9012), .A2(n9011), .ZN(n5218) );
  OAI21_X1 U6358 ( .B1(n8990), .B2(n5581), .A(n8991), .ZN(n5580) );
  INV_X1 U6359 ( .A(n5569), .ZN(n5568) );
  NAND2_X1 U6360 ( .A1(n5786), .A2(n5785), .ZN(n5219) );
  INV_X1 U6361 ( .A(n5737), .ZN(n5736) );
  NAND2_X1 U6362 ( .A1(n5738), .A2(n8446), .ZN(n5737) );
  INV_X1 U6363 ( .A(n5577), .ZN(n5576) );
  NAND2_X1 U6364 ( .A1(n9061), .A2(n8905), .ZN(n5577) );
  NOR2_X1 U6365 ( .A1(n9834), .A2(n5529), .ZN(n5528) );
  INV_X1 U6366 ( .A(n5352), .ZN(n5351) );
  AND2_X1 U6367 ( .A1(n8788), .A2(n8787), .ZN(n5352) );
  NOR2_X1 U6368 ( .A1(n6632), .A2(n5153), .ZN(n5220) );
  NAND2_X1 U6369 ( .A1(n8270), .A2(n5691), .ZN(n5688) );
  NAND2_X1 U6370 ( .A1(n8026), .A2(n8025), .ZN(n8110) );
  NAND2_X1 U6371 ( .A1(n9682), .A2(n8756), .ZN(n9656) );
  INV_X1 U6372 ( .A(n10679), .ZN(n5433) );
  NAND2_X1 U6373 ( .A1(n5739), .A2(n5736), .ZN(n8033) );
  INV_X1 U6374 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5838) );
  INV_X1 U6375 ( .A(n8475), .ZN(n5361) );
  NOR2_X1 U6376 ( .A1(n8310), .A2(n8311), .ZN(n8353) );
  OAI21_X1 U6377 ( .B1(n5717), .B2(n5720), .A(n5715), .ZN(n8753) );
  OAI21_X1 U6378 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9319) );
  INV_X1 U6379 ( .A(n8464), .ZN(n8695) );
  XNOR2_X1 U6380 ( .A(n6727), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7535) );
  OR2_X1 U6381 ( .A1(n6621), .A2(n6620), .ZN(n5221) );
  NAND2_X1 U6382 ( .A1(n8280), .A2(n8282), .ZN(n8281) );
  NAND2_X1 U6383 ( .A1(n5404), .A2(n5403), .ZN(n8813) );
  INV_X1 U6384 ( .A(n10346), .ZN(n10756) );
  NAND2_X1 U6385 ( .A1(n8664), .A2(n8663), .ZN(n9717) );
  INV_X1 U6386 ( .A(n9717), .ZN(n5459) );
  NAND2_X1 U6387 ( .A1(n8815), .A2(n5427), .ZN(n5428) );
  INV_X1 U6388 ( .A(n5439), .ZN(n10630) );
  NOR2_X1 U6389 ( .A1(n5429), .A2(n10806), .ZN(n5222) );
  AND2_X1 U6390 ( .A1(n5809), .A2(n10154), .ZN(n5223) );
  AOI21_X1 U6391 ( .B1(n9642), .B2(n5307), .A(n5146), .ZN(n5304) );
  AND2_X1 U6392 ( .A1(n5527), .A2(n5142), .ZN(n5224) );
  INV_X1 U6393 ( .A(n5156), .ZN(n5617) );
  OAI22_X1 U6394 ( .A1(n7789), .A2(n7788), .B1(n7787), .B2(n9391), .ZN(n7928)
         );
  INV_X1 U6395 ( .A(n9330), .ZN(n9370) );
  OAI21_X1 U6396 ( .B1(n6958), .B2(n6957), .A(n10659), .ZN(n10661) );
  OR2_X1 U6397 ( .A1(n8746), .A2(n8787), .ZN(n7299) );
  NAND2_X1 U6398 ( .A1(n9874), .A2(n6468), .ZN(n7399) );
  NAND2_X1 U6399 ( .A1(n6421), .A2(n6419), .ZN(n6423) );
  AND2_X1 U6400 ( .A1(n8318), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5225) );
  NOR2_X1 U6401 ( .A1(n8853), .A2(n9221), .ZN(n5226) );
  XNOR2_X1 U6402 ( .A(n6697), .B(P2_IR_REG_26__SCAN_IN), .ZN(n7173) );
  NAND2_X1 U6403 ( .A1(n6512), .A2(n7734), .ZN(n7812) );
  AND2_X1 U6404 ( .A1(n5574), .A2(n5575), .ZN(n5227) );
  AND2_X1 U6405 ( .A1(n6765), .A2(n7173), .ZN(n7172) );
  NAND2_X1 U6406 ( .A1(n6501), .A2(n6500), .ZN(n7863) );
  NAND3_X1 U6407 ( .A1(n6773), .A2(n6693), .A3(n5745), .ZN(n5228) );
  INV_X1 U6408 ( .A(n7159), .ZN(n7250) );
  NOR2_X1 U6409 ( .A1(n11079), .A2(n8197), .ZN(n5229) );
  AND2_X1 U6410 ( .A1(n5520), .A2(n5519), .ZN(n5230) );
  NAND2_X1 U6411 ( .A1(n6516), .A2(n6517), .ZN(n5231) );
  AND2_X1 U6412 ( .A1(n8386), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5232) );
  NOR2_X1 U6413 ( .A1(n7495), .A2(n5722), .ZN(n5233) );
  NOR2_X1 U6414 ( .A1(n7990), .A2(n7991), .ZN(n5234) );
  INV_X1 U6415 ( .A(n6421), .ZN(n10464) );
  INV_X1 U6416 ( .A(n7456), .ZN(n5434) );
  NAND3_X1 U6417 ( .A1(n5910), .A2(n5909), .A3(n5908), .ZN(n6875) );
  INV_X1 U6418 ( .A(n7014), .ZN(n5320) );
  INV_X1 U6419 ( .A(n11020), .ZN(n11086) );
  AND2_X2 U6420 ( .A1(n6371), .A2(n6651), .ZN(n11181) );
  AND2_X1 U6421 ( .A1(n5479), .A2(n5478), .ZN(n5235) );
  AND2_X1 U6422 ( .A1(n5481), .A2(n8401), .ZN(n5236) );
  NAND2_X1 U6423 ( .A1(n6880), .A2(n6874), .ZN(n6873) );
  NOR2_X1 U6424 ( .A1(n7608), .A2(n7609), .ZN(n5237) );
  NOR2_X1 U6425 ( .A1(n7613), .A2(n7614), .ZN(n5238) );
  NOR2_X1 U6426 ( .A1(n11026), .A2(n11025), .ZN(n5239) );
  AND2_X1 U6427 ( .A1(n5496), .A2(n5495), .ZN(n5240) );
  NOR2_X1 U6428 ( .A1(n11010), .A2(n7241), .ZN(n5241) );
  INV_X1 U6429 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5382) );
  AND2_X1 U6430 ( .A1(n7981), .A2(n7989), .ZN(n5260) );
  XNOR2_X1 U6431 ( .A(n7974), .B(n7989), .ZN(n7769) );
  AOI21_X1 U6432 ( .B1(n10484), .B2(n10746), .A(n5267), .ZN(n6372) );
  INV_X1 U6433 ( .A(n10746), .ZN(n10713) );
  NAND2_X1 U6434 ( .A1(n6868), .A2(n6866), .ZN(n6867) );
  NOR2_X1 U6435 ( .A1(n9424), .A2(n9425), .ZN(n9423) );
  OR2_X2 U6436 ( .A1(n5686), .A2(n5416), .ZN(n5412) );
  INV_X1 U6437 ( .A(n5593), .ZN(n5594) );
  OR2_X1 U6438 ( .A1(n9491), .A2(n11090), .ZN(n5263) );
  NAND2_X1 U6439 ( .A1(n7372), .A2(n7371), .ZN(n7370) );
  OAI21_X1 U6440 ( .B1(n7508), .B2(n10349), .A(n11160), .ZN(n5682) );
  NAND2_X1 U6441 ( .A1(n8140), .A2(n5750), .ZN(n8247) );
  NAND2_X1 U6442 ( .A1(n8802), .A2(n11178), .ZN(n5596) );
  NAND2_X1 U6443 ( .A1(n5402), .A2(n5401), .ZN(n5400) );
  NAND2_X1 U6444 ( .A1(n6970), .A2(n8917), .ZN(n6969) );
  NAND3_X1 U6445 ( .A1(n8986), .A2(n9028), .A3(n9027), .ZN(n8987) );
  NAND2_X1 U6446 ( .A1(n8966), .A2(n8967), .ZN(n8977) );
  NAND2_X1 U6447 ( .A1(n5242), .A2(n9079), .ZN(n8944) );
  NAND2_X1 U6448 ( .A1(n8941), .A2(n5209), .ZN(n5242) );
  NAND2_X1 U6449 ( .A1(n9013), .A2(n9039), .ZN(n5605) );
  NAND2_X1 U6450 ( .A1(n5273), .A2(n5270), .ZN(n9010) );
  AOI21_X1 U6451 ( .B1(n6043), .B2(n6042), .A(n5788), .ZN(n6055) );
  AOI21_X1 U6452 ( .B1(n8962), .B2(n9091), .A(n9051), .ZN(n8963) );
  OAI21_X1 U6453 ( .B1(n7210), .B2(n5515), .A(n5514), .ZN(n7768) );
  NAND2_X1 U6454 ( .A1(n5734), .A2(n5729), .ZN(n9544) );
  NAND3_X1 U6455 ( .A1(n5345), .A2(n5346), .A3(n5251), .ZN(P2_U3296) );
  NAND3_X1 U6456 ( .A1(n8783), .A2(n8782), .A3(n5256), .ZN(n5255) );
  AND2_X4 U6457 ( .A1(n6734), .A2(n6687), .ZN(n6773) );
  NAND3_X1 U6458 ( .A1(n5264), .A2(n5263), .A3(n5211), .ZN(P2_U3200) );
  NAND2_X1 U6459 ( .A1(n6315), .A2(n9084), .ZN(n8822) );
  NAND2_X1 U6460 ( .A1(n5564), .A2(n5568), .ZN(n6400) );
  NOR2_X1 U6461 ( .A1(n10525), .A2(n6321), .ZN(n10509) );
  NAND2_X1 U6462 ( .A1(n10509), .A2(n9019), .ZN(n5564) );
  NAND2_X1 U6463 ( .A1(n6336), .A2(n5845), .ZN(n6334) );
  NAND2_X1 U6464 ( .A1(n5589), .A2(n8870), .ZN(n7666) );
  INV_X1 U6465 ( .A(n10562), .ZN(n5586) );
  NOR2_X1 U6466 ( .A1(n10527), .A2(n10526), .ZN(n10525) );
  OAI21_X1 U6467 ( .B1(n9130), .B2(n9129), .A(n5269), .ZN(P1_U3242) );
  INV_X1 U6468 ( .A(n9005), .ZN(n5272) );
  NAND3_X1 U6469 ( .A1(n9001), .A2(n9000), .A3(n6401), .ZN(n5273) );
  AOI21_X1 U6470 ( .B1(n5605), .B2(n5218), .A(n9054), .ZN(n9016) );
  OAI21_X1 U6471 ( .B1(n5445), .B2(n6020), .A(n5219), .ZN(n5442) );
  NAND2_X1 U6472 ( .A1(n5443), .A2(n5441), .ZN(n6043) );
  NAND2_X1 U6473 ( .A1(n6055), .A2(n5790), .ZN(n6054) );
  OAI21_X1 U6474 ( .B1(n8989), .B2(n8990), .A(n5276), .ZN(n8993) );
  INV_X1 U6475 ( .A(n9686), .ZN(n5292) );
  OAI21_X1 U6476 ( .B1(n5292), .B2(n5154), .A(n5293), .ZN(n9653) );
  NAND2_X1 U6477 ( .A1(n5303), .A2(n5301), .ZN(n5463) );
  INV_X1 U6478 ( .A(n9197), .ZN(n9611) );
  INV_X1 U6479 ( .A(n5470), .ZN(n5313) );
  NAND2_X1 U6480 ( .A1(n5214), .A2(n8832), .ZN(n5316) );
  NAND2_X4 U6481 ( .A1(n6423), .A2(n5166), .ZN(n6624) );
  NAND2_X1 U6482 ( .A1(n6187), .A2(n5152), .ZN(n6203) );
  NAND3_X1 U6483 ( .A1(n6512), .A2(n5231), .A3(n7734), .ZN(n5325) );
  NAND2_X1 U6484 ( .A1(n8281), .A2(n5327), .ZN(n5326) );
  NOR2_X1 U6485 ( .A1(n9895), .A2(n5336), .ZN(n5335) );
  INV_X1 U6486 ( .A(n9897), .ZN(n5334) );
  NAND2_X1 U6487 ( .A1(n9853), .A2(n5341), .ZN(n5340) );
  NAND2_X1 U6488 ( .A1(n9853), .A2(n9854), .ZN(n9852) );
  NOR2_X2 U6489 ( .A1(n6295), .A2(n5344), .ZN(n6336) );
  OR2_X2 U6490 ( .A1(n6113), .A2(n5837), .ZN(n6295) );
  NAND3_X1 U6491 ( .A1(n5833), .A2(n5967), .A3(n5832), .ZN(n6113) );
  AOI21_X1 U6492 ( .B1(n8749), .B2(n5174), .A(n5347), .ZN(n5345) );
  NAND2_X1 U6493 ( .A1(n8750), .A2(n5174), .ZN(n5346) );
  NAND3_X1 U6494 ( .A1(n7232), .A2(n6686), .A3(n7133), .ZN(n6726) );
  AND3_X2 U6495 ( .A1(n7132), .A2(n6686), .A3(n5353), .ZN(n6734) );
  NAND2_X1 U6496 ( .A1(n5358), .A2(n5355), .ZN(n8484) );
  OAI211_X1 U6497 ( .C1(n5364), .C2(n5357), .A(n5356), .B(n8477), .ZN(n5355)
         );
  INV_X1 U6498 ( .A(n8480), .ZN(n5357) );
  NAND2_X1 U6499 ( .A1(n5359), .A2(n8695), .ZN(n5358) );
  NAND2_X1 U6500 ( .A1(n8471), .A2(n8730), .ZN(n5364) );
  NAND2_X1 U6501 ( .A1(n5365), .A2(n5366), .ZN(n8686) );
  NAND2_X1 U6502 ( .A1(n8624), .A2(n5368), .ZN(n5365) );
  AOI21_X1 U6503 ( .B1(n5371), .B2(n5369), .A(n5204), .ZN(n5368) );
  AND2_X1 U6504 ( .A1(n9582), .A2(n8622), .ZN(n5379) );
  INV_X2 U6505 ( .A(n7757), .ZN(n8037) );
  NAND3_X1 U6506 ( .A1(n6693), .A2(n5384), .A3(n6773), .ZN(n6698) );
  NAND3_X1 U6507 ( .A1(n6693), .A2(n6773), .A3(n5386), .ZN(n6700) );
  AND2_X1 U6508 ( .A1(n5745), .A2(n6694), .ZN(n5386) );
  AND2_X1 U6509 ( .A1(n5390), .A2(n5389), .ZN(n8494) );
  OAI21_X1 U6510 ( .B1(n8486), .B2(n5392), .A(n5391), .ZN(n5390) );
  NOR2_X2 U6511 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5911) );
  NAND2_X2 U6512 ( .A1(n8246), .A2(n5751), .ZN(n8270) );
  NAND2_X2 U6513 ( .A1(n8247), .A2(n8248), .ZN(n8246) );
  NOR2_X2 U6514 ( .A1(n6295), .A2(n5843), .ZN(n5864) );
  OAI211_X2 U6515 ( .C1(n8842), .C2(n6396), .A(n5394), .B(n5393), .ZN(n6869)
         );
  NAND2_X4 U6516 ( .A1(n6707), .A2(n8701), .ZN(n8853) );
  OR2_X1 U6517 ( .A1(n6707), .A2(n6931), .ZN(n5394) );
  NAND2_X4 U6518 ( .A1(n5138), .A2(n6406), .ZN(n6707) );
  OAI21_X2 U6519 ( .B1(n7026), .B2(n5397), .A(n5395), .ZN(n7347) );
  AND2_X2 U6520 ( .A1(n5400), .A2(n5399), .ZN(n10513) );
  NAND2_X1 U6521 ( .A1(n7662), .A2(n5406), .ZN(n5404) );
  NAND2_X1 U6522 ( .A1(n5412), .A2(n5413), .ZN(n6264) );
  INV_X1 U6523 ( .A(n5428), .ZN(n8251) );
  AND2_X1 U6524 ( .A1(n10514), .A2(n5430), .ZN(n10501) );
  NAND2_X1 U6525 ( .A1(n10514), .A2(n10517), .ZN(n10515) );
  NOR2_X2 U6526 ( .A1(n7386), .A2(n7744), .ZN(n7512) );
  NOR2_X2 U6527 ( .A1(n10630), .A2(n10725), .ZN(n10593) );
  NAND2_X1 U6528 ( .A1(n9653), .A2(n9660), .ZN(n5440) );
  NAND2_X1 U6529 ( .A1(n6005), .A2(n5444), .ZN(n5443) );
  INV_X1 U6530 ( .A(n5445), .ZN(n5444) );
  NAND2_X1 U6531 ( .A1(n5460), .A2(n5453), .ZN(n5452) );
  INV_X1 U6532 ( .A(n5175), .ZN(n5468) );
  NAND2_X1 U6533 ( .A1(n5471), .A2(n6054), .ZN(n8027) );
  NAND2_X1 U6534 ( .A1(n6057), .A2(n6056), .ZN(n5471) );
  OAI21_X1 U6535 ( .B1(n7241), .B2(P2_REG1_REG_3__SCAN_IN), .A(n5472), .ZN(
        n5473) );
  INV_X1 U6536 ( .A(n11028), .ZN(n5472) );
  NOR2_X1 U6537 ( .A1(n9472), .A2(n9471), .ZN(n9470) );
  NAND2_X1 U6538 ( .A1(n8401), .A2(n8362), .ZN(n5478) );
  NAND2_X1 U6539 ( .A1(n8353), .A2(n5489), .ZN(n5487) );
  XNOR2_X1 U6540 ( .A(n7244), .B(n7535), .ZN(n11043) );
  NAND2_X1 U6541 ( .A1(n5501), .A2(n5504), .ZN(n7207) );
  NAND2_X1 U6542 ( .A1(n5502), .A2(n5503), .ZN(n5501) );
  INV_X1 U6543 ( .A(n11008), .ZN(n5502) );
  NAND2_X1 U6544 ( .A1(n8375), .A2(n5505), .ZN(n5507) );
  NAND2_X1 U6545 ( .A1(n5510), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5508) );
  INV_X1 U6546 ( .A(n8375), .ZN(n5510) );
  XNOR2_X1 U6547 ( .A(n5506), .B(n5513), .ZN(n8378) );
  NAND3_X1 U6548 ( .A1(n5509), .A2(n5508), .A3(n5507), .ZN(n5506) );
  NAND2_X1 U6549 ( .A1(n7975), .A2(n7977), .ZN(n5517) );
  NAND2_X1 U6550 ( .A1(n8197), .A2(n5523), .ZN(n5521) );
  NAND3_X1 U6551 ( .A1(n5526), .A2(n5525), .A3(n5524), .ZN(n9394) );
  NAND2_X1 U6552 ( .A1(n8320), .A2(n5142), .ZN(n5526) );
  INV_X1 U6553 ( .A(n5527), .ZN(n8365) );
  AOI22_X1 U6554 ( .A1(n9537), .A2(n9536), .B1(n9362), .B2(n9541), .ZN(n9527)
         );
  NAND2_X1 U6555 ( .A1(n5773), .A2(n5774), .ZN(n5602) );
  NAND2_X1 U6556 ( .A1(n5624), .A2(n5627), .ZN(n6088) );
  NAND2_X1 U6557 ( .A1(n5956), .A2(n5770), .ZN(n5974) );
  AOI21_X1 U6558 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7243), .A(n11027), .ZN(
        n7244) );
  NOR2_X1 U6559 ( .A1(n8216), .A2(n11077), .ZN(n8219) );
  NOR2_X1 U6560 ( .A1(n10981), .A2(n10980), .ZN(n10983) );
  NOR2_X1 U6561 ( .A1(n8014), .A2(n11078), .ZN(n11077) );
  NOR2_X1 U6562 ( .A1(n10983), .A2(n7236), .ZN(n10999) );
  OAI21_X1 U6563 ( .B1(n7234), .B2(n7233), .A(n7235), .ZN(n10981) );
  NOR2_X1 U6564 ( .A1(n10999), .A2(n10998), .ZN(n10997) );
  NAND2_X1 U6565 ( .A1(n7399), .A2(n5193), .ZN(n5537) );
  NAND3_X1 U6566 ( .A1(n6481), .A2(n6482), .A3(n5145), .ZN(n5536) );
  NAND2_X1 U6567 ( .A1(n7863), .A2(n6505), .ZN(n6511) );
  NAND2_X1 U6568 ( .A1(n7863), .A2(n5550), .ZN(n7735) );
  NAND2_X1 U6569 ( .A1(n6837), .A2(n5553), .ZN(n6442) );
  NAND2_X1 U6570 ( .A1(n6433), .A2(n6645), .ZN(n5553) );
  NAND3_X1 U6571 ( .A1(n6837), .A2(n5553), .A3(n6438), .ZN(n6895) );
  NAND2_X1 U6572 ( .A1(n8822), .A2(n5558), .ZN(n5554) );
  NAND2_X1 U6573 ( .A1(n5554), .A2(n5555), .ZN(n8249) );
  NAND2_X1 U6574 ( .A1(n10525), .A2(n5568), .ZN(n5563) );
  INV_X1 U6575 ( .A(n8904), .ZN(n5579) );
  NAND3_X1 U6576 ( .A1(n5571), .A2(n5573), .A3(n8910), .ZN(n8908) );
  NAND2_X1 U6577 ( .A1(n9063), .A2(n5572), .ZN(n5571) );
  AND2_X1 U6578 ( .A1(n8904), .A2(n5575), .ZN(n5572) );
  NAND3_X1 U6579 ( .A1(n9063), .A2(n5575), .A3(n5577), .ZN(n5573) );
  AOI21_X1 U6580 ( .B1(n5586), .B2(n5582), .A(n5580), .ZN(n10527) );
  NAND2_X1 U6581 ( .A1(n10562), .A2(n8979), .ZN(n10549) );
  NAND2_X1 U6582 ( .A1(n7664), .A2(n8931), .ZN(n5589) );
  NAND2_X1 U6583 ( .A1(n6410), .A2(n10746), .ZN(n5595) );
  NAND2_X1 U6584 ( .A1(n5590), .A2(n5592), .ZN(n6418) );
  NAND2_X2 U6585 ( .A1(n8806), .A2(n5591), .ZN(n5593) );
  AOI21_X2 U6586 ( .B1(n5594), .B2(n10713), .A(n11180), .ZN(n5592) );
  AND2_X1 U6587 ( .A1(n5864), .A2(n10321), .ZN(n5865) );
  NAND2_X1 U6588 ( .A1(n5864), .A2(n5597), .ZN(n5868) );
  XNOR2_X2 U6589 ( .A(n6434), .B(n5941), .ZN(n6880) );
  NAND2_X1 U6590 ( .A1(n5599), .A2(n6282), .ZN(n6267) );
  INV_X1 U6591 ( .A(n6391), .ZN(n5601) );
  NAND2_X1 U6592 ( .A1(n5976), .A2(n5774), .ZN(n5990) );
  NAND2_X1 U6593 ( .A1(n5973), .A2(n5974), .ZN(n5976) );
  INV_X1 U6594 ( .A(n5774), .ZN(n5603) );
  INV_X1 U6595 ( .A(n5773), .ZN(n5973) );
  OR2_X1 U6596 ( .A1(n6171), .A2(n5614), .ZN(n5610) );
  NAND2_X1 U6597 ( .A1(n6171), .A2(n5608), .ZN(n5607) );
  NAND2_X1 U6598 ( .A1(n6171), .A2(n6170), .ZN(n5616) );
  OAI21_X1 U6599 ( .B1(n6054), .B2(n5621), .A(n5618), .ZN(n6108) );
  NAND2_X1 U6600 ( .A1(n6054), .A2(n5625), .ZN(n5624) );
  NAND2_X1 U6601 ( .A1(n6054), .A2(n5791), .ZN(n6082) );
  NAND2_X1 U6602 ( .A1(n5633), .A2(n5631), .ZN(n6142) );
  NAND2_X1 U6603 ( .A1(n6110), .A2(n5797), .ZN(n6126) );
  NOR2_X1 U6604 ( .A1(n6125), .A2(n5635), .ZN(n5634) );
  INV_X1 U6605 ( .A(n5797), .ZN(n5635) );
  INV_X1 U6606 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5757) );
  INV_X1 U6607 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5639) );
  INV_X1 U6608 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5638) );
  NAND3_X1 U6609 ( .A1(n5757), .A2(n5639), .A3(n5638), .ZN(n5637) );
  NAND2_X1 U6610 ( .A1(n5642), .A2(n5641), .ZN(n5644) );
  INV_X1 U6611 ( .A(n9356), .ZN(n5642) );
  NAND3_X1 U6612 ( .A1(n5644), .A2(n9172), .A3(n5643), .ZN(P2_U3160) );
  NAND3_X1 U6613 ( .A1(n5155), .A2(n9356), .A3(n9370), .ZN(n5643) );
  NAND2_X1 U6614 ( .A1(n9168), .A2(n5649), .ZN(n5647) );
  NAND2_X1 U6615 ( .A1(n9356), .A2(n9166), .ZN(n9225) );
  NAND2_X1 U6616 ( .A1(n9262), .A2(n5654), .ZN(n5652) );
  NAND2_X1 U6617 ( .A1(n5652), .A2(n5207), .ZN(n9303) );
  NAND2_X1 U6618 ( .A1(n7151), .A2(n5660), .ZN(n5658) );
  NAND2_X1 U6619 ( .A1(n7151), .A2(n7145), .ZN(n5659) );
  NAND2_X1 U6620 ( .A1(n5661), .A2(n5215), .ZN(n9291) );
  OAI21_X2 U6621 ( .B1(n8258), .B2(n5666), .A(n5663), .ZN(n9132) );
  NAND2_X1 U6622 ( .A1(n5672), .A2(n5671), .ZN(n5673) );
  NAND2_X1 U6623 ( .A1(n7705), .A2(n7530), .ZN(n5671) );
  INV_X1 U6624 ( .A(n5673), .ZN(n7581) );
  NAND2_X1 U6625 ( .A1(n5675), .A2(n5674), .ZN(n9310) );
  NAND2_X1 U6626 ( .A1(n5682), .A2(n5681), .ZN(n7662) );
  NAND2_X1 U6627 ( .A1(n7508), .A2(n10349), .ZN(n5681) );
  NAND2_X2 U6628 ( .A1(n7370), .A2(n6073), .ZN(n7508) );
  NAND3_X1 U6629 ( .A1(n5687), .A2(n10605), .A3(n5688), .ZN(n5686) );
  INV_X1 U6630 ( .A(n7899), .ZN(n5708) );
  INV_X1 U6631 ( .A(n5711), .ZN(n5710) );
  NAND2_X1 U6632 ( .A1(n10513), .A2(n10526), .ZN(n10512) );
  INV_X1 U6633 ( .A(n8122), .ZN(n5717) );
  NAND2_X1 U6634 ( .A1(n9623), .A2(n5726), .ZN(n5725) );
  OAI21_X1 U6635 ( .B1(n7942), .B2(n5737), .A(n5735), .ZN(n8034) );
  NAND2_X1 U6636 ( .A1(n8755), .A2(n5740), .ZN(n9682) );
  NAND2_X1 U6637 ( .A1(n9682), .A2(n5217), .ZN(n8760) );
  AND2_X1 U6638 ( .A1(n6696), .A2(n5742), .ZN(n7105) );
  NAND2_X1 U6639 ( .A1(n6696), .A2(n5213), .ZN(n9797) );
  NAND2_X1 U6640 ( .A1(n6696), .A2(n6695), .ZN(n7092) );
  NAND3_X1 U6641 ( .A1(n6773), .A2(n6693), .A3(n6688), .ZN(n7148) );
  NAND2_X1 U6642 ( .A1(n9061), .A2(n9057), .ZN(n8858) );
  MUX2_X1 U6643 ( .A(n8461), .B(n8460), .S(n8464), .Z(n8470) );
  NAND2_X1 U6644 ( .A1(n8719), .A2(n8718), .ZN(n8749) );
  XNOR2_X1 U6645 ( .A(n8406), .B(n8407), .ZN(n6392) );
  NAND2_X1 U6646 ( .A1(n6392), .A2(SI_29_), .ZN(n8410) );
  OR2_X1 U6647 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  OR2_X1 U6648 ( .A1(n6111), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6128) );
  CLKBUF_X1 U6649 ( .A(n6113), .Z(n6111) );
  NAND2_X1 U6650 ( .A1(n5771), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5758) );
  CLKBUF_X1 U6651 ( .A(n6406), .Z(n8349) );
  INV_X1 U6652 ( .A(n9235), .ZN(n9368) );
  XNOR2_X1 U6653 ( .A(n7096), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U6654 ( .A1(n9797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7096) );
  CLKBUF_X1 U6655 ( .A(n7942), .Z(n8081) );
  INV_X1 U6656 ( .A(n7395), .ZN(n7396) );
  NAND2_X1 U6657 ( .A1(n7395), .A2(n7143), .ZN(n7144) );
  NAND2_X1 U6658 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  XNOR2_X1 U6659 ( .A(n7094), .B(n7093), .ZN(n7098) );
  OR2_X1 U6660 ( .A1(n7132), .A2(n7131), .ZN(n7134) );
  NOR2_X1 U6661 ( .A1(n7308), .A2(n5753), .ZN(n7491) );
  NAND2_X1 U6662 ( .A1(n7287), .A2(n7283), .ZN(n7282) );
  INV_X1 U6663 ( .A(n7097), .ZN(n7099) );
  NAND2_X1 U6664 ( .A1(n7800), .A2(n7799), .ZN(n7942) );
  OR2_X1 U6665 ( .A1(n7299), .A2(n7189), .ZN(n7303) );
  OR2_X1 U6666 ( .A1(n7110), .A2(n7131), .ZN(n7112) );
  NAND2_X1 U6667 ( .A1(n7104), .A2(n7109), .ZN(n7158) );
  NAND2_X1 U6668 ( .A1(n7104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U6669 ( .A1(n7092), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U6670 ( .A1(n7830), .A2(n7829), .ZN(n5747) );
  INV_X1 U6671 ( .A(n10593), .ZN(n10608) );
  AND4_X1 U6672 ( .A1(n6844), .A2(n7363), .A3(n7138), .A4(n7146), .ZN(n5748)
         );
  AND2_X1 U6673 ( .A1(n9184), .A2(n9513), .ZN(n5749) );
  INV_X1 U6674 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8193) );
  OR2_X1 U6675 ( .A1(n9846), .A2(n9857), .ZN(n5750) );
  OR2_X1 U6676 ( .A1(n9862), .A2(n10740), .ZN(n5751) );
  AND2_X1 U6677 ( .A1(n6444), .A2(n6426), .ZN(n5752) );
  NAND2_X1 U6678 ( .A1(n11185), .A2(n11127), .ZN(n10806) );
  INV_X1 U6679 ( .A(n10806), .ZN(n6368) );
  XNOR2_X1 U6680 ( .A(n7562), .B(n7528), .ZN(n7521) );
  AND2_X1 U6681 ( .A1(n10464), .A2(n8088), .ZN(n9011) );
  NOR2_X1 U6682 ( .A1(n5429), .A2(n10739), .ZN(n6414) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5759) );
  OR2_X1 U6684 ( .A1(n10968), .A2(n7159), .ZN(n11081) );
  INV_X1 U6685 ( .A(n10579), .ZN(n10793) );
  AND2_X1 U6686 ( .A1(n7306), .A2(n7305), .ZN(n5753) );
  INV_X1 U6687 ( .A(n10514), .ZN(n10537) );
  NOR2_X1 U6688 ( .A1(n9366), .A2(n9367), .ZN(n5754) );
  AND2_X2 U6689 ( .A1(n7684), .A2(n11105), .ZN(n11124) );
  AND2_X1 U6690 ( .A1(n9671), .A2(n9658), .ZN(n5755) );
  NAND2_X1 U6691 ( .A1(n9565), .A2(n9582), .ZN(n5756) );
  NAND2_X1 U6692 ( .A1(n8988), .A2(n9002), .ZN(n8996) );
  INV_X1 U6693 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8370) );
  INV_X1 U6694 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6157) );
  INV_X1 U6695 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7106) );
  AND2_X1 U6696 ( .A1(n6381), .A2(n6380), .ZN(n6382) );
  INV_X1 U6697 ( .A(n7238), .ZN(n7239) );
  NOR2_X1 U6698 ( .A1(n8028), .A2(n7945), .ZN(n8212) );
  NAND2_X1 U6699 ( .A1(n8767), .A2(n5756), .ZN(n8769) );
  NAND2_X1 U6700 ( .A1(n6637), .A2(n7011), .ZN(n6436) );
  INV_X1 U6701 ( .A(n9008), .ZN(n9009) );
  INV_X1 U6702 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6066) );
  INV_X1 U6703 ( .A(n8630), .ZN(n8416) );
  INV_X1 U6704 ( .A(n8603), .ZN(n8414) );
  NOR2_X1 U6705 ( .A1(n10993), .A2(n7202), .ZN(n7203) );
  INV_X1 U6706 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U6707 ( .A1(n8028), .A2(n8193), .ZN(n8194) );
  AND2_X1 U6708 ( .A1(n8417), .A2(n10010), .ZN(n8643) );
  NOR2_X1 U6709 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n8413), .ZN(n8570) );
  INV_X1 U6710 ( .A(n6233), .ZN(n5858) );
  INV_X1 U6711 ( .A(n6075), .ZN(n5853) );
  INV_X1 U6712 ( .A(n6243), .ZN(n5859) );
  OR2_X1 U6713 ( .A1(n6257), .A2(n9866), .ZN(n5896) );
  OR2_X1 U6714 ( .A1(n6067), .A2(n6066), .ZN(n6075) );
  NOR2_X1 U6715 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5831) );
  NAND2_X1 U6716 ( .A1(n8416), .A2(n8415), .ZN(n8644) );
  OR2_X1 U6717 ( .A1(n9243), .A2(n9578), .ZN(n9157) );
  INV_X1 U6718 ( .A(n9312), .ZN(n9151) );
  XNOR2_X1 U6719 ( .A(n7528), .B(n7428), .ZN(n7310) );
  OR2_X1 U6720 ( .A1(n8615), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8630) );
  AND2_X1 U6721 ( .A1(n7758), .A2(n10196), .ZN(n7836) );
  INV_X1 U6722 ( .A(n11081), .ZN(n8377) );
  OR2_X1 U6723 ( .A1(n9732), .A2(n9593), .ZN(n9199) );
  INV_X1 U6724 ( .A(n7723), .ZN(n7787) );
  INV_X1 U6725 ( .A(n7274), .ZN(n7176) );
  INV_X1 U6726 ( .A(n9672), .ZN(n9667) );
  NAND2_X1 U6727 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6736) );
  INV_X1 U6728 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6163) );
  INV_X1 U6729 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U6730 ( .A1(n5859), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U6731 ( .A1(n5860), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5889) );
  OR2_X1 U6732 ( .A1(n6255), .A2(n9811), .ZN(n6257) );
  NAND2_X1 U6733 ( .A1(n5855), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6164) );
  OR2_X1 U6734 ( .A1(n10595), .A2(n10709), .ZN(n6250) );
  NAND2_X1 U6735 ( .A1(n5857), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6222) );
  INV_X1 U6736 ( .A(n6707), .ZN(n6205) );
  INV_X1 U6737 ( .A(SI_24_), .ZN(n10143) );
  INV_X1 U6738 ( .A(SI_20_), .ZN(n9956) );
  AND2_X1 U6739 ( .A1(n8828), .A2(n6763), .ZN(n6702) );
  NAND2_X1 U6740 ( .A1(n9147), .A2(n9613), .ZN(n9148) );
  NAND2_X1 U6741 ( .A1(n7521), .A2(n9393), .ZN(n7522) );
  AND2_X1 U6742 ( .A1(n9775), .A2(n8464), .ZN(n7319) );
  XNOR2_X1 U6743 ( .A(n7158), .B(n7250), .ZN(n7336) );
  INV_X1 U6744 ( .A(n9373), .ZN(n9361) );
  OR2_X1 U6745 ( .A1(n8037), .A2(n9213), .ZN(n8715) );
  AND2_X1 U6746 ( .A1(n8379), .A2(n9256), .ZN(n8380) );
  AND2_X1 U6747 ( .A1(n8653), .A2(n8645), .ZN(n9555) );
  INV_X1 U6748 ( .A(n9387), .ZN(n8181) );
  INV_X1 U6749 ( .A(n7299), .ZN(n7693) );
  INV_X1 U6750 ( .A(n9613), .ZN(n9757) );
  INV_X1 U6751 ( .A(n9384), .ZN(n9134) );
  INV_X1 U6752 ( .A(n9388), .ZN(n8078) );
  INV_X1 U6753 ( .A(n9775), .ZN(n9754) );
  INV_X1 U6754 ( .A(n9643), .ZN(n9689) );
  NAND2_X1 U6755 ( .A1(n6767), .A2(n6766), .ZN(n7678) );
  OR2_X1 U6756 ( .A1(n6951), .A2(n7131), .ZN(n6952) );
  OR2_X1 U6757 ( .A1(n6099), .A2(n6098), .ZN(n6118) );
  OR2_X1 U6758 ( .A1(n6164), .A2(n6163), .ZN(n6177) );
  NAND2_X1 U6759 ( .A1(n5856), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U6760 ( .A1(n5852), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6067) );
  OR2_X1 U6761 ( .A1(n6118), .A2(n6117), .ZN(n6134) );
  INV_X1 U6762 ( .A(n9932), .ZN(n9878) );
  OR2_X1 U6763 ( .A1(n6193), .A2(n6192), .ZN(n6212) );
  INV_X1 U6764 ( .A(n9917), .ZN(n9930) );
  OR2_X1 U6765 ( .A1(n10518), .A2(n6258), .ZN(n5878) );
  INV_X1 U6766 ( .A(n5139), .ZN(n6917) );
  INV_X1 U6767 ( .A(n9006), .ZN(n6401) );
  AND2_X1 U6768 ( .A1(n6278), .A2(n6277), .ZN(n10685) );
  OAI21_X1 U6769 ( .B1(n10693), .B2(n10789), .A(n6264), .ZN(n10535) );
  AND4_X1 U6770 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n9857)
         );
  AND2_X1 U6771 ( .A1(n10475), .A2(n10474), .ZN(n10671) );
  AND2_X1 U6772 ( .A1(n6917), .A2(n9040), .ZN(n11156) );
  AND2_X1 U6773 ( .A1(n8088), .A2(n9054), .ZN(n6655) );
  NAND2_X1 U6774 ( .A1(n7382), .A2(n8857), .ZN(n7381) );
  INV_X1 U6775 ( .A(n10672), .ZN(n10655) );
  NAND2_X1 U6776 ( .A1(n7173), .A2(n6702), .ZN(n7296) );
  AND2_X1 U6777 ( .A1(n7337), .A2(n7336), .ZN(n9373) );
  INV_X1 U6778 ( .A(n9375), .ZN(n9359) );
  INV_X1 U6779 ( .A(n9348), .ZN(n9377) );
  AND4_X1 U6780 ( .A1(n8715), .A2(n8425), .A3(n8424), .A4(n8423), .ZN(n8717)
         );
  AND4_X1 U6781 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n9337)
         );
  AND4_X1 U6782 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n9767)
         );
  NAND2_X1 U6783 ( .A1(n7254), .A2(n7253), .ZN(n11033) );
  INV_X1 U6784 ( .A(n11040), .ZN(n11076) );
  OR2_X1 U6785 ( .A1(n9775), .A2(n7693), .ZN(n11103) );
  INV_X1 U6786 ( .A(n9698), .ZN(n11120) );
  AOI21_X1 U6787 ( .B1(n7677), .B2(n7679), .A(n7176), .ZN(n7193) );
  NOR2_X1 U6788 ( .A1(n7299), .A2(n8800), .ZN(n9704) );
  OR2_X1 U6789 ( .A1(n9203), .A2(n9704), .ZN(n9779) );
  INV_X1 U6790 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6844) );
  INV_X1 U6791 ( .A(n9912), .ZN(n9928) );
  AND2_X1 U6792 ( .A1(n6671), .A2(n5139), .ZN(n9932) );
  INV_X1 U6793 ( .A(n8847), .ZN(n6405) );
  AND2_X1 U6794 ( .A1(n6249), .A2(n6248), .ZN(n9812) );
  AND4_X1 U6795 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n10764)
         );
  OR2_X1 U6796 ( .A1(n6755), .A2(n6917), .ZN(n10374) );
  OR2_X1 U6797 ( .A1(n6755), .A2(n6752), .ZN(n10956) );
  INV_X1 U6798 ( .A(n10422), .ZN(n10904) );
  INV_X1 U6799 ( .A(n10374), .ZN(n10962) );
  NAND2_X1 U6800 ( .A1(n9027), .A2(n8991), .ZN(n10536) );
  INV_X1 U6801 ( .A(n10576), .ZN(n10664) );
  NAND2_X1 U6802 ( .A1(n9015), .A2(n6323), .ZN(n10746) );
  AND2_X1 U6803 ( .A1(n6707), .A2(n7113), .ZN(n8854) );
  AND2_X1 U6804 ( .A1(n6420), .A2(n6655), .ZN(n11127) );
  OAI21_X1 U6805 ( .B1(n10812), .B2(P1_D_REG_0__SCAN_IN), .A(n10815), .ZN(
        n6955) );
  INV_X1 U6806 ( .A(n6365), .ZN(n10812) );
  AND2_X1 U6807 ( .A1(n6009), .A2(n6023), .ZN(n6852) );
  INV_X1 U6808 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10276) );
  OR2_X1 U6809 ( .A1(n7296), .A2(n8097), .ZN(n7252) );
  OR2_X1 U6810 ( .A1(n7321), .A2(n7320), .ZN(n9330) );
  INV_X1 U6811 ( .A(n9327), .ZN(n9380) );
  INV_X1 U6812 ( .A(n9531), .ZN(n9716) );
  INV_X1 U6813 ( .A(n9767), .ZN(n9645) );
  OR2_X1 U6814 ( .A1(P2_U3150), .A2(n7256), .ZN(n11040) );
  INV_X1 U6815 ( .A(n11033), .ZN(n11096) );
  OR2_X1 U6816 ( .A1(n10968), .A2(n7250), .ZN(n11090) );
  NAND2_X1 U6817 ( .A1(n9692), .A2(n7694), .ZN(n9698) );
  OR2_X1 U6818 ( .A1(n9751), .A2(n9750), .ZN(n9795) );
  AND2_X1 U6819 ( .A1(n7278), .A2(n7277), .ZN(n11192) );
  INV_X1 U6820 ( .A(n7338), .ZN(n7318) );
  INV_X1 U6821 ( .A(n8746), .ZN(n7732) );
  INV_X1 U6822 ( .A(n8028), .ZN(n8211) );
  NOR2_X1 U6823 ( .A1(n6685), .A2(n6684), .ZN(n6705) );
  AND2_X1 U6824 ( .A1(n6659), .A2(n10659), .ZN(n9936) );
  INV_X1 U6825 ( .A(n10676), .ZN(n9938) );
  NAND2_X1 U6826 ( .A1(n5894), .A2(n5893), .ZN(n10520) );
  INV_X1 U6827 ( .A(n10644), .ZN(n10344) );
  NAND2_X1 U6828 ( .A1(n6716), .A2(n6715), .ZN(n10967) );
  INV_X1 U6829 ( .A(n10580), .ZN(n10658) );
  INV_X1 U6830 ( .A(n10651), .ZN(n10638) );
  NOR2_X1 U6831 ( .A1(n6414), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U6832 ( .A1(n11181), .A2(n11127), .ZN(n10739) );
  INV_X1 U6833 ( .A(n11181), .ZN(n11180) );
  INV_X1 U6834 ( .A(n10472), .ZN(n10775) );
  NAND2_X1 U6835 ( .A1(n6371), .A2(n6955), .ZN(n11182) );
  INV_X2 U6836 ( .A(n11182), .ZN(n11185) );
  INV_X1 U6837 ( .A(n10826), .ZN(n10827) );
  NOR2_X2 U6838 ( .A1(n7252), .A2(P2_U3151), .ZN(P2_U3893) );
  INV_X1 U6839 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U6840 ( .A1(n5760), .A2(SI_1_), .ZN(n5764) );
  OAI21_X1 U6841 ( .B1(n5760), .B2(SI_1_), .A(n5764), .ZN(n5934) );
  INV_X1 U6842 ( .A(n5934), .ZN(n5763) );
  INV_X1 U6843 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5924) );
  INV_X1 U6844 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7123) );
  INV_X1 U6845 ( .A(SI_0_), .ZN(n5923) );
  NOR2_X1 U6846 ( .A1(n5762), .A2(n5923), .ZN(n5932) );
  NAND2_X1 U6847 ( .A1(n5763), .A2(n5932), .ZN(n5936) );
  NAND2_X1 U6848 ( .A1(n5936), .A2(n5764), .ZN(n5912) );
  MUX2_X1 U6849 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5771), .Z(n5765) );
  NAND2_X1 U6850 ( .A1(n5765), .A2(SI_2_), .ZN(n5767) );
  OAI21_X1 U6851 ( .B1(n5765), .B2(SI_2_), .A(n5767), .ZN(n5913) );
  INV_X1 U6852 ( .A(n5913), .ZN(n5766) );
  NAND2_X1 U6853 ( .A1(n5912), .A2(n5766), .ZN(n5915) );
  NAND2_X1 U6854 ( .A1(n5915), .A2(n5767), .ZN(n5954) );
  MUX2_X1 U6855 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n5771), .Z(n5768) );
  NAND2_X1 U6856 ( .A1(n5768), .A2(SI_3_), .ZN(n5770) );
  OAI21_X1 U6857 ( .B1(n5768), .B2(SI_3_), .A(n5770), .ZN(n5769) );
  INV_X1 U6858 ( .A(n5769), .ZN(n5953) );
  NAND2_X1 U6859 ( .A1(n5954), .A2(n5953), .ZN(n5956) );
  INV_X4 U6860 ( .A(n7113), .ZN(n8701) );
  MUX2_X1 U6861 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8701), .Z(n5772) );
  OAI21_X1 U6862 ( .B1(n5772), .B2(SI_4_), .A(n5774), .ZN(n5773) );
  MUX2_X1 U6863 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n5823), .Z(n5775) );
  NAND2_X1 U6864 ( .A1(n5775), .A2(SI_5_), .ZN(n5777) );
  OAI21_X1 U6865 ( .B1(n5775), .B2(SI_5_), .A(n5777), .ZN(n5776) );
  INV_X1 U6866 ( .A(n5776), .ZN(n5989) );
  NAND2_X1 U6867 ( .A1(n5992), .A2(n5777), .ZN(n6003) );
  MUX2_X1 U6868 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n5823), .Z(n5778) );
  NAND2_X1 U6869 ( .A1(n5778), .A2(SI_6_), .ZN(n5780) );
  OAI21_X1 U6870 ( .B1(n5778), .B2(SI_6_), .A(n5780), .ZN(n5779) );
  INV_X1 U6871 ( .A(n5779), .ZN(n6002) );
  NAND2_X1 U6872 ( .A1(n5781), .A2(SI_7_), .ZN(n5783) );
  OAI21_X1 U6873 ( .B1(n5781), .B2(SI_7_), .A(n5783), .ZN(n5782) );
  INV_X1 U6874 ( .A(n5782), .ZN(n6020) );
  MUX2_X1 U6875 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n5823), .Z(n5784) );
  XNOR2_X1 U6876 ( .A(n5784), .B(SI_8_), .ZN(n6027) );
  INV_X1 U6877 ( .A(n5784), .ZN(n5786) );
  INV_X1 U6878 ( .A(SI_8_), .ZN(n5785) );
  MUX2_X1 U6879 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n5823), .Z(n5787) );
  XNOR2_X1 U6880 ( .A(n5787), .B(n10170), .ZN(n6042) );
  NOR2_X1 U6881 ( .A1(n5787), .A2(SI_9_), .ZN(n5788) );
  MUX2_X1 U6882 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n5823), .Z(n5789) );
  NAND2_X1 U6883 ( .A1(n5789), .A2(SI_10_), .ZN(n5791) );
  OAI21_X1 U6884 ( .B1(n5789), .B2(SI_10_), .A(n5791), .ZN(n6056) );
  INV_X1 U6885 ( .A(n6056), .ZN(n5790) );
  MUX2_X1 U6886 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n5823), .Z(n5792) );
  XNOR2_X1 U6887 ( .A(n5792), .B(SI_11_), .ZN(n6081) );
  MUX2_X1 U6888 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n5823), .Z(n5793) );
  NAND2_X1 U6889 ( .A1(n5793), .A2(SI_12_), .ZN(n5794) );
  OAI21_X1 U6890 ( .B1(n5793), .B2(SI_12_), .A(n5794), .ZN(n6087) );
  MUX2_X1 U6891 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n5823), .Z(n5795) );
  NAND2_X1 U6892 ( .A1(n5795), .A2(SI_13_), .ZN(n5797) );
  OAI21_X1 U6893 ( .B1(n5795), .B2(SI_13_), .A(n5797), .ZN(n5796) );
  INV_X1 U6894 ( .A(n5796), .ZN(n6107) );
  NAND2_X1 U6895 ( .A1(n6108), .A2(n6107), .ZN(n6110) );
  MUX2_X1 U6896 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n5823), .Z(n5798) );
  XNOR2_X1 U6897 ( .A(n5798), .B(SI_14_), .ZN(n6125) );
  MUX2_X1 U6898 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n5823), .Z(n5799) );
  NAND2_X1 U6899 ( .A1(n5799), .A2(SI_15_), .ZN(n5800) );
  OAI21_X1 U6900 ( .B1(n5799), .B2(SI_15_), .A(n5800), .ZN(n6140) );
  MUX2_X1 U6901 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n5823), .Z(n5801) );
  XNOR2_X1 U6902 ( .A(n5801), .B(SI_16_), .ZN(n6154) );
  INV_X1 U6903 ( .A(n5801), .ZN(n5803) );
  INV_X1 U6904 ( .A(SI_16_), .ZN(n5802) );
  NAND2_X1 U6905 ( .A1(n5803), .A2(n5802), .ZN(n5804) );
  OAI21_X2 U6906 ( .B1(n6155), .B2(n6154), .A(n5804), .ZN(n6171) );
  MUX2_X1 U6907 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n5823), .Z(n5805) );
  MUX2_X1 U6908 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n5823), .Z(n5806) );
  NAND2_X1 U6909 ( .A1(n5806), .A2(SI_18_), .ZN(n5807) );
  OAI21_X1 U6910 ( .B1(n5806), .B2(SI_18_), .A(n5807), .ZN(n6183) );
  MUX2_X1 U6911 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n5823), .Z(n5808) );
  XNOR2_X1 U6912 ( .A(n5808), .B(SI_19_), .ZN(n6201) );
  INV_X1 U6913 ( .A(n5808), .ZN(n5809) );
  MUX2_X1 U6914 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n5823), .Z(n5810) );
  NOR2_X1 U6915 ( .A1(n5810), .A2(SI_20_), .ZN(n5811) );
  MUX2_X1 U6916 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n5823), .Z(n5812) );
  NAND2_X1 U6917 ( .A1(n5812), .A2(SI_21_), .ZN(n5814) );
  OAI21_X1 U6918 ( .B1(n5812), .B2(SI_21_), .A(n5814), .ZN(n5813) );
  INV_X1 U6919 ( .A(n5813), .ZN(n6228) );
  NAND2_X1 U6920 ( .A1(n6227), .A2(n6228), .ZN(n5815) );
  NAND2_X1 U6921 ( .A1(n5815), .A2(n5814), .ZN(n5817) );
  MUX2_X1 U6922 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n5823), .Z(n5816) );
  INV_X1 U6923 ( .A(SI_22_), .ZN(n10150) );
  MUX2_X1 U6924 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8701), .Z(n5819) );
  XNOR2_X1 U6925 ( .A(n5819), .B(n10142), .ZN(n6251) );
  NAND2_X1 U6926 ( .A1(n6252), .A2(n6251), .ZN(n5822) );
  INV_X1 U6927 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U6928 ( .A1(n5820), .A2(n10142), .ZN(n5821) );
  NAND2_X1 U6929 ( .A1(n5822), .A2(n5821), .ZN(n5903) );
  MUX2_X1 U6930 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8701), .Z(n5825) );
  XNOR2_X1 U6931 ( .A(n5825), .B(n10143), .ZN(n5902) );
  NAND2_X1 U6932 ( .A1(n5903), .A2(n5902), .ZN(n5880) );
  MUX2_X1 U6933 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n5823), .Z(n5824) );
  NAND2_X1 U6934 ( .A1(n5824), .A2(SI_25_), .ZN(n5829) );
  OAI21_X1 U6935 ( .B1(n5824), .B2(SI_25_), .A(n5829), .ZN(n5881) );
  INV_X1 U6936 ( .A(n5881), .ZN(n5827) );
  INV_X1 U6937 ( .A(n5825), .ZN(n5826) );
  NAND2_X1 U6938 ( .A1(n5826), .A2(n10143), .ZN(n5879) );
  MUX2_X1 U6939 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n8701), .Z(n6265) );
  XNOR2_X1 U6940 ( .A(n6265), .B(SI_26_), .ZN(n6384) );
  XNOR2_X1 U6941 ( .A(n6391), .B(n6384), .ZN(n8662) );
  AND4_X2 U6943 ( .A1(n5830), .A2(n10288), .A3(n10283), .A4(n10079), .ZN(n5833) );
  AND2_X2 U6944 ( .A1(n5911), .A2(n5831), .ZN(n5967) );
  INV_X2 U6945 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10284) );
  INV_X2 U6946 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6058) );
  NOR2_X1 U6947 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5836) );
  NOR2_X1 U6948 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5835) );
  NOR2_X1 U6949 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5834) );
  NAND4_X1 U6950 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n10096), .ZN(n5837)
         );
  AND2_X1 U6951 ( .A1(n10316), .A2(n5845), .ZN(n5842) );
  NAND2_X1 U6952 ( .A1(n10311), .A2(n10312), .ZN(n6342) );
  NAND2_X1 U6953 ( .A1(n5842), .A2(n5198), .ZN(n5843) );
  XNOR2_X2 U6954 ( .A(n5846), .B(n10316), .ZN(n6406) );
  NAND2_X1 U6955 ( .A1(n8662), .A2(n8854), .ZN(n5848) );
  INV_X1 U6956 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8306) );
  OR2_X1 U6957 ( .A1(n8853), .A2(n8306), .ZN(n5847) );
  INV_X1 U6958 ( .A(n10688), .ZN(n10517) );
  NAND2_X1 U6959 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5982) );
  INV_X1 U6960 ( .A(n5982), .ZN(n5849) );
  NAND2_X1 U6961 ( .A1(n5849), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5996) );
  INV_X1 U6962 ( .A(n5996), .ZN(n5850) );
  NAND2_X1 U6963 ( .A1(n5850), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6014) );
  INV_X1 U6964 ( .A(n6014), .ZN(n5851) );
  NAND2_X1 U6965 ( .A1(n5851), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6035) );
  INV_X1 U6966 ( .A(n6147), .ZN(n5855) );
  INV_X1 U6967 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6192) );
  INV_X1 U6968 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6221) );
  INV_X1 U6969 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9811) );
  INV_X1 U6970 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9866) );
  INV_X1 U6971 ( .A(n5896), .ZN(n5860) );
  INV_X1 U6972 ( .A(n5889), .ZN(n5861) );
  NAND2_X1 U6973 ( .A1(n5861), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6271) );
  INV_X1 U6974 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6975 ( .A1(n5889), .A2(n5862), .ZN(n5863) );
  NAND2_X1 U6976 ( .A1(n6271), .A2(n5863), .ZN(n10518) );
  OAI21_X1 U6977 ( .B1(n5865), .B2(n5969), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5867) );
  INV_X2 U6978 ( .A(n5872), .ZN(n5870) );
  INV_X1 U6979 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5875) );
  AND2_X2 U6980 ( .A1(n5871), .A2(n5872), .ZN(n5926) );
  NAND2_X1 U6981 ( .A1(n8848), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5874) );
  AND2_X2 U6982 ( .A1(n9223), .A2(n5872), .ZN(n5944) );
  NAND2_X1 U6983 ( .A1(n5960), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5873) );
  OAI211_X1 U6984 ( .C1(n6405), .C2(n5875), .A(n5874), .B(n5873), .ZN(n5876)
         );
  INV_X1 U6985 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U6986 ( .A1(n5880), .A2(n5879), .ZN(n5882) );
  NAND2_X1 U6987 ( .A1(n5882), .A2(n5881), .ZN(n5884) );
  NAND2_X1 U6988 ( .A1(n5884), .A2(n5883), .ZN(n8830) );
  INV_X1 U6989 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8268) );
  OR2_X1 U6990 ( .A1(n8853), .A2(n8268), .ZN(n5885) );
  INV_X1 U6991 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U6992 ( .A1(n5896), .A2(n5887), .ZN(n5888) );
  NAND2_X1 U6993 ( .A1(n5889), .A2(n5888), .ZN(n10540) );
  INV_X1 U6994 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U6995 ( .A1(n8848), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6996 ( .A1(n5960), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5890) );
  OAI211_X1 U6997 ( .C1(n6405), .C2(n10701), .A(n5891), .B(n5890), .ZN(n5892)
         );
  INV_X1 U6998 ( .A(n5892), .ZN(n5893) );
  NAND2_X1 U6999 ( .A1(n6257), .A2(n9866), .ZN(n5895) );
  AND2_X1 U7000 ( .A1(n5896), .A2(n5895), .ZN(n10555) );
  NAND2_X1 U7001 ( .A1(n10555), .A2(n6289), .ZN(n5901) );
  INV_X1 U7002 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10707) );
  NAND2_X1 U7003 ( .A1(n8848), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7004 ( .A1(n5960), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U7005 ( .C1(n6405), .C2(n10707), .A(n5898), .B(n5897), .ZN(n5899)
         );
  INV_X1 U7006 ( .A(n5899), .ZN(n5900) );
  XNOR2_X1 U7007 ( .A(n5903), .B(n5902), .ZN(n8639) );
  NAND2_X1 U7008 ( .A1(n8639), .A2(n8854), .ZN(n5905) );
  INV_X1 U7009 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8243) );
  OR2_X1 U7010 ( .A1(n8853), .A2(n8243), .ZN(n5904) );
  NAND2_X1 U7011 ( .A1(n5944), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7012 ( .A1(n5926), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5906) );
  AND2_X1 U7013 ( .A1(n5907), .A2(n5906), .ZN(n5910) );
  NAND2_X1 U7014 ( .A1(n8847), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7015 ( .A1(n5134), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5908) );
  OR2_X1 U7016 ( .A1(n5911), .A2(n5969), .ZN(n5949) );
  INV_X1 U7017 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6731) );
  INV_X1 U7018 ( .A(n5912), .ZN(n5914) );
  NAND2_X1 U7019 ( .A1(n5914), .A2(n5913), .ZN(n5916) );
  NAND2_X1 U7020 ( .A1(n5916), .A2(n5915), .ZN(n8842) );
  INV_X1 U7021 ( .A(n6869), .ZN(n5917) );
  NAND2_X1 U7022 ( .A1(n7014), .A2(n6869), .ZN(n8905) );
  NAND2_X1 U7023 ( .A1(n5137), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7024 ( .A1(n5135), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7025 ( .A1(n5944), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5918) );
  AND3_X1 U7026 ( .A1(n5920), .A2(n5919), .A3(n5918), .ZN(n5922) );
  NAND2_X1 U7027 ( .A1(n5926), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5921) );
  NOR2_X1 U7028 ( .A1(n8701), .A2(n5923), .ZN(n5925) );
  XNOR2_X1 U7029 ( .A(n5925), .B(n5924), .ZN(n10823) );
  MUX2_X1 U7030 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10823), .S(n6707), .Z(n6964)
         );
  NAND2_X1 U7031 ( .A1(n6426), .A2(n6964), .ZN(n6874) );
  NAND2_X1 U7032 ( .A1(n5944), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7033 ( .A1(n5926), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5927) );
  AND2_X2 U7034 ( .A1(n5928), .A2(n5927), .ZN(n5931) );
  NAND2_X1 U7035 ( .A1(n5136), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7036 ( .A1(n6195), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5929) );
  INV_X1 U7037 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7038 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  AND2_X1 U7039 ( .A1(n5936), .A2(n5935), .ZN(n7114) );
  INV_X1 U7040 ( .A(n7114), .ZN(n6739) );
  NAND2_X1 U7041 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5937) );
  MUX2_X1 U7042 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5937), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5939) );
  INV_X1 U7043 ( .A(n5911), .ZN(n5938) );
  NAND2_X1 U7044 ( .A1(n5939), .A2(n5938), .ZN(n6784) );
  OR2_X1 U7045 ( .A1(n6707), .A2(n6784), .ZN(n5940) );
  INV_X1 U7046 ( .A(n6434), .ZN(n6967) );
  NAND2_X1 U7047 ( .A1(n6967), .A2(n5941), .ZN(n5942) );
  NAND2_X1 U7048 ( .A1(n6873), .A2(n5942), .ZN(n6868) );
  INV_X1 U7049 ( .A(n6869), .ZN(n7086) );
  NAND2_X1 U7050 ( .A1(n7014), .A2(n7086), .ZN(n5943) );
  INV_X1 U7051 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7031) );
  NAND2_X1 U7052 ( .A1(n5135), .A2(n7031), .ZN(n5948) );
  NAND2_X1 U7053 ( .A1(n5926), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7054 ( .A1(n8847), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7055 ( .A1(n5944), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7056 ( .A1(n5949), .A2(n10276), .ZN(n5950) );
  NAND2_X1 U7057 ( .A1(n5950), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5952) );
  INV_X1 U7058 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7059 ( .A(n5952), .B(n5951), .ZN(n10358) );
  INV_X1 U7060 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6723) );
  OR2_X1 U7061 ( .A1(n8853), .A2(n6723), .ZN(n5958) );
  OR2_X1 U7062 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7063 ( .A1(n5956), .A2(n5955), .ZN(n7316) );
  OR2_X1 U7064 ( .A1(n6396), .A2(n7316), .ZN(n5957) );
  OAI211_X1 U7065 ( .C1(n6707), .C2(n10358), .A(n5958), .B(n5957), .ZN(n6985)
         );
  NAND2_X1 U7066 ( .A1(n6997), .A2(n6985), .ZN(n9061) );
  NAND2_X1 U7067 ( .A1(n6889), .A2(n8858), .ZN(n6888) );
  NAND2_X1 U7068 ( .A1(n6997), .A2(n7034), .ZN(n5959) );
  NAND2_X1 U7069 ( .A1(n6888), .A2(n5959), .ZN(n6992) );
  NAND2_X1 U7070 ( .A1(n5960), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5966) );
  INV_X1 U7071 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7072 ( .A1(n7031), .A2(n5961), .ZN(n5962) );
  AND2_X1 U7073 ( .A1(n5962), .A2(n5982), .ZN(n9880) );
  NAND2_X1 U7074 ( .A1(n6289), .A2(n9880), .ZN(n5965) );
  NAND2_X1 U7075 ( .A1(n5926), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7076 ( .A1(n8847), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5963) );
  AND4_X2 U7077 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n7420)
         );
  NOR2_X1 U7078 ( .A1(n5967), .A2(n5969), .ZN(n5968) );
  MUX2_X1 U7079 ( .A(n5969), .B(n5968), .S(P1_IR_REG_4__SCAN_IN), .Z(n5970) );
  INV_X1 U7080 ( .A(n5970), .ZN(n5972) );
  NAND2_X1 U7081 ( .A1(n5967), .A2(n5971), .ZN(n6006) );
  NAND2_X1 U7082 ( .A1(n5972), .A2(n6006), .ZN(n10373) );
  OR2_X1 U7083 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U7084 ( .A1(n5976), .A2(n5975), .ZN(n7527) );
  OR2_X1 U7085 ( .A1(n6396), .A2(n7527), .ZN(n5978) );
  INV_X1 U7086 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6724) );
  OR2_X1 U7087 ( .A1(n8853), .A2(n6724), .ZN(n5977) );
  OAI211_X1 U7088 ( .C1(n6707), .C2(n10373), .A(n5978), .B(n5977), .ZN(n5979)
         );
  NAND2_X1 U7089 ( .A1(n7420), .A2(n5979), .ZN(n8910) );
  INV_X2 U7090 ( .A(n7420), .ZN(n10355) );
  INV_X1 U7091 ( .A(n5979), .ZN(n7000) );
  NAND2_X1 U7092 ( .A1(n10355), .A2(n7000), .ZN(n9063) );
  NAND2_X1 U7093 ( .A1(n8910), .A2(n9063), .ZN(n8861) );
  NAND2_X1 U7094 ( .A1(n6992), .A2(n8861), .ZN(n6991) );
  NAND2_X1 U7095 ( .A1(n7420), .A2(n7000), .ZN(n5980) );
  NAND2_X1 U7096 ( .A1(n6991), .A2(n5980), .ZN(n6970) );
  NAND2_X1 U7097 ( .A1(n8847), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7098 ( .A1(n5960), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5986) );
  INV_X1 U7099 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7100 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  AND2_X1 U7101 ( .A1(n5996), .A2(n5983), .ZN(n7423) );
  NAND2_X1 U7102 ( .A1(n5134), .A2(n7423), .ZN(n5985) );
  NAND2_X1 U7103 ( .A1(n5926), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7104 ( .A1(n6006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7105 ( .A(n5988), .B(n10079), .ZN(n6801) );
  OR2_X1 U7106 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  AND2_X1 U7107 ( .A1(n5992), .A2(n5991), .ZN(n7533) );
  INV_X1 U7108 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6725) );
  OR2_X1 U7109 ( .A1(n8853), .A2(n6725), .ZN(n5993) );
  NAND2_X1 U7110 ( .A1(n9877), .A2(n7418), .ZN(n8911) );
  INV_X1 U7111 ( .A(n9877), .ZN(n10354) );
  NAND2_X1 U7112 ( .A1(n8911), .A2(n9064), .ZN(n8917) );
  NAND2_X1 U7113 ( .A1(n9877), .A2(n11129), .ZN(n5994) );
  NAND2_X1 U7114 ( .A1(n5960), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7115 ( .A1(n8847), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6000) );
  INV_X1 U7116 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7117 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  AND2_X1 U7118 ( .A1(n6014), .A2(n5997), .ZN(n7409) );
  NAND2_X1 U7119 ( .A1(n6289), .A2(n7409), .ZN(n5999) );
  NAND2_X1 U7120 ( .A1(n5926), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7121 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7122 ( .A1(n6005), .A2(n6004), .ZN(n7578) );
  OR2_X1 U7123 ( .A1(n7578), .A2(n6396), .ZN(n6011) );
  AND2_X1 U7124 ( .A1(n6030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7125 ( .A1(n6007), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6009) );
  INV_X1 U7126 ( .A(n6007), .ZN(n6008) );
  NAND2_X1 U7127 ( .A1(n6008), .A2(n10283), .ZN(n6023) );
  AOI22_X1 U7128 ( .A1(n6206), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6205), .B2(
        n6852), .ZN(n6010) );
  NAND2_X1 U7129 ( .A1(n6011), .A2(n6010), .ZN(n7405) );
  NAND2_X1 U7130 ( .A1(n7042), .A2(n7405), .ZN(n9067) );
  INV_X1 U7131 ( .A(n7042), .ZN(n10353) );
  NAND2_X1 U7132 ( .A1(n10353), .A2(n7064), .ZN(n9070) );
  NAND2_X1 U7133 ( .A1(n9067), .A2(n9070), .ZN(n8914) );
  NAND2_X1 U7134 ( .A1(n7042), .A2(n7064), .ZN(n6012) );
  NAND2_X1 U7135 ( .A1(n8847), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7136 ( .A1(n5960), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6018) );
  INV_X1 U7137 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7138 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  AND2_X1 U7139 ( .A1(n6035), .A2(n6015), .ZN(n7443) );
  NAND2_X1 U7140 ( .A1(n6289), .A2(n7443), .ZN(n6017) );
  NAND2_X1 U7141 ( .A1(n5926), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7142 ( .A1(n7750), .A2(n6396), .ZN(n6026) );
  NAND2_X1 U7143 ( .A1(n6023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6024) );
  XNOR2_X1 U7144 ( .A(n6024), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7145 ( .A1(n6206), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6205), .B2(
        n6909), .ZN(n6025) );
  NAND2_X1 U7146 ( .A1(n6026), .A2(n6025), .ZN(n7049) );
  OR2_X1 U7147 ( .A1(n7353), .A2(n7049), .ZN(n8922) );
  NAND2_X1 U7148 ( .A1(n7353), .A2(n7049), .ZN(n8921) );
  NAND2_X1 U7149 ( .A1(n8922), .A2(n8921), .ZN(n8868) );
  INV_X1 U7150 ( .A(n7353), .ZN(n10352) );
  NAND2_X1 U7151 ( .A1(n7825), .A2(n8854), .ZN(n6033) );
  NAND2_X1 U7152 ( .A1(n10283), .A2(n10284), .ZN(n6029) );
  NOR2_X1 U7153 ( .A1(n6030), .A2(n6029), .ZN(n6044) );
  OR2_X1 U7154 ( .A1(n6044), .A2(n5969), .ZN(n6031) );
  XNOR2_X1 U7155 ( .A(n6031), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7638) );
  AOI22_X1 U7156 ( .A1(n6206), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6205), .B2(
        n7638), .ZN(n6032) );
  NAND2_X1 U7157 ( .A1(n5960), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7158 ( .A1(n8847), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7159 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  AND2_X1 U7160 ( .A1(n6047), .A2(n6036), .ZN(n7999) );
  NAND2_X1 U7161 ( .A1(n5135), .A2(n7999), .ZN(n6038) );
  NAND2_X1 U7162 ( .A1(n5926), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7163 ( .A1(n8009), .A2(n7868), .ZN(n8901) );
  NAND2_X1 U7164 ( .A1(n8009), .A2(n7868), .ZN(n8926) );
  NAND2_X1 U7165 ( .A1(n8901), .A2(n8926), .ZN(n8866) );
  NAND2_X1 U7166 ( .A1(n7347), .A2(n8866), .ZN(n7346) );
  INV_X1 U7167 ( .A(n7868), .ZN(n10351) );
  OR2_X1 U7168 ( .A1(n8009), .A2(n10351), .ZN(n6041) );
  NAND2_X1 U7169 ( .A1(n7346), .A2(n6041), .ZN(n7382) );
  XNOR2_X1 U7170 ( .A(n6043), .B(n6042), .ZN(n7934) );
  NAND2_X1 U7171 ( .A1(n7934), .A2(n8854), .ZN(n6046) );
  NAND2_X1 U7172 ( .A1(n6044), .A2(n10288), .ZN(n6093) );
  NAND2_X1 U7173 ( .A1(n6093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6059) );
  XNOR2_X1 U7174 ( .A(n6059), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U7175 ( .A1(n6206), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6205), .B2(
        n10397), .ZN(n6045) );
  NAND2_X1 U7176 ( .A1(n6046), .A2(n6045), .ZN(n7456) );
  NAND2_X1 U7177 ( .A1(n5960), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7178 ( .A1(n8847), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6051) );
  INV_X1 U7179 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U7180 ( .A1(n6047), .A2(n7866), .ZN(n6048) );
  AND2_X1 U7181 ( .A1(n6067), .A2(n6048), .ZN(n7870) );
  NAND2_X1 U7182 ( .A1(n6289), .A2(n7870), .ZN(n6050) );
  NAND2_X1 U7183 ( .A1(n8848), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6049) );
  OR2_X1 U7184 ( .A1(n7456), .A2(n8002), .ZN(n8891) );
  NAND2_X1 U7185 ( .A1(n7456), .A2(n8002), .ZN(n8896) );
  NAND2_X1 U7186 ( .A1(n8891), .A2(n8896), .ZN(n8857) );
  INV_X1 U7187 ( .A(n8002), .ZN(n7739) );
  OR2_X1 U7188 ( .A1(n7456), .A2(n7739), .ZN(n6053) );
  NAND2_X1 U7189 ( .A1(n7381), .A2(n6053), .ZN(n7372) );
  INV_X1 U7190 ( .A(n6055), .ZN(n6057) );
  NAND2_X1 U7191 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NAND2_X1 U7192 ( .A1(n6060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7193 ( .A1(n6062), .A2(n6061), .ZN(n6083) );
  OR2_X1 U7194 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  AOI22_X1 U7195 ( .A1(n6206), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6205), .B2(
        n10963), .ZN(n6064) );
  NAND2_X1 U7196 ( .A1(n8847), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7197 ( .A1(n5960), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7198 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  AND2_X1 U7199 ( .A1(n6075), .A2(n6068), .ZN(n7740) );
  NAND2_X1 U7200 ( .A1(n6289), .A2(n7740), .ZN(n6070) );
  NAND2_X1 U7201 ( .A1(n8848), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7202 ( .A1(n7744), .A2(n7515), .ZN(n9077) );
  NAND2_X1 U7203 ( .A1(n7744), .A2(n7515), .ZN(n8894) );
  NAND2_X1 U7204 ( .A1(n9077), .A2(n8894), .ZN(n7371) );
  INV_X1 U7205 ( .A(n7515), .ZN(n11157) );
  OR2_X1 U7206 ( .A1(n7744), .A2(n11157), .ZN(n6073) );
  NAND2_X1 U7207 ( .A1(n8847), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7208 ( .A1(n5960), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6079) );
  INV_X1 U7209 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7210 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  AND2_X1 U7211 ( .A1(n6099), .A2(n6076), .ZN(n7816) );
  NAND2_X1 U7212 ( .A1(n6289), .A2(n7816), .ZN(n6078) );
  NAND2_X1 U7213 ( .A1(n8848), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7214 ( .A1(n8011), .A2(n8854), .ZN(n6086) );
  NAND2_X1 U7215 ( .A1(n6083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7216 ( .A(n6084), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U7217 ( .A1(n6206), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6205), .B2(
        n10891), .ZN(n6085) );
  NAND2_X1 U7218 ( .A1(n6088), .A2(n6087), .ZN(n6090) );
  NAND2_X1 U7219 ( .A1(n6090), .A2(n6089), .ZN(n8106) );
  OR2_X1 U7220 ( .A1(n8106), .A2(n6396), .ZN(n6097) );
  INV_X1 U7221 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6091) );
  NAND3_X1 U7222 ( .A1(n6091), .A2(n6058), .A3(n6061), .ZN(n6092) );
  OAI21_X1 U7223 ( .B1(n6093), .B2(n6092), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6094) );
  MUX2_X1 U7224 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6094), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6095) );
  AND2_X1 U7225 ( .A1(n6111), .A2(n6095), .ZN(n10412) );
  AOI22_X1 U7226 ( .A1(n6206), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6205), .B2(
        n10412), .ZN(n6096) );
  NAND2_X1 U7227 ( .A1(n5960), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7228 ( .A1(n8847), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7229 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  AND2_X1 U7230 ( .A1(n6118), .A2(n6100), .ZN(n8073) );
  NAND2_X1 U7231 ( .A1(n5135), .A2(n8073), .ZN(n6102) );
  NAND2_X1 U7232 ( .A1(n8848), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6101) );
  NAND4_X1 U7233 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n11154)
         );
  NOR2_X1 U7234 ( .A1(n7671), .A2(n11154), .ZN(n6106) );
  NAND2_X1 U7235 ( .A1(n7671), .A2(n11154), .ZN(n6105) );
  OR2_X1 U7236 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  NAND2_X1 U7237 ( .A1(n6110), .A2(n6109), .ZN(n8161) );
  OR2_X1 U7238 ( .A1(n8161), .A2(n6396), .ZN(n6116) );
  NAND2_X1 U7239 ( .A1(n6111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6112) );
  MUX2_X1 U7240 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6112), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6114) );
  AOI22_X1 U7241 ( .A1(n6206), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6205), .B2(
        n10948), .ZN(n6115) );
  NAND2_X1 U7242 ( .A1(n8847), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7243 ( .A1(n5960), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7244 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  AND2_X1 U7245 ( .A1(n6134), .A2(n6119), .ZN(n8156) );
  NAND2_X1 U7246 ( .A1(n6289), .A2(n8156), .ZN(n6121) );
  NAND2_X1 U7247 ( .A1(n8848), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6120) );
  NAND4_X1 U7248 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n10348)
         );
  INV_X1 U7249 ( .A(n10348), .ZN(n8285) );
  NAND2_X1 U7250 ( .A1(n8159), .A2(n8285), .ZN(n6124) );
  XNOR2_X1 U7251 ( .A(n6126), .B(n6125), .ZN(n8517) );
  NAND2_X1 U7252 ( .A1(n8517), .A2(n8854), .ZN(n6132) );
  NAND2_X1 U7253 ( .A1(n6128), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6127) );
  MUX2_X1 U7254 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6127), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6130) );
  INV_X1 U7255 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U7256 ( .A1(n6129), .A2(n10296), .ZN(n6156) );
  NAND2_X1 U7257 ( .A1(n6130), .A2(n6156), .ZN(n10422) );
  AOI22_X1 U7258 ( .A1(n6206), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6205), .B2(
        n10904), .ZN(n6131) );
  NAND2_X1 U7259 ( .A1(n5960), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7260 ( .A1(n8847), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6138) );
  INV_X1 U7261 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7262 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  AND2_X1 U7263 ( .A1(n6147), .A2(n6135), .ZN(n8287) );
  NAND2_X1 U7264 ( .A1(n5134), .A2(n8287), .ZN(n6137) );
  NAND2_X1 U7265 ( .A1(n8848), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7266 ( .A1(n6540), .A2(n10764), .ZN(n8942) );
  NAND2_X1 U7267 ( .A1(n6141), .A2(n6140), .ZN(n6143) );
  NAND2_X1 U7268 ( .A1(n6143), .A2(n6142), .ZN(n8508) );
  OR2_X1 U7269 ( .A1(n8508), .A2(n6396), .ZN(n6146) );
  NAND2_X1 U7270 ( .A1(n6156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U7271 ( .A(n6144), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U7272 ( .A1(n6206), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6205), .B2(
        n10917), .ZN(n6145) );
  NAND2_X1 U7273 ( .A1(n5960), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7274 ( .A1(n8848), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6151) );
  INV_X1 U7275 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U7276 ( .A1(n6147), .A2(n8339), .ZN(n6148) );
  AND2_X1 U7277 ( .A1(n6164), .A2(n6148), .ZN(n8819) );
  NAND2_X1 U7278 ( .A1(n5134), .A2(n8819), .ZN(n6150) );
  NAND2_X1 U7279 ( .A1(n8847), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6149) );
  NAND4_X1 U7280 ( .A1(n6152), .A2(n6151), .A3(n6150), .A4(n6149), .ZN(n10346)
         );
  NAND2_X1 U7281 ( .A1(n6546), .A2(n10346), .ZN(n8948) );
  NAND2_X1 U7282 ( .A1(n10767), .A2(n10756), .ZN(n8947) );
  NAND2_X1 U7283 ( .A1(n8948), .A2(n8947), .ZN(n8874) );
  NAND2_X1 U7284 ( .A1(n10767), .A2(n10346), .ZN(n6153) );
  NAND2_X1 U7285 ( .A1(n8813), .A2(n6153), .ZN(n8141) );
  XNOR2_X1 U7286 ( .A(n6155), .B(n6154), .ZN(n8531) );
  NAND2_X1 U7287 ( .A1(n8531), .A2(n8854), .ZN(n6162) );
  INV_X1 U7288 ( .A(n6156), .ZN(n6158) );
  NAND2_X1 U7289 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  NAND2_X1 U7290 ( .A1(n6187), .A2(n10096), .ZN(n6172) );
  OR2_X1 U7291 ( .A1(n6187), .A2(n10096), .ZN(n6160) );
  AOI22_X1 U7292 ( .A1(n6206), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6205), .B2(
        n10441), .ZN(n6161) );
  NAND2_X1 U7293 ( .A1(n5960), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7294 ( .A1(n8848), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7295 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  AND2_X1 U7296 ( .A1(n6177), .A2(n6165), .ZN(n9849) );
  NAND2_X1 U7297 ( .A1(n6289), .A2(n9849), .ZN(n6167) );
  NAND2_X1 U7298 ( .A1(n8847), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7299 ( .A1(n10759), .A2(n9857), .ZN(n9087) );
  NAND2_X1 U7300 ( .A1(n8950), .A2(n9087), .ZN(n8144) );
  NAND2_X1 U7301 ( .A1(n8141), .A2(n8144), .ZN(n8140) );
  INV_X1 U7302 ( .A(n10759), .ZN(n9846) );
  XNOR2_X1 U7303 ( .A(n6171), .B(n6170), .ZN(n8547) );
  NAND2_X1 U7304 ( .A1(n8547), .A2(n8854), .ZN(n6175) );
  NAND2_X1 U7305 ( .A1(n6172), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6173) );
  XNOR2_X1 U7306 ( .A(n6173), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U7307 ( .A1(n6206), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6205), .B2(
        n10457), .ZN(n6174) );
  NAND2_X1 U7308 ( .A1(n5960), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7309 ( .A1(n8848), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6181) );
  INV_X1 U7310 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7311 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  AND2_X1 U7312 ( .A1(n6193), .A2(n6178), .ZN(n9859) );
  NAND2_X1 U7313 ( .A1(n5135), .A2(n9859), .ZN(n6180) );
  NAND2_X1 U7314 ( .A1(n8847), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7315 ( .A1(n10753), .A2(n10740), .ZN(n8890) );
  NAND2_X1 U7316 ( .A1(n10753), .A2(n10740), .ZN(n8960) );
  NAND2_X1 U7317 ( .A1(n8890), .A2(n8960), .ZN(n8248) );
  NAND2_X1 U7318 ( .A1(n5141), .A2(n6183), .ZN(n6184) );
  NAND2_X1 U7319 ( .A1(n6185), .A2(n6184), .ZN(n8555) );
  OR2_X1 U7320 ( .A1(n8555), .A2(n6396), .ZN(n6191) );
  OAI21_X1 U7321 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7322 ( .A1(n6188), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6189) );
  AND2_X1 U7323 ( .A1(n6203), .A2(n6189), .ZN(n10934) );
  AOI22_X1 U7324 ( .A1(n6206), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6205), .B2(
        n10934), .ZN(n6190) );
  NAND2_X1 U7325 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  AND2_X1 U7326 ( .A1(n6212), .A2(n6194), .ZN(n9916) );
  NAND2_X1 U7327 ( .A1(n5134), .A2(n9916), .ZN(n6199) );
  NAND2_X1 U7328 ( .A1(n5960), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7329 ( .A1(n8847), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7330 ( .A1(n8848), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7331 ( .A1(n9913), .A2(n10644), .ZN(n6200) );
  XNOR2_X1 U7332 ( .A(n6202), .B(n6201), .ZN(n8577) );
  NAND2_X1 U7333 ( .A1(n8577), .A2(n8854), .ZN(n6208) );
  XNOR2_X2 U7334 ( .A(n6204), .B(n10303), .ZN(n6421) );
  AOI22_X1 U7335 ( .A1(n6206), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10464), 
        .B2(n6205), .ZN(n6207) );
  NAND2_X1 U7336 ( .A1(n5960), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7337 ( .A1(n8847), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6209) );
  AND2_X1 U7338 ( .A1(n6210), .A2(n6209), .ZN(n6216) );
  INV_X1 U7339 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7340 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  NAND2_X1 U7341 ( .A1(n6222), .A2(n6213), .ZN(n10660) );
  OR2_X1 U7342 ( .A1(n10660), .A2(n6258), .ZN(n6215) );
  NAND2_X1 U7343 ( .A1(n8848), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7344 ( .A1(n10657), .A2(n10742), .ZN(n8959) );
  NAND2_X1 U7345 ( .A1(n10657), .A2(n10742), .ZN(n9094) );
  XNOR2_X1 U7346 ( .A(n6218), .B(n6217), .ZN(n8587) );
  NAND2_X1 U7347 ( .A1(n8587), .A2(n8854), .ZN(n6220) );
  INV_X1 U7348 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10054) );
  OR2_X1 U7349 ( .A1(n8853), .A2(n10054), .ZN(n6219) );
  NAND2_X1 U7350 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  AND2_X1 U7351 ( .A1(n6233), .A2(n6223), .ZN(n10633) );
  NAND2_X1 U7352 ( .A1(n10633), .A2(n6289), .ZN(n6226) );
  AOI22_X1 U7353 ( .A1(n8848), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n5960), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7354 ( .A1(n8847), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7355 ( .A1(n10631), .A2(n10645), .ZN(n8973) );
  NAND2_X1 U7356 ( .A1(n10631), .A2(n10645), .ZN(n8886) );
  INV_X1 U7357 ( .A(n10645), .ZN(n10616) );
  INV_X1 U7358 ( .A(n6227), .ZN(n6229) );
  XNOR2_X1 U7359 ( .A(n6229), .B(n6228), .ZN(n8599) );
  NAND2_X1 U7360 ( .A1(n8599), .A2(n8854), .ZN(n6231) );
  INV_X1 U7361 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7873) );
  OR2_X1 U7362 ( .A1(n8853), .A2(n7873), .ZN(n6230) );
  INV_X1 U7363 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7364 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  NAND2_X1 U7365 ( .A1(n6243), .A2(n6234), .ZN(n10609) );
  OR2_X1 U7366 ( .A1(n10609), .A2(n6258), .ZN(n6237) );
  AOI22_X1 U7367 ( .A1(n8847), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5960), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7368 ( .A1(n8848), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7369 ( .A1(n10725), .A2(n10626), .ZN(n8974) );
  NAND2_X1 U7370 ( .A1(n10725), .A2(n10626), .ZN(n8975) );
  NAND2_X1 U7371 ( .A1(n8974), .A2(n8975), .ZN(n10605) );
  XNOR2_X1 U7372 ( .A(n6239), .B(SI_22_), .ZN(n8612) );
  NAND2_X1 U7373 ( .A1(n8612), .A2(n8854), .ZN(n6241) );
  INV_X1 U7374 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8086) );
  OR2_X1 U7375 ( .A1(n8853), .A2(n8086), .ZN(n6240) );
  INV_X1 U7376 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7377 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  NAND2_X1 U7378 ( .A1(n6255), .A2(n6244), .ZN(n10596) );
  OR2_X1 U7379 ( .A1(n10596), .A2(n6258), .ZN(n6249) );
  INV_X1 U7380 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U7381 ( .A1(n8848), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7382 ( .A1(n5960), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6245) );
  OAI211_X1 U7383 ( .C1(n6405), .C2(n10722), .A(n6246), .B(n6245), .ZN(n6247)
         );
  INV_X1 U7384 ( .A(n6247), .ZN(n6248) );
  OR2_X1 U7385 ( .A1(n10595), .A2(n9812), .ZN(n8969) );
  NAND2_X1 U7386 ( .A1(n10595), .A2(n9812), .ZN(n8978) );
  NAND2_X1 U7387 ( .A1(n8969), .A2(n8978), .ZN(n10586) );
  XNOR2_X1 U7388 ( .A(n6252), .B(n6251), .ZN(n8626) );
  NAND2_X1 U7389 ( .A1(n8626), .A2(n8854), .ZN(n6254) );
  INV_X1 U7390 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8130) );
  OR2_X1 U7391 ( .A1(n8853), .A2(n8130), .ZN(n6253) );
  NAND2_X1 U7392 ( .A1(n6255), .A2(n9811), .ZN(n6256) );
  NAND2_X1 U7393 ( .A1(n6257), .A2(n6256), .ZN(n10567) );
  OR2_X1 U7394 ( .A1(n10567), .A2(n6258), .ZN(n6263) );
  INV_X1 U7395 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U7396 ( .A1(n5960), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7397 ( .A1(n8848), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6259) );
  OAI211_X1 U7398 ( .C1(n6405), .C2(n10717), .A(n6260), .B(n6259), .ZN(n6261)
         );
  INV_X1 U7399 ( .A(n6261), .ZN(n6262) );
  NAND2_X1 U7400 ( .A1(n6263), .A2(n6262), .ZN(n10590) );
  OR2_X1 U7401 ( .A1(n10688), .A2(n10694), .ZN(n9028) );
  NAND2_X1 U7402 ( .A1(n10688), .A2(n10694), .ZN(n8992) );
  NAND2_X1 U7403 ( .A1(n9028), .A2(n8992), .ZN(n10526) );
  INV_X1 U7404 ( .A(n6265), .ZN(n6266) );
  INV_X1 U7405 ( .A(SI_26_), .ZN(n10141) );
  NAND2_X1 U7406 ( .A1(n6266), .A2(n10141), .ZN(n6282) );
  MUX2_X1 U7407 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n8701), .Z(n6279) );
  INV_X1 U7408 ( .A(SI_27_), .ZN(n6280) );
  XNOR2_X1 U7409 ( .A(n6279), .B(n6280), .ZN(n6284) );
  NAND2_X1 U7410 ( .A1(n8674), .A2(n8854), .ZN(n6269) );
  INV_X1 U7411 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8347) );
  OR2_X1 U7412 ( .A1(n8853), .A2(n8347), .ZN(n6268) );
  NAND2_X2 U7413 ( .A1(n6269), .A2(n6268), .ZN(n10679) );
  INV_X1 U7414 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7415 ( .A1(n6271), .A2(n6270), .ZN(n6272) );
  NAND2_X1 U7416 ( .A1(n10502), .A2(n6289), .ZN(n6278) );
  INV_X1 U7417 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7418 ( .A1(n5960), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7419 ( .A1(n8848), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6273) );
  OAI211_X1 U7420 ( .C1(n6405), .C2(n6275), .A(n6274), .B(n6273), .ZN(n6276)
         );
  INV_X1 U7421 ( .A(n6276), .ZN(n6277) );
  OR2_X1 U7422 ( .A1(n10679), .A2(n10685), .ZN(n9029) );
  INV_X1 U7423 ( .A(n6279), .ZN(n6281) );
  NAND2_X1 U7424 ( .A1(n6281), .A2(n6280), .ZN(n6283) );
  AND2_X1 U7425 ( .A1(n6282), .A2(n6283), .ZN(n6386) );
  INV_X1 U7426 ( .A(n6283), .ZN(n6285) );
  OR2_X1 U7427 ( .A1(n6285), .A2(n6284), .ZN(n6380) );
  MUX2_X1 U7428 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8701), .Z(n6378) );
  INV_X1 U7429 ( .A(SI_28_), .ZN(n10137) );
  XNOR2_X1 U7430 ( .A(n6378), .B(n10137), .ZN(n6381) );
  INV_X1 U7431 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8345) );
  OR2_X1 U7432 ( .A1(n8853), .A2(n8345), .ZN(n6288) );
  XNOR2_X1 U7433 ( .A(n6326), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n10491) );
  NAND2_X1 U7434 ( .A1(n10491), .A2(n6289), .ZN(n6294) );
  INV_X1 U7435 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7436 ( .A1(n8848), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7437 ( .A1(n5960), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6290) );
  OAI211_X1 U7438 ( .C1(n6405), .C2(n6373), .A(n6291), .B(n6290), .ZN(n6292)
         );
  INV_X1 U7439 ( .A(n6292), .ZN(n6293) );
  NAND2_X1 U7440 ( .A1(n6680), .A2(n10676), .ZN(n9020) );
  XNOR2_X1 U7441 ( .A(n6377), .B(n8998), .ZN(n10485) );
  NAND2_X1 U7442 ( .A1(n6299), .A2(n6341), .ZN(n6296) );
  NAND2_X1 U7443 ( .A1(n6297), .A2(n10312), .ZN(n6348) );
  MUX2_X1 U7444 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6300), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6301) );
  NAND2_X1 U7445 ( .A1(n8860), .A2(n9120), .ZN(n6424) );
  OR2_X1 U7446 ( .A1(n6423), .A2(n6424), .ZN(n6660) );
  INV_X1 U7447 ( .A(n6655), .ZN(n6827) );
  AND2_X1 U7448 ( .A1(n6660), .A2(n6827), .ZN(n6960) );
  NAND2_X1 U7449 ( .A1(n6421), .A2(n9120), .ZN(n6420) );
  NAND2_X1 U7450 ( .A1(n6420), .A2(n6423), .ZN(n6303) );
  NAND2_X1 U7451 ( .A1(n6960), .A2(n6303), .ZN(n11166) );
  INV_X1 U7452 ( .A(n11164), .ZN(n8233) );
  INV_X1 U7453 ( .A(n6880), .ZN(n8865) );
  NOR2_X1 U7454 ( .A1(n6426), .A2(n6877), .ZN(n6879) );
  NAND2_X1 U7455 ( .A1(n8865), .A2(n6879), .ZN(n6305) );
  NAND2_X1 U7456 ( .A1(n6967), .A2(n7011), .ZN(n6304) );
  NAND2_X1 U7457 ( .A1(n6305), .A2(n6304), .ZN(n8904) );
  NAND2_X1 U7458 ( .A1(n8908), .A2(n9064), .ZN(n6306) );
  NAND2_X1 U7459 ( .A1(n6306), .A2(n8911), .ZN(n7020) );
  NAND2_X1 U7460 ( .A1(n7020), .A2(n9070), .ZN(n6307) );
  NAND2_X1 U7461 ( .A1(n6307), .A2(n9067), .ZN(n7349) );
  AND2_X1 U7462 ( .A1(n8901), .A2(n8922), .ZN(n6308) );
  AND2_X1 U7463 ( .A1(n8891), .A2(n6308), .ZN(n9071) );
  NAND2_X1 U7464 ( .A1(n7349), .A2(n9071), .ZN(n6311) );
  NAND2_X1 U7465 ( .A1(n8926), .A2(n8921), .ZN(n6309) );
  NAND3_X1 U7466 ( .A1(n8891), .A2(n8901), .A3(n6309), .ZN(n6310) );
  AND2_X1 U7467 ( .A1(n6310), .A2(n8896), .ZN(n9073) );
  NAND2_X1 U7468 ( .A1(n6311), .A2(n9073), .ZN(n7369) );
  INV_X1 U7469 ( .A(n7371), .ZN(n8928) );
  NAND2_X1 U7470 ( .A1(n7369), .A2(n8928), .ZN(n6312) );
  NAND2_X1 U7471 ( .A1(n7821), .A2(n10349), .ZN(n8895) );
  INV_X1 U7472 ( .A(n11154), .ZN(n7819) );
  OR2_X1 U7473 ( .A1(n7671), .A2(n7819), .ZN(n8940) );
  NAND2_X1 U7474 ( .A1(n7671), .A2(n7819), .ZN(n9078) );
  NAND2_X1 U7475 ( .A1(n7666), .A2(n8940), .ZN(n7898) );
  OR2_X1 U7476 ( .A1(n7907), .A2(n8285), .ZN(n9083) );
  NAND2_X1 U7477 ( .A1(n7907), .A2(n8285), .ZN(n9079) );
  NAND2_X1 U7478 ( .A1(n9083), .A2(n9079), .ZN(n8873) );
  INV_X1 U7479 ( .A(n8943), .ZN(n6314) );
  INV_X1 U7480 ( .A(n9079), .ZN(n6313) );
  NOR2_X1 U7481 ( .A1(n6314), .A2(n6313), .ZN(n8938) );
  NAND2_X1 U7482 ( .A1(n8051), .A2(n8938), .ZN(n6315) );
  INV_X1 U7483 ( .A(n8874), .ZN(n6316) );
  INV_X1 U7484 ( .A(n8144), .ZN(n8876) );
  NAND2_X1 U7485 ( .A1(n8249), .A2(n8960), .ZN(n6317) );
  NOR2_X1 U7486 ( .A1(n10745), .A2(n10644), .ZN(n8957) );
  NAND2_X1 U7487 ( .A1(n10745), .A2(n10644), .ZN(n8961) );
  NAND2_X1 U7488 ( .A1(n10640), .A2(n9094), .ZN(n10623) );
  NAND2_X1 U7489 ( .A1(n10623), .A2(n10624), .ZN(n10622) );
  NAND2_X1 U7490 ( .A1(n10622), .A2(n8886), .ZN(n10614) );
  INV_X1 U7491 ( .A(n10605), .ZN(n10615) );
  NAND2_X1 U7492 ( .A1(n10614), .A2(n10615), .ZN(n10613) );
  INV_X1 U7493 ( .A(n8886), .ZN(n6318) );
  NAND2_X1 U7494 ( .A1(n8974), .A2(n6318), .ZN(n6319) );
  AND2_X1 U7495 ( .A1(n6319), .A2(n8975), .ZN(n8884) );
  INV_X1 U7496 ( .A(n8969), .ZN(n8981) );
  OR2_X1 U7497 ( .A1(n10579), .A2(n10551), .ZN(n8982) );
  NAND2_X1 U7498 ( .A1(n10579), .A2(n10551), .ZN(n8979) );
  NAND2_X1 U7499 ( .A1(n10563), .A2(n10566), .ZN(n10562) );
  NAND2_X1 U7500 ( .A1(n10556), .A2(n10693), .ZN(n9024) );
  NAND2_X1 U7501 ( .A1(n10532), .A2(n9024), .ZN(n10550) );
  INV_X1 U7502 ( .A(n10536), .ZN(n6320) );
  INV_X1 U7503 ( .A(n8992), .ZN(n6321) );
  OAI21_X1 U7504 ( .B1(n6322), .B2(n8998), .A(n6400), .ZN(n10484) );
  NAND2_X1 U7505 ( .A1(n10464), .A2(n6419), .ZN(n9015) );
  INV_X1 U7506 ( .A(n9120), .ZN(n6663) );
  NAND2_X1 U7507 ( .A1(n8860), .A2(n6663), .ZN(n6323) );
  INV_X1 U7508 ( .A(n7049), .ZN(n11139) );
  NAND2_X1 U7509 ( .A1(n7048), .A2(n11139), .ZN(n7356) );
  NAND2_X1 U7510 ( .A1(n10807), .A2(n10652), .ZN(n10653) );
  NAND2_X1 U7511 ( .A1(n10789), .A2(n10574), .ZN(n10554) );
  NOR2_X2 U7512 ( .A1(n10554), .A2(n10538), .ZN(n10514) );
  INV_X1 U7513 ( .A(n10501), .ZN(n6324) );
  AND2_X1 U7514 ( .A1(n6419), .A2(n8860), .ZN(n9040) );
  INV_X1 U7515 ( .A(n6326), .ZN(n8803) );
  INV_X1 U7516 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6672) );
  NOR2_X1 U7517 ( .A1(n6258), .A2(n6672), .ZN(n6330) );
  INV_X1 U7518 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U7519 ( .A1(n8848), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7520 ( .A1(n5960), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6327) );
  OAI211_X1 U7521 ( .C1(n6405), .C2(n6415), .A(n6328), .B(n6327), .ZN(n6329)
         );
  AOI21_X1 U7522 ( .B1(n8803), .B2(n6330), .A(n6329), .ZN(n10487) );
  OAI22_X1 U7523 ( .A1(n10685), .A2(n10763), .B1(n10487), .B2(n10741), .ZN(
        n6331) );
  INV_X1 U7524 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7525 ( .A1(n6336), .A2(n6332), .ZN(n6339) );
  NAND2_X1 U7526 ( .A1(n6339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6333) );
  MUX2_X1 U7527 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6333), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6335) );
  INV_X1 U7528 ( .A(n6336), .ZN(n6337) );
  NAND2_X1 U7529 ( .A1(n6337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6338) );
  MUX2_X1 U7530 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6338), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6340) );
  NAND2_X1 U7531 ( .A1(n6348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7532 ( .A1(n8269), .A2(P1_B_REG_SCAN_IN), .ZN(n6351) );
  INV_X1 U7533 ( .A(n8245), .ZN(n6350) );
  MUX2_X1 U7534 ( .A(n6351), .B(P1_B_REG_SCAN_IN), .S(n6350), .Z(n6352) );
  INV_X1 U7535 ( .A(n6352), .ZN(n6354) );
  NOR4_X1 U7536 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6363) );
  NOR4_X1 U7537 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6362) );
  OR4_X1 U7538 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6360) );
  NOR4_X1 U7539 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6358) );
  NOR4_X1 U7540 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6357) );
  NOR4_X1 U7541 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6356) );
  NOR4_X1 U7542 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6355) );
  NAND4_X1 U7543 ( .A1(n6358), .A2(n6357), .A3(n6356), .A4(n6355), .ZN(n6359)
         );
  NOR4_X1 U7544 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        n6360), .A4(n6359), .ZN(n6361) );
  NAND3_X1 U7545 ( .A1(n6363), .A2(n6362), .A3(n6361), .ZN(n6364) );
  NAND2_X1 U7546 ( .A1(n6365), .A2(n6364), .ZN(n6650) );
  NAND2_X1 U7547 ( .A1(n6420), .A2(n9040), .ZN(n6665) );
  NAND3_X1 U7548 ( .A1(n10813), .A2(n6650), .A3(n6665), .ZN(n6958) );
  NAND2_X1 U7549 ( .A1(n8308), .A2(n8269), .ZN(n10814) );
  OAI21_X1 U7550 ( .B1(n10812), .B2(P1_D_REG_1__SCAN_IN), .A(n10814), .ZN(
        n6649) );
  NAND2_X1 U7551 ( .A1(n11164), .A2(n9054), .ZN(n6657) );
  NAND2_X1 U7552 ( .A1(n6649), .A2(n6657), .ZN(n6366) );
  NAND2_X1 U7553 ( .A1(n8308), .A2(n8245), .ZN(n10815) );
  MUX2_X1 U7554 ( .A(n6367), .B(n6372), .S(n11185), .Z(n6370) );
  NAND2_X1 U7555 ( .A1(n6370), .A2(n6369), .ZN(P1_U3518) );
  INV_X1 U7556 ( .A(n6955), .ZN(n6651) );
  MUX2_X1 U7557 ( .A(n6373), .B(n6372), .S(n11181), .Z(n6375) );
  NAND2_X1 U7558 ( .A1(n6375), .A2(n6374), .ZN(P1_U3550) );
  NAND2_X1 U7559 ( .A1(n10493), .A2(n10676), .ZN(n6376) );
  AOI22_X2 U7560 ( .A1(n6377), .A2(n6376), .B1(n6680), .B2(n9938), .ZN(n6399)
         );
  INV_X1 U7561 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7562 ( .A1(n6379), .A2(n10137), .ZN(n6385) );
  INV_X1 U7563 ( .A(n6385), .ZN(n6383) );
  NOR2_X1 U7564 ( .A1(n6383), .A2(n6382), .ZN(n6388) );
  OR2_X1 U7565 ( .A1(n6384), .A2(n6388), .ZN(n6390) );
  AND2_X1 U7566 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  OR2_X1 U7567 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  MUX2_X1 U7568 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8701), .Z(n8407) );
  INV_X1 U7569 ( .A(n6392), .ZN(n6394) );
  INV_X1 U7570 ( .A(SI_29_), .ZN(n6393) );
  NAND2_X1 U7571 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  NAND2_X1 U7572 ( .A1(n8410), .A2(n6395), .ZN(n8841) );
  INV_X1 U7573 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8350) );
  OR2_X1 U7574 ( .A1(n8853), .A2(n8350), .ZN(n6397) );
  OR2_X1 U7575 ( .A1(n8809), .A2(n10487), .ZN(n9032) );
  NAND2_X1 U7576 ( .A1(n8809), .A2(n10487), .ZN(n9111) );
  NAND2_X1 U7577 ( .A1(n9032), .A2(n9111), .ZN(n9006) );
  INV_X1 U7578 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U7579 ( .A1(n8848), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U7580 ( .A1(n5960), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6403) );
  OAI211_X1 U7581 ( .C1(n6405), .C2(n10674), .A(n6404), .B(n6403), .ZN(n9937)
         );
  INV_X1 U7582 ( .A(n8349), .ZN(n6752) );
  NAND2_X1 U7583 ( .A1(n6752), .A2(P1_B_REG_SCAN_IN), .ZN(n6407) );
  AND2_X1 U7584 ( .A1(n11155), .A2(n6407), .ZN(n10474) );
  NAND2_X1 U7585 ( .A1(n9937), .A2(n10474), .ZN(n6408) );
  OAI211_X1 U7586 ( .C1(n5429), .C2(n5159), .A(n10672), .B(n10479), .ZN(n8806)
         );
  INV_X1 U7587 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6411) );
  NOR2_X1 U7588 ( .A1(n11185), .A2(n6411), .ZN(n6412) );
  NOR2_X1 U7589 ( .A1(n11181), .A2(n6415), .ZN(n6416) );
  NAND2_X1 U7590 ( .A1(n6418), .A2(n6417), .ZN(P1_U3551) );
  OR2_X1 U7591 ( .A1(n6420), .A2(n6419), .ZN(n6422) );
  OR2_X1 U7592 ( .A1(n6421), .A2(n6424), .ZN(n7005) );
  INV_X1 U7593 ( .A(n6424), .ZN(n6425) );
  AND2_X2 U7594 ( .A1(n6685), .A2(n6425), .ZN(n6444) );
  INV_X1 U7595 ( .A(n6685), .ZN(n6430) );
  NAND2_X1 U7596 ( .A1(n6430), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U7597 ( .A1(n6433), .A2(n6428), .ZN(n6839) );
  INV_X1 U7598 ( .A(n6429), .ZN(n6605) );
  NAND2_X1 U7599 ( .A1(n6426), .A2(n6605), .ZN(n6432) );
  AOI22_X1 U7600 ( .A1(n6964), .A2(n6444), .B1(n6430), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U7601 ( .A1(n6432), .A2(n6431), .ZN(n6838) );
  INV_X2 U7602 ( .A(n6624), .ZN(n6645) );
  NAND2_X1 U7603 ( .A1(n6434), .A2(n6444), .ZN(n6435) );
  NAND2_X1 U7604 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  XNOR2_X1 U7605 ( .A(n6437), .B(n6624), .ZN(n6441) );
  INV_X1 U7606 ( .A(n6441), .ZN(n6438) );
  NAND2_X1 U7607 ( .A1(n6434), .A2(n6605), .ZN(n6440) );
  OR2_X1 U7608 ( .A1(n5941), .A2(n6579), .ZN(n6439) );
  NAND2_X1 U7609 ( .A1(n6440), .A2(n6439), .ZN(n6898) );
  NAND2_X1 U7610 ( .A1(n6895), .A2(n6898), .ZN(n6443) );
  NAND2_X1 U7611 ( .A1(n6442), .A2(n6441), .ZN(n6896) );
  NAND2_X1 U7612 ( .A1(n6443), .A2(n6896), .ZN(n8831) );
  INV_X1 U7613 ( .A(n8831), .ZN(n6449) );
  XNOR2_X1 U7614 ( .A(n6445), .B(n6624), .ZN(n6450) );
  OR2_X1 U7615 ( .A1(n7014), .A2(n6644), .ZN(n6447) );
  NAND2_X1 U7616 ( .A1(n6869), .A2(n6444), .ZN(n6446) );
  NAND2_X1 U7617 ( .A1(n6447), .A2(n6446), .ZN(n6451) );
  XNOR2_X1 U7618 ( .A(n6450), .B(n6451), .ZN(n8834) );
  INV_X1 U7619 ( .A(n8834), .ZN(n6448) );
  INV_X1 U7620 ( .A(n6450), .ZN(n6453) );
  INV_X1 U7621 ( .A(n6451), .ZN(n6452) );
  NAND2_X1 U7622 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  OAI22_X1 U7623 ( .A1(n6997), .A2(n6579), .B1(n7034), .B2(n6455), .ZN(n6456)
         );
  XNOR2_X1 U7624 ( .A(n6456), .B(n6645), .ZN(n6461) );
  INV_X2 U7625 ( .A(n6605), .ZN(n6644) );
  OR2_X1 U7626 ( .A1(n6997), .A2(n6644), .ZN(n6458) );
  NAND2_X1 U7627 ( .A1(n6985), .A2(n6444), .ZN(n6457) );
  NAND2_X1 U7628 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  XNOR2_X1 U7629 ( .A(n6461), .B(n6459), .ZN(n6983) );
  INV_X1 U7630 ( .A(n6459), .ZN(n6460) );
  OAI22_X1 U7631 ( .A1(n7420), .A2(n6579), .B1(n7000), .B2(n6455), .ZN(n6462)
         );
  XNOR2_X1 U7632 ( .A(n6462), .B(n6645), .ZN(n6465) );
  OR2_X1 U7633 ( .A1(n7420), .A2(n6644), .ZN(n6464) );
  NAND2_X1 U7634 ( .A1(n5979), .A2(n6444), .ZN(n6463) );
  NAND2_X1 U7635 ( .A1(n6464), .A2(n6463), .ZN(n6466) );
  XNOR2_X1 U7636 ( .A(n6465), .B(n6466), .ZN(n9875) );
  INV_X1 U7637 ( .A(n6465), .ZN(n6467) );
  NAND2_X1 U7638 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  OAI22_X1 U7639 ( .A1(n9877), .A2(n6579), .B1(n11129), .B2(n6455), .ZN(n6469)
         );
  XNOR2_X1 U7640 ( .A(n6469), .B(n6645), .ZN(n6479) );
  OR2_X1 U7641 ( .A1(n9877), .A2(n6644), .ZN(n6471) );
  NAND2_X1 U7642 ( .A1(n7418), .A2(n6444), .ZN(n6470) );
  AND2_X1 U7643 ( .A1(n6471), .A2(n6470), .ZN(n7416) );
  OAI22_X1 U7644 ( .A1(n7042), .A2(n6579), .B1(n7064), .B2(n6455), .ZN(n6472)
         );
  XNOR2_X1 U7645 ( .A(n6472), .B(n6624), .ZN(n6476) );
  OR2_X1 U7646 ( .A1(n7042), .A2(n6644), .ZN(n6474) );
  NAND2_X1 U7647 ( .A1(n7405), .A2(n6444), .ZN(n6473) );
  NAND2_X1 U7648 ( .A1(n6474), .A2(n6473), .ZN(n7401) );
  NAND2_X1 U7649 ( .A1(n6476), .A2(n7401), .ZN(n6475) );
  OAI21_X1 U7650 ( .B1(n6479), .B2(n7416), .A(n6475), .ZN(n6482) );
  INV_X1 U7651 ( .A(n6479), .ZN(n7400) );
  INV_X1 U7652 ( .A(n7416), .ZN(n6477) );
  OAI21_X1 U7653 ( .B1(n7400), .B2(n6477), .A(n7401), .ZN(n6480) );
  INV_X1 U7654 ( .A(n6476), .ZN(n7402) );
  NOR2_X1 U7655 ( .A1(n6477), .A2(n7401), .ZN(n6478) );
  AOI22_X1 U7656 ( .A1(n6480), .A2(n7402), .B1(n6479), .B2(n6478), .ZN(n6481)
         );
  OR2_X1 U7657 ( .A1(n7353), .A2(n6644), .ZN(n6484) );
  NAND2_X1 U7658 ( .A1(n7049), .A2(n6444), .ZN(n6483) );
  AND2_X1 U7659 ( .A1(n6484), .A2(n6483), .ZN(n7437) );
  NAND2_X1 U7660 ( .A1(n7049), .A2(n6637), .ZN(n6485) );
  OAI21_X1 U7661 ( .B1(n7353), .B2(n6579), .A(n6485), .ZN(n6486) );
  XNOR2_X1 U7662 ( .A(n6486), .B(n6624), .ZN(n7438) );
  NAND2_X1 U7663 ( .A1(n8009), .A2(n6637), .ZN(n6488) );
  OR2_X1 U7664 ( .A1(n7868), .A2(n6579), .ZN(n6487) );
  NAND2_X1 U7665 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  XNOR2_X1 U7666 ( .A(n6489), .B(n6645), .ZN(n7858) );
  NAND2_X1 U7667 ( .A1(n8009), .A2(n6444), .ZN(n6491) );
  OR2_X1 U7668 ( .A1(n7868), .A2(n6644), .ZN(n6490) );
  AND2_X1 U7669 ( .A1(n6491), .A2(n6490), .ZN(n6497) );
  NAND2_X1 U7670 ( .A1(n7858), .A2(n6497), .ZN(n6492) );
  NAND2_X1 U7671 ( .A1(n7857), .A2(n6492), .ZN(n6501) );
  NAND2_X1 U7672 ( .A1(n7456), .A2(n6637), .ZN(n6494) );
  OR2_X1 U7673 ( .A1(n8002), .A2(n6579), .ZN(n6493) );
  NAND2_X1 U7674 ( .A1(n6494), .A2(n6493), .ZN(n6495) );
  XNOR2_X1 U7675 ( .A(n6495), .B(n6624), .ZN(n6502) );
  NOR2_X1 U7676 ( .A1(n8002), .A2(n6644), .ZN(n6496) );
  AOI21_X1 U7677 ( .B1(n7456), .B2(n6444), .A(n6496), .ZN(n6503) );
  XNOR2_X1 U7678 ( .A(n6502), .B(n6503), .ZN(n7862) );
  INV_X1 U7679 ( .A(n7858), .ZN(n6498) );
  INV_X1 U7680 ( .A(n6497), .ZN(n8005) );
  NAND2_X1 U7681 ( .A1(n6498), .A2(n8005), .ZN(n6499) );
  AND2_X1 U7682 ( .A1(n7862), .A2(n6499), .ZN(n6500) );
  INV_X1 U7683 ( .A(n6502), .ZN(n6504) );
  NAND2_X1 U7684 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  NAND2_X1 U7685 ( .A1(n7744), .A2(n6637), .ZN(n6507) );
  OR2_X1 U7686 ( .A1(n7515), .A2(n6579), .ZN(n6506) );
  NAND2_X1 U7687 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  XNOR2_X1 U7688 ( .A(n6508), .B(n6645), .ZN(n6510) );
  NOR2_X1 U7689 ( .A1(n7515), .A2(n6644), .ZN(n6509) );
  AOI21_X1 U7690 ( .B1(n7744), .B2(n6444), .A(n6509), .ZN(n7736) );
  NAND2_X1 U7691 ( .A1(n7735), .A2(n7736), .ZN(n6512) );
  NAND2_X1 U7692 ( .A1(n6511), .A2(n6510), .ZN(n7734) );
  OAI22_X1 U7693 ( .A1(n11160), .A2(n6455), .B1(n10349), .B2(n6579), .ZN(n6513) );
  XNOR2_X1 U7694 ( .A(n6513), .B(n6645), .ZN(n6516) );
  OR2_X1 U7695 ( .A1(n11160), .A2(n6579), .ZN(n6515) );
  OR2_X1 U7696 ( .A1(n10349), .A2(n6644), .ZN(n6514) );
  AND2_X1 U7697 ( .A1(n6515), .A2(n6514), .ZN(n6517) );
  INV_X1 U7698 ( .A(n6516), .ZN(n6519) );
  INV_X1 U7699 ( .A(n6517), .ZN(n6518) );
  NAND2_X1 U7700 ( .A1(n6519), .A2(n6518), .ZN(n7813) );
  NAND2_X1 U7701 ( .A1(n7671), .A2(n6637), .ZN(n6521) );
  NAND2_X1 U7702 ( .A1(n11154), .A2(n6444), .ZN(n6520) );
  NAND2_X1 U7703 ( .A1(n6521), .A2(n6520), .ZN(n6522) );
  XNOR2_X1 U7704 ( .A(n6522), .B(n6624), .ZN(n6524) );
  AND2_X1 U7705 ( .A1(n11154), .A2(n6605), .ZN(n6523) );
  AOI21_X1 U7706 ( .B1(n7671), .B2(n6444), .A(n6523), .ZN(n6525) );
  XNOR2_X1 U7707 ( .A(n6524), .B(n6525), .ZN(n8068) );
  INV_X1 U7708 ( .A(n6524), .ZN(n6526) );
  NAND2_X1 U7709 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  NAND2_X1 U7710 ( .A1(n7907), .A2(n6637), .ZN(n6529) );
  NAND2_X1 U7711 ( .A1(n10348), .A2(n6444), .ZN(n6528) );
  NAND2_X1 U7712 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  XNOR2_X1 U7713 ( .A(n6530), .B(n6624), .ZN(n6534) );
  AND2_X1 U7714 ( .A1(n10348), .A2(n6605), .ZN(n6531) );
  AOI21_X1 U7715 ( .B1(n7907), .B2(n6444), .A(n6531), .ZN(n6532) );
  XNOR2_X1 U7716 ( .A(n6534), .B(n6532), .ZN(n8151) );
  INV_X1 U7717 ( .A(n6532), .ZN(n6533) );
  NAND2_X1 U7718 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  NAND2_X1 U7719 ( .A1(n6540), .A2(n6637), .ZN(n6537) );
  OR2_X1 U7720 ( .A1(n10764), .A2(n6579), .ZN(n6536) );
  NAND2_X1 U7721 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  XNOR2_X1 U7722 ( .A(n6538), .B(n6645), .ZN(n6542) );
  NOR2_X1 U7723 ( .A1(n10764), .A2(n6644), .ZN(n6539) );
  AOI21_X1 U7724 ( .B1(n6540), .B2(n6444), .A(n6539), .ZN(n8282) );
  INV_X1 U7725 ( .A(n6541), .ZN(n6543) );
  NAND2_X1 U7726 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  OAI22_X1 U7727 ( .A1(n6546), .A2(n6455), .B1(n10756), .B2(n6579), .ZN(n6545)
         );
  XNOR2_X1 U7728 ( .A(n6545), .B(n6645), .ZN(n6547) );
  OAI22_X1 U7729 ( .A1(n6546), .A2(n6579), .B1(n10756), .B2(n6644), .ZN(n8338)
         );
  INV_X1 U7730 ( .A(n6547), .ZN(n6548) );
  NAND2_X1 U7731 ( .A1(n10759), .A2(n6637), .ZN(n6550) );
  OR2_X1 U7732 ( .A1(n9857), .A2(n6579), .ZN(n6549) );
  NAND2_X1 U7733 ( .A1(n6550), .A2(n6549), .ZN(n6551) );
  XNOR2_X1 U7734 ( .A(n6551), .B(n6645), .ZN(n6555) );
  NOR2_X1 U7735 ( .A1(n9857), .A2(n6644), .ZN(n6552) );
  AOI21_X1 U7736 ( .B1(n10759), .B2(n6444), .A(n6552), .ZN(n6554) );
  XNOR2_X1 U7737 ( .A(n6555), .B(n6554), .ZN(n9844) );
  INV_X1 U7738 ( .A(n9844), .ZN(n6553) );
  NAND2_X1 U7739 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  NAND2_X1 U7740 ( .A1(n9841), .A2(n6556), .ZN(n9853) );
  NAND2_X1 U7741 ( .A1(n10753), .A2(n6637), .ZN(n6558) );
  OR2_X1 U7742 ( .A1(n10740), .A2(n6579), .ZN(n6557) );
  NAND2_X1 U7743 ( .A1(n6558), .A2(n6557), .ZN(n6559) );
  XNOR2_X1 U7744 ( .A(n6559), .B(n6624), .ZN(n6561) );
  NOR2_X1 U7745 ( .A1(n10740), .A2(n6644), .ZN(n6560) );
  AOI21_X1 U7746 ( .B1(n10753), .B2(n6444), .A(n6560), .ZN(n6562) );
  XNOR2_X1 U7747 ( .A(n6561), .B(n6562), .ZN(n9854) );
  INV_X1 U7748 ( .A(n6561), .ZN(n6563) );
  NAND2_X1 U7749 ( .A1(n6563), .A2(n6562), .ZN(n6564) );
  OAI22_X1 U7750 ( .A1(n9913), .A2(n6455), .B1(n10644), .B2(n6579), .ZN(n6565)
         );
  XNOR2_X1 U7751 ( .A(n6565), .B(n6645), .ZN(n9908) );
  OR2_X1 U7752 ( .A1(n9913), .A2(n6579), .ZN(n6567) );
  OR2_X1 U7753 ( .A1(n10644), .A2(n6644), .ZN(n6566) );
  AND2_X1 U7754 ( .A1(n6567), .A2(n6566), .ZN(n9907) );
  NAND2_X1 U7755 ( .A1(n10657), .A2(n6637), .ZN(n6569) );
  INV_X1 U7756 ( .A(n10742), .ZN(n10343) );
  NAND2_X1 U7757 ( .A1(n10343), .A2(n6444), .ZN(n6568) );
  NAND2_X1 U7758 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  XNOR2_X1 U7759 ( .A(n6570), .B(n6624), .ZN(n6592) );
  NOR2_X1 U7760 ( .A1(n10742), .A2(n6644), .ZN(n6571) );
  AOI21_X1 U7761 ( .B1(n10657), .B2(n6444), .A(n6571), .ZN(n6593) );
  XNOR2_X1 U7762 ( .A(n6592), .B(n6593), .ZN(n9884) );
  NAND2_X1 U7763 ( .A1(n10631), .A2(n6637), .ZN(n6573) );
  OR2_X1 U7764 ( .A1(n10645), .A2(n6579), .ZN(n6572) );
  NAND2_X1 U7765 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  XNOR2_X1 U7766 ( .A(n6574), .B(n6624), .ZN(n6596) );
  NOR2_X1 U7767 ( .A1(n10645), .A2(n6644), .ZN(n6575) );
  AOI21_X1 U7768 ( .B1(n10631), .B2(n6444), .A(n6575), .ZN(n6597) );
  XNOR2_X1 U7769 ( .A(n6596), .B(n6597), .ZN(n9888) );
  AND2_X1 U7770 ( .A1(n9884), .A2(n9888), .ZN(n6606) );
  NAND2_X1 U7771 ( .A1(n10595), .A2(n6637), .ZN(n6577) );
  OR2_X1 U7772 ( .A1(n9812), .A2(n6579), .ZN(n6576) );
  NAND2_X1 U7773 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  XNOR2_X1 U7774 ( .A(n6578), .B(n6645), .ZN(n6608) );
  NAND2_X1 U7775 ( .A1(n10725), .A2(n6637), .ZN(n6581) );
  OR2_X1 U7776 ( .A1(n10626), .A2(n6579), .ZN(n6580) );
  NAND2_X1 U7777 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  XNOR2_X1 U7778 ( .A(n6582), .B(n6624), .ZN(n6587) );
  NAND2_X1 U7779 ( .A1(n10725), .A2(n6444), .ZN(n6584) );
  OR2_X1 U7780 ( .A1(n10626), .A2(n6644), .ZN(n6583) );
  NAND2_X1 U7781 ( .A1(n6584), .A2(n6583), .ZN(n6588) );
  NAND2_X1 U7782 ( .A1(n6587), .A2(n6588), .ZN(n6609) );
  AND2_X1 U7783 ( .A1(n6608), .A2(n6609), .ZN(n6586) );
  AND2_X1 U7784 ( .A1(n6606), .A2(n6586), .ZN(n6585) );
  NAND2_X1 U7785 ( .A1(n9817), .A2(n6585), .ZN(n6604) );
  INV_X1 U7786 ( .A(n6586), .ZN(n6602) );
  INV_X1 U7787 ( .A(n6587), .ZN(n6590) );
  INV_X1 U7788 ( .A(n6588), .ZN(n6589) );
  NAND2_X1 U7789 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  NAND2_X1 U7790 ( .A1(n6609), .A2(n6591), .ZN(n9829) );
  INV_X1 U7791 ( .A(n9829), .ZN(n6601) );
  INV_X1 U7792 ( .A(n9888), .ZN(n6595) );
  INV_X1 U7793 ( .A(n6592), .ZN(n6594) );
  NAND2_X1 U7794 ( .A1(n6594), .A2(n6593), .ZN(n9885) );
  OR2_X1 U7795 ( .A1(n6595), .A2(n9885), .ZN(n6600) );
  INV_X1 U7796 ( .A(n6596), .ZN(n6598) );
  NAND2_X1 U7797 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  AND2_X1 U7798 ( .A1(n6600), .A2(n6599), .ZN(n9825) );
  AND2_X1 U7799 ( .A1(n6601), .A2(n9825), .ZN(n6607) );
  OR2_X1 U7800 ( .A1(n6602), .A2(n6607), .ZN(n6603) );
  NAND2_X1 U7801 ( .A1(n6604), .A2(n6603), .ZN(n9894) );
  AOI22_X1 U7802 ( .A1(n10595), .A2(n6444), .B1(n6605), .B2(n10709), .ZN(n9896) );
  NOR2_X1 U7803 ( .A1(n9894), .A2(n9896), .ZN(n9897) );
  AOI21_X1 U7804 ( .B1(n9827), .B2(n6609), .A(n6608), .ZN(n9895) );
  AOI22_X1 U7805 ( .A1(n10579), .A2(n6637), .B1(n6444), .B2(n10590), .ZN(n6610) );
  XNOR2_X1 U7806 ( .A(n6610), .B(n6624), .ZN(n6611) );
  OAI22_X1 U7807 ( .A1(n10793), .A2(n6579), .B1(n10551), .B2(n6644), .ZN(n6612) );
  XNOR2_X1 U7808 ( .A(n6611), .B(n6612), .ZN(n9809) );
  NAND2_X1 U7809 ( .A1(n6611), .A2(n6613), .ZN(n6614) );
  NAND2_X1 U7810 ( .A1(n10556), .A2(n6637), .ZN(n6616) );
  NAND2_X1 U7811 ( .A1(n10710), .A2(n6444), .ZN(n6615) );
  NAND2_X1 U7812 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  XNOR2_X1 U7813 ( .A(n6617), .B(n6624), .ZN(n6621) );
  NAND2_X1 U7814 ( .A1(n10556), .A2(n6444), .ZN(n6619) );
  NAND2_X1 U7815 ( .A1(n10710), .A2(n6605), .ZN(n6618) );
  NAND2_X1 U7816 ( .A1(n6619), .A2(n6618), .ZN(n6620) );
  NAND2_X1 U7817 ( .A1(n6621), .A2(n6620), .ZN(n9863) );
  NAND2_X1 U7818 ( .A1(n10538), .A2(n6637), .ZN(n6623) );
  NAND2_X1 U7819 ( .A1(n10520), .A2(n6444), .ZN(n6622) );
  NAND2_X1 U7820 ( .A1(n6623), .A2(n6622), .ZN(n6625) );
  XNOR2_X1 U7821 ( .A(n6625), .B(n6624), .ZN(n6631) );
  OAI22_X1 U7822 ( .A1(n10785), .A2(n6579), .B1(n10684), .B2(n6644), .ZN(n6630) );
  XNOR2_X1 U7823 ( .A(n6631), .B(n6630), .ZN(n9834) );
  NAND2_X1 U7824 ( .A1(n10688), .A2(n6637), .ZN(n6627) );
  NAND2_X1 U7825 ( .A1(n10503), .A2(n6444), .ZN(n6626) );
  NAND2_X1 U7826 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  XNOR2_X1 U7827 ( .A(n6628), .B(n6645), .ZN(n6633) );
  NOR2_X1 U7828 ( .A1(n10694), .A2(n6644), .ZN(n6629) );
  AOI21_X1 U7829 ( .B1(n10688), .B2(n6444), .A(n6629), .ZN(n6634) );
  XNOR2_X1 U7830 ( .A(n6633), .B(n6634), .ZN(n9922) );
  NOR2_X1 U7831 ( .A1(n6631), .A2(n6630), .ZN(n9923) );
  INV_X1 U7832 ( .A(n6633), .ZN(n6636) );
  INV_X1 U7833 ( .A(n6634), .ZN(n6635) );
  NAND2_X1 U7834 ( .A1(n10679), .A2(n6637), .ZN(n6639) );
  NAND2_X1 U7835 ( .A1(n9933), .A2(n6444), .ZN(n6638) );
  NAND2_X1 U7836 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  XNOR2_X1 U7837 ( .A(n6640), .B(n6645), .ZN(n6643) );
  NOR2_X1 U7838 ( .A1(n10685), .A2(n6644), .ZN(n6641) );
  AOI21_X1 U7839 ( .B1(n10679), .B2(n6444), .A(n6641), .ZN(n6642) );
  NAND2_X1 U7840 ( .A1(n6643), .A2(n6642), .ZN(n6676) );
  OAI21_X1 U7841 ( .B1(n6643), .B2(n6642), .A(n6676), .ZN(n9174) );
  OAI22_X1 U7842 ( .A1(n10493), .A2(n6579), .B1(n10676), .B2(n6644), .ZN(n6646) );
  XNOR2_X1 U7843 ( .A(n6646), .B(n6645), .ZN(n6648) );
  OAI22_X1 U7844 ( .A1(n10493), .A2(n6455), .B1(n10676), .B2(n6579), .ZN(n6647) );
  XNOR2_X1 U7845 ( .A(n6648), .B(n6647), .ZN(n6654) );
  INV_X1 U7846 ( .A(n6654), .ZN(n6677) );
  INV_X1 U7847 ( .A(n6649), .ZN(n6956) );
  NAND3_X1 U7848 ( .A1(n6651), .A2(n6956), .A3(n6650), .ZN(n6670) );
  INV_X1 U7849 ( .A(n10813), .ZN(n6652) );
  NOR2_X1 U7850 ( .A1(n6670), .A2(n6652), .ZN(n6656) );
  NOR2_X1 U7851 ( .A1(n11127), .A2(n9040), .ZN(n6662) );
  NAND3_X1 U7852 ( .A1(n6677), .A2(n9926), .A3(n6676), .ZN(n6653) );
  NAND3_X1 U7853 ( .A1(n9177), .A2(n6654), .A3(n9926), .ZN(n6682) );
  AND2_X1 U7854 ( .A1(n6655), .A2(n6663), .ZN(n6963) );
  NAND2_X1 U7855 ( .A1(n6656), .A2(n6963), .ZN(n6659) );
  INV_X1 U7856 ( .A(n6657), .ZN(n6658) );
  INV_X1 U7857 ( .A(n10491), .ZN(n6675) );
  INV_X1 U7858 ( .A(n6660), .ZN(n6661) );
  NAND2_X1 U7859 ( .A1(n10813), .A2(n6661), .ZN(n9125) );
  INV_X1 U7860 ( .A(n6662), .ZN(n6664) );
  NAND2_X1 U7861 ( .A1(n6663), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7729) );
  NAND3_X1 U7862 ( .A1(n9125), .A2(n6664), .A3(n7729), .ZN(n6667) );
  INV_X1 U7863 ( .A(n6665), .ZN(n6666) );
  AOI21_X1 U7864 ( .B1(n6670), .B2(n6667), .A(n6666), .ZN(n6840) );
  NAND2_X1 U7865 ( .A1(n6840), .A2(n6668), .ZN(n6669) );
  NOR2_X1 U7866 ( .A1(n6670), .A2(n9125), .ZN(n6671) );
  NAND2_X1 U7867 ( .A1(n6671), .A2(n6917), .ZN(n9912) );
  OAI22_X1 U7868 ( .A1(n10487), .A2(n9878), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6672), .ZN(n6673) );
  AOI21_X1 U7869 ( .B1(n9928), .B2(n9933), .A(n6673), .ZN(n6674) );
  OAI21_X1 U7870 ( .B1(n6675), .B2(n9930), .A(n6674), .ZN(n6679) );
  NOR3_X1 U7871 ( .A1(n6677), .A2(n9919), .A3(n6676), .ZN(n6678) );
  AOI211_X1 U7872 ( .C1(n6680), .C2(n9904), .A(n6679), .B(n6678), .ZN(n6681)
         );
  NAND3_X1 U7873 ( .A1(n6683), .A2(n6682), .A3(n6681), .ZN(P1_U3220) );
  INV_X1 U7874 ( .A(n8128), .ZN(n6684) );
  NOR3_X1 U7875 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n6691) );
  NOR2_X1 U7876 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6690) );
  NOR2_X1 U7877 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6689) );
  AND2_X2 U7878 ( .A1(n6692), .A2(n6832), .ZN(n6693) );
  INV_X1 U7879 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U7880 ( .A1(n6698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U7881 ( .A1(n6700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U7882 ( .A1(n5228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6703) );
  INV_X2 U7883 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7884 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6710) );
  INV_X1 U7885 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6704) );
  XNOR2_X1 U7886 ( .A(n6784), .B(n6704), .ZN(n6709) );
  INV_X1 U7887 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6959) );
  INV_X1 U7888 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6712) );
  NOR3_X1 U7889 ( .A1(n6709), .A2(n6959), .A3(n6712), .ZN(n6793) );
  NOR2_X1 U7890 ( .A1(n6705), .A2(P1_U3086), .ZN(n6716) );
  NAND2_X1 U7891 ( .A1(n8128), .A2(n9040), .ZN(n6706) );
  NAND2_X1 U7892 ( .A1(n6707), .A2(n6706), .ZN(n6715) );
  INV_X1 U7893 ( .A(n6715), .ZN(n6708) );
  NAND2_X1 U7894 ( .A1(n6716), .A2(n6708), .ZN(n6755) );
  OR2_X1 U7895 ( .A1(n5139), .A2(n8349), .ZN(n9124) );
  AOI211_X1 U7896 ( .C1(n6710), .C2(n6709), .A(n6793), .B(n10952), .ZN(n6722)
         );
  NAND2_X1 U7897 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6714) );
  INV_X1 U7898 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6711) );
  XNOR2_X1 U7899 ( .A(n6784), .B(n6711), .ZN(n6713) );
  INV_X1 U7900 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6829) );
  NOR3_X1 U7901 ( .A1(n6713), .A2(n6829), .A3(n6712), .ZN(n6785) );
  AOI211_X1 U7902 ( .C1(n6714), .C2(n6713), .A(n6785), .B(n10956), .ZN(n6721)
         );
  NOR2_X1 U7903 ( .A1(n10374), .A2(n6784), .ZN(n6720) );
  INV_X1 U7904 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6718) );
  INV_X1 U7905 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6717) );
  OAI22_X1 U7906 ( .A1(n10967), .A2(n6718), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6717), .ZN(n6719) );
  OR4_X1 U7907 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(P1_U3244)
         );
  NAND2_X1 U7908 ( .A1(n8701), .A2(P1_U3086), .ZN(n9220) );
  NOR2_X1 U7909 ( .A1(n8701), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10820) );
  INV_X2 U7910 ( .A(n10820), .ZN(n9222) );
  OAI222_X1 U7911 ( .A1(n9220), .A2(n5759), .B1(n9222), .B2(n6739), .C1(
        P1_U3086), .C2(n6784), .ZN(P1_U3354) );
  OAI222_X1 U7912 ( .A1(n9220), .A2(n6723), .B1(n9222), .B2(n7316), .C1(
        P1_U3086), .C2(n10358), .ZN(P1_U3352) );
  OAI222_X1 U7913 ( .A1(P1_U3086), .A2(n10373), .B1(n9222), .B2(n7527), .C1(
        n6724), .C2(n9220), .ZN(P1_U3351) );
  INV_X1 U7914 ( .A(n7533), .ZN(n6728) );
  OAI222_X1 U7915 ( .A1(P1_U3086), .A2(n6801), .B1(n9222), .B2(n6728), .C1(
        n6725), .C2(n9220), .ZN(P1_U3350) );
  NOR2_X2 U7916 ( .A1(n8701), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9802) );
  INV_X1 U7917 ( .A(n9802), .ZN(n8844) );
  INV_X1 U7918 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U7919 ( .A1(n6726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6727) );
  INV_X1 U7920 ( .A(n7535), .ZN(n11046) );
  NAND2_X1 U7921 ( .A1(n8701), .A2(P2_U3151), .ZN(n9800) );
  OAI222_X1 U7922 ( .A1(n8844), .A2(n6729), .B1(n11046), .B2(P2_U3151), .C1(
        n9800), .C2(n6728), .ZN(P2_U3290) );
  INV_X1 U7923 ( .A(n9220), .ZN(n7068) );
  AOI22_X1 U7924 ( .A1(n6852), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7068), .ZN(n6730) );
  OAI21_X1 U7925 ( .B1(n7578), .B2(n9222), .A(n6730), .ZN(P1_U3349) );
  OAI222_X1 U7926 ( .A1(n9220), .A2(n6731), .B1(n9222), .B2(n8842), .C1(
        P1_U3086), .C2(n6931), .ZN(P1_U3353) );
  INV_X1 U7927 ( .A(n9800), .ZN(n8329) );
  INV_X1 U7928 ( .A(n8329), .ZN(n9804) );
  NAND2_X1 U7929 ( .A1(n6732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7930 ( .A1(n11016), .A2(P2_STATE_REG_SCAN_IN), .B1(n9802), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n6733) );
  OAI21_X1 U7931 ( .B1(n7316), .B2(n9804), .A(n6733), .ZN(P2_U3292) );
  OR2_X1 U7932 ( .A1(n6734), .A2(n7131), .ZN(n6748) );
  XNOR2_X1 U7933 ( .A(n6748), .B(n6747), .ZN(n11061) );
  INV_X1 U7934 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6735) );
  OAI222_X1 U7935 ( .A1(n9804), .A2(n7578), .B1(n11061), .B2(P2_U3151), .C1(
        n6735), .C2(n8844), .ZN(P2_U3289) );
  INV_X1 U7936 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6740) );
  MUX2_X1 U7937 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6736), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6738) );
  INV_X1 U7938 ( .A(n7132), .ZN(n6737) );
  NAND2_X1 U7939 ( .A1(n6738), .A2(n6737), .ZN(n7234) );
  OAI222_X1 U7940 ( .A1(n8844), .A2(n6740), .B1(n7234), .B2(P2_U3151), .C1(
        n9804), .C2(n6739), .ZN(P2_U3294) );
  INV_X1 U7941 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6745) );
  INV_X1 U7942 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U7943 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  NAND2_X1 U7944 ( .A1(n6743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6744) );
  XNOR2_X1 U7945 ( .A(n6744), .B(P2_IR_REG_4__SCAN_IN), .ZN(n11034) );
  OAI222_X1 U7946 ( .A1(n8844), .A2(n6745), .B1(n7243), .B2(P2_U3151), .C1(
        n9804), .C2(n7527), .ZN(P2_U3291) );
  AOI22_X1 U7947 ( .A1(n6909), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7068), .ZN(n6746) );
  OAI21_X1 U7948 ( .B1(n7750), .B2(n9222), .A(n6746), .ZN(P1_U3348) );
  NAND2_X1 U7949 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  NAND2_X1 U7950 ( .A1(n6749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6758) );
  XNOR2_X1 U7951 ( .A(n6758), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7747) );
  INV_X1 U7952 ( .A(n7747), .ZN(n7227) );
  INV_X1 U7953 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6750) );
  OAI222_X1 U7954 ( .A1(n9804), .A2(n7750), .B1(n7227), .B2(P2_U3151), .C1(
        n6750), .C2(n8844), .ZN(P2_U3288) );
  INV_X1 U7955 ( .A(n7825), .ZN(n6761) );
  AOI22_X1 U7956 ( .A1(n7638), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7068), .ZN(n6751) );
  OAI21_X1 U7957 ( .B1(n6761), .B2(n9222), .A(n6751), .ZN(P1_U3347) );
  OR2_X1 U7958 ( .A1(n5139), .A2(n6752), .ZN(n6923) );
  OAI22_X1 U7959 ( .A1(n6829), .A2(n6923), .B1(n9124), .B2(n6959), .ZN(n6753)
         );
  XNOR2_X1 U7960 ( .A(n6753), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6756) );
  INV_X1 U7961 ( .A(n10967), .ZN(n10396) );
  AOI22_X1 U7962 ( .A1(n10396), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6754) );
  OAI21_X1 U7963 ( .B1(n6756), .B2(n6755), .A(n6754), .ZN(P1_U3243) );
  INV_X1 U7964 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6762) );
  INV_X1 U7965 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U7966 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NAND2_X1 U7967 ( .A1(n6759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6760) );
  XNOR2_X1 U7968 ( .A(n6760), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7824) );
  OAI222_X1 U7969 ( .A1(n8844), .A2(n6762), .B1(n9800), .B2(n6761), .C1(
        P2_U3151), .C2(n7771), .ZN(P2_U3287) );
  INV_X1 U7970 ( .A(n8097), .ZN(n7295) );
  INV_X1 U7971 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6769) );
  INV_X1 U7972 ( .A(n8828), .ZN(n6764) );
  NAND2_X1 U7973 ( .A1(n7172), .A2(n6769), .ZN(n6767) );
  OR2_X1 U7974 ( .A1(n7173), .A2(n8828), .ZN(n6766) );
  INV_X1 U7975 ( .A(n7678), .ZN(n7177) );
  NAND2_X1 U7976 ( .A1(n7177), .A2(n7318), .ZN(n6768) );
  OAI21_X1 U7977 ( .B1(n7318), .B2(n6769), .A(n6768), .ZN(P2_U3377) );
  INV_X1 U7978 ( .A(n7934), .ZN(n6776) );
  AOI22_X1 U7979 ( .A1(n10397), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7068), .ZN(n6770) );
  OAI21_X1 U7980 ( .B1(n6776), .B2(n9222), .A(n6770), .ZN(P1_U3346) );
  OR2_X1 U7981 ( .A1(n6833), .A2(n7131), .ZN(n6771) );
  XNOR2_X1 U7982 ( .A(n6771), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8028) );
  INV_X1 U7983 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6772) );
  OAI222_X1 U7984 ( .A1(n9804), .A2(n8027), .B1(n8211), .B2(P2_U3151), .C1(
        n6772), .C2(n8844), .ZN(P2_U3285) );
  INV_X1 U7985 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6822) );
  OR2_X1 U7986 ( .A1(n6773), .A2(n7131), .ZN(n6774) );
  XNOR2_X1 U7987 ( .A(n6774), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7989) );
  INV_X1 U7988 ( .A(n7989), .ZN(n6775) );
  OAI222_X1 U7989 ( .A1(n9804), .A2(n6776), .B1(n8844), .B2(n6822), .C1(
        P2_U3151), .C2(n6775), .ZN(P2_U3286) );
  INV_X1 U7990 ( .A(n10963), .ZN(n7640) );
  INV_X1 U7991 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6777) );
  OAI222_X1 U7992 ( .A1(P1_U3086), .A2(n7640), .B1(n9222), .B2(n8027), .C1(
        n6777), .C2(n9220), .ZN(P1_U3345) );
  INV_X1 U7993 ( .A(n7172), .ZN(n6778) );
  INV_X1 U7994 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6782) );
  INV_X1 U7995 ( .A(n6779), .ZN(n6780) );
  NOR3_X1 U7996 ( .A1(n7173), .A2(n6763), .A3(n6780), .ZN(n6781) );
  AOI21_X1 U7997 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(P2_U3376) );
  AND2_X1 U7998 ( .A1(n6783), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7999 ( .A1(n6783), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8000 ( .A1(n6783), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8001 ( .A1(n6783), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8002 ( .A1(n6783), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8003 ( .A1(n6783), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8004 ( .A1(n6783), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8005 ( .A1(n6783), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8006 ( .A1(n6783), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8007 ( .A1(n6783), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8008 ( .A1(n6783), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8009 ( .A1(n6783), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8010 ( .A1(n6783), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8011 ( .A1(n6783), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8012 ( .A1(n6783), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8013 ( .A1(n6783), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8014 ( .A1(n6783), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8015 ( .A1(n6783), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8016 ( .A1(n6783), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8017 ( .A1(n6783), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8018 ( .A1(n6783), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8019 ( .A1(n6783), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8020 ( .A1(n6783), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8021 ( .A1(n6783), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8022 ( .A1(n6783), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8023 ( .A1(n6783), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8024 ( .A1(n6783), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8025 ( .A1(n6783), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8026 ( .A1(n6783), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8027 ( .A1(n6783), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U8028 ( .A(n10373), .ZN(n6800) );
  INV_X1 U8029 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6788) );
  INV_X1 U8030 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6787) );
  INV_X1 U8031 ( .A(n6784), .ZN(n6794) );
  AOI21_X1 U8032 ( .B1(n6794), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6785), .ZN(
        n6926) );
  XOR2_X1 U8033 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6931), .Z(n6925) );
  NOR2_X1 U8034 ( .A1(n6926), .A2(n6925), .ZN(n6924) );
  INV_X1 U8035 ( .A(n6924), .ZN(n6786) );
  OAI21_X1 U8036 ( .B1(n6931), .B2(n6787), .A(n6786), .ZN(n10364) );
  XNOR2_X1 U8037 ( .A(n10358), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U8038 ( .A1(n10364), .A2(n10365), .ZN(n10363) );
  OAI21_X1 U8039 ( .B1(n10358), .B2(n6788), .A(n10363), .ZN(n10381) );
  INV_X1 U8040 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6789) );
  MUX2_X1 U8041 ( .A(n6789), .B(P1_REG1_REG_4__SCAN_IN), .S(n10373), .Z(n10382) );
  NAND2_X1 U8042 ( .A1(n10381), .A2(n10382), .ZN(n10380) );
  INV_X1 U8043 ( .A(n10380), .ZN(n6790) );
  AOI21_X1 U8044 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6800), .A(n6790), .ZN(
        n6792) );
  XOR2_X1 U8045 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6801), .Z(n6791) );
  NOR2_X1 U8046 ( .A1(n6792), .A2(n6791), .ZN(n6809) );
  AOI211_X1 U8047 ( .C1(n6792), .C2(n6791), .A(n10956), .B(n6809), .ZN(n6808)
         );
  INV_X1 U8048 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6797) );
  INV_X1 U8049 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6796) );
  XOR2_X1 U8050 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6931), .Z(n6928) );
  NOR2_X1 U8051 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  INV_X1 U8052 ( .A(n6927), .ZN(n6795) );
  OAI21_X1 U8053 ( .B1(n6931), .B2(n6796), .A(n6795), .ZN(n10367) );
  XNOR2_X1 U8054 ( .A(n10358), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U8055 ( .A1(n10367), .A2(n10368), .ZN(n10366) );
  OAI21_X1 U8056 ( .B1(n10358), .B2(n6797), .A(n10366), .ZN(n10378) );
  INV_X1 U8057 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6798) );
  MUX2_X1 U8058 ( .A(n6798), .B(P1_REG2_REG_4__SCAN_IN), .S(n10373), .Z(n10379) );
  NAND2_X1 U8059 ( .A1(n10378), .A2(n10379), .ZN(n10377) );
  INV_X1 U8060 ( .A(n10377), .ZN(n6799) );
  INV_X1 U8061 ( .A(n6801), .ZN(n6813) );
  XNOR2_X1 U8062 ( .A(n6813), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6802) );
  NOR2_X1 U8063 ( .A1(n6803), .A2(n6802), .ZN(n6812) );
  AOI211_X1 U8064 ( .C1(n6803), .C2(n6802), .A(n10952), .B(n6812), .ZN(n6807)
         );
  INV_X1 U8065 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8066 ( .A1(n10962), .A2(n6813), .ZN(n6804) );
  NAND2_X1 U8067 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7419) );
  OAI211_X1 U8068 ( .C1(n6805), .C2(n10967), .A(n6804), .B(n7419), .ZN(n6806)
         );
  OR3_X1 U8069 ( .A1(n6808), .A2(n6807), .A3(n6806), .ZN(P1_U3248) );
  AOI21_X1 U8070 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6813), .A(n6809), .ZN(
        n6811) );
  XNOR2_X1 U8071 ( .A(n6852), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U8072 ( .A1(n6811), .A2(n6810), .ZN(n6851) );
  AOI211_X1 U8073 ( .C1(n6811), .C2(n6810), .A(n10956), .B(n6851), .ZN(n6820)
         );
  AOI21_X1 U8074 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6813), .A(n6812), .ZN(
        n6815) );
  XNOR2_X1 U8075 ( .A(n6852), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6814) );
  NOR2_X1 U8076 ( .A1(n6815), .A2(n6814), .ZN(n6848) );
  AOI211_X1 U8077 ( .C1(n6815), .C2(n6814), .A(n10952), .B(n6848), .ZN(n6819)
         );
  INV_X1 U8078 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8079 ( .A1(n10962), .A2(n6852), .ZN(n6816) );
  NAND2_X1 U8080 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7406) );
  OAI211_X1 U8081 ( .C1(n6817), .C2(n10967), .A(n6816), .B(n7406), .ZN(n6818)
         );
  OR3_X1 U8082 ( .A1(n6820), .A2(n6819), .A3(n6818), .ZN(P1_U3249) );
  NOR2_X1 U8083 ( .A1(n10396), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8084 ( .A1(n7739), .A2(P1_U3973), .ZN(n6821) );
  OAI21_X1 U8085 ( .B1(P1_U3973), .B2(n6822), .A(n6821), .ZN(P1_U3563) );
  NAND2_X1 U8086 ( .A1(n6426), .A2(P1_U3973), .ZN(n6823) );
  OAI21_X1 U8087 ( .B1(P1_U3973), .B2(n7123), .A(n6823), .ZN(P1_U3554) );
  INV_X1 U8088 ( .A(n6879), .ZN(n6824) );
  NAND2_X1 U8089 ( .A1(n6426), .A2(n6877), .ZN(n9055) );
  NAND2_X1 U8090 ( .A1(n6824), .A2(n9055), .ZN(n8859) );
  INV_X1 U8091 ( .A(n8859), .ZN(n6826) );
  NOR2_X1 U8092 ( .A1(n11178), .A2(n10746), .ZN(n6825) );
  OAI222_X1 U8093 ( .A1(n6877), .A2(n6827), .B1(n6826), .B2(n6825), .C1(n10741), .C2(n6967), .ZN(n6860) );
  NAND2_X1 U8094 ( .A1(n6860), .A2(n11181), .ZN(n6828) );
  OAI21_X1 U8095 ( .B1(n11181), .B2(n6829), .A(n6828), .ZN(P1_U3522) );
  AOI22_X1 U8096 ( .A1(n10412), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7068), .ZN(n6830) );
  OAI21_X1 U8097 ( .B1(n8106), .B2(n9222), .A(n6830), .ZN(P1_U3343) );
  INV_X1 U8098 ( .A(n10891), .ZN(n7643) );
  INV_X1 U8099 ( .A(n8011), .ZN(n6835) );
  INV_X1 U8100 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U8101 ( .A1(n7643), .A2(P1_U3086), .B1(n9222), .B2(n6835), .C1(
        n6831), .C2(n9220), .ZN(P1_U3344) );
  INV_X1 U8102 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U8103 ( .A1(n6843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U8104 ( .A(n6834), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8214) );
  INV_X1 U8105 ( .A(n8214), .ZN(n11095) );
  OAI222_X1 U8106 ( .A1(n8844), .A2(n6836), .B1(n9800), .B2(n6835), .C1(
        P2_U3151), .C2(n11095), .ZN(P2_U3284) );
  OAI21_X1 U8107 ( .B1(n6839), .B2(n6838), .A(n6837), .ZN(n6919) );
  NAND2_X1 U8108 ( .A1(n6840), .A2(n10813), .ZN(n8835) );
  AOI22_X1 U8109 ( .A1(n9932), .A2(n6434), .B1(n8835), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U8110 ( .A1(n9904), .A2(n6964), .ZN(n6841) );
  OAI211_X1 U8111 ( .C1(n6919), .C2(n9919), .A(n6842), .B(n6841), .ZN(P1_U3232) );
  NAND2_X1 U8112 ( .A1(n7142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6845) );
  XNOR2_X1 U8113 ( .A(n6845), .B(n6844), .ZN(n8318) );
  INV_X1 U8114 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6846) );
  OAI222_X1 U8115 ( .A1(n9804), .A2(n8106), .B1(n8318), .B2(P2_U3151), .C1(
        n6846), .C2(n8844), .ZN(P2_U3283) );
  INV_X1 U8116 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7080) );
  INV_X1 U8117 ( .A(n9857), .ZN(n8823) );
  NAND2_X1 U8118 ( .A1(n8823), .A2(P1_U3973), .ZN(n6847) );
  OAI21_X1 U8119 ( .B1(P1_U3973), .B2(n7080), .A(n6847), .ZN(P1_U3570) );
  XNOR2_X1 U8120 ( .A(n6909), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6849) );
  NOR2_X1 U8121 ( .A1(n6850), .A2(n6849), .ZN(n6902) );
  AOI211_X1 U8122 ( .C1(n6850), .C2(n6849), .A(n10952), .B(n6902), .ZN(n6859)
         );
  AOI21_X1 U8123 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6852), .A(n6851), .ZN(
        n6854) );
  XNOR2_X1 U8124 ( .A(n6909), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6853) );
  NOR2_X1 U8125 ( .A1(n6854), .A2(n6853), .ZN(n6908) );
  AOI211_X1 U8126 ( .C1(n6854), .C2(n6853), .A(n10956), .B(n6908), .ZN(n6858)
         );
  INV_X1 U8127 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8128 ( .A1(n10962), .A2(n6909), .ZN(n6855) );
  NAND2_X1 U8129 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7441) );
  OAI211_X1 U8130 ( .C1(n6856), .C2(n10967), .A(n6855), .B(n7441), .ZN(n6857)
         );
  OR3_X1 U8131 ( .A1(n6859), .A2(n6858), .A3(n6857), .ZN(P1_U3250) );
  INV_X1 U8132 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6862) );
  NAND2_X1 U8133 ( .A1(n6860), .A2(n11185), .ZN(n6861) );
  OAI21_X1 U8134 ( .B1(n11185), .B2(n6862), .A(n6861), .ZN(P1_U3453) );
  NOR2_X1 U8135 ( .A1(n7142), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6950) );
  OR2_X1 U8136 ( .A1(n6950), .A2(n7131), .ZN(n6863) );
  XNOR2_X1 U8137 ( .A(n6863), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8390) );
  AOI22_X1 U8138 ( .A1(n8390), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9802), .ZN(n6864) );
  OAI21_X1 U8139 ( .B1(n8161), .B2(n9800), .A(n6864), .ZN(P2_U3282) );
  AOI22_X1 U8140 ( .A1(n10948), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7068), .ZN(n6865) );
  OAI21_X1 U8141 ( .B1(n8161), .B2(n9222), .A(n6865), .ZN(P1_U3342) );
  INV_X1 U8142 ( .A(n6866), .ZN(n8863) );
  OAI21_X1 U8143 ( .B1(n6868), .B2(n6866), .A(n6867), .ZN(n7088) );
  AOI211_X1 U8144 ( .C1(n6869), .C2(n6876), .A(n10655), .B(n6890), .ZN(n7083)
         );
  XNOR2_X1 U8145 ( .A(n8904), .B(n6866), .ZN(n6870) );
  OAI222_X1 U8146 ( .A1(n10763), .A2(n6967), .B1(n10741), .B2(n6997), .C1(
        n6870), .C2(n10713), .ZN(n7082) );
  AOI211_X1 U8147 ( .C1(n11178), .C2(n7088), .A(n7083), .B(n7082), .ZN(n6943)
         );
  OAI22_X1 U8148 ( .A1(n10739), .A2(n7086), .B1(n11181), .B2(n6787), .ZN(n6871) );
  INV_X1 U8149 ( .A(n6871), .ZN(n6872) );
  OAI21_X1 U8150 ( .B1(n6943), .B2(n11180), .A(n6872), .ZN(P1_U3524) );
  OAI21_X1 U8151 ( .B1(n6880), .B2(n6874), .A(n6873), .ZN(n7017) );
  AOI22_X1 U8152 ( .A1(n5320), .A2(n11155), .B1(n11156), .B2(n6426), .ZN(n6878) );
  OAI211_X1 U8153 ( .C1(n6877), .C2(n5941), .A(n10672), .B(n6876), .ZN(n7009)
         );
  NAND2_X1 U8154 ( .A1(n6878), .A2(n7009), .ZN(n6882) );
  XNOR2_X1 U8155 ( .A(n6880), .B(n6879), .ZN(n6881) );
  NOR2_X1 U8156 ( .A1(n6881), .A2(n10713), .ZN(n7004) );
  AOI211_X1 U8157 ( .C1(n11178), .C2(n7017), .A(n6882), .B(n7004), .ZN(n6947)
         );
  INV_X1 U8158 ( .A(n10739), .ZN(n7604) );
  AOI22_X1 U8159 ( .A1(n7604), .A2(n7011), .B1(P1_REG1_REG_1__SCAN_IN), .B2(
        n11180), .ZN(n6883) );
  OAI21_X1 U8160 ( .B1(n6947), .B2(n11180), .A(n6883), .ZN(P1_U3523) );
  INV_X1 U8161 ( .A(n8858), .ZN(n6885) );
  NAND2_X1 U8162 ( .A1(n6886), .A2(n6885), .ZN(n6884) );
  OAI21_X1 U8163 ( .B1(n6886), .B2(n6885), .A(n6884), .ZN(n6887) );
  NAND2_X1 U8164 ( .A1(n6887), .A2(n10746), .ZN(n7040) );
  AOI22_X1 U8165 ( .A1(n11155), .A2(n10355), .B1(n5320), .B2(n11156), .ZN(
        n6892) );
  OAI21_X1 U8166 ( .B1(n6889), .B2(n8858), .A(n6888), .ZN(n7038) );
  NAND2_X1 U8167 ( .A1(n7038), .A2(n11178), .ZN(n6891) );
  OAI211_X1 U8168 ( .C1(n6890), .C2(n7034), .A(n6993), .B(n10672), .ZN(n7030)
         );
  NAND4_X1 U8169 ( .A1(n7040), .A2(n6892), .A3(n6891), .A4(n7030), .ZN(n6981)
         );
  OAI22_X1 U8170 ( .A1(n10739), .A2(n7034), .B1(n11181), .B2(n6788), .ZN(n6893) );
  AOI21_X1 U8171 ( .B1(n6981), .B2(n11181), .A(n6893), .ZN(n6894) );
  INV_X1 U8172 ( .A(n6894), .ZN(P1_U3525) );
  NAND2_X1 U8173 ( .A1(n6895), .A2(n6896), .ZN(n6897) );
  XOR2_X1 U8174 ( .A(n6898), .B(n6897), .Z(n6901) );
  AOI22_X1 U8175 ( .A1(n5320), .A2(n9932), .B1(n9928), .B2(n6426), .ZN(n6900)
         );
  AOI22_X1 U8176 ( .A1(n9904), .A2(n7011), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8835), .ZN(n6899) );
  OAI211_X1 U8177 ( .C1(n6901), .C2(n9919), .A(n6900), .B(n6899), .ZN(P1_U3222) );
  AOI21_X1 U8178 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6909), .A(n6902), .ZN(
        n6903) );
  XNOR2_X1 U8179 ( .A(n7638), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6904) );
  NOR2_X1 U8180 ( .A1(n6903), .A2(n6904), .ZN(n7637) );
  INV_X1 U8181 ( .A(n6903), .ZN(n6906) );
  INV_X1 U8182 ( .A(n6904), .ZN(n6905) );
  INV_X1 U8183 ( .A(n10952), .ZN(n10916) );
  OAI21_X1 U8184 ( .B1(n6906), .B2(n6905), .A(n10916), .ZN(n6916) );
  INV_X1 U8185 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U8186 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7997) );
  OAI21_X1 U8187 ( .B1(n10967), .B2(n6907), .A(n7997), .ZN(n6914) );
  AOI21_X1 U8188 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6909), .A(n6908), .ZN(
        n6912) );
  INV_X1 U8189 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6910) );
  MUX2_X1 U8190 ( .A(n6910), .B(P1_REG1_REG_8__SCAN_IN), .S(n7638), .Z(n6911)
         );
  NOR2_X1 U8191 ( .A1(n6912), .A2(n6911), .ZN(n7631) );
  AOI211_X1 U8192 ( .C1(n6912), .C2(n6911), .A(n10956), .B(n7631), .ZN(n6913)
         );
  AOI211_X1 U8193 ( .C1(n10962), .C2(n7638), .A(n6914), .B(n6913), .ZN(n6915)
         );
  OAI21_X1 U8194 ( .B1(n7637), .B2(n6916), .A(n6915), .ZN(P1_U3251) );
  NAND2_X1 U8195 ( .A1(n6917), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6918) );
  XOR2_X1 U8196 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6918), .Z(n6922) );
  INV_X1 U8197 ( .A(P1_U3973), .ZN(n10357) );
  INV_X1 U8198 ( .A(n6919), .ZN(n6920) );
  NOR2_X1 U8199 ( .A1(n6920), .A2(n6923), .ZN(n6921) );
  AOI211_X1 U8200 ( .C1(n6923), .C2(n6922), .A(n10357), .B(n6921), .ZN(n10372)
         );
  AOI211_X1 U8201 ( .C1(n6926), .C2(n6925), .A(n6924), .B(n10956), .ZN(n6934)
         );
  AOI211_X1 U8202 ( .C1(n6929), .C2(n6928), .A(n6927), .B(n10952), .ZN(n6933)
         );
  AOI22_X1 U8203 ( .A1(n10396), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6930) );
  OAI21_X1 U8204 ( .B1(n6931), .B2(n10374), .A(n6930), .ZN(n6932) );
  OR4_X1 U8205 ( .A1(n10372), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(P1_U3245) );
  NAND2_X1 U8206 ( .A1(n6935), .A2(n6949), .ZN(n6936) );
  OR2_X1 U8207 ( .A1(n7142), .A2(n7140), .ZN(n6937) );
  NAND2_X1 U8208 ( .A1(n6937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7078) );
  XNOR2_X1 U8209 ( .A(n7078), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9420) );
  AOI22_X1 U8210 ( .A1(n9420), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n9802), .ZN(n6938) );
  OAI21_X1 U8211 ( .B1(n8508), .B2(n9804), .A(n6938), .ZN(P2_U3280) );
  AOI22_X1 U8212 ( .A1(n10917), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7068), .ZN(n6939) );
  OAI21_X1 U8213 ( .B1(n8508), .B2(n9222), .A(n6939), .ZN(P1_U3340) );
  INV_X1 U8214 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6940) );
  OAI22_X1 U8215 ( .A1(n10806), .A2(n7086), .B1(n11185), .B2(n6940), .ZN(n6941) );
  INV_X1 U8216 ( .A(n6941), .ZN(n6942) );
  OAI21_X1 U8217 ( .B1(n6943), .B2(n11182), .A(n6942), .ZN(P1_U3459) );
  INV_X1 U8218 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6944) );
  OAI22_X1 U8219 ( .A1(n10806), .A2(n5941), .B1(n11185), .B2(n6944), .ZN(n6945) );
  INV_X1 U8220 ( .A(n6945), .ZN(n6946) );
  OAI21_X1 U8221 ( .B1(n6947), .B2(n11182), .A(n6946), .ZN(P1_U3456) );
  INV_X1 U8222 ( .A(n8517), .ZN(n6953) );
  INV_X1 U8223 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6948) );
  OAI222_X1 U8224 ( .A1(n10422), .A2(P1_U3086), .B1(n9222), .B2(n6953), .C1(
        n6948), .C2(n9220), .ZN(P1_U3341) );
  INV_X1 U8225 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6954) );
  AND2_X1 U8226 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  XNOR2_X1 U8227 ( .A(n6952), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9401) );
  INV_X1 U8228 ( .A(n9401), .ZN(n8386) );
  OAI222_X1 U8229 ( .A1(n8844), .A2(n6954), .B1(n9800), .B2(n6953), .C1(
        P2_U3151), .C2(n8386), .ZN(P2_U3281) );
  NAND2_X1 U8230 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  INV_X2 U8231 ( .A(n10661), .ZN(n7511) );
  NAND2_X1 U8232 ( .A1(n10601), .A2(n11155), .ZN(n10572) );
  NOR2_X1 U8233 ( .A1(n10601), .A2(n6959), .ZN(n6962) );
  AND3_X1 U8234 ( .A1(n8859), .A2(n6960), .A3(n10661), .ZN(n6961) );
  AOI211_X1 U8235 ( .C1(n10632), .C2(P1_REG3_REG_0__SCAN_IN), .A(n6962), .B(
        n6961), .ZN(n6966) );
  NOR2_X1 U8236 ( .A1(n10576), .A2(n10655), .ZN(n10480) );
  OAI21_X1 U8237 ( .B1(n10480), .B2(n10580), .A(n6964), .ZN(n6965) );
  OAI211_X1 U8238 ( .C1(n6967), .C2(n10572), .A(n6966), .B(n6965), .ZN(
        P1_U3293) );
  XNOR2_X1 U8239 ( .A(n8917), .B(n8908), .ZN(n6968) );
  OAI222_X1 U8240 ( .A1(n10763), .A2(n7420), .B1(n10741), .B2(n7042), .C1(
        n6968), .C2(n10713), .ZN(n11130) );
  INV_X1 U8241 ( .A(n11130), .ZN(n6978) );
  OAI21_X1 U8242 ( .B1(n6970), .B2(n8917), .A(n6969), .ZN(n11132) );
  NAND2_X1 U8243 ( .A1(n11166), .A2(n7005), .ZN(n6971) );
  INV_X1 U8244 ( .A(n6994), .ZN(n6973) );
  INV_X1 U8245 ( .A(n6972), .ZN(n7022) );
  OAI211_X1 U8246 ( .C1(n11129), .C2(n6973), .A(n7022), .B(n10672), .ZN(n11128) );
  AOI22_X1 U8247 ( .A1(n7511), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7423), .B2(
        n10632), .ZN(n6975) );
  NAND2_X1 U8248 ( .A1(n10580), .A2(n7418), .ZN(n6974) );
  OAI211_X1 U8249 ( .C1(n11128), .C2(n10576), .A(n6975), .B(n6974), .ZN(n6976)
         );
  AOI21_X1 U8250 ( .B1(n11132), .B2(n10651), .A(n6976), .ZN(n6977) );
  OAI21_X1 U8251 ( .B1(n6978), .B2(n7511), .A(n6977), .ZN(P1_U3288) );
  INV_X1 U8252 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6979) );
  OAI22_X1 U8253 ( .A1(n10806), .A2(n7034), .B1(n11185), .B2(n6979), .ZN(n6980) );
  AOI21_X1 U8254 ( .B1(n6981), .B2(n11185), .A(n6980), .ZN(n6982) );
  INV_X1 U8255 ( .A(n6982), .ZN(P1_U3462) );
  XOR2_X1 U8256 ( .A(n6984), .B(n6983), .Z(n6990) );
  AOI22_X1 U8257 ( .A1(n9904), .A2(n6985), .B1(n10355), .B2(n9932), .ZN(n6989)
         );
  NAND2_X1 U8258 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10359) );
  INV_X1 U8259 ( .A(n10359), .ZN(n6987) );
  NOR2_X1 U8260 ( .A1(n7014), .A2(n9912), .ZN(n6986) );
  AOI211_X1 U8261 ( .C1(n9917), .C2(n7031), .A(n6987), .B(n6986), .ZN(n6988)
         );
  OAI211_X1 U8262 ( .C1(n6990), .C2(n9919), .A(n6989), .B(n6988), .ZN(P1_U3218) );
  OAI21_X1 U8263 ( .B1(n6992), .B2(n8861), .A(n6991), .ZN(n7076) );
  AOI21_X1 U8264 ( .B1(n6993), .B2(n5979), .A(n10655), .ZN(n6995) );
  AND2_X1 U8265 ( .A1(n6995), .A2(n6994), .ZN(n7070) );
  XNOR2_X1 U8266 ( .A(n5227), .B(n8861), .ZN(n6996) );
  OAI222_X1 U8267 ( .A1(n10741), .A2(n9877), .B1(n10763), .B2(n6997), .C1(
        n6996), .C2(n10713), .ZN(n7073) );
  AOI211_X1 U8268 ( .C1(n11178), .C2(n7076), .A(n7070), .B(n7073), .ZN(n7003)
         );
  AOI22_X1 U8269 ( .A1(n7604), .A2(n5979), .B1(n11180), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6998) );
  OAI21_X1 U8270 ( .B1(n7003), .B2(n11180), .A(n6998), .ZN(P1_U3526) );
  INV_X1 U8271 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6999) );
  OAI22_X1 U8272 ( .A1(n10806), .A2(n7000), .B1(n11185), .B2(n6999), .ZN(n7001) );
  INV_X1 U8273 ( .A(n7001), .ZN(n7002) );
  OAI21_X1 U8274 ( .B1(n7003), .B2(n11182), .A(n7002), .ZN(P1_U3465) );
  INV_X1 U8275 ( .A(n7004), .ZN(n7019) );
  INV_X1 U8276 ( .A(n11166), .ZN(n7008) );
  INV_X1 U8277 ( .A(n7005), .ZN(n7006) );
  NAND2_X1 U8278 ( .A1(n10661), .A2(n7006), .ZN(n8065) );
  INV_X1 U8279 ( .A(n8065), .ZN(n7007) );
  AOI21_X1 U8280 ( .B1(n7008), .B2(n10661), .A(n7007), .ZN(n7520) );
  INV_X1 U8281 ( .A(n7520), .ZN(n7037) );
  INV_X1 U8282 ( .A(n6426), .ZN(n7010) );
  NAND2_X1 U8283 ( .A1(n10601), .A2(n11156), .ZN(n10488) );
  OAI22_X1 U8284 ( .A1(n7010), .A2(n10488), .B1(n7009), .B2(n10576), .ZN(n7016) );
  AOI22_X1 U8285 ( .A1(n7511), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10632), .ZN(n7013) );
  NAND2_X1 U8286 ( .A1(n10580), .A2(n7011), .ZN(n7012) );
  OAI211_X1 U8287 ( .C1(n7014), .C2(n10572), .A(n7013), .B(n7012), .ZN(n7015)
         );
  AOI211_X1 U8288 ( .C1(n7017), .C2(n7037), .A(n7016), .B(n7015), .ZN(n7018)
         );
  OAI21_X1 U8289 ( .B1(n7019), .B2(n7511), .A(n7018), .ZN(P1_U3292) );
  XOR2_X1 U8290 ( .A(n7020), .B(n8914), .Z(n7021) );
  NAND2_X1 U8291 ( .A1(n7021), .A2(n10746), .ZN(n7058) );
  AOI211_X1 U8292 ( .C1(n7405), .C2(n7022), .A(n10655), .B(n7048), .ZN(n7056)
         );
  INV_X1 U8293 ( .A(n10572), .ZN(n8272) );
  AOI22_X1 U8294 ( .A1(n10352), .A2(n8272), .B1(n10580), .B2(n7405), .ZN(n7024) );
  AOI22_X1 U8295 ( .A1(n7511), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7409), .B2(
        n10632), .ZN(n7023) );
  OAI211_X1 U8296 ( .C1(n9877), .C2(n10488), .A(n7024), .B(n7023), .ZN(n7025)
         );
  AOI21_X1 U8297 ( .B1(n7056), .B2(n10664), .A(n7025), .ZN(n7029) );
  OAI21_X1 U8298 ( .B1(n7027), .B2(n8914), .A(n7026), .ZN(n7057) );
  NAND2_X1 U8299 ( .A1(n7057), .A2(n7037), .ZN(n7028) );
  OAI211_X1 U8300 ( .C1(n7058), .C2(n7511), .A(n7029), .B(n7028), .ZN(P1_U3287) );
  NOR2_X1 U8301 ( .A1(n7030), .A2(n10576), .ZN(n7036) );
  INV_X1 U8302 ( .A(n10488), .ZN(n10569) );
  AOI22_X1 U8303 ( .A1(n8272), .A2(n10355), .B1(n5320), .B2(n10569), .ZN(n7033) );
  AOI22_X1 U8304 ( .A1(n7511), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10632), .B2(
        n7031), .ZN(n7032) );
  OAI211_X1 U8305 ( .C1(n7034), .C2(n10658), .A(n7033), .B(n7032), .ZN(n7035)
         );
  AOI211_X1 U8306 ( .C1(n7038), .C2(n7037), .A(n7036), .B(n7035), .ZN(n7039)
         );
  OAI21_X1 U8307 ( .B1(n7511), .B2(n7040), .A(n7039), .ZN(P1_U3290) );
  XNOR2_X1 U8308 ( .A(n7349), .B(n5397), .ZN(n7041) );
  NAND2_X1 U8309 ( .A1(n7041), .A2(n10746), .ZN(n7045) );
  OAI22_X1 U8310 ( .A1(n7042), .A2(n10763), .B1(n7868), .B2(n10741), .ZN(n7043) );
  INV_X1 U8311 ( .A(n7043), .ZN(n7044) );
  NAND2_X1 U8312 ( .A1(n7045), .A2(n7044), .ZN(n11140) );
  INV_X1 U8313 ( .A(n11140), .ZN(n7054) );
  OAI21_X1 U8314 ( .B1(n7047), .B2(n8868), .A(n7046), .ZN(n11142) );
  OAI211_X1 U8315 ( .C1(n7048), .C2(n11139), .A(n10672), .B(n7356), .ZN(n11138) );
  AOI22_X1 U8316 ( .A1(n7511), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7443), .B2(
        n10632), .ZN(n7051) );
  NAND2_X1 U8317 ( .A1(n7049), .A2(n10580), .ZN(n7050) );
  OAI211_X1 U8318 ( .C1(n11138), .C2(n10576), .A(n7051), .B(n7050), .ZN(n7052)
         );
  AOI21_X1 U8319 ( .B1(n11142), .B2(n10651), .A(n7052), .ZN(n7053) );
  OAI21_X1 U8320 ( .B1(n7054), .B2(n7511), .A(n7053), .ZN(P1_U3286) );
  OAI22_X1 U8321 ( .A1(n7353), .A2(n10741), .B1(n9877), .B2(n10763), .ZN(n7055) );
  AOI211_X1 U8322 ( .C1(n7057), .C2(n11178), .A(n7056), .B(n7055), .ZN(n7059)
         );
  NAND2_X1 U8323 ( .A1(n7059), .A2(n7058), .ZN(n7066) );
  INV_X1 U8324 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7060) );
  OAI22_X1 U8325 ( .A1(n10739), .A2(n7064), .B1(n11181), .B2(n7060), .ZN(n7061) );
  AOI21_X1 U8326 ( .B1(n7066), .B2(n11181), .A(n7061), .ZN(n7062) );
  INV_X1 U8327 ( .A(n7062), .ZN(P1_U3528) );
  INV_X1 U8328 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7063) );
  OAI22_X1 U8329 ( .A1(n10806), .A2(n7064), .B1(n11185), .B2(n7063), .ZN(n7065) );
  AOI21_X1 U8330 ( .B1(n7066), .B2(n11185), .A(n7065), .ZN(n7067) );
  INV_X1 U8331 ( .A(n7067), .ZN(P1_U3471) );
  INV_X1 U8332 ( .A(n8531), .ZN(n7081) );
  AOI22_X1 U8333 ( .A1(n10441), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7068), .ZN(n7069) );
  OAI21_X1 U8334 ( .B1(n7081), .B2(n9222), .A(n7069), .ZN(P1_U3339) );
  INV_X1 U8335 ( .A(n7070), .ZN(n7072) );
  AOI22_X1 U8336 ( .A1(n10580), .A2(n5979), .B1(n10632), .B2(n9880), .ZN(n7071) );
  OAI21_X1 U8337 ( .B1(n7072), .B2(n10576), .A(n7071), .ZN(n7075) );
  MUX2_X1 U8338 ( .A(n7073), .B(P1_REG2_REG_4__SCAN_IN), .S(n7511), .Z(n7074)
         );
  AOI211_X1 U8339 ( .C1(n10651), .C2(n7076), .A(n7075), .B(n7074), .ZN(n7077)
         );
  INV_X1 U8340 ( .A(n7077), .ZN(P1_U3289) );
  NAND2_X1 U8341 ( .A1(n7078), .A2(n7138), .ZN(n7079) );
  NAND2_X1 U8342 ( .A1(n7079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7364) );
  XNOR2_X1 U8343 ( .A(n7364), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9439) );
  INV_X1 U8344 ( .A(n9439), .ZN(n8382) );
  OAI222_X1 U8345 ( .A1(n8382), .A2(P2_U3151), .B1(n9800), .B2(n7081), .C1(
        n8844), .C2(n7080), .ZN(P2_U3279) );
  INV_X1 U8346 ( .A(n7082), .ZN(n7090) );
  NAND2_X1 U8347 ( .A1(n7083), .A2(n10664), .ZN(n7085) );
  AOI22_X1 U8348 ( .A1(n7511), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10632), .ZN(n7084) );
  OAI211_X1 U8349 ( .C1(n7086), .C2(n10658), .A(n7085), .B(n7084), .ZN(n7087)
         );
  AOI21_X1 U8350 ( .B1(n10651), .B2(n7088), .A(n7087), .ZN(n7089) );
  OAI21_X1 U8351 ( .B1(n7090), .B2(n7511), .A(n7089), .ZN(P1_U3291) );
  NAND2_X1 U8352 ( .A1(n10357), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7091) );
  OAI21_X1 U8353 ( .B1(n10487), .B2(n10357), .A(n7091), .ZN(P1_U3583) );
  NAND2_X1 U8354 ( .A1(n7105), .A2(n7106), .ZN(n7104) );
  NOR2_X1 U8355 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7095) );
  NAND2_X1 U8356 ( .A1(n7155), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7103) );
  INV_X1 U8357 ( .A(n7098), .ZN(n8839) );
  NAND2_X1 U8358 ( .A1(n7757), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U8359 ( .A1(n7539), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7101) );
  AND2_X2 U8360 ( .A1(n8839), .A2(n7099), .ZN(n7156) );
  OAI21_X1 U8361 ( .B1(n7105), .B2(n7131), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n7108) );
  NAND2_X1 U8362 ( .A1(n7313), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U8363 ( .A1(n7532), .A2(n7114), .ZN(n7117) );
  INV_X1 U8364 ( .A(n7234), .ZN(n7115) );
  NAND2_X1 U8365 ( .A1(n7534), .A2(n7115), .ZN(n7116) );
  OR2_X1 U8366 ( .A1(n7305), .A2(n7304), .ZN(n8456) );
  NAND2_X1 U8367 ( .A1(n7305), .A2(n7304), .ZN(n8458) );
  NAND2_X1 U8368 ( .A1(n7757), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U8369 ( .A1(n7156), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U8370 ( .A1(n7155), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8371 ( .A1(n7539), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7119) );
  NAND4_X1 U8372 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n7164)
         );
  INV_X1 U8373 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U8374 ( .A1(n8701), .A2(SI_0_), .ZN(n7124) );
  XNOR2_X1 U8375 ( .A(n7124), .B(n7123), .ZN(n9806) );
  OR2_X1 U8376 ( .A1(n7164), .A2(n7686), .ZN(n8455) );
  INV_X1 U8377 ( .A(n8455), .ZN(n7283) );
  NAND2_X1 U8378 ( .A1(n7282), .A2(n8456), .ZN(n7427) );
  INV_X1 U8379 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11106) );
  OR2_X1 U8380 ( .A1(n8037), .A2(n11106), .ZN(n7129) );
  NAND2_X1 U8381 ( .A1(n7155), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7128) );
  INV_X1 U8382 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7125) );
  NAND2_X1 U8383 ( .A1(n7156), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7126) );
  NAND2_X1 U8384 ( .A1(n7313), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7136) );
  XNOR2_X2 U8385 ( .A(n7134), .B(n7133), .ZN(n7237) );
  INV_X1 U8386 ( .A(n7237), .ZN(n7219) );
  NAND2_X1 U8387 ( .A1(n7534), .A2(n7219), .ZN(n7135) );
  XNOR2_X1 U8388 ( .A(n7427), .B(n8469), .ZN(n11102) );
  NAND3_X1 U8389 ( .A1(n7363), .A2(n7138), .A3(n7137), .ZN(n7139) );
  NAND2_X1 U8390 ( .A1(n7148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7149) );
  INV_X1 U8391 ( .A(n8800), .ZN(n8084) );
  AOI21_X1 U8392 ( .B1(n8746), .B2(n8084), .A(n7153), .ZN(n7152) );
  AND2_X1 U8393 ( .A1(n9775), .A2(n7152), .ZN(n7154) );
  NAND2_X2 U8394 ( .A1(n7189), .A2(n8800), .ZN(n8464) );
  NAND2_X1 U8395 ( .A1(n7732), .A2(n8787), .ZN(n7191) );
  INV_X1 U8396 ( .A(n9203), .ZN(n7654) );
  NAND2_X1 U8397 ( .A1(n7155), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7157) );
  INV_X1 U8398 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7697) );
  INV_X1 U8399 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7212) );
  INV_X1 U8400 ( .A(n7336), .ZN(n7161) );
  AOI22_X1 U8401 ( .A1(n9393), .A2(n7160), .B1(n7162), .B2(n7305), .ZN(n7169)
         );
  INV_X1 U8402 ( .A(n7686), .ZN(n7163) );
  NAND2_X1 U8403 ( .A1(n7164), .A2(n7163), .ZN(n7284) );
  NAND2_X1 U8404 ( .A1(n8725), .A2(n7284), .ZN(n7285) );
  INV_X1 U8405 ( .A(n7304), .ZN(n7715) );
  OR2_X1 U8406 ( .A1(n7305), .A2(n7715), .ZN(n7165) );
  NAND2_X1 U8407 ( .A1(n7285), .A2(n7165), .ZN(n7166) );
  NAND2_X1 U8408 ( .A1(n7166), .A2(n8469), .ZN(n7432) );
  OAI21_X1 U8409 ( .B1(n8469), .B2(n7166), .A(n7432), .ZN(n7167) );
  AND2_X1 U8410 ( .A1(n7189), .A2(n8746), .ZN(n8785) );
  AND2_X1 U8411 ( .A1(n7153), .A2(n8800), .ZN(n7268) );
  NAND2_X1 U8412 ( .A1(n7167), .A2(n9643), .ZN(n7168) );
  OAI211_X1 U8413 ( .C1(n11102), .C2(n7654), .A(n7169), .B(n7168), .ZN(n11107)
         );
  INV_X1 U8414 ( .A(n9704), .ZN(n7653) );
  OAI22_X1 U8415 ( .A1(n11102), .A2(n7653), .B1(n11104), .B2(n9775), .ZN(n7170) );
  NOR2_X1 U8416 ( .A1(n11107), .A2(n7170), .ZN(n11101) );
  NAND3_X1 U8417 ( .A1(n8746), .A2(n8800), .A3(n8787), .ZN(n7171) );
  NAND2_X1 U8418 ( .A1(n7679), .A2(n7678), .ZN(n7681) );
  NAND2_X1 U8419 ( .A1(n7172), .A2(n6782), .ZN(n7175) );
  OR2_X1 U8420 ( .A1(n7173), .A2(n6763), .ZN(n7174) );
  NAND2_X1 U8421 ( .A1(n7176), .A2(n7177), .ZN(n7270) );
  NOR2_X1 U8422 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n7181) );
  NOR4_X1 U8423 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n7180) );
  NOR4_X1 U8424 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n7179) );
  NOR4_X1 U8425 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n7178) );
  NAND4_X1 U8426 ( .A1(n7181), .A2(n7180), .A3(n7179), .A4(n7178), .ZN(n7187)
         );
  NOR4_X1 U8427 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n7185) );
  NOR4_X1 U8428 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n7184) );
  NOR4_X1 U8429 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n7183) );
  NOR4_X1 U8430 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n7182) );
  NAND4_X1 U8431 ( .A1(n7185), .A2(n7184), .A3(n7183), .A4(n7182), .ZN(n7186)
         );
  OAI21_X1 U8432 ( .B1(n7187), .B2(n7186), .A(n7172), .ZN(n7273) );
  AND2_X1 U8433 ( .A1(n7318), .A2(n7273), .ZN(n7188) );
  NOR2_X1 U8434 ( .A1(n7274), .A2(n7189), .ZN(n7300) );
  NAND2_X1 U8435 ( .A1(n7300), .A2(n9704), .ZN(n7190) );
  NAND3_X1 U8436 ( .A1(n7681), .A2(n7682), .A3(n7190), .ZN(n7194) );
  INV_X1 U8437 ( .A(n7191), .ZN(n7192) );
  INV_X1 U8438 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7217) );
  OR2_X1 U8439 ( .A1(n8232), .A2(n7217), .ZN(n7195) );
  OAI21_X1 U8440 ( .B1(n11101), .B2(n5132), .A(n7195), .ZN(P2_U3461) );
  OR2_X1 U8441 ( .A1(n8464), .A2(n8097), .ZN(n7196) );
  NAND2_X1 U8442 ( .A1(n7196), .A2(n7252), .ZN(n7251) );
  OR2_X1 U8443 ( .A1(n7251), .A2(n7534), .ZN(n7197) );
  NAND2_X1 U8444 ( .A1(n7197), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8445 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U8446 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n7237), .ZN(n7201) );
  OAI21_X1 U8447 ( .B1(n7237), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7201), .ZN(
        n10994) );
  AND2_X1 U8448 ( .A1(n10974), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U8449 ( .A1(n7232), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7199) );
  OAI21_X1 U8450 ( .B1(n7234), .B2(n7198), .A(n7199), .ZN(n10977) );
  INV_X1 U8451 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10976) );
  INV_X1 U8452 ( .A(n7199), .ZN(n7200) );
  NOR2_X1 U8453 ( .A1(n10975), .A2(n7200), .ZN(n10995) );
  NOR2_X1 U8454 ( .A1(n10994), .A2(n10995), .ZN(n10993) );
  INV_X1 U8455 ( .A(n7201), .ZN(n7202) );
  XNOR2_X1 U8456 ( .A(n7203), .B(n11016), .ZN(n11009) );
  NOR2_X1 U8457 ( .A1(n11016), .A2(n7203), .ZN(n7204) );
  NAND2_X1 U8458 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n7243), .ZN(n7205) );
  OAI21_X1 U8459 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n7243), .A(n7205), .ZN(
        n11025) );
  INV_X1 U8460 ( .A(n7205), .ZN(n7206) );
  NOR2_X1 U8461 ( .A1(n7535), .A2(n7207), .ZN(n7208) );
  INV_X1 U8462 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U8463 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n11061), .ZN(n7209) );
  OAI21_X1 U8464 ( .B1(n11061), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7209), .ZN(
        n11069) );
  NOR2_X1 U8465 ( .A1(n11070), .A2(n11069), .ZN(n11068) );
  AOI21_X1 U8466 ( .B1(n7803), .B2(n7210), .A(n7608), .ZN(n7264) );
  NOR2_X1 U8467 ( .A1(n7158), .A2(P2_U3151), .ZN(n8333) );
  INV_X1 U8468 ( .A(n8333), .ZN(n7211) );
  OR2_X1 U8469 ( .A1(n7251), .A2(n7211), .ZN(n10968) );
  MUX2_X1 U8470 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8795), .Z(n7221) );
  INV_X1 U8471 ( .A(n7221), .ZN(n7222) );
  MUX2_X1 U8472 ( .A(n7697), .B(n7212), .S(n7159), .Z(n7220) );
  INV_X1 U8473 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10980) );
  MUX2_X1 U8474 ( .A(n10976), .B(n10980), .S(n7159), .Z(n7215) );
  XNOR2_X1 U8475 ( .A(n7215), .B(n7234), .ZN(n10987) );
  INV_X1 U8476 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7214) );
  INV_X1 U8477 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7213) );
  MUX2_X1 U8478 ( .A(n7214), .B(n7213), .S(n7159), .Z(n10969) );
  NAND2_X1 U8479 ( .A1(n10969), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10988) );
  INV_X1 U8480 ( .A(n7215), .ZN(n7216) );
  AOI22_X1 U8481 ( .A1(n10987), .A2(n10988), .B1(n7234), .B2(n7216), .ZN(
        n11003) );
  MUX2_X1 U8482 ( .A(n7125), .B(n7217), .S(n7159), .Z(n7218) );
  XNOR2_X1 U8483 ( .A(n7218), .B(n7219), .ZN(n11004) );
  OAI22_X1 U8484 ( .A1(n11003), .A2(n11004), .B1(n7219), .B2(n7218), .ZN(
        n11018) );
  XNOR2_X1 U8485 ( .A(n7220), .B(n11016), .ZN(n11019) );
  NOR2_X1 U8486 ( .A1(n11018), .A2(n11019), .ZN(n11017) );
  AOI21_X1 U8487 ( .B1(n11016), .B2(n7220), .A(n11017), .ZN(n11037) );
  XNOR2_X1 U8488 ( .A(n11034), .B(n7221), .ZN(n11036) );
  NAND2_X1 U8489 ( .A1(n11037), .A2(n11036), .ZN(n11035) );
  MUX2_X1 U8490 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8795), .Z(n7223) );
  XNOR2_X1 U8491 ( .A(n7223), .B(n7535), .ZN(n11049) );
  MUX2_X1 U8492 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8795), .Z(n7224) );
  NOR2_X1 U8493 ( .A1(n7224), .A2(n11061), .ZN(n7225) );
  AOI21_X1 U8494 ( .B1(n7224), .B2(n11061), .A(n7225), .ZN(n11065) );
  NAND2_X1 U8495 ( .A1(n11066), .A2(n11065), .ZN(n11064) );
  INV_X1 U8496 ( .A(n7225), .ZN(n7226) );
  NAND2_X1 U8497 ( .A1(n11064), .A2(n7226), .ZN(n7230) );
  MUX2_X1 U8498 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8795), .Z(n7228) );
  NOR2_X1 U8499 ( .A1(n7228), .A2(n7227), .ZN(n7620) );
  AOI21_X1 U8500 ( .B1(n7228), .B2(n7227), .A(n7620), .ZN(n7229) );
  NOR2_X1 U8501 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  NAND2_X1 U8502 ( .A1(P2_U3893), .A2(n7158), .ZN(n11020) );
  OAI21_X1 U8503 ( .B1(n7619), .B2(n7231), .A(n11086), .ZN(n7263) );
  INV_X1 U8504 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7249) );
  AND2_X1 U8505 ( .A1(n10974), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U8506 ( .A1(n7232), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7235) );
  INV_X1 U8507 ( .A(n7235), .ZN(n7236) );
  NAND2_X1 U8508 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(n7237), .ZN(n7238) );
  NOR2_X1 U8509 ( .A1(n10997), .A2(n7239), .ZN(n7240) );
  NOR2_X1 U8510 ( .A1(n11016), .A2(n7240), .ZN(n7241) );
  NAND2_X1 U8511 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n7243), .ZN(n7242) );
  NOR2_X1 U8512 ( .A1(n7535), .A2(n7244), .ZN(n7245) );
  INV_X1 U8513 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U8514 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n11061), .ZN(n7246) );
  OAI21_X1 U8515 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n11061), .A(n7246), .ZN(
        n11060) );
  INV_X1 U8516 ( .A(n7246), .ZN(n7247) );
  AOI21_X1 U8517 ( .B1(n7249), .B2(n7248), .A(n7613), .ZN(n7260) );
  INV_X1 U8518 ( .A(n7158), .ZN(n8796) );
  OR2_X1 U8519 ( .A1(n7159), .A2(P2_U3151), .ZN(n8330) );
  OR3_X1 U8520 ( .A1(n7251), .A2(n8796), .A3(n8330), .ZN(n7254) );
  INV_X1 U8521 ( .A(n7252), .ZN(n7256) );
  NAND2_X1 U8522 ( .A1(n8333), .A2(n7256), .ZN(n7253) );
  INV_X1 U8523 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7255) );
  NOR2_X1 U8524 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7255), .ZN(n7765) );
  INV_X1 U8525 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7257) );
  NOR2_X1 U8526 ( .A1(n11040), .A2(n7257), .ZN(n7258) );
  AOI211_X1 U8527 ( .C1(n7747), .C2(n11033), .A(n7765), .B(n7258), .ZN(n7259)
         );
  OAI21_X1 U8528 ( .B1(n7260), .B2(n11090), .A(n7259), .ZN(n7261) );
  INV_X1 U8529 ( .A(n7261), .ZN(n7262) );
  OAI211_X1 U8530 ( .C1(n7264), .C2(n11081), .A(n7263), .B(n7262), .ZN(
        P2_U3189) );
  NAND2_X1 U8531 ( .A1(n7164), .A2(n7686), .ZN(n8454) );
  NAND2_X1 U8532 ( .A1(n8455), .A2(n8454), .ZN(n8728) );
  INV_X1 U8533 ( .A(n8728), .ZN(n7266) );
  NOR2_X1 U8534 ( .A1(n9779), .A2(n9643), .ZN(n7265) );
  INV_X1 U8535 ( .A(n7305), .ZN(n7486) );
  OAI222_X1 U8536 ( .A1(n7686), .A2(n9775), .B1(n7266), .B2(n7265), .C1(n9773), 
        .C2(n7486), .ZN(n7279) );
  NAND2_X1 U8537 ( .A1(n7279), .A2(n8232), .ZN(n7267) );
  OAI21_X1 U8538 ( .B1(n8232), .B2(n7213), .A(n7267), .ZN(P2_U3459) );
  INV_X1 U8539 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7281) );
  INV_X1 U8540 ( .A(n7268), .ZN(n7269) );
  OR3_X1 U8541 ( .A1(n7189), .A2(n7269), .A3(n7732), .ZN(n7291) );
  INV_X1 U8542 ( .A(n7270), .ZN(n7271) );
  NAND2_X1 U8543 ( .A1(n7271), .A2(n7273), .ZN(n7293) );
  NAND2_X1 U8544 ( .A1(n7319), .A2(n7291), .ZN(n7272) );
  NAND2_X1 U8545 ( .A1(n7272), .A2(n11103), .ZN(n7294) );
  NAND2_X1 U8546 ( .A1(n7294), .A2(n7327), .ZN(n7275) );
  OAI21_X1 U8547 ( .B1(n7291), .B2(n7293), .A(n7275), .ZN(n7276) );
  NAND2_X1 U8548 ( .A1(n7276), .A2(n7318), .ZN(n7278) );
  INV_X1 U8549 ( .A(n7293), .ZN(n7340) );
  NAND2_X1 U8550 ( .A1(n8797), .A2(n7340), .ZN(n7277) );
  NAND2_X1 U8551 ( .A1(n7279), .A2(n11195), .ZN(n7280) );
  OAI21_X1 U8552 ( .B1(n7281), .B2(n11195), .A(n7280), .ZN(P2_U3390) );
  OAI21_X1 U8553 ( .B1(n7287), .B2(n7283), .A(n7282), .ZN(n7718) );
  NOR2_X1 U8554 ( .A1(n7304), .A2(n9775), .ZN(n7289) );
  INV_X1 U8555 ( .A(n7164), .ZN(n7494) );
  INV_X1 U8556 ( .A(n7284), .ZN(n7307) );
  INV_X1 U8557 ( .A(n7285), .ZN(n7286) );
  AOI21_X1 U8558 ( .B1(n7307), .B2(n7287), .A(n7286), .ZN(n7288) );
  OAI222_X1 U8559 ( .A1(n9773), .A2(n7311), .B1(n9687), .B2(n7494), .C1(n9689), 
        .C2(n7288), .ZN(n7714) );
  AOI211_X1 U8560 ( .C1(n9779), .C2(n7718), .A(n7289), .B(n7714), .ZN(n11099)
         );
  OR2_X1 U8561 ( .A1(n11099), .A2(n5132), .ZN(n7290) );
  OAI21_X1 U8562 ( .B1(n8232), .B2(n10980), .A(n7290), .ZN(P2_U3460) );
  NOR2_X1 U8563 ( .A1(n7327), .A2(n7291), .ZN(n7292) );
  AOI21_X1 U8564 ( .B1(n7294), .B2(n7293), .A(n7292), .ZN(n7317) );
  NAND4_X1 U8565 ( .A1(n7317), .A2(n7296), .A3(n7295), .A4(n7677), .ZN(n7298)
         );
  INV_X1 U8566 ( .A(n7327), .ZN(n7297) );
  AOI22_X2 U8567 ( .A1(n7298), .A2(P2_STATE_REG_SCAN_IN), .B1(n8797), .B2(
        n7297), .ZN(n9348) );
  INV_X1 U8568 ( .A(n7300), .ZN(n7301) );
  NAND2_X1 U8569 ( .A1(n7301), .A2(n8746), .ZN(n7302) );
  XNOR2_X1 U8570 ( .A(n9158), .B(n7304), .ZN(n7306) );
  NOR2_X1 U8571 ( .A1(n7306), .A2(n7305), .ZN(n7308) );
  NAND2_X1 U8572 ( .A1(n7491), .A2(n7492), .ZN(n7490) );
  INV_X1 U8573 ( .A(n7308), .ZN(n7309) );
  NAND2_X1 U8574 ( .A1(n7490), .A2(n7309), .ZN(n7483) );
  XNOR2_X1 U8575 ( .A(n7310), .B(n7311), .ZN(n7484) );
  NAND2_X1 U8576 ( .A1(n7483), .A2(n7484), .ZN(n7323) );
  INV_X1 U8577 ( .A(n7310), .ZN(n7312) );
  NAND2_X1 U8578 ( .A1(n7312), .A2(n7311), .ZN(n7322) );
  AND2_X1 U8579 ( .A1(n7323), .A2(n7322), .ZN(n7326) );
  NAND2_X1 U8580 ( .A1(n7313), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7315) );
  NAND2_X1 U8581 ( .A1(n7534), .A2(n11016), .ZN(n7314) );
  XNOR2_X1 U8582 ( .A(n7521), .B(n7565), .ZN(n7325) );
  INV_X1 U8583 ( .A(n7317), .ZN(n7321) );
  NAND2_X1 U8584 ( .A1(n7319), .A2(n7318), .ZN(n7320) );
  AND2_X1 U8585 ( .A1(n7325), .A2(n7322), .ZN(n7324) );
  NAND2_X1 U8586 ( .A1(n7324), .A2(n7323), .ZN(n7523) );
  OAI211_X1 U8587 ( .C1(n7326), .C2(n7325), .A(n9370), .B(n7523), .ZN(n7345)
         );
  AND2_X1 U8588 ( .A1(n8797), .A2(n7327), .ZN(n7337) );
  INV_X1 U8589 ( .A(n7337), .ZN(n7328) );
  NAND2_X1 U8590 ( .A1(n7155), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7335) );
  INV_X1 U8591 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7329) );
  OR2_X1 U8592 ( .A1(n7548), .A2(n7329), .ZN(n7334) );
  NOR2_X1 U8593 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7540) );
  AND2_X1 U8594 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7330) );
  NOR2_X1 U8595 ( .A1(n7540), .A2(n7330), .ZN(n7706) );
  OR2_X1 U8596 ( .A1(n8037), .A2(n7706), .ZN(n7333) );
  INV_X1 U8597 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7331) );
  OR2_X1 U8598 ( .A1(n8711), .A2(n7331), .ZN(n7332) );
  NAND2_X1 U8599 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  NOR2_X1 U8600 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5382), .ZN(n11015) );
  AOI21_X1 U8601 ( .B1(n9327), .B2(n7562), .A(n11015), .ZN(n7342) );
  OAI21_X1 U8602 ( .B1(n9361), .B2(n7311), .A(n7342), .ZN(n7343) );
  AOI21_X1 U8603 ( .B1(n9359), .B2(n9392), .A(n7343), .ZN(n7344) );
  OAI211_X1 U8604 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9348), .A(n7345), .B(
        n7344), .ZN(P2_U3158) );
  OAI21_X1 U8605 ( .B1(n7347), .B2(n8866), .A(n7346), .ZN(n7348) );
  INV_X1 U8606 ( .A(n7348), .ZN(n7506) );
  NAND2_X1 U8607 ( .A1(n7349), .A2(n8922), .ZN(n7350) );
  INV_X1 U8608 ( .A(n8866), .ZN(n8924) );
  NAND3_X1 U8609 ( .A1(n7350), .A2(n8924), .A3(n8921), .ZN(n7383) );
  INV_X1 U8610 ( .A(n7383), .ZN(n7352) );
  AOI21_X1 U8611 ( .B1(n7350), .B2(n8921), .A(n8924), .ZN(n7351) );
  NOR3_X1 U8612 ( .A1(n7352), .A2(n7351), .A3(n10713), .ZN(n7355) );
  OAI22_X1 U8613 ( .A1(n7353), .A2(n10763), .B1(n8002), .B2(n10741), .ZN(n7354) );
  NOR2_X1 U8614 ( .A1(n7355), .A2(n7354), .ZN(n7501) );
  NAND2_X1 U8615 ( .A1(n7356), .A2(n8009), .ZN(n7357) );
  AND2_X1 U8616 ( .A1(n7385), .A2(n7357), .ZN(n7504) );
  AOI22_X1 U8617 ( .A1(n7504), .A2(n10672), .B1(n11127), .B2(n8009), .ZN(n7358) );
  OAI211_X1 U8618 ( .C1(n10770), .C2(n7506), .A(n7501), .B(n7358), .ZN(n7360)
         );
  NAND2_X1 U8619 ( .A1(n7360), .A2(n11181), .ZN(n7359) );
  OAI21_X1 U8620 ( .B1(n11181), .B2(n6910), .A(n7359), .ZN(P1_U3530) );
  INV_X1 U8621 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U8622 ( .A1(n7360), .A2(n11185), .ZN(n7361) );
  OAI21_X1 U8623 ( .B1(n11185), .B2(n7362), .A(n7361), .ZN(P1_U3477) );
  INV_X1 U8624 ( .A(n8547), .ZN(n7394) );
  NAND2_X1 U8625 ( .A1(n7364), .A2(n7363), .ZN(n7365) );
  NAND2_X1 U8626 ( .A1(n7365), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7366) );
  XNOR2_X1 U8627 ( .A(n7366), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9457) );
  INV_X1 U8628 ( .A(n9457), .ZN(n8396) );
  INV_X1 U8629 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7367) );
  OAI222_X1 U8630 ( .A1(n9804), .A2(n7394), .B1(n8396), .B2(P2_U3151), .C1(
        n7367), .C2(n8844), .ZN(P2_U3278) );
  INV_X1 U8631 ( .A(n10934), .ZN(n7368) );
  INV_X1 U8632 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10051) );
  OAI222_X1 U8633 ( .A1(P1_U3086), .A2(n7368), .B1(n9222), .B2(n8555), .C1(
        n10051), .C2(n9220), .ZN(P1_U3337) );
  XNOR2_X1 U8634 ( .A(n7369), .B(n8928), .ZN(n7597) );
  INV_X1 U8635 ( .A(n7597), .ZN(n7380) );
  NAND2_X1 U8636 ( .A1(n10661), .A2(n10746), .ZN(n10583) );
  OAI21_X1 U8637 ( .B1(n7372), .B2(n7371), .A(n7370), .ZN(n7600) );
  NAND2_X1 U8638 ( .A1(n7600), .A2(n10651), .ZN(n7379) );
  AOI211_X1 U8639 ( .C1(n7744), .C2(n7386), .A(n10655), .B(n7512), .ZN(n7595)
         );
  INV_X1 U8640 ( .A(n7744), .ZN(n7373) );
  NOR2_X1 U8641 ( .A1(n7373), .A2(n10658), .ZN(n7377) );
  NAND2_X1 U8642 ( .A1(n7739), .A2(n10569), .ZN(n7375) );
  AOI22_X1 U8643 ( .A1(n7511), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7740), .B2(
        n10632), .ZN(n7374) );
  OAI211_X1 U8644 ( .C1(n10349), .C2(n10572), .A(n7375), .B(n7374), .ZN(n7376)
         );
  AOI211_X1 U8645 ( .C1(n7595), .C2(n10664), .A(n7377), .B(n7376), .ZN(n7378)
         );
  OAI211_X1 U8646 ( .C1(n7380), .C2(n10583), .A(n7379), .B(n7378), .ZN(
        P1_U3283) );
  OAI21_X1 U8647 ( .B1(n7382), .B2(n8857), .A(n7381), .ZN(n7454) );
  INV_X1 U8648 ( .A(n7454), .ZN(n7393) );
  NAND2_X1 U8649 ( .A1(n7383), .A2(n8901), .ZN(n7384) );
  XNOR2_X1 U8650 ( .A(n7384), .B(n8857), .ZN(n7450) );
  INV_X1 U8651 ( .A(n10583), .ZN(n10529) );
  AOI21_X1 U8652 ( .B1(n7385), .B2(n7456), .A(n10655), .ZN(n7387) );
  AOI22_X1 U8653 ( .A1(n7387), .A2(n7386), .B1(n11155), .B2(n11157), .ZN(n7451) );
  AOI22_X1 U8654 ( .A1(n7511), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7870), .B2(
        n10632), .ZN(n7388) );
  OAI21_X1 U8655 ( .B1(n7868), .B2(n10488), .A(n7388), .ZN(n7389) );
  AOI21_X1 U8656 ( .B1(n7456), .B2(n10580), .A(n7389), .ZN(n7390) );
  OAI21_X1 U8657 ( .B1(n7451), .B2(n10576), .A(n7390), .ZN(n7391) );
  AOI21_X1 U8658 ( .B1(n7450), .B2(n10529), .A(n7391), .ZN(n7392) );
  OAI21_X1 U8659 ( .B1(n7393), .B2(n10638), .A(n7392), .ZN(P1_U3284) );
  INV_X1 U8660 ( .A(n10457), .ZN(n10439) );
  INV_X1 U8661 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10052) );
  OAI222_X1 U8662 ( .A1(P1_U3086), .A2(n10439), .B1(n9222), .B2(n7394), .C1(
        n10052), .C2(n9220), .ZN(P1_U3338) );
  INV_X1 U8663 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7398) );
  NAND2_X1 U8664 ( .A1(n7396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7397) );
  XNOR2_X1 U8665 ( .A(n7397), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8556) );
  OAI222_X1 U8666 ( .A1(n8844), .A2(n7398), .B1(n9486), .B2(P2_U3151), .C1(
        n9804), .C2(n8555), .ZN(P2_U3277) );
  NOR2_X1 U8667 ( .A1(n7399), .A2(n7400), .ZN(n7413) );
  NAND2_X1 U8668 ( .A1(n7399), .A2(n7400), .ZN(n7414) );
  OAI21_X1 U8669 ( .B1(n7413), .B2(n7416), .A(n7414), .ZN(n7404) );
  XNOR2_X1 U8670 ( .A(n7402), .B(n7401), .ZN(n7403) );
  XNOR2_X1 U8671 ( .A(n7404), .B(n7403), .ZN(n7412) );
  AOI22_X1 U8672 ( .A1(n9904), .A2(n7405), .B1(n10352), .B2(n9932), .ZN(n7411)
         );
  INV_X1 U8673 ( .A(n7406), .ZN(n7408) );
  NOR2_X1 U8674 ( .A1(n9877), .A2(n9912), .ZN(n7407) );
  AOI211_X1 U8675 ( .C1(n9917), .C2(n7409), .A(n7408), .B(n7407), .ZN(n7410)
         );
  OAI211_X1 U8676 ( .C1(n7412), .C2(n9919), .A(n7411), .B(n7410), .ZN(P1_U3239) );
  INV_X1 U8677 ( .A(n7413), .ZN(n7415) );
  NAND2_X1 U8678 ( .A1(n7415), .A2(n7414), .ZN(n7417) );
  XNOR2_X1 U8679 ( .A(n7417), .B(n7416), .ZN(n7426) );
  AOI22_X1 U8680 ( .A1(n9904), .A2(n7418), .B1(n10353), .B2(n9932), .ZN(n7425)
         );
  INV_X1 U8681 ( .A(n7419), .ZN(n7422) );
  NOR2_X1 U8682 ( .A1(n7420), .A2(n9912), .ZN(n7421) );
  AOI211_X1 U8683 ( .C1(n9917), .C2(n7423), .A(n7422), .B(n7421), .ZN(n7424)
         );
  OAI211_X1 U8684 ( .C1(n7426), .C2(n9919), .A(n7425), .B(n7424), .ZN(P1_U3227) );
  INV_X1 U8685 ( .A(n8469), .ZN(n8729) );
  NAND2_X1 U8686 ( .A1(n8729), .A2(n7427), .ZN(n7429) );
  NAND2_X1 U8687 ( .A1(n7311), .A2(n7428), .ZN(n8463) );
  NAND2_X1 U8688 ( .A1(n7565), .A2(n7562), .ZN(n8472) );
  INV_X1 U8689 ( .A(n7562), .ZN(n7698) );
  NAND2_X1 U8690 ( .A1(n9393), .A2(n7698), .ZN(n8480) );
  NAND2_X1 U8691 ( .A1(n8472), .A2(n8480), .ZN(n8724) );
  INV_X1 U8692 ( .A(n8724), .ZN(n7433) );
  NAND2_X1 U8693 ( .A1(n7430), .A2(n7433), .ZN(n7569) );
  OAI21_X1 U8694 ( .B1(n7430), .B2(n7433), .A(n7569), .ZN(n7692) );
  OAI22_X1 U8695 ( .A1(n8474), .A2(n9773), .B1(n7698), .B2(n9775), .ZN(n7435)
         );
  NAND2_X1 U8696 ( .A1(n7311), .A2(n11104), .ZN(n7431) );
  NAND2_X1 U8697 ( .A1(n7432), .A2(n7431), .ZN(n7564) );
  XNOR2_X1 U8698 ( .A(n7564), .B(n7433), .ZN(n7434) );
  OAI22_X1 U8699 ( .A1(n7434), .A2(n9689), .B1(n7311), .B2(n9687), .ZN(n7695)
         );
  AOI211_X1 U8700 ( .C1(n9779), .C2(n7692), .A(n7435), .B(n7695), .ZN(n11113)
         );
  NAND2_X1 U8701 ( .A1(n5132), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7436) );
  OAI21_X1 U8702 ( .B1(n11113), .B2(n5132), .A(n7436), .ZN(P2_U3462) );
  XNOR2_X1 U8703 ( .A(n7438), .B(n7437), .ZN(n7439) );
  XNOR2_X1 U8704 ( .A(n7440), .B(n7439), .ZN(n7448) );
  NOR2_X1 U8705 ( .A1(n11139), .A2(n9936), .ZN(n7447) );
  INV_X1 U8706 ( .A(n7441), .ZN(n7442) );
  AOI21_X1 U8707 ( .B1(n10353), .B2(n9928), .A(n7442), .ZN(n7445) );
  NAND2_X1 U8708 ( .A1(n9917), .A2(n7443), .ZN(n7444) );
  OAI211_X1 U8709 ( .C1(n7868), .C2(n9878), .A(n7445), .B(n7444), .ZN(n7446)
         );
  AOI211_X1 U8710 ( .C1(n7448), .C2(n9926), .A(n7447), .B(n7446), .ZN(n7449)
         );
  INV_X1 U8711 ( .A(n7449), .ZN(P1_U3213) );
  NAND2_X1 U8712 ( .A1(n7450), .A2(n10746), .ZN(n7452) );
  OAI211_X1 U8713 ( .C1(n7868), .C2(n10763), .A(n7452), .B(n7451), .ZN(n7453)
         );
  AOI21_X1 U8714 ( .B1(n11178), .B2(n7454), .A(n7453), .ZN(n7460) );
  INV_X1 U8715 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7632) );
  AOI22_X1 U8716 ( .A1(n7456), .A2(n7604), .B1(n11180), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7455) );
  OAI21_X1 U8717 ( .B1(n7460), .B2(n11180), .A(n7455), .ZN(P1_U3531) );
  INV_X1 U8718 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7457) );
  OAI22_X1 U8719 ( .A1(n5434), .A2(n10806), .B1(n11185), .B2(n7457), .ZN(n7458) );
  INV_X1 U8720 ( .A(n7458), .ZN(n7459) );
  OAI21_X1 U8721 ( .B1(n7460), .B2(n11182), .A(n7459), .ZN(P1_U3480) );
  NOR2_X1 U8722 ( .A1(n9377), .A2(P2_U3151), .ZN(n7498) );
  INV_X1 U8723 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7685) );
  OAI22_X1 U8724 ( .A1(n9375), .A2(n7486), .B1(n9380), .B2(n7686), .ZN(n7461)
         );
  AOI21_X1 U8725 ( .B1(n9370), .B2(n8728), .A(n7461), .ZN(n7462) );
  OAI21_X1 U8726 ( .B1(n7498), .B2(n7685), .A(n7462), .ZN(P2_U3172) );
  NOR2_X1 U8727 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7463) );
  AOI21_X1 U8728 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7463), .ZN(n10882) );
  NOR2_X1 U8729 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7464) );
  AOI21_X1 U8730 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7464), .ZN(n10879) );
  NOR2_X1 U8731 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7465) );
  AOI21_X1 U8732 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7465), .ZN(n10876) );
  NOR2_X1 U8733 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7466) );
  AOI21_X1 U8734 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7466), .ZN(n10873) );
  NOR2_X1 U8735 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7467) );
  AOI21_X1 U8736 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7467), .ZN(n10870) );
  NOR2_X1 U8737 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7468) );
  AOI21_X1 U8738 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7468), .ZN(n10867) );
  NOR2_X1 U8739 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7469) );
  AOI21_X1 U8740 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7469), .ZN(n10864) );
  NOR2_X1 U8741 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7470) );
  AOI21_X1 U8742 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7470), .ZN(n10861) );
  NOR2_X1 U8743 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7471) );
  AOI21_X1 U8744 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7471), .ZN(n10858) );
  NOR2_X1 U8745 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7472) );
  AOI21_X1 U8746 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7472), .ZN(n10855) );
  NOR2_X1 U8747 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7473) );
  AOI21_X1 U8748 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7473), .ZN(n10852) );
  NOR2_X1 U8749 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7474) );
  AOI21_X1 U8750 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7474), .ZN(n10849) );
  NOR2_X1 U8751 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7475) );
  AOI21_X1 U8752 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7475), .ZN(n10846) );
  NOR2_X1 U8753 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7476) );
  AOI21_X1 U8754 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7476), .ZN(n10843) );
  AND2_X1 U8755 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7477) );
  NOR2_X1 U8756 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7477), .ZN(n10829) );
  INV_X1 U8757 ( .A(n10829), .ZN(n10830) );
  INV_X1 U8758 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10992) );
  NAND3_X1 U8759 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U8760 ( .A1(n10992), .A2(n10831), .ZN(n10828) );
  NAND2_X1 U8761 ( .A1(n10830), .A2(n10828), .ZN(n10834) );
  NAND2_X1 U8762 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7478) );
  OAI21_X1 U8763 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7478), .ZN(n10833) );
  NOR2_X1 U8764 ( .A1(n10834), .A2(n10833), .ZN(n10832) );
  AOI21_X1 U8765 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10832), .ZN(n10837) );
  NAND2_X1 U8766 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7479) );
  OAI21_X1 U8767 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7479), .ZN(n10836) );
  NOR2_X1 U8768 ( .A1(n10837), .A2(n10836), .ZN(n10835) );
  AOI21_X1 U8769 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10835), .ZN(n10840) );
  NOR2_X1 U8770 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7480) );
  AOI21_X1 U8771 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7480), .ZN(n10839) );
  NAND2_X1 U8772 ( .A1(n10840), .A2(n10839), .ZN(n10838) );
  OAI21_X1 U8773 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10838), .ZN(n10842) );
  NAND2_X1 U8774 ( .A1(n10843), .A2(n10842), .ZN(n10841) );
  OAI21_X1 U8775 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10841), .ZN(n10845) );
  NAND2_X1 U8776 ( .A1(n10846), .A2(n10845), .ZN(n10844) );
  OAI21_X1 U8777 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10844), .ZN(n10848) );
  NAND2_X1 U8778 ( .A1(n10849), .A2(n10848), .ZN(n10847) );
  OAI21_X1 U8779 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10847), .ZN(n10851) );
  NAND2_X1 U8780 ( .A1(n10852), .A2(n10851), .ZN(n10850) );
  OAI21_X1 U8781 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10850), .ZN(n10854) );
  NAND2_X1 U8782 ( .A1(n10855), .A2(n10854), .ZN(n10853) );
  OAI21_X1 U8783 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10853), .ZN(n10857) );
  NAND2_X1 U8784 ( .A1(n10858), .A2(n10857), .ZN(n10856) );
  OAI21_X1 U8785 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10856), .ZN(n10860) );
  NAND2_X1 U8786 ( .A1(n10861), .A2(n10860), .ZN(n10859) );
  OAI21_X1 U8787 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10859), .ZN(n10863) );
  NAND2_X1 U8788 ( .A1(n10864), .A2(n10863), .ZN(n10862) );
  OAI21_X1 U8789 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10862), .ZN(n10866) );
  NAND2_X1 U8790 ( .A1(n10867), .A2(n10866), .ZN(n10865) );
  OAI21_X1 U8791 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10865), .ZN(n10869) );
  NAND2_X1 U8792 ( .A1(n10870), .A2(n10869), .ZN(n10868) );
  OAI21_X1 U8793 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10868), .ZN(n10872) );
  NAND2_X1 U8794 ( .A1(n10873), .A2(n10872), .ZN(n10871) );
  OAI21_X1 U8795 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10871), .ZN(n10875) );
  NAND2_X1 U8796 ( .A1(n10876), .A2(n10875), .ZN(n10874) );
  OAI21_X1 U8797 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10874), .ZN(n10878) );
  NAND2_X1 U8798 ( .A1(n10879), .A2(n10878), .ZN(n10877) );
  OAI21_X1 U8799 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10877), .ZN(n10881) );
  NAND2_X1 U8800 ( .A1(n10882), .A2(n10881), .ZN(n10880) );
  OAI21_X1 U8801 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10880), .ZN(n7482) );
  XNOR2_X1 U8802 ( .A(n5639), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7481) );
  XNOR2_X1 U8803 ( .A(n7482), .B(n7481), .ZN(ADD_1068_U4) );
  OAI21_X1 U8804 ( .B1(n7484), .B2(n7483), .A(n7323), .ZN(n7485) );
  NAND2_X1 U8805 ( .A1(n7485), .A2(n9370), .ZN(n7489) );
  OAI22_X1 U8806 ( .A1(n9361), .A2(n7486), .B1(n11104), .B2(n9380), .ZN(n7487)
         );
  AOI21_X1 U8807 ( .B1(n9359), .B2(n9393), .A(n7487), .ZN(n7488) );
  OAI211_X1 U8808 ( .C1(n7498), .C2(n11106), .A(n7489), .B(n7488), .ZN(
        P2_U3177) );
  INV_X1 U8809 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7497) );
  OAI21_X1 U8810 ( .B1(n7492), .B2(n7491), .A(n7490), .ZN(n7493) );
  NAND2_X1 U8811 ( .A1(n7493), .A2(n9370), .ZN(n7496) );
  OAI22_X1 U8812 ( .A1(n9361), .A2(n7494), .B1(n7304), .B2(n9380), .ZN(n7495)
         );
  OAI211_X1 U8813 ( .C1(n7498), .C2(n7497), .A(n7496), .B(n5233), .ZN(P2_U3162) );
  INV_X1 U8814 ( .A(n8009), .ZN(n7500) );
  AOI22_X1 U8815 ( .A1(n7511), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7999), .B2(
        n10632), .ZN(n7499) );
  OAI21_X1 U8816 ( .B1(n7500), .B2(n10658), .A(n7499), .ZN(n7503) );
  NOR2_X1 U8817 ( .A1(n7501), .A2(n7511), .ZN(n7502) );
  AOI211_X1 U8818 ( .C1(n7504), .C2(n10480), .A(n7503), .B(n7502), .ZN(n7505)
         );
  OAI21_X1 U8819 ( .B1(n7506), .B2(n10638), .A(n7505), .ZN(P1_U3285) );
  INV_X1 U8820 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U8821 ( .A1(n9933), .A2(P1_U3973), .ZN(n7507) );
  OAI21_X1 U8822 ( .B1(n8332), .B2(P1_U3973), .A(n7507), .ZN(P1_U3581) );
  XNOR2_X1 U8823 ( .A(n7508), .B(n8872), .ZN(n11163) );
  INV_X1 U8824 ( .A(n11163), .ZN(n11167) );
  INV_X1 U8825 ( .A(n7664), .ZN(n7509) );
  AOI211_X1 U8826 ( .C1(n8872), .C2(n7510), .A(n10713), .B(n7509), .ZN(n11161)
         );
  INV_X1 U8827 ( .A(n7511), .ZN(n10601) );
  OAI211_X1 U8828 ( .C1(n7512), .C2(n11160), .A(n10672), .B(n7669), .ZN(n11159) );
  AOI22_X1 U8829 ( .A1(n7511), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7816), .B2(
        n10632), .ZN(n7514) );
  NAND2_X1 U8830 ( .A1(n8272), .A2(n11154), .ZN(n7513) );
  OAI211_X1 U8831 ( .C1(n7515), .C2(n10488), .A(n7514), .B(n7513), .ZN(n7516)
         );
  AOI21_X1 U8832 ( .B1(n7821), .B2(n10580), .A(n7516), .ZN(n7517) );
  OAI21_X1 U8833 ( .B1(n11159), .B2(n10576), .A(n7517), .ZN(n7518) );
  AOI21_X1 U8834 ( .B1(n11161), .B2(n10601), .A(n7518), .ZN(n7519) );
  OAI21_X1 U8835 ( .B1(n11167), .B2(n7520), .A(n7519), .ZN(P1_U3282) );
  NAND2_X1 U8836 ( .A1(n7523), .A2(n7522), .ZN(n7705) );
  NAND2_X1 U8837 ( .A1(n7313), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7526) );
  NAND2_X1 U8838 ( .A1(n7534), .A2(n11034), .ZN(n7525) );
  INV_X1 U8839 ( .A(n11117), .ZN(n7708) );
  XNOR2_X1 U8840 ( .A(n7708), .B(n7528), .ZN(n7529) );
  NAND2_X1 U8841 ( .A1(n7529), .A2(n8474), .ZN(n7530) );
  OAI21_X1 U8842 ( .B1(n7529), .B2(n8474), .A(n7530), .ZN(n7704) );
  INV_X1 U8843 ( .A(n7530), .ZN(n7531) );
  NAND2_X1 U8844 ( .A1(n7313), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7538) );
  NAND2_X1 U8845 ( .A1(n5140), .A2(n7533), .ZN(n7537) );
  NAND2_X1 U8846 ( .A1(n7534), .A2(n7535), .ZN(n7536) );
  XNOR2_X1 U8847 ( .A(n7528), .B(n7723), .ZN(n7573) );
  NAND2_X1 U8848 ( .A1(n7155), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7545) );
  NAND2_X1 U8849 ( .A1(n7539), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U8850 ( .A1(n7156), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7543) );
  NAND2_X1 U8851 ( .A1(n7540), .A2(n10210), .ZN(n7550) );
  OR2_X1 U8852 ( .A1(n10210), .A2(n7540), .ZN(n7541) );
  AND2_X1 U8853 ( .A1(n7550), .A2(n7541), .ZN(n7722) );
  OR2_X1 U8854 ( .A1(n8037), .A2(n7722), .ZN(n7542) );
  NAND4_X1 U8855 ( .A1(n7545), .A2(n7544), .A3(n7543), .A4(n7542), .ZN(n9391)
         );
  XNOR2_X1 U8856 ( .A(n7573), .B(n7848), .ZN(n7546) );
  AOI21_X1 U8857 ( .B1(n7547), .B2(n7546), .A(n7581), .ZN(n7561) );
  NAND2_X1 U8858 ( .A1(n7155), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7555) );
  INV_X1 U8859 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7549) );
  OR2_X1 U8860 ( .A1(n7548), .A2(n7549), .ZN(n7554) );
  NAND2_X1 U8861 ( .A1(n7550), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7551) );
  AND2_X1 U8862 ( .A1(n7584), .A2(n7551), .ZN(n7852) );
  OR2_X1 U8863 ( .A1(n8037), .A2(n7852), .ZN(n7553) );
  INV_X1 U8864 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7851) );
  OR2_X1 U8865 ( .A1(n8711), .A2(n7851), .ZN(n7552) );
  NAND2_X1 U8866 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n11057) );
  INV_X1 U8867 ( .A(n11057), .ZN(n7556) );
  AOI21_X1 U8868 ( .B1(n9327), .B2(n7787), .A(n7556), .ZN(n7557) );
  OAI21_X1 U8869 ( .B1(n9361), .B2(n8474), .A(n7557), .ZN(n7559) );
  NOR2_X1 U8870 ( .A1(n9348), .A2(n7722), .ZN(n7558) );
  AOI211_X1 U8871 ( .C1(n9359), .C2(n9390), .A(n7559), .B(n7558), .ZN(n7560)
         );
  OAI21_X1 U8872 ( .B1(n7561), .B2(n9330), .A(n7560), .ZN(P2_U3167) );
  XNOR2_X1 U8873 ( .A(n9392), .B(n11117), .ZN(n8730) );
  NAND2_X1 U8874 ( .A1(n9393), .A2(n7562), .ZN(n7563) );
  NAND2_X1 U8875 ( .A1(n7564), .A2(n7563), .ZN(n7567) );
  NAND2_X1 U8876 ( .A1(n7565), .A2(n7698), .ZN(n7566) );
  NAND2_X1 U8877 ( .A1(n7567), .A2(n7566), .ZN(n7657) );
  XOR2_X1 U8878 ( .A(n8730), .B(n7657), .Z(n7568) );
  AOI222_X1 U8879 ( .A1(n9643), .A2(n7568), .B1(n9391), .B2(n7160), .C1(n9393), 
        .C2(n7162), .ZN(n11123) );
  NAND2_X1 U8880 ( .A1(n7569), .A2(n8472), .ZN(n7650) );
  XNOR2_X1 U8881 ( .A(n7650), .B(n8730), .ZN(n11121) );
  AOI22_X1 U8882 ( .A1(n11121), .A2(n9779), .B1(n9754), .B2(n11117), .ZN(n7570) );
  AND2_X1 U8883 ( .A1(n11123), .A2(n7570), .ZN(n11115) );
  OR2_X1 U8884 ( .A1(n8232), .A2(n7329), .ZN(n7571) );
  OAI21_X1 U8885 ( .B1(n11115), .B2(n5132), .A(n7571), .ZN(P2_U3463) );
  INV_X1 U8886 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7572) );
  INV_X1 U8887 ( .A(n8577), .ZN(n9218) );
  OAI222_X1 U8888 ( .A1(n8844), .A2(n7572), .B1(n9800), .B2(n9218), .C1(
        P2_U3151), .C2(n8787), .ZN(P2_U3276) );
  INV_X1 U8889 ( .A(n7573), .ZN(n7574) );
  NOR2_X1 U8890 ( .A1(n7574), .A2(n9391), .ZN(n7580) );
  NAND2_X1 U8891 ( .A1(n7313), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7577) );
  INV_X1 U8892 ( .A(n11061), .ZN(n7575) );
  NAND2_X1 U8893 ( .A1(n7534), .A2(n7575), .ZN(n7576) );
  OAI211_X1 U8894 ( .C1(n7524), .C2(n7578), .A(n7577), .B(n7576), .ZN(n7790)
         );
  INV_X1 U8895 ( .A(n7790), .ZN(n7910) );
  XNOR2_X1 U8896 ( .A(n7910), .B(n7528), .ZN(n7751) );
  XNOR2_X1 U8897 ( .A(n7751), .B(n7793), .ZN(n7579) );
  INV_X1 U8898 ( .A(n7752), .ZN(n7583) );
  OAI21_X1 U8899 ( .B1(n7581), .B2(n7580), .A(n7579), .ZN(n7582) );
  NAND3_X1 U8900 ( .A1(n7583), .A2(n9370), .A3(n7582), .ZN(n7594) );
  NAND2_X1 U8901 ( .A1(n7155), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7589) );
  OR2_X1 U8902 ( .A1(n7548), .A2(n7249), .ZN(n7588) );
  AND2_X1 U8903 ( .A1(n7584), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7585) );
  NOR2_X1 U8904 ( .A1(n7758), .A2(n7585), .ZN(n7804) );
  OR2_X1 U8905 ( .A1(n8037), .A2(n7804), .ZN(n7587) );
  OR2_X1 U8906 ( .A1(n8711), .A2(n7803), .ZN(n7586) );
  NAND2_X1 U8907 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n11074) );
  INV_X1 U8908 ( .A(n11074), .ZN(n7590) );
  AOI21_X1 U8909 ( .B1(n9327), .B2(n7790), .A(n7590), .ZN(n7591) );
  OAI21_X1 U8910 ( .B1(n9361), .B2(n7848), .A(n7591), .ZN(n7592) );
  AOI21_X1 U8911 ( .B1(n9359), .B2(n9389), .A(n7592), .ZN(n7593) );
  OAI211_X1 U8912 ( .C1(n7852), .C2(n9348), .A(n7594), .B(n7593), .ZN(P2_U3179) );
  OAI22_X1 U8913 ( .A1(n10349), .A2(n10741), .B1(n8002), .B2(n10763), .ZN(
        n7596) );
  AOI211_X1 U8914 ( .C1(n7597), .C2(n10746), .A(n7596), .B(n7595), .ZN(n7598)
         );
  INV_X1 U8915 ( .A(n7598), .ZN(n7599) );
  AOI21_X1 U8916 ( .B1(n7600), .B2(n11178), .A(n7599), .ZN(n7606) );
  INV_X1 U8917 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7601) );
  NOR2_X1 U8918 ( .A1(n11185), .A2(n7601), .ZN(n7602) );
  AOI21_X1 U8919 ( .B1(n7744), .B2(n6368), .A(n7602), .ZN(n7603) );
  OAI21_X1 U8920 ( .B1(n7606), .B2(n11182), .A(n7603), .ZN(P1_U3483) );
  INV_X1 U8921 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7630) );
  AOI22_X1 U8922 ( .A1(n7744), .A2(n7604), .B1(n11180), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7605) );
  OAI21_X1 U8923 ( .B1(n7606), .B2(n11180), .A(n7605), .ZN(P1_U3532) );
  NOR2_X1 U8924 ( .A1(n7747), .A2(n7607), .ZN(n7609) );
  INV_X1 U8925 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7610) );
  AOI22_X1 U8926 ( .A1(n7824), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7610), .B2(
        n7771), .ZN(n7611) );
  AOI21_X1 U8927 ( .B1(n5237), .B2(n7611), .A(n7768), .ZN(n7629) );
  NOR2_X1 U8928 ( .A1(n7747), .A2(n7612), .ZN(n7614) );
  INV_X1 U8929 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7896) );
  AOI22_X1 U8930 ( .A1(n7824), .A2(P2_REG1_REG_8__SCAN_IN), .B1(n7896), .B2(
        n7771), .ZN(n7615) );
  AOI21_X1 U8931 ( .B1(n5238), .B2(n7615), .A(n7770), .ZN(n7616) );
  NOR2_X1 U8932 ( .A1(n7616), .A2(n11090), .ZN(n7627) );
  MUX2_X1 U8933 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8795), .Z(n7617) );
  NOR2_X1 U8934 ( .A1(n7617), .A2(n7771), .ZN(n7776) );
  AOI21_X1 U8935 ( .B1(n7617), .B2(n7771), .A(n7776), .ZN(n7618) );
  INV_X1 U8936 ( .A(n7618), .ZN(n7622) );
  NOR2_X1 U8937 ( .A1(n7620), .A2(n7619), .ZN(n7621) );
  NOR2_X1 U8938 ( .A1(n7621), .A2(n7622), .ZN(n7775) );
  AOI21_X1 U8939 ( .B1(n7622), .B2(n7621), .A(n7775), .ZN(n7625) );
  AOI22_X1 U8940 ( .A1(n11033), .A2(n7824), .B1(n11076), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n7624) );
  NOR2_X1 U8941 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10196), .ZN(n7882) );
  INV_X1 U8942 ( .A(n7882), .ZN(n7623) );
  OAI211_X1 U8943 ( .C1(n7625), .C2(n11020), .A(n7624), .B(n7623), .ZN(n7626)
         );
  NOR2_X1 U8944 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  OAI21_X1 U8945 ( .B1(n7629), .B2(n11081), .A(n7628), .ZN(P2_U3190) );
  MUX2_X1 U8946 ( .A(n7630), .B(P1_REG1_REG_10__SCAN_IN), .S(n10963), .Z(
        n10958) );
  AOI21_X1 U8947 ( .B1(n7638), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7631), .ZN(
        n10393) );
  MUX2_X1 U8948 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7632), .S(n10397), .Z(n10392) );
  NAND2_X1 U8949 ( .A1(n10393), .A2(n10392), .ZN(n10391) );
  OAI21_X1 U8950 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10397), .A(n10391), .ZN(
        n10959) );
  NOR2_X1 U8951 ( .A1(n10958), .A2(n10959), .ZN(n10957) );
  AOI21_X1 U8952 ( .B1(n10963), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10957), .ZN(
        n10888) );
  INV_X1 U8953 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7633) );
  MUX2_X1 U8954 ( .A(n7633), .B(P1_REG1_REG_11__SCAN_IN), .S(n10891), .Z(
        n10887) );
  NOR2_X1 U8955 ( .A1(n10888), .A2(n10887), .ZN(n10886) );
  AOI21_X1 U8956 ( .B1(n10891), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10886), .ZN(
        n7636) );
  INV_X1 U8957 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7634) );
  MUX2_X1 U8958 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7634), .S(n10412), .Z(n7635) );
  NAND2_X1 U8959 ( .A1(n7635), .A2(n7636), .ZN(n10403) );
  OAI21_X1 U8960 ( .B1(n7636), .B2(n7635), .A(n10403), .ZN(n7645) );
  XOR2_X1 U8961 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10412), .Z(n10416) );
  NOR2_X1 U8962 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n10397), .ZN(n7639) );
  AOI21_X1 U8963 ( .B1(n10397), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7639), .ZN(
        n10389) );
  NAND2_X1 U8964 ( .A1(n10388), .A2(n10389), .ZN(n10387) );
  OAI21_X1 U8965 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n10397), .A(n10387), .ZN(
        n10955) );
  INV_X1 U8966 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7641) );
  AOI22_X1 U8967 ( .A1(n10963), .A2(n7641), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7640), .ZN(n10954) );
  NOR2_X1 U8968 ( .A1(n10955), .A2(n10954), .ZN(n10953) );
  INV_X1 U8969 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7642) );
  AOI22_X1 U8970 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7643), .B1(n10891), .B2(
        n7642), .ZN(n10884) );
  NOR2_X1 U8971 ( .A1(n10885), .A2(n10884), .ZN(n10883) );
  XNOR2_X1 U8972 ( .A(n10416), .B(n10415), .ZN(n7644) );
  AOI22_X1 U8973 ( .A1(n10910), .A2(n7645), .B1(n10916), .B2(n7644), .ZN(n7649) );
  INV_X1 U8974 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7646) );
  NAND2_X1 U8975 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8071) );
  OAI21_X1 U8976 ( .B1(n10967), .B2(n7646), .A(n8071), .ZN(n7647) );
  AOI21_X1 U8977 ( .B1(n10412), .B2(n10962), .A(n7647), .ZN(n7648) );
  NAND2_X1 U8978 ( .A1(n7649), .A2(n7648), .ZN(P1_U3255) );
  NAND2_X1 U8979 ( .A1(n7650), .A2(n8730), .ZN(n7652) );
  NOR2_X1 U8980 ( .A1(n9392), .A2(n7708), .ZN(n8479) );
  INV_X1 U8981 ( .A(n8479), .ZN(n7651) );
  NAND2_X1 U8982 ( .A1(n7652), .A2(n7651), .ZN(n7796) );
  NAND2_X1 U8983 ( .A1(n7848), .A2(n7787), .ZN(n8477) );
  NAND2_X1 U8984 ( .A1(n9391), .A2(n7723), .ZN(n8481) );
  NAND2_X1 U8985 ( .A1(n8477), .A2(n8481), .ZN(n8723) );
  XNOR2_X1 U8986 ( .A(n7796), .B(n8723), .ZN(n7728) );
  AOI21_X1 U8987 ( .B1(n7654), .B2(n7653), .A(n7728), .ZN(n7660) );
  NOR2_X1 U8988 ( .A1(n9392), .A2(n11117), .ZN(n7656) );
  NAND2_X1 U8989 ( .A1(n9392), .A2(n11117), .ZN(n7655) );
  XNOR2_X1 U8990 ( .A(n7789), .B(n8723), .ZN(n7658) );
  OAI22_X1 U8991 ( .A1(n7658), .A2(n9689), .B1(n8474), .B2(n9687), .ZN(n7721)
         );
  OAI22_X1 U8992 ( .A1(n7793), .A2(n9773), .B1(n7723), .B2(n9775), .ZN(n7659)
         );
  NOR3_X1 U8993 ( .A1(n7660), .A2(n7721), .A3(n7659), .ZN(n11126) );
  NAND2_X1 U8994 ( .A1(n5132), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7661) );
  OAI21_X1 U8995 ( .B1(n11126), .B2(n5132), .A(n7661), .ZN(P2_U3464) );
  XOR2_X1 U8996 ( .A(n8870), .B(n7662), .Z(n11179) );
  INV_X1 U8997 ( .A(n11179), .ZN(n7676) );
  INV_X1 U8998 ( .A(n8870), .ZN(n7663) );
  NAND3_X1 U8999 ( .A1(n7664), .A2(n8931), .A3(n7663), .ZN(n7665) );
  NAND3_X1 U9000 ( .A1(n7666), .A2(n10746), .A3(n7665), .ZN(n7668) );
  NAND2_X1 U9001 ( .A1(n10348), .A2(n11155), .ZN(n7667) );
  OAI211_X1 U9002 ( .C1(n10349), .C2(n10763), .A(n7668), .B(n7667), .ZN(n11177) );
  INV_X1 U9003 ( .A(n7669), .ZN(n7670) );
  INV_X1 U9004 ( .A(n7671), .ZN(n11175) );
  OAI211_X1 U9005 ( .C1(n7670), .C2(n11175), .A(n10672), .B(n7902), .ZN(n11173) );
  AOI22_X1 U9006 ( .A1(n7511), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8073), .B2(
        n10632), .ZN(n7673) );
  NAND2_X1 U9007 ( .A1(n7671), .A2(n10580), .ZN(n7672) );
  OAI211_X1 U9008 ( .C1(n11173), .C2(n10576), .A(n7673), .B(n7672), .ZN(n7674)
         );
  AOI21_X1 U9009 ( .B1(n11177), .B2(n10661), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9010 ( .B1(n7676), .B2(n10638), .A(n7675), .ZN(P1_U3281) );
  NAND2_X1 U9011 ( .A1(n7677), .A2(n7176), .ZN(n7680) );
  OAI22_X1 U9012 ( .A1(n7681), .A2(n7680), .B1(n7679), .B2(n7678), .ZN(n7683)
         );
  NAND2_X1 U9013 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  INV_X2 U9014 ( .A(n11124), .ZN(n9692) );
  NAND2_X1 U9015 ( .A1(n9692), .A2(n7160), .ZN(n9678) );
  OAI22_X1 U9016 ( .A1(n9662), .A2(n7686), .B1(n7685), .B2(n11105), .ZN(n7690)
         );
  NAND4_X1 U9017 ( .A1(n8728), .A2(n7687), .A3(n9775), .A4(n9692), .ZN(n7688)
         );
  OAI21_X1 U9018 ( .B1(n7214), .B2(n9692), .A(n7688), .ZN(n7689) );
  AOI211_X1 U9019 ( .C1(n9695), .C2(n7305), .A(n7690), .B(n7689), .ZN(n7691)
         );
  INV_X1 U9020 ( .A(n7691), .ZN(P2_U3233) );
  INV_X1 U9021 ( .A(n7692), .ZN(n7702) );
  NAND2_X1 U9022 ( .A1(n7693), .A2(n7189), .ZN(n9210) );
  INV_X1 U9023 ( .A(n9210), .ZN(n11110) );
  OR2_X1 U9024 ( .A1(n9203), .A2(n11110), .ZN(n7694) );
  INV_X1 U9025 ( .A(n7695), .ZN(n7696) );
  MUX2_X1 U9026 ( .A(n7697), .B(n7696), .S(n9692), .Z(n7701) );
  OAI22_X1 U9027 ( .A1(n9662), .A2(n7698), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n11105), .ZN(n7699) );
  AOI21_X1 U9028 ( .B1(n9695), .B2(n9392), .A(n7699), .ZN(n7700) );
  OAI211_X1 U9029 ( .C1(n7702), .C2(n9698), .A(n7701), .B(n7700), .ZN(P2_U3230) );
  AOI21_X1 U9030 ( .B1(n7705), .B2(n7704), .A(n7703), .ZN(n7713) );
  INV_X1 U9031 ( .A(n7706), .ZN(n11119) );
  INV_X1 U9032 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7707) );
  NOR2_X1 U9033 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7707), .ZN(n11032) );
  NOR2_X1 U9034 ( .A1(n9380), .A2(n7708), .ZN(n7709) );
  AOI211_X1 U9035 ( .C1(n9373), .C2(n9393), .A(n11032), .B(n7709), .ZN(n7710)
         );
  OAI21_X1 U9036 ( .B1(n7848), .B2(n9375), .A(n7710), .ZN(n7711) );
  AOI21_X1 U9037 ( .B1(n11119), .B2(n9377), .A(n7711), .ZN(n7712) );
  OAI21_X1 U9038 ( .B1(n7713), .B2(n9330), .A(n7712), .ZN(P2_U3170) );
  INV_X1 U9039 ( .A(n7714), .ZN(n7720) );
  AOI22_X1 U9040 ( .A1(n11116), .A2(n7715), .B1(n11118), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7716) );
  OAI21_X1 U9041 ( .B1(n10976), .B2(n9692), .A(n7716), .ZN(n7717) );
  AOI21_X1 U9042 ( .B1(n11120), .B2(n7718), .A(n7717), .ZN(n7719) );
  OAI21_X1 U9043 ( .B1(n7720), .B2(n11124), .A(n7719), .ZN(P2_U3232) );
  NAND2_X1 U9044 ( .A1(n7721), .A2(n9692), .ZN(n7727) );
  NOR2_X1 U9045 ( .A1(n9692), .A2(n11052), .ZN(n7725) );
  OAI22_X1 U9046 ( .A1(n9662), .A2(n7723), .B1(n7722), .B2(n11105), .ZN(n7724)
         );
  AOI211_X1 U9047 ( .C1(n9695), .C2(n9390), .A(n7725), .B(n7724), .ZN(n7726)
         );
  OAI211_X1 U9048 ( .C1(n7728), .C2(n9698), .A(n7727), .B(n7726), .ZN(P2_U3228) );
  NAND2_X1 U9049 ( .A1(n8587), .A2(n10820), .ZN(n7730) );
  OAI211_X1 U9050 ( .C1(n10054), .C2(n9220), .A(n7730), .B(n7729), .ZN(
        P1_U3335) );
  INV_X1 U9051 ( .A(n8587), .ZN(n7733) );
  INV_X1 U9052 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7731) );
  OAI222_X1 U9053 ( .A1(n9804), .A2(n7733), .B1(n7732), .B2(P2_U3151), .C1(
        n7731), .C2(n8844), .ZN(P2_U3275) );
  NAND2_X1 U9054 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  XNOR2_X1 U9055 ( .A(n7737), .B(n7736), .ZN(n7746) );
  NAND2_X1 U9056 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10964) );
  INV_X1 U9057 ( .A(n10964), .ZN(n7738) );
  AOI21_X1 U9058 ( .B1(n7739), .B2(n9928), .A(n7738), .ZN(n7742) );
  NAND2_X1 U9059 ( .A1(n9917), .A2(n7740), .ZN(n7741) );
  OAI211_X1 U9060 ( .C1(n10349), .C2(n9878), .A(n7742), .B(n7741), .ZN(n7743)
         );
  AOI21_X1 U9061 ( .B1(n7744), .B2(n9904), .A(n7743), .ZN(n7745) );
  OAI21_X1 U9062 ( .B1(n7746), .B2(n9919), .A(n7745), .ZN(P1_U3217) );
  NAND2_X1 U9063 ( .A1(n7313), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U9064 ( .A1(n7534), .A2(n7747), .ZN(n7748) );
  OAI211_X1 U9065 ( .C1(n7524), .C2(n7750), .A(n7749), .B(n7748), .ZN(n7786)
         );
  XNOR2_X1 U9066 ( .A(n7528), .B(n7786), .ZN(n7875) );
  XNOR2_X1 U9067 ( .A(n7875), .B(n7911), .ZN(n7755) );
  INV_X1 U9068 ( .A(n7751), .ZN(n7753) );
  AOI21_X1 U9069 ( .B1(n9390), .B2(n7753), .A(n7752), .ZN(n7754) );
  NAND2_X1 U9070 ( .A1(n7754), .A2(n7755), .ZN(n7877) );
  OAI21_X1 U9071 ( .B1(n7755), .B2(n7754), .A(n7877), .ZN(n7756) );
  NAND2_X1 U9072 ( .A1(n7756), .A2(n9370), .ZN(n7767) );
  OR2_X1 U9073 ( .A1(n7548), .A2(n7896), .ZN(n7763) );
  NAND2_X1 U9074 ( .A1(n7155), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7762) );
  NOR2_X1 U9075 ( .A1(n7758), .A2(n10196), .ZN(n7759) );
  OR2_X1 U9076 ( .A1(n7836), .A2(n7759), .ZN(n7842) );
  NAND2_X1 U9077 ( .A1(n7757), .A2(n7842), .ZN(n7761) );
  OR2_X1 U9078 ( .A1(n8711), .A2(n7610), .ZN(n7760) );
  NAND4_X1 U9079 ( .A1(n7763), .A2(n7762), .A3(n7761), .A4(n7760), .ZN(n9388)
         );
  OAI22_X1 U9080 ( .A1(n9361), .A2(n7793), .B1(n8078), .B2(n9375), .ZN(n7764)
         );
  AOI211_X1 U9081 ( .C1(n7786), .C2(n9327), .A(n7765), .B(n7764), .ZN(n7766)
         );
  OAI211_X1 U9082 ( .C1(n7804), .C2(n9348), .A(n7767), .B(n7766), .ZN(P2_U3153) );
  INV_X1 U9083 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7952) );
  AOI21_X1 U9084 ( .B1(n7952), .B2(n7769), .A(n7976), .ZN(n7785) );
  INV_X1 U9085 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7773) );
  XNOR2_X1 U9086 ( .A(n7988), .B(n7989), .ZN(n7772) );
  AOI21_X1 U9087 ( .B1(n7773), .B2(n7772), .A(n7990), .ZN(n7774) );
  NOR2_X1 U9088 ( .A1(n7774), .A2(n11090), .ZN(n7783) );
  MUX2_X1 U9089 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8795), .Z(n7979) );
  XOR2_X1 U9090 ( .A(n7989), .B(n7979), .Z(n7778) );
  NOR2_X1 U9091 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  NOR2_X1 U9092 ( .A1(n7777), .A2(n7778), .ZN(n7980) );
  AOI21_X1 U9093 ( .B1(n7778), .B2(n7777), .A(n7980), .ZN(n7781) );
  AOI22_X1 U9094 ( .A1(n11033), .A2(n7989), .B1(n11076), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n7780) );
  NOR2_X1 U9095 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7835), .ZN(n7964) );
  INV_X1 U9096 ( .A(n7964), .ZN(n7779) );
  OAI211_X1 U9097 ( .C1(n7781), .C2(n11020), .A(n7780), .B(n7779), .ZN(n7782)
         );
  NOR2_X1 U9098 ( .A1(n7783), .A2(n7782), .ZN(n7784) );
  OAI21_X1 U9099 ( .B1(n7785), .B2(n11081), .A(n7784), .ZN(P2_U3191) );
  NAND2_X1 U9100 ( .A1(n7911), .A2(n7786), .ZN(n8443) );
  INV_X1 U9101 ( .A(n7786), .ZN(n8077) );
  AND2_X1 U9102 ( .A1(n9391), .A2(n7787), .ZN(n7788) );
  NAND2_X1 U9103 ( .A1(n7793), .A2(n7790), .ZN(n8475) );
  NAND2_X1 U9104 ( .A1(n9390), .A2(n7910), .ZN(n8483) );
  NAND2_X1 U9105 ( .A1(n8475), .A2(n8483), .ZN(n8726) );
  NAND2_X1 U9106 ( .A1(n7928), .A2(n8726), .ZN(n7791) );
  NAND2_X1 U9107 ( .A1(n7793), .A2(n7910), .ZN(n7830) );
  NAND2_X1 U9108 ( .A1(n7791), .A2(n7830), .ZN(n7792) );
  XOR2_X1 U9109 ( .A(n8727), .B(n7792), .Z(n7794) );
  OAI22_X1 U9110 ( .A1(n7794), .A2(n9689), .B1(n7793), .B2(n9687), .ZN(n8079)
         );
  INV_X1 U9111 ( .A(n8079), .ZN(n7810) );
  INV_X1 U9112 ( .A(n8723), .ZN(n7795) );
  NAND2_X1 U9113 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  NAND2_X1 U9114 ( .A1(n7797), .A2(n8477), .ZN(n7846) );
  NAND2_X1 U9115 ( .A1(n7846), .A2(n7847), .ZN(n7800) );
  AND2_X1 U9116 ( .A1(n7798), .A2(n8475), .ZN(n7799) );
  INV_X1 U9117 ( .A(n8081), .ZN(n7802) );
  NAND2_X1 U9118 ( .A1(n7800), .A2(n8475), .ZN(n7801) );
  AND2_X1 U9119 ( .A1(n7801), .A2(n8727), .ZN(n8076) );
  NOR3_X1 U9120 ( .A1(n7802), .A2(n8076), .A3(n9698), .ZN(n7808) );
  NOR2_X1 U9121 ( .A1(n9678), .A2(n8078), .ZN(n7807) );
  NOR2_X1 U9122 ( .A1(n9692), .A2(n7803), .ZN(n7806) );
  OAI22_X1 U9123 ( .A1(n9662), .A2(n8077), .B1(n7804), .B2(n11105), .ZN(n7805)
         );
  NOR4_X1 U9124 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n7809)
         );
  OAI21_X1 U9125 ( .B1(n11124), .B2(n7810), .A(n7809), .ZN(P2_U3226) );
  INV_X1 U9126 ( .A(n8599), .ZN(n7874) );
  AOI22_X1 U9127 ( .A1(n7189), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9802), .ZN(n7811) );
  OAI21_X1 U9128 ( .B1(n7874), .B2(n9800), .A(n7811), .ZN(P2_U3274) );
  NAND2_X1 U9129 ( .A1(n5231), .A2(n7813), .ZN(n7814) );
  XNOR2_X1 U9130 ( .A(n7812), .B(n7814), .ZN(n7823) );
  NAND2_X1 U9131 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10892) );
  INV_X1 U9132 ( .A(n10892), .ZN(n7815) );
  AOI21_X1 U9133 ( .B1(n11157), .B2(n9928), .A(n7815), .ZN(n7818) );
  NAND2_X1 U9134 ( .A1(n9917), .A2(n7816), .ZN(n7817) );
  OAI211_X1 U9135 ( .C1(n7819), .C2(n9878), .A(n7818), .B(n7817), .ZN(n7820)
         );
  AOI21_X1 U9136 ( .B1(n7821), .B2(n9904), .A(n7820), .ZN(n7822) );
  OAI21_X1 U9137 ( .B1(n7823), .B2(n9919), .A(n7822), .ZN(P1_U3236) );
  AOI22_X1 U9138 ( .A1(n7313), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7534), .B2(
        n7824), .ZN(n7827) );
  NAND2_X1 U9139 ( .A1(n7825), .A2(n5140), .ZN(n7826) );
  NAND2_X1 U9140 ( .A1(n8078), .A2(n7888), .ZN(n8446) );
  AND2_X1 U9141 ( .A1(n9388), .A2(n7931), .ZN(n8444) );
  INV_X1 U9142 ( .A(n8444), .ZN(n7939) );
  NAND2_X1 U9143 ( .A1(n8446), .A2(n7939), .ZN(n8733) );
  NAND2_X1 U9144 ( .A1(n8081), .A2(n7940), .ZN(n7828) );
  XOR2_X1 U9145 ( .A(n8733), .B(n7828), .Z(n7891) );
  NAND2_X1 U9146 ( .A1(n7911), .A2(n8077), .ZN(n7829) );
  AND2_X1 U9147 ( .A1(n8726), .A2(n7831), .ZN(n7926) );
  NAND2_X1 U9148 ( .A1(n7928), .A2(n7926), .ZN(n7832) );
  NAND2_X1 U9149 ( .A1(n7832), .A2(n7929), .ZN(n7833) );
  XNOR2_X1 U9150 ( .A(n7833), .B(n8733), .ZN(n7834) );
  AOI22_X1 U9151 ( .A1(n7834), .A2(n9643), .B1(n7162), .B2(n9389), .ZN(n7890)
         );
  MUX2_X1 U9152 ( .A(n7610), .B(n7890), .S(n9692), .Z(n7845) );
  NAND2_X1 U9153 ( .A1(n7155), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U9154 ( .A1(n7156), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U9155 ( .A1(n7539), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U9156 ( .A1(n7836), .A2(n7835), .ZN(n7946) );
  OR2_X1 U9157 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  AND2_X1 U9158 ( .A1(n7946), .A2(n7837), .ZN(n7963) );
  OR2_X1 U9159 ( .A1(n8037), .A2(n7963), .ZN(n7838) );
  NAND4_X1 U9160 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n9387)
         );
  INV_X1 U9161 ( .A(n7842), .ZN(n7884) );
  OAI22_X1 U9162 ( .A1(n9678), .A2(n8181), .B1(n7884), .B2(n11105), .ZN(n7843)
         );
  AOI21_X1 U9163 ( .B1(n11116), .B2(n7888), .A(n7843), .ZN(n7844) );
  OAI211_X1 U9164 ( .C1(n7891), .C2(n9698), .A(n7845), .B(n7844), .ZN(P2_U3225) );
  XNOR2_X1 U9165 ( .A(n7846), .B(n7847), .ZN(n7914) );
  INV_X1 U9166 ( .A(n7914), .ZN(n7856) );
  XNOR2_X1 U9167 ( .A(n7928), .B(n7847), .ZN(n7849) );
  OAI22_X1 U9168 ( .A1(n7849), .A2(n9689), .B1(n7848), .B2(n9687), .ZN(n7912)
         );
  INV_X1 U9169 ( .A(n7912), .ZN(n7850) );
  MUX2_X1 U9170 ( .A(n7851), .B(n7850), .S(n9692), .Z(n7855) );
  OAI22_X1 U9171 ( .A1(n9662), .A2(n7910), .B1(n7852), .B2(n11105), .ZN(n7853)
         );
  AOI21_X1 U9172 ( .B1(n9695), .B2(n9389), .A(n7853), .ZN(n7854) );
  OAI211_X1 U9173 ( .C1(n9698), .C2(n7856), .A(n7855), .B(n7854), .ZN(P2_U3227) );
  INV_X1 U9174 ( .A(n7857), .ZN(n7859) );
  NAND2_X1 U9175 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  OAI21_X1 U9176 ( .B1(n7859), .B2(n7858), .A(n7860), .ZN(n8004) );
  NOR2_X1 U9177 ( .A1(n8004), .A2(n8005), .ZN(n8003) );
  INV_X1 U9178 ( .A(n7860), .ZN(n7861) );
  NOR3_X1 U9179 ( .A1(n8003), .A2(n7862), .A3(n7861), .ZN(n7865) );
  INV_X1 U9180 ( .A(n7863), .ZN(n7864) );
  OAI21_X1 U9181 ( .B1(n7865), .B2(n7864), .A(n9926), .ZN(n7872) );
  NOR2_X1 U9182 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7866), .ZN(n10395) );
  AOI21_X1 U9183 ( .B1(n11157), .B2(n9932), .A(n10395), .ZN(n7867) );
  OAI21_X1 U9184 ( .B1(n7868), .B2(n9912), .A(n7867), .ZN(n7869) );
  AOI21_X1 U9185 ( .B1(n7870), .B2(n9917), .A(n7869), .ZN(n7871) );
  OAI211_X1 U9186 ( .C1(n5434), .C2(n9936), .A(n7872), .B(n7871), .ZN(P1_U3231) );
  OAI222_X1 U9187 ( .A1(P1_U3086), .A2(n9054), .B1(n9222), .B2(n7874), .C1(
        n7873), .C2(n9220), .ZN(P1_U3334) );
  NAND2_X1 U9188 ( .A1(n7877), .A2(n7876), .ZN(n7960) );
  XNOR2_X1 U9189 ( .A(n9158), .B(n7931), .ZN(n7878) );
  NOR2_X1 U9190 ( .A1(n7878), .A2(n9388), .ZN(n7959) );
  INV_X1 U9191 ( .A(n7959), .ZN(n7879) );
  NAND2_X1 U9192 ( .A1(n7878), .A2(n9388), .ZN(n7958) );
  NAND2_X1 U9193 ( .A1(n7879), .A2(n7958), .ZN(n7880) );
  XNOR2_X1 U9194 ( .A(n7960), .B(n7880), .ZN(n7887) );
  NOR2_X1 U9195 ( .A1(n9375), .A2(n8181), .ZN(n7881) );
  AOI211_X1 U9196 ( .C1(n9373), .C2(n9389), .A(n7882), .B(n7881), .ZN(n7883)
         );
  OAI21_X1 U9197 ( .B1(n7884), .B2(n9348), .A(n7883), .ZN(n7885) );
  AOI21_X1 U9198 ( .B1(n7888), .B2(n9327), .A(n7885), .ZN(n7886) );
  OAI21_X1 U9199 ( .B1(n7887), .B2(n9330), .A(n7886), .ZN(P2_U3161) );
  INV_X1 U9200 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7893) );
  AOI22_X1 U9201 ( .A1(n9754), .A2(n7888), .B1(n9387), .B2(n7160), .ZN(n7889)
         );
  OAI211_X1 U9202 ( .C1(n7891), .C2(n9752), .A(n7890), .B(n7889), .ZN(n7894)
         );
  NAND2_X1 U9203 ( .A1(n7894), .A2(n11195), .ZN(n7892) );
  OAI21_X1 U9204 ( .B1(n7893), .B2(n11195), .A(n7892), .ZN(P2_U3414) );
  NAND2_X1 U9205 ( .A1(n7894), .A2(n8232), .ZN(n7895) );
  OAI21_X1 U9206 ( .B1(n8232), .B2(n7896), .A(n7895), .ZN(P2_U3467) );
  INV_X1 U9207 ( .A(n8051), .ZN(n7897) );
  AOI21_X1 U9208 ( .B1(n8873), .B2(n7898), .A(n7897), .ZN(n7918) );
  XOR2_X1 U9209 ( .A(n7899), .B(n8873), .Z(n7920) );
  NAND2_X1 U9210 ( .A1(n7920), .A2(n10651), .ZN(n7909) );
  AOI22_X1 U9211 ( .A1(n7511), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8156), .B2(
        n10632), .ZN(n7901) );
  NAND2_X1 U9212 ( .A1(n10569), .A2(n11154), .ZN(n7900) );
  OAI211_X1 U9213 ( .C1(n10764), .C2(n10572), .A(n7901), .B(n7900), .ZN(n7906)
         );
  INV_X1 U9214 ( .A(n7902), .ZN(n7904) );
  INV_X1 U9215 ( .A(n8059), .ZN(n7903) );
  OAI211_X1 U9216 ( .C1(n8159), .C2(n7904), .A(n7903), .B(n10672), .ZN(n7916)
         );
  NOR2_X1 U9217 ( .A1(n7916), .A2(n10576), .ZN(n7905) );
  AOI211_X1 U9218 ( .C1(n10580), .C2(n7907), .A(n7906), .B(n7905), .ZN(n7908)
         );
  OAI211_X1 U9219 ( .C1(n7918), .C2(n10583), .A(n7909), .B(n7908), .ZN(
        P1_U3280) );
  OAI22_X1 U9220 ( .A1(n7911), .A2(n9773), .B1(n7910), .B2(n9775), .ZN(n7913)
         );
  AOI211_X1 U9221 ( .C1(n7914), .C2(n9779), .A(n7913), .B(n7912), .ZN(n11137)
         );
  OR2_X1 U9222 ( .A1(n11137), .A2(n5132), .ZN(n7915) );
  OAI21_X1 U9223 ( .B1(n8232), .B2(n7549), .A(n7915), .ZN(P2_U3465) );
  INV_X1 U9224 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7921) );
  INV_X1 U9225 ( .A(n10764), .ZN(n10347) );
  AOI22_X1 U9226 ( .A1(n10347), .A2(n11155), .B1(n11156), .B2(n11154), .ZN(
        n7917) );
  OAI211_X1 U9227 ( .C1(n7918), .C2(n10713), .A(n7917), .B(n7916), .ZN(n7919)
         );
  AOI21_X1 U9228 ( .B1(n7920), .B2(n11178), .A(n7919), .ZN(n7923) );
  MUX2_X1 U9229 ( .A(n7921), .B(n7923), .S(n11181), .Z(n7922) );
  OAI21_X1 U9230 ( .B1(n8159), .B2(n10739), .A(n7922), .ZN(P1_U3535) );
  INV_X1 U9231 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7924) );
  MUX2_X1 U9232 ( .A(n7924), .B(n7923), .S(n11185), .Z(n7925) );
  OAI21_X1 U9233 ( .B1(n8159), .B2(n10806), .A(n7925), .ZN(P1_U3492) );
  AND2_X1 U9234 ( .A1(n7926), .A2(n8733), .ZN(n7927) );
  NAND2_X1 U9235 ( .A1(n7928), .A2(n7927), .ZN(n7933) );
  INV_X1 U9236 ( .A(n8733), .ZN(n7930) );
  NAND2_X1 U9237 ( .A1(n8078), .A2(n7931), .ZN(n7932) );
  NAND2_X1 U9238 ( .A1(n7934), .A2(n5140), .ZN(n7936) );
  AOI22_X1 U9239 ( .A1(n7313), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7534), .B2(
        n7989), .ZN(n7935) );
  AND2_X1 U9240 ( .A1(n8024), .A2(n9387), .ZN(n8445) );
  INV_X1 U9241 ( .A(n8445), .ZN(n8089) );
  INV_X1 U9242 ( .A(n8024), .ZN(n7937) );
  NAND2_X1 U9243 ( .A1(n8181), .A2(n7937), .ZN(n8451) );
  NAND2_X1 U9244 ( .A1(n8089), .A2(n8451), .ZN(n8735) );
  XOR2_X1 U9245 ( .A(n8023), .B(n8735), .Z(n7938) );
  OAI22_X1 U9246 ( .A1(n7938), .A2(n9689), .B1(n8078), .B2(n9687), .ZN(n7970)
         );
  INV_X1 U9247 ( .A(n7970), .ZN(n7957) );
  NAND2_X1 U9248 ( .A1(n7940), .A2(n7939), .ZN(n8496) );
  INV_X1 U9249 ( .A(n8496), .ZN(n7941) );
  INV_X1 U9250 ( .A(n8033), .ZN(n7943) );
  AOI21_X1 U9251 ( .B1(n8735), .B2(n7944), .A(n7943), .ZN(n7972) );
  NAND2_X1 U9252 ( .A1(n7155), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7951) );
  INV_X1 U9253 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7945) );
  OR2_X1 U9254 ( .A1(n7548), .A2(n7945), .ZN(n7950) );
  NAND2_X1 U9255 ( .A1(n7946), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7947) );
  AND2_X1 U9256 ( .A1(n8015), .A2(n7947), .ZN(n8184) );
  OR2_X1 U9257 ( .A1(n8037), .A2(n8184), .ZN(n7949) );
  OR2_X1 U9258 ( .A1(n8711), .A2(n8193), .ZN(n7948) );
  INV_X1 U9259 ( .A(n8260), .ZN(n9386) );
  OAI22_X1 U9260 ( .A1(n9692), .A2(n7952), .B1(n7963), .B2(n11105), .ZN(n7953)
         );
  AOI21_X1 U9261 ( .B1(n9695), .B2(n9386), .A(n7953), .ZN(n7954) );
  OAI21_X1 U9262 ( .B1(n8024), .B2(n9662), .A(n7954), .ZN(n7955) );
  AOI21_X1 U9263 ( .B1(n7972), .B2(n11120), .A(n7955), .ZN(n7956) );
  OAI21_X1 U9264 ( .B1(n7957), .B2(n11124), .A(n7956), .ZN(P2_U3224) );
  OAI21_X1 U9265 ( .B1(n7960), .B2(n7959), .A(n7958), .ZN(n7962) );
  XNOR2_X1 U9266 ( .A(n8024), .B(n7528), .ZN(n8177) );
  XNOR2_X1 U9267 ( .A(n8177), .B(n9387), .ZN(n7961) );
  NAND2_X1 U9268 ( .A1(n7962), .A2(n7961), .ZN(n8179) );
  OAI211_X1 U9269 ( .C1(n7962), .C2(n7961), .A(n8179), .B(n9370), .ZN(n7969)
         );
  INV_X1 U9270 ( .A(n7963), .ZN(n7967) );
  AOI21_X1 U9271 ( .B1(n9373), .B2(n9388), .A(n7964), .ZN(n7965) );
  OAI21_X1 U9272 ( .B1(n8260), .B2(n9375), .A(n7965), .ZN(n7966) );
  AOI21_X1 U9273 ( .B1(n9377), .B2(n7967), .A(n7966), .ZN(n7968) );
  OAI211_X1 U9274 ( .C1(n8024), .C2(n9380), .A(n7969), .B(n7968), .ZN(P2_U3171) );
  OAI22_X1 U9275 ( .A1(n8024), .A2(n9775), .B1(n8260), .B2(n9773), .ZN(n7971)
         );
  AOI211_X1 U9276 ( .C1(n7972), .C2(n9779), .A(n7971), .B(n7970), .ZN(n11149)
         );
  NAND2_X1 U9277 ( .A1(n5132), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7973) );
  OAI21_X1 U9278 ( .B1(n11149), .B2(n5132), .A(n7973), .ZN(P2_U3468) );
  NOR2_X1 U9279 ( .A1(n7989), .A2(n7974), .ZN(n7975) );
  MUX2_X1 U9280 ( .A(n8193), .B(P2_REG2_REG_10__SCAN_IN), .S(n8028), .Z(n7977)
         );
  INV_X1 U9281 ( .A(n7977), .ZN(n7978) );
  AOI21_X1 U9282 ( .B1(n5230), .B2(n7978), .A(n8195), .ZN(n7996) );
  INV_X1 U9283 ( .A(n7979), .ZN(n7981) );
  MUX2_X1 U9284 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8795), .Z(n7982) );
  AND2_X1 U9285 ( .A1(n7982), .A2(n8211), .ZN(n8200) );
  OR2_X1 U9286 ( .A1(n7982), .A2(n8211), .ZN(n8201) );
  INV_X1 U9287 ( .A(n8201), .ZN(n7983) );
  NOR2_X1 U9288 ( .A1(n8200), .A2(n7983), .ZN(n7985) );
  OAI21_X1 U9289 ( .B1(n8202), .B2(n7985), .A(n11086), .ZN(n7984) );
  AOI21_X1 U9290 ( .B1(n8202), .B2(n7985), .A(n7984), .ZN(n7987) );
  INV_X1 U9291 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8180) );
  OAI22_X1 U9292 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8180), .B1(n11096), .B2(
        n8211), .ZN(n7986) );
  AOI211_X1 U9293 ( .C1(n11076), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7987), .B(
        n7986), .ZN(n7995) );
  NOR2_X1 U9294 ( .A1(n7989), .A2(n7988), .ZN(n7991) );
  AOI22_X1 U9295 ( .A1(n8028), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n7945), .B2(
        n8211), .ZN(n7992) );
  AOI21_X1 U9296 ( .B1(n5234), .B2(n7992), .A(n8213), .ZN(n7993) );
  OR2_X1 U9297 ( .A1(n7993), .A2(n11090), .ZN(n7994) );
  OAI211_X1 U9298 ( .C1(n7996), .C2(n11081), .A(n7995), .B(n7994), .ZN(
        P2_U3192) );
  INV_X1 U9299 ( .A(n7997), .ZN(n7998) );
  AOI21_X1 U9300 ( .B1(n10352), .B2(n9928), .A(n7998), .ZN(n8001) );
  NAND2_X1 U9301 ( .A1(n9917), .A2(n7999), .ZN(n8000) );
  OAI211_X1 U9302 ( .C1(n8002), .C2(n9878), .A(n8001), .B(n8000), .ZN(n8008)
         );
  AOI21_X1 U9303 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8006) );
  NOR2_X1 U9304 ( .A1(n8006), .A2(n9919), .ZN(n8007) );
  AOI211_X1 U9305 ( .C1(n8009), .C2(n9904), .A(n8008), .B(n8007), .ZN(n8010)
         );
  INV_X1 U9306 ( .A(n8010), .ZN(P1_U3221) );
  NAND2_X1 U9307 ( .A1(n8011), .A2(n5140), .ZN(n8013) );
  AOI22_X1 U9308 ( .A1(n7313), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7534), .B2(
        n8214), .ZN(n8012) );
  NAND2_X1 U9309 ( .A1(n7155), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8021) );
  INV_X1 U9310 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8014) );
  OR2_X1 U9311 ( .A1(n7548), .A2(n8014), .ZN(n8020) );
  NAND2_X1 U9312 ( .A1(n8015), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8016) );
  AND2_X1 U9313 ( .A1(n8035), .A2(n8016), .ZN(n8263) );
  OR2_X1 U9314 ( .A1(n8037), .A2(n8263), .ZN(n8019) );
  INV_X1 U9315 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8017) );
  OR2_X1 U9316 ( .A1(n8711), .A2(n8017), .ZN(n8018) );
  NOR2_X1 U9317 ( .A1(n8265), .A2(n8293), .ZN(n8502) );
  INV_X1 U9318 ( .A(n8502), .ZN(n8022) );
  NAND2_X1 U9319 ( .A1(n8181), .A2(n8024), .ZN(n8025) );
  AOI22_X1 U9320 ( .A1(n7313), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7534), .B2(
        n8028), .ZN(n8029) );
  NOR2_X1 U9321 ( .A1(n8226), .A2(n9386), .ZN(n8101) );
  OR2_X1 U9322 ( .A1(n8110), .A2(n8101), .ZN(n8030) );
  NAND2_X1 U9323 ( .A1(n8226), .A2(n9386), .ZN(n8102) );
  NAND2_X1 U9324 ( .A1(n8030), .A2(n8102), .ZN(n8031) );
  XOR2_X1 U9325 ( .A(n8739), .B(n8031), .Z(n8032) );
  OAI22_X1 U9326 ( .A1(n8032), .A2(n9689), .B1(n8260), .B2(n9687), .ZN(n8132)
         );
  INV_X1 U9327 ( .A(n8132), .ZN(n8047) );
  OR2_X1 U9328 ( .A1(n8226), .A2(n8260), .ZN(n8488) );
  NAND2_X1 U9329 ( .A1(n8488), .A2(n8089), .ZN(n8495) );
  NAND2_X1 U9330 ( .A1(n8226), .A2(n8260), .ZN(n8498) );
  XNOR2_X1 U9331 ( .A(n8122), .B(n8739), .ZN(n8134) );
  INV_X1 U9332 ( .A(n8265), .ZN(n8131) );
  NAND2_X1 U9333 ( .A1(n7155), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8042) );
  INV_X1 U9334 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8124) );
  OR2_X1 U9335 ( .A1(n8711), .A2(n8124), .ZN(n8041) );
  AND2_X1 U9336 ( .A1(n8035), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8036) );
  NOR2_X1 U9337 ( .A1(n8113), .A2(n8036), .ZN(n8100) );
  OR2_X1 U9338 ( .A1(n8037), .A2(n8100), .ZN(n8040) );
  INV_X1 U9339 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8038) );
  OR2_X1 U9340 ( .A1(n7548), .A2(n8038), .ZN(n8039) );
  NAND4_X1 U9341 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n9384)
         );
  OAI22_X1 U9342 ( .A1(n9692), .A2(n8017), .B1(n8263), .B2(n11105), .ZN(n8043)
         );
  AOI21_X1 U9343 ( .B1(n9695), .B2(n9384), .A(n8043), .ZN(n8044) );
  OAI21_X1 U9344 ( .B1(n8131), .B2(n9662), .A(n8044), .ZN(n8045) );
  AOI21_X1 U9345 ( .B1(n8134), .B2(n11120), .A(n8045), .ZN(n8046) );
  OAI21_X1 U9346 ( .B1(n8047), .B2(n11124), .A(n8046), .ZN(P2_U3222) );
  NAND2_X1 U9347 ( .A1(n8048), .A2(n8943), .ZN(n8049) );
  NAND2_X1 U9348 ( .A1(n8050), .A2(n8049), .ZN(n8234) );
  OR2_X1 U9349 ( .A1(n8234), .A2(n11166), .ZN(n8058) );
  NAND2_X1 U9350 ( .A1(n8051), .A2(n9079), .ZN(n8052) );
  XNOR2_X1 U9351 ( .A(n8052), .B(n8943), .ZN(n8056) );
  NAND2_X1 U9352 ( .A1(n10346), .A2(n11155), .ZN(n8054) );
  NAND2_X1 U9353 ( .A1(n10348), .A2(n11156), .ZN(n8053) );
  NAND2_X1 U9354 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  AOI21_X1 U9355 ( .B1(n8056), .B2(n10746), .A(n8055), .ZN(n8057) );
  NAND2_X1 U9356 ( .A1(n8058), .A2(n8057), .ZN(n8237) );
  NAND2_X1 U9357 ( .A1(n8237), .A2(n10601), .ZN(n8064) );
  OAI21_X1 U9358 ( .B1(n8059), .B2(n8290), .A(n10672), .ZN(n8060) );
  NOR2_X1 U9359 ( .A1(n8060), .A2(n8815), .ZN(n8235) );
  AOI22_X1 U9360 ( .A1(n7511), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8287), .B2(
        n10632), .ZN(n8061) );
  OAI21_X1 U9361 ( .B1(n8290), .B2(n10658), .A(n8061), .ZN(n8062) );
  AOI21_X1 U9362 ( .B1(n8235), .B2(n10664), .A(n8062), .ZN(n8063) );
  OAI211_X1 U9363 ( .C1(n8234), .C2(n8065), .A(n8064), .B(n8063), .ZN(P1_U3279) );
  OAI21_X1 U9364 ( .B1(n8068), .B2(n8067), .A(n8066), .ZN(n8069) );
  NAND2_X1 U9365 ( .A1(n8069), .A2(n9926), .ZN(n8075) );
  NAND2_X1 U9366 ( .A1(n9932), .A2(n10348), .ZN(n8070) );
  OAI211_X1 U9367 ( .C1(n10349), .C2(n9912), .A(n8071), .B(n8070), .ZN(n8072)
         );
  AOI21_X1 U9368 ( .B1(n8073), .B2(n9917), .A(n8072), .ZN(n8074) );
  OAI211_X1 U9369 ( .C1(n11175), .C2(n9936), .A(n8075), .B(n8074), .ZN(
        P1_U3224) );
  NOR2_X1 U9370 ( .A1(n8076), .A2(n9752), .ZN(n8082) );
  OAI22_X1 U9371 ( .A1(n8078), .A2(n9773), .B1(n8077), .B2(n9775), .ZN(n8080)
         );
  AOI211_X1 U9372 ( .C1(n8082), .C2(n8081), .A(n8080), .B(n8079), .ZN(n11147)
         );
  NAND2_X1 U9373 ( .A1(n5132), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8083) );
  OAI21_X1 U9374 ( .B1(n11147), .B2(n5132), .A(n8083), .ZN(P2_U3466) );
  INV_X1 U9375 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8085) );
  INV_X1 U9376 ( .A(n8612), .ZN(n8087) );
  OAI222_X1 U9377 ( .A1(n8844), .A2(n8085), .B1(n9800), .B2(n8087), .C1(
        P2_U3151), .C2(n8084), .ZN(P2_U3273) );
  OAI222_X1 U9378 ( .A1(n8088), .A2(P1_U3086), .B1(n9222), .B2(n8087), .C1(
        n8086), .C2(n9220), .ZN(P1_U3333) );
  NAND2_X1 U9379 ( .A1(n8033), .A2(n8089), .ZN(n8090) );
  XNOR2_X1 U9380 ( .A(n8226), .B(n8260), .ZN(n8736) );
  XNOR2_X1 U9381 ( .A(n8090), .B(n8736), .ZN(n8230) );
  XOR2_X1 U9382 ( .A(n8110), .B(n8736), .Z(n8093) );
  INV_X1 U9383 ( .A(n8293), .ZN(n9385) );
  AOI22_X1 U9384 ( .A1(n9385), .A2(n7160), .B1(n7162), .B2(n9387), .ZN(n8092)
         );
  NAND2_X1 U9385 ( .A1(n8230), .A2(n9203), .ZN(n8091) );
  OAI211_X1 U9386 ( .C1(n8093), .C2(n9689), .A(n8092), .B(n8091), .ZN(n8228)
         );
  AOI21_X1 U9387 ( .B1(n11110), .B2(n8230), .A(n8228), .ZN(n8096) );
  OAI22_X1 U9388 ( .A1(n9692), .A2(n8193), .B1(n8184), .B2(n11105), .ZN(n8094)
         );
  AOI21_X1 U9389 ( .B1(n11116), .B2(n8226), .A(n8094), .ZN(n8095) );
  OAI21_X1 U9390 ( .B1(n8096), .B2(n11124), .A(n8095), .ZN(P2_U3223) );
  INV_X1 U9391 ( .A(n8626), .ZN(n8099) );
  NAND2_X1 U9392 ( .A1(n8097), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8799) );
  NAND2_X1 U9393 ( .A1(n9802), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8098) );
  OAI211_X1 U9394 ( .C1(n8099), .C2(n9804), .A(n8799), .B(n8098), .ZN(P2_U3272) );
  INV_X1 U9395 ( .A(n8100), .ZN(n8302) );
  NOR2_X1 U9396 ( .A1(n8265), .A2(n9385), .ZN(n8104) );
  OR2_X1 U9397 ( .A1(n8101), .A2(n8104), .ZN(n8111) );
  OR2_X1 U9398 ( .A1(n8110), .A2(n8111), .ZN(n8105) );
  AND2_X1 U9399 ( .A1(n5212), .A2(n8102), .ZN(n8103) );
  AND2_X1 U9400 ( .A1(n8105), .A2(n8112), .ZN(n8109) );
  INV_X1 U9401 ( .A(n8318), .ZN(n8208) );
  AOI22_X1 U9402 ( .A1(n7313), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7534), .B2(
        n8208), .ZN(n8107) );
  NAND2_X1 U9403 ( .A1(n8108), .A2(n8107), .ZN(n8505) );
  AOI21_X1 U9404 ( .B1(n8109), .B2(n8737), .A(n9689), .ZN(n8120) );
  NAND2_X1 U9405 ( .A1(n7155), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U9406 ( .A1(n7539), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8117) );
  NOR2_X1 U9407 ( .A1(n8113), .A2(n8321), .ZN(n8114) );
  OR2_X1 U9408 ( .A1(n8168), .A2(n8114), .ZN(n9322) );
  NAND2_X1 U9409 ( .A1(n7757), .A2(n9322), .ZN(n8116) );
  NAND2_X1 U9410 ( .A1(n7156), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8115) );
  NAND4_X1 U9411 ( .A1(n8118), .A2(n8117), .A3(n8116), .A4(n8115), .ZN(n9383)
         );
  OAI22_X1 U9412 ( .A1(n9688), .A2(n9773), .B1(n8293), .B2(n9687), .ZN(n8119)
         );
  AOI21_X1 U9413 ( .B1(n8120), .B2(n8164), .A(n8119), .ZN(n8136) );
  INV_X1 U9414 ( .A(n8136), .ZN(n8121) );
  AOI21_X1 U9415 ( .B1(n11118), .B2(n8302), .A(n8121), .ZN(n8127) );
  XNOR2_X1 U9416 ( .A(n8160), .B(n8737), .ZN(n8138) );
  INV_X1 U9417 ( .A(n8505), .ZN(n8305) );
  OAI22_X1 U9418 ( .A1(n8305), .A2(n9662), .B1(n8124), .B2(n9692), .ZN(n8125)
         );
  AOI21_X1 U9419 ( .B1(n8138), .B2(n11120), .A(n8125), .ZN(n8126) );
  OAI21_X1 U9420 ( .B1(n8127), .B2(n11124), .A(n8126), .ZN(P2_U3221) );
  NAND2_X1 U9421 ( .A1(n8626), .A2(n10820), .ZN(n8129) );
  OR2_X1 U9422 ( .A1(n8128), .A2(P1_U3086), .ZN(n9126) );
  OAI211_X1 U9423 ( .C1(n8130), .C2(n9220), .A(n8129), .B(n9126), .ZN(P1_U3332) );
  OAI22_X1 U9424 ( .A1(n8131), .A2(n9775), .B1(n9134), .B2(n9773), .ZN(n8133)
         );
  AOI211_X1 U9425 ( .C1(n8134), .C2(n9779), .A(n8133), .B(n8132), .ZN(n11153)
         );
  NAND2_X1 U9426 ( .A1(n5132), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8135) );
  OAI21_X1 U9427 ( .B1(n11153), .B2(n5132), .A(n8135), .ZN(P2_U3470) );
  OAI21_X1 U9428 ( .B1(n8305), .B2(n9775), .A(n8136), .ZN(n8137) );
  AOI21_X1 U9429 ( .B1(n9779), .B2(n8138), .A(n8137), .ZN(n11172) );
  OR2_X1 U9430 ( .A1(n8232), .A2(n8038), .ZN(n8139) );
  OAI21_X1 U9431 ( .B1(n11172), .B2(n5132), .A(n8139), .ZN(P2_U3471) );
  OAI21_X1 U9432 ( .B1(n8141), .B2(n8144), .A(n8140), .ZN(n10762) );
  AOI211_X1 U9433 ( .C1(n10759), .C2(n8816), .A(n10655), .B(n8251), .ZN(n10757) );
  NAND2_X1 U9434 ( .A1(n10759), .A2(n10580), .ZN(n8143) );
  AOI22_X1 U9435 ( .A1(n7511), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9849), .B2(
        n10632), .ZN(n8142) );
  OAI211_X1 U9436 ( .C1(n10756), .C2(n10488), .A(n8143), .B(n8142), .ZN(n8148)
         );
  XNOR2_X1 U9437 ( .A(n8145), .B(n8144), .ZN(n8146) );
  INV_X1 U9438 ( .A(n10740), .ZN(n10345) );
  AOI22_X1 U9439 ( .A1(n8146), .A2(n10746), .B1(n11155), .B2(n10345), .ZN(
        n10761) );
  NOR2_X1 U9440 ( .A1(n10761), .A2(n7511), .ZN(n8147) );
  AOI211_X1 U9441 ( .C1(n10757), .C2(n10664), .A(n8148), .B(n8147), .ZN(n8149)
         );
  OAI21_X1 U9442 ( .B1(n10762), .B2(n10638), .A(n8149), .ZN(P1_U3277) );
  OAI211_X1 U9443 ( .C1(n8152), .C2(n8151), .A(n8150), .B(n9926), .ZN(n8158)
         );
  NAND2_X1 U9444 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10949) );
  INV_X1 U9445 ( .A(n10949), .ZN(n8153) );
  AOI21_X1 U9446 ( .B1(n9928), .B2(n11154), .A(n8153), .ZN(n8154) );
  OAI21_X1 U9447 ( .B1(n10764), .B2(n9878), .A(n8154), .ZN(n8155) );
  AOI21_X1 U9448 ( .B1(n8156), .B2(n9917), .A(n8155), .ZN(n8157) );
  OAI211_X1 U9449 ( .C1(n8159), .C2(n9936), .A(n8158), .B(n8157), .ZN(P1_U3234) );
  NAND2_X1 U9450 ( .A1(n8505), .A2(n9134), .ZN(n8491) );
  OR2_X1 U9451 ( .A1(n8161), .A2(n7524), .ZN(n8163) );
  AOI22_X1 U9452 ( .A1(n7313), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7534), .B2(
        n8390), .ZN(n8162) );
  XNOR2_X1 U9453 ( .A(n9328), .B(n9688), .ZN(n8525) );
  INV_X1 U9454 ( .A(n8525), .ZN(n8752) );
  XNOR2_X1 U9455 ( .A(n8753), .B(n8752), .ZN(n8190) );
  INV_X1 U9456 ( .A(n8190), .ZN(n8176) );
  XNOR2_X1 U9457 ( .A(n9191), .B(n8525), .ZN(n8165) );
  OAI22_X1 U9458 ( .A1(n8165), .A2(n9689), .B1(n9134), .B2(n9687), .ZN(n8188)
         );
  INV_X1 U9459 ( .A(n9322), .ZN(n8166) );
  OAI22_X1 U9460 ( .A1(n9190), .A2(n11103), .B1(n8166), .B2(n11105), .ZN(n8167) );
  OAI21_X1 U9461 ( .B1(n8188), .B2(n8167), .A(n9692), .ZN(n8175) );
  NAND2_X1 U9462 ( .A1(n7156), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U9463 ( .A1(n7155), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U9464 ( .A1(n7539), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8171) );
  OR2_X1 U9465 ( .A1(n8168), .A2(n9237), .ZN(n8169) );
  AND2_X1 U9466 ( .A1(n8169), .A2(n8511), .ZN(n9691) );
  OR2_X1 U9467 ( .A1(n8037), .A2(n9691), .ZN(n8170) );
  NAND4_X1 U9468 ( .A1(n8173), .A2(n8172), .A3(n8171), .A4(n8170), .ZN(n9382)
         );
  AOI22_X1 U9469 ( .A1(n9695), .A2(n9382), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n11124), .ZN(n8174) );
  OAI211_X1 U9470 ( .C1(n8176), .C2(n9698), .A(n8175), .B(n8174), .ZN(P2_U3220) );
  OR2_X1 U9471 ( .A1(n8177), .A2(n8181), .ZN(n8178) );
  NAND2_X1 U9472 ( .A1(n8179), .A2(n8178), .ZN(n8258) );
  XNOR2_X1 U9473 ( .A(n8226), .B(n7528), .ZN(n8257) );
  XNOR2_X1 U9474 ( .A(n8259), .B(n8260), .ZN(n8187) );
  OAI22_X1 U9475 ( .A1(n9361), .A2(n8181), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8180), .ZN(n8182) );
  AOI21_X1 U9476 ( .B1(n9359), .B2(n9385), .A(n8182), .ZN(n8183) );
  OAI21_X1 U9477 ( .B1(n8184), .B2(n9348), .A(n8183), .ZN(n8185) );
  AOI21_X1 U9478 ( .B1(n8226), .B2(n9327), .A(n8185), .ZN(n8186) );
  OAI21_X1 U9479 ( .B1(n8187), .B2(n9330), .A(n8186), .ZN(P2_U3157) );
  OAI22_X1 U9480 ( .A1(n9190), .A2(n9775), .B1(n9669), .B2(n9773), .ZN(n8189)
         );
  AOI211_X1 U9481 ( .C1(n9779), .C2(n8190), .A(n8189), .B(n8188), .ZN(n11187)
         );
  NAND2_X1 U9482 ( .A1(n5132), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8191) );
  OAI21_X1 U9483 ( .B1(n11187), .B2(n5132), .A(n8191), .ZN(P2_U3472) );
  INV_X1 U9484 ( .A(n8639), .ZN(n8244) );
  AOI22_X1 U9485 ( .A1(n6763), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9802), .ZN(n8192) );
  OAI21_X1 U9486 ( .B1(n8244), .B2(n9800), .A(n8192), .ZN(P2_U3271) );
  NOR2_X1 U9487 ( .A1(n8214), .A2(n8196), .ZN(n8197) );
  NAND2_X1 U9488 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8318), .ZN(n8198) );
  OAI21_X1 U9489 ( .B1(n8318), .B2(P2_REG2_REG_12__SCAN_IN), .A(n8198), .ZN(
        n8199) );
  AOI21_X1 U9490 ( .B1(n5229), .B2(n8199), .A(n8317), .ZN(n8225) );
  MUX2_X1 U9491 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8795), .Z(n8312) );
  XNOR2_X1 U9492 ( .A(n8312), .B(n8208), .ZN(n8206) );
  MUX2_X1 U9493 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8795), .Z(n8203) );
  OR2_X1 U9494 ( .A1(n8203), .A2(n11095), .ZN(n8204) );
  XNOR2_X1 U9495 ( .A(n8203), .B(n8214), .ZN(n11085) );
  NAND2_X1 U9496 ( .A1(n11084), .A2(n11085), .ZN(n11083) );
  NAND2_X1 U9497 ( .A1(n8204), .A2(n11083), .ZN(n8205) );
  NAND2_X1 U9498 ( .A1(n8206), .A2(n8205), .ZN(n8313) );
  OAI21_X1 U9499 ( .B1(n8206), .B2(n8205), .A(n8313), .ZN(n8223) );
  INV_X1 U9500 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8210) );
  INV_X1 U9501 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8207) );
  NOR2_X1 U9502 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8207), .ZN(n8299) );
  AOI21_X1 U9503 ( .B1(n11033), .B2(n8208), .A(n8299), .ZN(n8209) );
  OAI21_X1 U9504 ( .B1(n11040), .B2(n8210), .A(n8209), .ZN(n8222) );
  NOR2_X1 U9505 ( .A1(n8214), .A2(n8215), .ZN(n8216) );
  XNOR2_X1 U9506 ( .A(n8215), .B(n8214), .ZN(n11078) );
  NAND2_X1 U9507 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8318), .ZN(n8217) );
  OAI21_X1 U9508 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8318), .A(n8217), .ZN(
        n8218) );
  AOI21_X1 U9509 ( .B1(n8219), .B2(n8218), .A(n8309), .ZN(n8220) );
  NOR2_X1 U9510 ( .A1(n8220), .A2(n11090), .ZN(n8221) );
  AOI211_X1 U9511 ( .C1(n11086), .C2(n8223), .A(n8222), .B(n8221), .ZN(n8224)
         );
  OAI21_X1 U9512 ( .B1(n8225), .B2(n11081), .A(n8224), .ZN(P2_U3194) );
  INV_X1 U9513 ( .A(n8226), .ZN(n8227) );
  NOR2_X1 U9514 ( .A1(n8227), .A2(n9775), .ZN(n8229) );
  AOI211_X1 U9515 ( .C1(n8230), .C2(n9704), .A(n8229), .B(n8228), .ZN(n11151)
         );
  OR2_X1 U9516 ( .A1(n11151), .A2(n5132), .ZN(n8231) );
  OAI21_X1 U9517 ( .B1(n8232), .B2(n7945), .A(n8231), .ZN(P2_U3469) );
  NOR2_X1 U9518 ( .A1(n8234), .A2(n8233), .ZN(n8236) );
  OR3_X1 U9519 ( .A1(n8237), .A2(n8236), .A3(n8235), .ZN(n8240) );
  MUX2_X1 U9520 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n8240), .S(n11185), .Z(n8238) );
  INV_X1 U9521 ( .A(n8238), .ZN(n8239) );
  OAI21_X1 U9522 ( .B1(n8290), .B2(n10806), .A(n8239), .ZN(P1_U3495) );
  MUX2_X1 U9523 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n8240), .S(n11181), .Z(n8241) );
  INV_X1 U9524 ( .A(n8241), .ZN(n8242) );
  OAI21_X1 U9525 ( .B1(n8290), .B2(n10739), .A(n8242), .ZN(P1_U3536) );
  OAI222_X1 U9526 ( .A1(P1_U3086), .A2(n8245), .B1(n9222), .B2(n8244), .C1(
        n8243), .C2(n9220), .ZN(P1_U3331) );
  OAI21_X1 U9527 ( .B1(n8247), .B2(n8248), .A(n8246), .ZN(n10755) );
  INV_X1 U9528 ( .A(n8248), .ZN(n8952) );
  XNOR2_X1 U9529 ( .A(n8249), .B(n8952), .ZN(n8250) );
  OAI222_X1 U9530 ( .A1(n10763), .A2(n9857), .B1(n10741), .B2(n10644), .C1(
        n10713), .C2(n8250), .ZN(n10751) );
  INV_X1 U9531 ( .A(n8271), .ZN(n8252) );
  AOI211_X1 U9532 ( .C1(n10753), .C2(n5428), .A(n10655), .B(n8252), .ZN(n10752) );
  NAND2_X1 U9533 ( .A1(n10752), .A2(n10664), .ZN(n8254) );
  AOI22_X1 U9534 ( .A1(n7511), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9859), .B2(
        n10632), .ZN(n8253) );
  OAI211_X1 U9535 ( .C1(n9862), .C2(n10658), .A(n8254), .B(n8253), .ZN(n8255)
         );
  AOI21_X1 U9536 ( .B1(n10751), .B2(n10661), .A(n8255), .ZN(n8256) );
  OAI21_X1 U9537 ( .B1(n10755), .B2(n10638), .A(n8256), .ZN(P1_U3276) );
  XNOR2_X1 U9538 ( .A(n8265), .B(n7528), .ZN(n8292) );
  XNOR2_X1 U9539 ( .A(n8292), .B(n8293), .ZN(n8295) );
  XOR2_X1 U9540 ( .A(n8296), .B(n8295), .Z(n8267) );
  INV_X1 U9541 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10223) );
  OAI22_X1 U9542 ( .A1(n9361), .A2(n8260), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10223), .ZN(n8261) );
  AOI21_X1 U9543 ( .B1(n9359), .B2(n9384), .A(n8261), .ZN(n8262) );
  OAI21_X1 U9544 ( .B1(n8263), .B2(n9348), .A(n8262), .ZN(n8264) );
  AOI21_X1 U9545 ( .B1(n8265), .B2(n9327), .A(n8264), .ZN(n8266) );
  OAI21_X1 U9546 ( .B1(n8267), .B2(n9330), .A(n8266), .ZN(P2_U3176) );
  OAI222_X1 U9547 ( .A1(P1_U3086), .A2(n8269), .B1(n9222), .B2(n8830), .C1(
        n8268), .C2(n9220), .ZN(P1_U3330) );
  XNOR2_X1 U9548 ( .A(n9913), .B(n10344), .ZN(n8878) );
  XNOR2_X1 U9549 ( .A(n8270), .B(n8878), .ZN(n10750) );
  AOI211_X1 U9550 ( .C1(n10745), .C2(n8271), .A(n10655), .B(n10652), .ZN(
        n10743) );
  NOR2_X1 U9551 ( .A1(n9913), .A2(n10658), .ZN(n8276) );
  NAND2_X1 U9552 ( .A1(n10343), .A2(n8272), .ZN(n8274) );
  AOI22_X1 U9553 ( .A1(n7511), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9916), .B2(
        n10632), .ZN(n8273) );
  OAI211_X1 U9554 ( .C1(n10740), .C2(n10488), .A(n8274), .B(n8273), .ZN(n8275)
         );
  AOI211_X1 U9555 ( .C1(n10743), .C2(n10664), .A(n8276), .B(n8275), .ZN(n8279)
         );
  XNOR2_X1 U9556 ( .A(n8277), .B(n8878), .ZN(n10747) );
  NAND2_X1 U9557 ( .A1(n10747), .A2(n10529), .ZN(n8278) );
  OAI211_X1 U9558 ( .C1(n10750), .C2(n10638), .A(n8279), .B(n8278), .ZN(
        P1_U3275) );
  OAI21_X1 U9559 ( .B1(n8280), .B2(n8282), .A(n8281), .ZN(n8283) );
  NAND2_X1 U9560 ( .A1(n8283), .A2(n9926), .ZN(n8289) );
  AOI22_X1 U9561 ( .A1(n9932), .A2(n10346), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8284) );
  OAI21_X1 U9562 ( .B1(n8285), .B2(n9912), .A(n8284), .ZN(n8286) );
  AOI21_X1 U9563 ( .B1(n8287), .B2(n9917), .A(n8286), .ZN(n8288) );
  OAI211_X1 U9564 ( .C1(n8290), .C2(n9936), .A(n8289), .B(n8288), .ZN(P1_U3215) );
  INV_X1 U9565 ( .A(n8662), .ZN(n8307) );
  AOI22_X1 U9566 ( .A1(n7173), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9802), .ZN(n8291) );
  OAI21_X1 U9567 ( .B1(n8307), .B2(n9800), .A(n8291), .ZN(P2_U3269) );
  INV_X1 U9568 ( .A(n8292), .ZN(n8294) );
  XNOR2_X1 U9569 ( .A(n8505), .B(n7528), .ZN(n9131) );
  XNOR2_X1 U9570 ( .A(n9131), .B(n9134), .ZN(n8297) );
  OAI211_X1 U9571 ( .C1(n8298), .C2(n8297), .A(n9132), .B(n9370), .ZN(n8304)
         );
  AOI21_X1 U9572 ( .B1(n9373), .B2(n9385), .A(n8299), .ZN(n8300) );
  OAI21_X1 U9573 ( .B1(n9688), .B2(n9375), .A(n8300), .ZN(n8301) );
  AOI21_X1 U9574 ( .B1(n9377), .B2(n8302), .A(n8301), .ZN(n8303) );
  OAI211_X1 U9575 ( .C1(n8305), .C2(n9380), .A(n8304), .B(n8303), .ZN(P2_U3164) );
  OAI222_X1 U9576 ( .A1(n8308), .A2(P1_U3086), .B1(n9222), .B2(n8307), .C1(
        n8306), .C2(n9220), .ZN(P1_U3329) );
  INV_X1 U9577 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8311) );
  XNOR2_X1 U9578 ( .A(n8351), .B(n8390), .ZN(n8310) );
  AOI21_X1 U9579 ( .B1(n8311), .B2(n8310), .A(n8353), .ZN(n8328) );
  MUX2_X1 U9580 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8795), .Z(n8388) );
  XNOR2_X1 U9581 ( .A(n8388), .B(n8390), .ZN(n8316) );
  OR2_X1 U9582 ( .A1(n8312), .A2(n8318), .ZN(n8314) );
  NAND2_X1 U9583 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U9584 ( .A1(n8316), .A2(n8315), .ZN(n8391) );
  OAI21_X1 U9585 ( .B1(n8316), .B2(n8315), .A(n8391), .ZN(n8326) );
  XNOR2_X1 U9586 ( .A(n8364), .B(n8390), .ZN(n8320) );
  INV_X1 U9587 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8319) );
  AOI21_X1 U9588 ( .B1(n8320), .B2(n8319), .A(n8365), .ZN(n8324) );
  NAND2_X1 U9589 ( .A1(n11076), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8323) );
  NOR2_X1 U9590 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8321), .ZN(n9323) );
  AOI21_X1 U9591 ( .B1(n11033), .B2(n8390), .A(n9323), .ZN(n8322) );
  OAI211_X1 U9592 ( .C1(n8324), .C2(n11081), .A(n8323), .B(n8322), .ZN(n8325)
         );
  AOI21_X1 U9593 ( .B1(n11086), .B2(n8326), .A(n8325), .ZN(n8327) );
  OAI21_X1 U9594 ( .B1(n8328), .B2(n11090), .A(n8327), .ZN(P2_U3195) );
  NAND2_X1 U9595 ( .A1(n8674), .A2(n8329), .ZN(n8331) );
  OAI211_X1 U9596 ( .C1(n8332), .C2(n8844), .A(n8331), .B(n8330), .ZN(P2_U3268) );
  INV_X1 U9597 ( .A(n8435), .ZN(n8346) );
  AOI21_X1 U9598 ( .B1(n9802), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8333), .ZN(
        n8334) );
  OAI21_X1 U9599 ( .B1(n8346), .B2(n9800), .A(n8334), .ZN(P2_U3267) );
  NAND2_X1 U9600 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  XOR2_X1 U9601 ( .A(n8338), .B(n8337), .Z(n8344) );
  NOR2_X1 U9602 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8339), .ZN(n10922) );
  AOI21_X1 U9603 ( .B1(n8823), .B2(n9932), .A(n10922), .ZN(n8341) );
  NAND2_X1 U9604 ( .A1(n9917), .A2(n8819), .ZN(n8340) );
  OAI211_X1 U9605 ( .C1(n10764), .C2(n9912), .A(n8341), .B(n8340), .ZN(n8342)
         );
  AOI21_X1 U9606 ( .B1(n10767), .B2(n9904), .A(n8342), .ZN(n8343) );
  OAI21_X1 U9607 ( .B1(n8344), .B2(n9919), .A(n8343), .ZN(P1_U3241) );
  OAI222_X1 U9608 ( .A1(P1_U3086), .A2(n5139), .B1(n9222), .B2(n8346), .C1(
        n8345), .C2(n9220), .ZN(P1_U3327) );
  INV_X1 U9609 ( .A(n8674), .ZN(n8348) );
  OAI222_X1 U9610 ( .A1(P1_U3086), .A2(n8349), .B1(n9222), .B2(n8348), .C1(
        n8347), .C2(n9220), .ZN(P1_U3328) );
  OAI222_X1 U9611 ( .A1(P1_U3086), .A2(n5872), .B1(n9222), .B2(n8841), .C1(
        n8350), .C2(n9220), .ZN(P1_U3326) );
  NOR2_X1 U9612 ( .A1(n8390), .A2(n8351), .ZN(n8352) );
  INV_X1 U9613 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8354) );
  MUX2_X1 U9614 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8354), .S(n9401), .Z(n9404)
         );
  NOR2_X1 U9615 ( .A1(n9420), .A2(n8355), .ZN(n8358) );
  INV_X1 U9616 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9425) );
  INV_X1 U9617 ( .A(n9420), .ZN(n8356) );
  INV_X1 U9618 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8359) );
  AOI22_X1 U9619 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9439), .B1(n8382), .B2(
        n8359), .ZN(n9443) );
  NOR2_X1 U9620 ( .A1(n9457), .A2(n8360), .ZN(n8361) );
  INV_X1 U9621 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9453) );
  NOR2_X1 U9622 ( .A1(n9453), .A2(n9452), .ZN(n9451) );
  NAND2_X1 U9623 ( .A1(n9486), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8362) );
  OAI21_X1 U9624 ( .B1(n9486), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8362), .ZN(
        n9471) );
  INV_X1 U9625 ( .A(n8362), .ZN(n8363) );
  XNOR2_X1 U9626 ( .A(n7153), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8401) );
  INV_X1 U9627 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9414) );
  INV_X1 U9628 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8366) );
  MUX2_X1 U9629 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n8366), .S(n9401), .Z(n9396)
         );
  NAND2_X1 U9630 ( .A1(n8386), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8367) );
  NOR2_X1 U9631 ( .A1(n9420), .A2(n8368), .ZN(n8369) );
  MUX2_X1 U9632 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n8370), .S(n9439), .Z(n9433)
         );
  NAND2_X1 U9633 ( .A1(n9457), .A2(n8372), .ZN(n8373) );
  INV_X1 U9634 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9455) );
  XNOR2_X1 U9635 ( .A(n8556), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n9474) );
  INV_X1 U9636 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U9637 ( .A1(n8375), .A2(n9633), .ZN(n8374) );
  INV_X1 U9638 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8376) );
  MUX2_X1 U9639 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8376), .S(n7153), .Z(n8403)
         );
  NAND2_X1 U9640 ( .A1(n8378), .A2(n8377), .ZN(n8381) );
  NAND2_X1 U9641 ( .A1(n11033), .A2(n7153), .ZN(n8379) );
  NAND2_X1 U9642 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9256) );
  MUX2_X1 U9643 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n7159), .Z(n8397) );
  XNOR2_X1 U9644 ( .A(n8397), .B(n9457), .ZN(n9465) );
  MUX2_X1 U9645 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8795), .Z(n8383) );
  OR2_X1 U9646 ( .A1(n8383), .A2(n8382), .ZN(n8395) );
  XNOR2_X1 U9647 ( .A(n8383), .B(n9439), .ZN(n9437) );
  MUX2_X1 U9648 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8795), .Z(n8385) );
  INV_X1 U9649 ( .A(n8385), .ZN(n8384) );
  NAND2_X1 U9650 ( .A1(n9420), .A2(n8384), .ZN(n8394) );
  XNOR2_X1 U9651 ( .A(n8385), .B(n9420), .ZN(n9418) );
  MUX2_X1 U9652 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8795), .Z(n8387) );
  OR2_X1 U9653 ( .A1(n8387), .A2(n8386), .ZN(n8393) );
  XNOR2_X1 U9654 ( .A(n8387), .B(n9401), .ZN(n9399) );
  INV_X1 U9655 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U9656 ( .A1(n8390), .A2(n8389), .ZN(n8392) );
  NAND2_X1 U9657 ( .A1(n8392), .A2(n8391), .ZN(n9398) );
  NAND2_X1 U9658 ( .A1(n9399), .A2(n9398), .ZN(n9397) );
  NAND2_X1 U9659 ( .A1(n8393), .A2(n9397), .ZN(n9417) );
  NAND2_X1 U9660 ( .A1(n9418), .A2(n9417), .ZN(n9416) );
  NAND2_X1 U9661 ( .A1(n8394), .A2(n9416), .ZN(n9436) );
  NAND2_X1 U9662 ( .A1(n9437), .A2(n9436), .ZN(n9435) );
  NAND2_X1 U9663 ( .A1(n8395), .A2(n9435), .ZN(n9464) );
  NAND2_X1 U9664 ( .A1(n9465), .A2(n9464), .ZN(n9463) );
  OAI21_X1 U9665 ( .B1(n8397), .B2(n8396), .A(n9463), .ZN(n8400) );
  INV_X1 U9666 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8398) );
  MUX2_X1 U9667 ( .A(n9633), .B(n8398), .S(n7159), .Z(n8399) );
  NAND2_X1 U9668 ( .A1(n8400), .A2(n8399), .ZN(n9480) );
  NOR2_X1 U9669 ( .A1(n8400), .A2(n8399), .ZN(n9482) );
  AOI21_X1 U9670 ( .B1(n9486), .B2(n9480), .A(n9482), .ZN(n8405) );
  INV_X1 U9671 ( .A(n8401), .ZN(n8402) );
  MUX2_X1 U9672 ( .A(n8403), .B(n8402), .S(n7159), .Z(n8404) );
  INV_X1 U9673 ( .A(n8406), .ZN(n8408) );
  NAND2_X1 U9674 ( .A1(n8408), .A2(n8407), .ZN(n8409) );
  MUX2_X1 U9675 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8701), .Z(n8698) );
  XNOR2_X1 U9676 ( .A(n8698), .B(SI_30_), .ZN(n8699) );
  XNOR2_X2 U9677 ( .A(n8700), .B(n8699), .ZN(n9219) );
  NAND2_X1 U9678 ( .A1(n9219), .A2(n5140), .ZN(n8412) );
  NAND2_X1 U9679 ( .A1(n7313), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U9680 ( .A1(n8412), .A2(n8411), .ZN(n8716) );
  INV_X1 U9681 ( .A(n8559), .ZN(n8413) );
  NAND2_X1 U9682 ( .A1(n8570), .A2(n10195), .ZN(n8591) );
  INV_X1 U9683 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10002) );
  INV_X1 U9684 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8415) );
  INV_X1 U9685 ( .A(n8644), .ZN(n8417) );
  INV_X1 U9686 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10010) );
  INV_X1 U9687 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U9688 ( .A1(n8643), .A2(n10001), .ZN(n8667) );
  INV_X1 U9689 ( .A(n8667), .ZN(n8418) );
  INV_X1 U9690 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10232) );
  AND2_X2 U9691 ( .A1(n8418), .A2(n10232), .ZN(n8666) );
  INV_X1 U9692 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U9693 ( .A1(n8666), .A2(n8419), .ZN(n8680) );
  OR2_X2 U9694 ( .A1(n8680), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9213) );
  INV_X1 U9695 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8420) );
  OR2_X1 U9696 ( .A1(n7548), .A2(n8420), .ZN(n8425) );
  INV_X1 U9697 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8421) );
  OR2_X1 U9698 ( .A1(n8708), .A2(n8421), .ZN(n8424) );
  INV_X1 U9699 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8422) );
  OR2_X1 U9700 ( .A1(n8711), .A2(n8422), .ZN(n8423) );
  OR2_X1 U9701 ( .A1(n8716), .A2(n8717), .ZN(n8786) );
  OR2_X1 U9702 ( .A1(n8841), .A2(n7524), .ZN(n8427) );
  NAND2_X1 U9703 ( .A1(n7313), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U9704 ( .A1(n8427), .A2(n8426), .ZN(n9703) );
  INV_X1 U9705 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8428) );
  OR2_X1 U9706 ( .A1(n8708), .A2(n8428), .ZN(n8433) );
  INV_X1 U9707 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8429) );
  OR2_X1 U9708 ( .A1(n7548), .A2(n8429), .ZN(n8432) );
  INV_X1 U9709 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8430) );
  OR2_X1 U9710 ( .A1(n8711), .A2(n8430), .ZN(n8431) );
  AND2_X1 U9711 ( .A1(n8779), .A2(n8695), .ZN(n8434) );
  AND2_X1 U9712 ( .A1(n8786), .A2(n8434), .ZN(n8696) );
  NAND2_X1 U9713 ( .A1(n8435), .A2(n5140), .ZN(n8437) );
  NAND2_X1 U9714 ( .A1(n7313), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U9715 ( .A1(n7155), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U9716 ( .A1(n7156), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U9717 ( .A1(n7539), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U9718 ( .A1(n8680), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8438) );
  OR2_X2 U9719 ( .A1(n8037), .A2(n9502), .ZN(n8439) );
  NAND4_X1 U9720 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n9517)
         );
  AOI22_X1 U9721 ( .A1(n8696), .A2(n9708), .B1(n8464), .B2(n9517), .ZN(n8693)
         );
  INV_X1 U9722 ( .A(n8443), .ZN(n8450) );
  INV_X1 U9723 ( .A(n8446), .ZN(n8449) );
  NOR2_X1 U9724 ( .A1(n8445), .A2(n8444), .ZN(n8447) );
  MUX2_X1 U9725 ( .A(n8447), .B(n8446), .S(n8464), .Z(n8448) );
  NAND2_X1 U9726 ( .A1(n8448), .A2(n8451), .ZN(n8485) );
  INV_X1 U9727 ( .A(n8485), .ZN(n8497) );
  OAI21_X1 U9728 ( .B1(n8450), .B2(n8449), .A(n8497), .ZN(n8452) );
  NAND3_X1 U9729 ( .A1(n8452), .A2(n8451), .A3(n8498), .ZN(n8487) );
  NAND2_X1 U9730 ( .A1(n8454), .A2(n8458), .ZN(n8453) );
  NAND2_X1 U9731 ( .A1(n8453), .A2(n8456), .ZN(n8461) );
  NAND2_X1 U9732 ( .A1(n8454), .A2(n7189), .ZN(n8457) );
  NAND3_X1 U9733 ( .A1(n8457), .A2(n8456), .A3(n8455), .ZN(n8459) );
  NAND2_X1 U9734 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  NAND2_X1 U9735 ( .A1(n8480), .A2(n8462), .ZN(n8466) );
  NAND2_X1 U9736 ( .A1(n8472), .A2(n8463), .ZN(n8465) );
  MUX2_X1 U9737 ( .A(n8466), .B(n8465), .S(n8464), .Z(n8467) );
  INV_X1 U9738 ( .A(n8467), .ZN(n8468) );
  OAI21_X1 U9739 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8471) );
  INV_X1 U9740 ( .A(n8472), .ZN(n8473) );
  OAI21_X1 U9741 ( .B1(n8474), .B2(n11117), .A(n8481), .ZN(n8476) );
  INV_X1 U9742 ( .A(n8477), .ZN(n8478) );
  NAND2_X1 U9743 ( .A1(n8481), .A2(n8483), .ZN(n8482) );
  AOI22_X1 U9744 ( .A1(n8484), .A2(n8483), .B1(n8464), .B2(n8482), .ZN(n8486)
         );
  INV_X1 U9745 ( .A(n8488), .ZN(n8489) );
  NOR2_X1 U9746 ( .A1(n8502), .A2(n8489), .ZN(n8490) );
  AOI21_X1 U9747 ( .B1(n8494), .B2(n8490), .A(n8499), .ZN(n8493) );
  INV_X1 U9748 ( .A(n8737), .ZN(n8492) );
  OAI21_X1 U9749 ( .B1(n8493), .B2(n8492), .A(n8491), .ZN(n8507) );
  INV_X1 U9750 ( .A(n8498), .ZN(n8500) );
  NOR3_X1 U9751 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(n8503) );
  OAI21_X1 U9752 ( .B1(n8503), .B2(n8502), .A(n8737), .ZN(n8504) );
  OAI21_X1 U9753 ( .B1(n9134), .B2(n8505), .A(n8504), .ZN(n8506) );
  MUX2_X1 U9754 ( .A(n8507), .B(n8506), .S(n8464), .Z(n8526) );
  OR2_X1 U9755 ( .A1(n8508), .A2(n7524), .ZN(n8510) );
  AOI22_X1 U9756 ( .A1(n7313), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7534), .B2(
        n9420), .ZN(n8509) );
  NAND2_X1 U9757 ( .A1(n7155), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U9758 ( .A1(n7539), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U9759 ( .A1(n7156), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8513) );
  AOI21_X1 U9760 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n8511), .A(n8534), .ZN(
        n9372) );
  OR2_X1 U9761 ( .A1(n8037), .A2(n9372), .ZN(n8512) );
  NAND4_X1 U9762 ( .A1(n8515), .A2(n8514), .A3(n8513), .A4(n8512), .ZN(n9694)
         );
  NAND2_X1 U9763 ( .A1(n9768), .A2(n9694), .ZN(n8516) );
  NAND2_X1 U9764 ( .A1(n9674), .A2(n9774), .ZN(n9657) );
  NAND2_X1 U9765 ( .A1(n8517), .A2(n5140), .ZN(n8519) );
  AOI22_X1 U9766 ( .A1(n7313), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7534), .B2(
        n9401), .ZN(n8518) );
  NAND2_X1 U9767 ( .A1(n8519), .A2(n8518), .ZN(n9232) );
  NAND2_X1 U9768 ( .A1(n9232), .A2(n9382), .ZN(n9194) );
  AND2_X1 U9769 ( .A1(n9382), .A2(n8695), .ZN(n8520) );
  AOI21_X1 U9770 ( .B1(n9232), .B2(n8464), .A(n8520), .ZN(n8521) );
  NAND2_X1 U9771 ( .A1(n9672), .A2(n8521), .ZN(n8527) );
  OAI21_X1 U9772 ( .B1(n9667), .B2(n9194), .A(n8527), .ZN(n8524) );
  NAND2_X1 U9773 ( .A1(n9190), .A2(n9383), .ZN(n8522) );
  NAND2_X1 U9774 ( .A1(n9328), .A2(n9688), .ZN(n8754) );
  MUX2_X1 U9775 ( .A(n8522), .B(n8754), .S(n8464), .Z(n8523) );
  OAI211_X1 U9776 ( .C1(n8526), .C2(n8525), .A(n8524), .B(n8523), .ZN(n8546)
         );
  INV_X1 U9777 ( .A(n8527), .ZN(n8540) );
  OR2_X1 U9778 ( .A1(n9232), .A2(n9382), .ZN(n8528) );
  NOR2_X1 U9779 ( .A1(n9774), .A2(n8695), .ZN(n8530) );
  NOR2_X1 U9780 ( .A1(n9694), .A2(n8464), .ZN(n8529) );
  MUX2_X1 U9781 ( .A(n8530), .B(n8529), .S(n9674), .Z(n8539) );
  NAND2_X1 U9782 ( .A1(n8531), .A2(n5140), .ZN(n8533) );
  AOI22_X1 U9783 ( .A1(n7313), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7534), .B2(
        n9439), .ZN(n8532) );
  NAND2_X1 U9784 ( .A1(n8533), .A2(n8532), .ZN(n9661) );
  NAND2_X1 U9785 ( .A1(n7155), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8538) );
  OAI21_X1 U9786 ( .B1(n9284), .B2(n8534), .A(n8550), .ZN(n9655) );
  INV_X1 U9787 ( .A(n9655), .ZN(n9287) );
  OR2_X1 U9788 ( .A1(n8037), .A2(n9287), .ZN(n8537) );
  OR2_X1 U9789 ( .A1(n8711), .A2(n8370), .ZN(n8536) );
  OR2_X1 U9790 ( .A1(n7548), .A2(n8359), .ZN(n8535) );
  OR2_X1 U9791 ( .A1(n9661), .A2(n9767), .ZN(n8541) );
  NAND2_X1 U9792 ( .A1(n9661), .A2(n9767), .ZN(n8542) );
  NAND2_X1 U9793 ( .A1(n8541), .A2(n8542), .ZN(n9660) );
  AOI211_X1 U9794 ( .C1(n8540), .C2(n9685), .A(n8539), .B(n9660), .ZN(n8545)
         );
  INV_X1 U9795 ( .A(n8541), .ZN(n8758) );
  INV_X1 U9796 ( .A(n8542), .ZN(n8543) );
  MUX2_X1 U9797 ( .A(n8758), .B(n8543), .S(n8464), .Z(n8544) );
  AOI21_X1 U9798 ( .B1(n8546), .B2(n8545), .A(n8544), .ZN(n8582) );
  NAND2_X1 U9799 ( .A1(n8547), .A2(n5140), .ZN(n8549) );
  AOI22_X1 U9800 ( .A1(n7313), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7534), .B2(
        n9457), .ZN(n8548) );
  OR2_X1 U9801 ( .A1(n7548), .A2(n9453), .ZN(n8554) );
  NAND2_X1 U9802 ( .A1(n7155), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U9803 ( .A1(n7539), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8552) );
  AOI21_X1 U9804 ( .B1(n8550), .B2(P2_REG3_REG_17__SCAN_IN), .A(n8559), .ZN(
        n9648) );
  OR2_X1 U9805 ( .A1(n8037), .A2(n9648), .ZN(n8551) );
  NAND4_X1 U9806 ( .A1(n8554), .A2(n8553), .A3(n8552), .A4(n8551), .ZN(n9628)
         );
  MUX2_X1 U9807 ( .A(n9755), .B(n9628), .S(n8464), .Z(n8581) );
  NAND2_X1 U9808 ( .A1(n8582), .A2(n8581), .ZN(n8565) );
  OR2_X1 U9809 ( .A1(n8555), .A2(n7524), .ZN(n8558) );
  AOI22_X1 U9810 ( .A1(n7313), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7534), .B2(
        n8556), .ZN(n8557) );
  INV_X1 U9811 ( .A(n9748), .ZN(n9635) );
  NAND2_X1 U9812 ( .A1(n7155), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U9813 ( .A1(n7539), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U9814 ( .A1(n7156), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8561) );
  XNOR2_X1 U9815 ( .A(P2_REG3_REG_18__SCAN_IN), .B(n8559), .ZN(n9632) );
  OR2_X1 U9816 ( .A1(n8037), .A2(n9632), .ZN(n8560) );
  NAND4_X1 U9817 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8560), .ZN(n9613)
         );
  NAND2_X1 U9818 ( .A1(n9635), .A2(n9757), .ZN(n8580) );
  NAND3_X1 U9819 ( .A1(n8565), .A2(n8580), .A3(n9628), .ZN(n8564) );
  AND2_X1 U9820 ( .A1(n9748), .A2(n9613), .ZN(n8566) );
  NAND2_X1 U9821 ( .A1(n8564), .A2(n8762), .ZN(n8569) );
  NAND2_X1 U9822 ( .A1(n8565), .A2(n9755), .ZN(n8567) );
  AOI21_X1 U9823 ( .B1(n8567), .B2(n8580), .A(n8566), .ZN(n8568) );
  MUX2_X1 U9824 ( .A(n8569), .B(n8568), .S(n8464), .Z(n8584) );
  NAND2_X1 U9825 ( .A1(n7156), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U9826 ( .A1(n7155), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U9827 ( .A1(n7539), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8574) );
  INV_X1 U9828 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U9829 ( .A1(n8571), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8572) );
  AND2_X1 U9830 ( .A1(n8591), .A2(n8572), .ZN(n9618) );
  OR2_X1 U9831 ( .A1(n8037), .A2(n9618), .ZN(n8573) );
  NAND4_X1 U9832 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n9629)
         );
  NAND2_X1 U9833 ( .A1(n8577), .A2(n5140), .ZN(n8579) );
  AOI22_X1 U9834 ( .A1(n7313), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7534), .B2(
        n7153), .ZN(n8578) );
  XOR2_X1 U9835 ( .A(n9629), .B(n9744), .Z(n9616) );
  NAND2_X1 U9836 ( .A1(n8762), .A2(n8580), .ZN(n9626) );
  NOR3_X1 U9837 ( .A1(n8582), .A2(n8581), .A3(n9626), .ZN(n8583) );
  NOR3_X1 U9838 ( .A1(n8584), .A2(n9616), .A3(n8583), .ZN(n8598) );
  INV_X1 U9839 ( .A(n9744), .ZN(n9617) );
  NOR2_X1 U9840 ( .A1(n9617), .A2(n8464), .ZN(n8586) );
  NOR2_X1 U9841 ( .A1(n9744), .A2(n8695), .ZN(n8585) );
  MUX2_X1 U9842 ( .A(n8586), .B(n8585), .S(n9629), .Z(n8597) );
  NAND2_X1 U9843 ( .A1(n8587), .A2(n5140), .ZN(n8589) );
  NAND2_X1 U9844 ( .A1(n7313), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U9845 ( .A1(n7156), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8596) );
  INV_X1 U9846 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8590) );
  OR2_X1 U9847 ( .A1(n8708), .A2(n8590), .ZN(n8595) );
  NAND2_X1 U9848 ( .A1(n8591), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8592) );
  AND2_X1 U9849 ( .A1(n8603), .A2(n8592), .ZN(n9604) );
  OR2_X1 U9850 ( .A1(n8037), .A2(n9604), .ZN(n8594) );
  INV_X1 U9851 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9605) );
  OR2_X1 U9852 ( .A1(n8711), .A2(n9605), .ZN(n8593) );
  NAND2_X1 U9853 ( .A1(n9740), .A2(n9268), .ZN(n8610) );
  NAND2_X1 U9854 ( .A1(n8764), .A2(n8610), .ZN(n9607) );
  NOR3_X1 U9855 ( .A1(n8598), .A2(n8597), .A3(n9607), .ZN(n8624) );
  NAND2_X1 U9856 ( .A1(n8599), .A2(n5140), .ZN(n8601) );
  NAND2_X1 U9857 ( .A1(n7313), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U9858 ( .A1(n7156), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8609) );
  INV_X1 U9859 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8602) );
  OR2_X1 U9860 ( .A1(n8708), .A2(n8602), .ZN(n8608) );
  NAND2_X1 U9861 ( .A1(n8603), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8604) );
  AND2_X1 U9862 ( .A1(n8615), .A2(n8604), .ZN(n9266) );
  OR2_X1 U9863 ( .A1(n8037), .A2(n9266), .ZN(n8607) );
  INV_X1 U9864 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8605) );
  OR2_X1 U9865 ( .A1(n8711), .A2(n8605), .ZN(n8606) );
  NAND2_X1 U9866 ( .A1(n9736), .A2(n9337), .ZN(n8621) );
  MUX2_X1 U9867 ( .A(n8764), .B(n8610), .S(n8464), .Z(n8611) );
  NAND2_X1 U9868 ( .A1(n9564), .A2(n8611), .ZN(n8623) );
  NAND2_X1 U9869 ( .A1(n8612), .A2(n5140), .ZN(n8614) );
  NAND2_X1 U9870 ( .A1(n7313), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U9871 ( .A1(n7156), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U9872 ( .A1(n7155), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U9873 ( .A1(n7539), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U9874 ( .A1(n8615), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8616) );
  AND2_X1 U9875 ( .A1(n8630), .A2(n8616), .ZN(n9584) );
  OR2_X1 U9876 ( .A1(n8037), .A2(n9584), .ZN(n8617) );
  XNOR2_X1 U9877 ( .A(n9732), .B(n9593), .ZN(n9582) );
  MUX2_X1 U9878 ( .A(n8621), .B(n9565), .S(n8464), .Z(n8622) );
  INV_X1 U9879 ( .A(n9732), .ZN(n9587) );
  NAND2_X1 U9880 ( .A1(n9587), .A2(n9593), .ZN(n8625) );
  INV_X1 U9881 ( .A(n9593), .ZN(n9250) );
  NAND2_X1 U9882 ( .A1(n9732), .A2(n9250), .ZN(n9567) );
  MUX2_X1 U9883 ( .A(n8625), .B(n9567), .S(n8464), .Z(n8638) );
  NAND2_X1 U9884 ( .A1(n8626), .A2(n5140), .ZN(n8628) );
  NAND2_X1 U9885 ( .A1(n7313), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U9886 ( .A1(n7156), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8636) );
  INV_X1 U9887 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8629) );
  OR2_X1 U9888 ( .A1(n8708), .A2(n8629), .ZN(n8635) );
  NAND2_X1 U9889 ( .A1(n8630), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8631) );
  AND2_X1 U9890 ( .A1(n8644), .A2(n8631), .ZN(n9248) );
  OR2_X1 U9891 ( .A1(n8037), .A2(n9248), .ZN(n8634) );
  INV_X1 U9892 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8632) );
  OR2_X1 U9893 ( .A1(n8711), .A2(n8632), .ZN(n8633) );
  OR2_X1 U9894 ( .A1(n8637), .A2(n9246), .ZN(n8768) );
  NAND2_X1 U9895 ( .A1(n8637), .A2(n9246), .ZN(n8766) );
  NAND2_X1 U9896 ( .A1(n8768), .A2(n8766), .ZN(n9569) );
  NAND2_X1 U9897 ( .A1(n8639), .A2(n5140), .ZN(n8641) );
  NAND2_X1 U9898 ( .A1(n7313), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U9899 ( .A1(n7156), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8649) );
  INV_X1 U9900 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8642) );
  OR2_X1 U9901 ( .A1(n8708), .A2(n8642), .ZN(n8648) );
  INV_X1 U9902 ( .A(n8643), .ZN(n8653) );
  NAND2_X1 U9903 ( .A1(n8644), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8645) );
  OR2_X1 U9904 ( .A1(n8037), .A2(n9555), .ZN(n8647) );
  INV_X1 U9905 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9556) );
  OR2_X1 U9906 ( .A1(n8711), .A2(n9556), .ZN(n8646) );
  NAND2_X1 U9907 ( .A1(n9725), .A2(n9277), .ZN(n8772) );
  MUX2_X1 U9908 ( .A(n8768), .B(n8766), .S(n8464), .Z(n8650) );
  MUX2_X1 U9909 ( .A(n8772), .B(n8773), .S(n8464), .Z(n8659) );
  NAND2_X1 U9910 ( .A1(n7313), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U9911 ( .A1(n7156), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U9912 ( .A1(n7155), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U9913 ( .A1(n7539), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U9914 ( .A1(n8653), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8654) );
  AND2_X1 U9915 ( .A1(n8667), .A2(n8654), .ZN(n9540) );
  OR2_X1 U9916 ( .A1(n8037), .A2(n9540), .ZN(n8655) );
  NAND2_X1 U9917 ( .A1(n9541), .A2(n9549), .ZN(n8660) );
  INV_X1 U9918 ( .A(n9549), .ZN(n9362) );
  NAND2_X1 U9919 ( .A1(n9721), .A2(n9362), .ZN(n8774) );
  MUX2_X1 U9920 ( .A(n8660), .B(n8774), .S(n8464), .Z(n8661) );
  NAND2_X1 U9921 ( .A1(n8662), .A2(n5140), .ZN(n8664) );
  NAND2_X1 U9922 ( .A1(n7313), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U9923 ( .A1(n7156), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8673) );
  INV_X1 U9924 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8665) );
  OR2_X1 U9925 ( .A1(n8708), .A2(n8665), .ZN(n8672) );
  INV_X1 U9926 ( .A(n8666), .ZN(n8678) );
  NAND2_X1 U9927 ( .A1(n8667), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8668) );
  AND2_X1 U9928 ( .A1(n8678), .A2(n8668), .ZN(n9358) );
  OR2_X1 U9929 ( .A1(n8037), .A2(n9358), .ZN(n8671) );
  INV_X1 U9930 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8669) );
  OR2_X1 U9931 ( .A1(n8711), .A2(n8669), .ZN(n8670) );
  NAND2_X1 U9932 ( .A1(n9717), .A2(n9162), .ZN(n9513) );
  NAND2_X1 U9933 ( .A1(n9182), .A2(n9513), .ZN(n9532) );
  NAND2_X1 U9934 ( .A1(n8674), .A2(n5140), .ZN(n8676) );
  NAND2_X1 U9935 ( .A1(n7313), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U9936 ( .A1(n7156), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8684) );
  INV_X1 U9937 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8677) );
  OR2_X1 U9938 ( .A1(n8708), .A2(n8677), .ZN(n8683) );
  NAND2_X1 U9939 ( .A1(n8678), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8679) );
  INV_X1 U9940 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9522) );
  OR2_X1 U9941 ( .A1(n8711), .A2(n9522), .ZN(n8681) );
  NAND2_X1 U9942 ( .A1(n9713), .A2(n9531), .ZN(n9184) );
  MUX2_X1 U9943 ( .A(n9513), .B(n9182), .S(n8464), .Z(n8685) );
  OAI211_X1 U9944 ( .C1(n8686), .C2(n9532), .A(n9200), .B(n8685), .ZN(n8688)
         );
  MUX2_X1 U9945 ( .A(n9185), .B(n9184), .S(n8464), .Z(n8687) );
  NAND2_X1 U9946 ( .A1(n8688), .A2(n8687), .ZN(n8692) );
  MUX2_X1 U9947 ( .A(n9517), .B(n9708), .S(n8464), .Z(n8689) );
  AOI21_X1 U9948 ( .B1(n8692), .B2(n8693), .A(n8689), .ZN(n8690) );
  INV_X1 U9949 ( .A(n8690), .ZN(n8691) );
  NAND2_X1 U9950 ( .A1(n9703), .A2(n9505), .ZN(n8720) );
  OAI211_X1 U9951 ( .C1(n8693), .C2(n8692), .A(n8691), .B(n9201), .ZN(n8697)
         );
  INV_X1 U9952 ( .A(n8786), .ZN(n8694) );
  AOI211_X1 U9953 ( .C1(n8697), .C2(n8720), .A(n8695), .B(n8694), .ZN(n8750)
         );
  NAND2_X1 U9954 ( .A1(n8697), .A2(n8696), .ZN(n8719) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8701), .Z(n8702) );
  INV_X1 U9956 ( .A(SI_31_), .ZN(n9939) );
  XNOR2_X1 U9957 ( .A(n8702), .B(n9939), .ZN(n8703) );
  NAND2_X1 U9958 ( .A1(n10821), .A2(n5140), .ZN(n8706) );
  NAND2_X1 U9959 ( .A1(n7313), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U9960 ( .A1(n8706), .A2(n8705), .ZN(n8784) );
  INV_X1 U9961 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8707) );
  OR2_X1 U9962 ( .A1(n8708), .A2(n8707), .ZN(n8714) );
  INV_X1 U9963 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8709) );
  OR2_X1 U9964 ( .A1(n7548), .A2(n8709), .ZN(n8713) );
  INV_X1 U9965 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8710) );
  OR2_X1 U9966 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  INV_X1 U9967 ( .A(n8717), .ZN(n9381) );
  OAI22_X1 U9968 ( .A1(n8784), .A2(n8751), .B1(n9702), .B2(n9381), .ZN(n8722)
         );
  NOR2_X1 U9969 ( .A1(n8722), .A2(n8746), .ZN(n8718) );
  INV_X1 U9970 ( .A(n8720), .ZN(n8721) );
  NOR2_X1 U9971 ( .A1(n8722), .A2(n8721), .ZN(n8782) );
  NAND2_X1 U9972 ( .A1(n9708), .A2(n9227), .ZN(n8778) );
  NAND2_X1 U9973 ( .A1(n9187), .A2(n8778), .ZN(n9499) );
  INV_X1 U9974 ( .A(n9607), .ZN(n9198) );
  INV_X1 U9975 ( .A(n9626), .ZN(n9622) );
  NOR4_X1 U9976 ( .A1(n8725), .A2(n7189), .A3(n8724), .A4(n8723), .ZN(n8732)
         );
  NOR3_X1 U9977 ( .A1(n8728), .A2(n8727), .A3(n8726), .ZN(n8731) );
  NAND4_X1 U9978 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n8734)
         );
  NOR4_X1 U9979 ( .A1(n8736), .A2(n8735), .A3(n8734), .A4(n8733), .ZN(n8738)
         );
  NAND4_X1 U9980 ( .A1(n8752), .A2(n8739), .A3(n8738), .A4(n8737), .ZN(n8740)
         );
  NOR4_X1 U9981 ( .A1(n9660), .A2(n9685), .A3(n9667), .A4(n8740), .ZN(n8741)
         );
  XNOR2_X1 U9982 ( .A(n9755), .B(n9628), .ZN(n9641) );
  NAND4_X1 U9983 ( .A1(n9198), .A2(n9622), .A3(n8741), .A4(n9641), .ZN(n8742)
         );
  NOR4_X1 U9984 ( .A1(n9569), .A2(n9616), .A3(n9595), .A4(n8742), .ZN(n8743)
         );
  NAND4_X1 U9985 ( .A1(n9545), .A2(n9553), .A3(n8743), .A4(n9582), .ZN(n8744)
         );
  NOR4_X1 U9986 ( .A1(n9499), .A2(n9516), .A3(n9532), .A4(n8744), .ZN(n8745)
         );
  NAND4_X1 U9987 ( .A1(n8782), .A2(n8745), .A3(n8786), .A4(n8779), .ZN(n8747)
         );
  NAND2_X1 U9988 ( .A1(n8747), .A2(n8746), .ZN(n8748) );
  NOR2_X1 U9989 ( .A1(n9700), .A2(n9493), .ZN(n8789) );
  NOR2_X1 U9990 ( .A1(n8789), .A2(n8787), .ZN(n8792) );
  NAND2_X1 U9991 ( .A1(n8753), .A2(n8752), .ZN(n8755) );
  OR2_X1 U9992 ( .A1(n9232), .A2(n9669), .ZN(n8756) );
  INV_X1 U9993 ( .A(n9657), .ZN(n8757) );
  NOR2_X1 U9994 ( .A1(n9660), .A2(n8757), .ZN(n9658) );
  OR2_X1 U9995 ( .A1(n8758), .A2(n9658), .ZN(n8759) );
  NAND2_X1 U9996 ( .A1(n9638), .A2(n9641), .ZN(n9640) );
  INV_X1 U9997 ( .A(n9628), .ZN(n9761) );
  OR2_X1 U9998 ( .A1(n9755), .A2(n9761), .ZN(n8761) );
  NAND2_X1 U9999 ( .A1(n9640), .A2(n8761), .ZN(n9623) );
  INV_X1 U10000 ( .A(n9629), .ZN(n9347) );
  NAND2_X1 U10001 ( .A1(n9744), .A2(n9347), .ZN(n8763) );
  NAND2_X1 U10002 ( .A1(n9608), .A2(n9198), .ZN(n8765) );
  AND2_X1 U10003 ( .A1(n9567), .A2(n8766), .ZN(n8767) );
  AND2_X1 U10004 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  INV_X1 U10005 ( .A(n8770), .ZN(n8771) );
  INV_X1 U10006 ( .A(n9513), .ZN(n8775) );
  OAI211_X1 U10007 ( .C1(n9183), .C2(n8775), .A(n9182), .B(n9185), .ZN(n8777)
         );
  INV_X1 U10008 ( .A(n9187), .ZN(n8776) );
  AOI21_X1 U10009 ( .B1(n8777), .B2(n9184), .A(n8776), .ZN(n8781) );
  INV_X1 U10010 ( .A(n8778), .ZN(n8780) );
  OAI21_X1 U10011 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8783) );
  INV_X1 U10012 ( .A(n8788), .ZN(n8793) );
  INV_X1 U10013 ( .A(n8789), .ZN(n8790) );
  NOR2_X1 U10014 ( .A1(n8790), .A2(n7153), .ZN(n8791) );
  AOI211_X1 U10015 ( .C1(n8793), .C2(n8792), .A(n8791), .B(n8799), .ZN(n8794)
         );
  NAND3_X1 U10016 ( .A1(n8797), .A2(n8796), .A3(n7159), .ZN(n8798) );
  OAI211_X1 U10017 ( .C1(n8800), .C2(n8799), .A(n8798), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8801) );
  NAND2_X1 U10018 ( .A1(n8802), .A2(n10651), .ZN(n8811) );
  INV_X1 U10019 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8805) );
  NAND3_X1 U10020 ( .A1(n8803), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n10632), 
        .ZN(n8804) );
  OAI21_X1 U10021 ( .B1(n10601), .B2(n8805), .A(n8804), .ZN(n8808) );
  NOR2_X1 U10022 ( .A1(n8806), .A2(n10576), .ZN(n8807) );
  AOI211_X1 U10023 ( .C1(n10580), .C2(n8809), .A(n8808), .B(n8807), .ZN(n8810)
         );
  OAI211_X1 U10024 ( .C1(n8812), .C2(n7511), .A(n8811), .B(n8810), .ZN(
        P1_U3356) );
  OAI21_X1 U10025 ( .B1(n8814), .B2(n8874), .A(n8813), .ZN(n10771) );
  INV_X1 U10026 ( .A(n8815), .ZN(n8818) );
  INV_X1 U10027 ( .A(n8816), .ZN(n8817) );
  AOI211_X1 U10028 ( .C1(n10767), .C2(n8818), .A(n10655), .B(n8817), .ZN(
        n10765) );
  NAND2_X1 U10029 ( .A1(n10767), .A2(n10580), .ZN(n8821) );
  AOI22_X1 U10030 ( .A1(n7511), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8819), .B2(
        n10632), .ZN(n8820) );
  OAI211_X1 U10031 ( .C1(n10764), .C2(n10488), .A(n8821), .B(n8820), .ZN(n8826) );
  XNOR2_X1 U10032 ( .A(n8822), .B(n8874), .ZN(n8824) );
  AOI22_X1 U10033 ( .A1(n8824), .A2(n10746), .B1(n11155), .B2(n8823), .ZN(
        n10769) );
  NOR2_X1 U10034 ( .A1(n10769), .A2(n7511), .ZN(n8825) );
  AOI211_X1 U10035 ( .C1(n10765), .C2(n10664), .A(n8826), .B(n8825), .ZN(n8827) );
  OAI21_X1 U10036 ( .B1(n10638), .B2(n10771), .A(n8827), .ZN(P1_U3278) );
  AOI22_X1 U10037 ( .A1(n8828), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9802), .ZN(n8829) );
  OAI21_X1 U10038 ( .B1(n8830), .B2(n9804), .A(n8829), .ZN(P2_U3270) );
  INV_X1 U10039 ( .A(n8832), .ZN(n8833) );
  AOI21_X1 U10040 ( .B1(n8834), .B2(n8831), .A(n8833), .ZN(n8838) );
  AOI22_X1 U10041 ( .A1(n10356), .A2(n9932), .B1(n9928), .B2(n6434), .ZN(n8837) );
  AOI22_X1 U10042 ( .A1(n9904), .A2(n6869), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8835), .ZN(n8836) );
  OAI211_X1 U10043 ( .C1(n8838), .C2(n9919), .A(n8837), .B(n8836), .ZN(
        P1_U3237) );
  AOI22_X1 U10044 ( .A1(n8839), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9802), .ZN(n8840) );
  OAI21_X1 U10045 ( .B1(n8841), .B2(n9800), .A(n8840), .ZN(P2_U3266) );
  INV_X1 U10046 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8843) );
  OAI222_X1 U10047 ( .A1(n8844), .A2(n8843), .B1(n7237), .B2(P2_U3151), .C1(
        n9800), .C2(n8842), .ZN(P2_U3293) );
  NAND2_X1 U10048 ( .A1(n10464), .A2(n9054), .ZN(n9014) );
  NAND2_X1 U10049 ( .A1(n10821), .A2(n8854), .ZN(n8846) );
  INV_X1 U10050 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10817) );
  OR2_X1 U10051 ( .A1(n8853), .A2(n10817), .ZN(n8845) );
  NAND2_X1 U10052 ( .A1(n8847), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U10053 ( .A1(n8848), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U10054 ( .A1(n5960), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8849) );
  NAND3_X1 U10055 ( .A1(n8851), .A2(n8850), .A3(n8849), .ZN(n10475) );
  INV_X1 U10056 ( .A(n10475), .ZN(n8852) );
  OR2_X1 U10057 ( .A1(n10472), .A2(n8852), .ZN(n9118) );
  INV_X1 U10058 ( .A(n9118), .ZN(n9017) );
  NAND2_X1 U10059 ( .A1(n10472), .A2(n8852), .ZN(n9039) );
  INV_X1 U10060 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9221) );
  INV_X1 U10061 ( .A(n10779), .ZN(n10471) );
  INV_X1 U10062 ( .A(n9937), .ZN(n8856) );
  NOR2_X1 U10063 ( .A1(n10471), .A2(n8856), .ZN(n9004) );
  INV_X1 U10064 ( .A(n9004), .ZN(n8855) );
  NAND2_X1 U10065 ( .A1(n9039), .A2(n8855), .ZN(n9117) );
  AND2_X1 U10066 ( .A1(n10471), .A2(n8856), .ZN(n9110) );
  INV_X1 U10067 ( .A(n10624), .ZN(n8879) );
  INV_X1 U10068 ( .A(n10642), .ZN(n10649) );
  INV_X1 U10069 ( .A(n8857), .ZN(n8929) );
  INV_X1 U10070 ( .A(n8917), .ZN(n8864) );
  NOR4_X1 U10071 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n8862)
         );
  NAND4_X1 U10072 ( .A1(n8865), .A2(n8864), .A3(n8863), .A4(n8862), .ZN(n8867)
         );
  NOR4_X1 U10073 ( .A1(n8914), .A2(n8868), .A3(n8867), .A4(n8866), .ZN(n8869)
         );
  NAND4_X1 U10074 ( .A1(n8870), .A2(n8929), .A3(n8928), .A4(n8869), .ZN(n8871)
         );
  NOR4_X1 U10075 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8871), .ZN(n8875)
         );
  NAND4_X1 U10076 ( .A1(n8952), .A2(n8943), .A3(n8876), .A4(n8875), .ZN(n8877)
         );
  NOR4_X1 U10077 ( .A1(n8879), .A2(n8878), .A3(n10649), .A4(n8877), .ZN(n8880)
         );
  NAND4_X1 U10078 ( .A1(n10566), .A2(n5418), .A3(n10615), .A4(n8880), .ZN(
        n8881) );
  NOR4_X1 U10079 ( .A1(n10526), .A2(n10550), .A3(n10536), .A4(n8881), .ZN(
        n8882) );
  NAND4_X1 U10080 ( .A1(n6401), .A2(n10500), .A3(n8998), .A4(n8882), .ZN(n8883) );
  NOR4_X1 U10081 ( .A1(n9017), .A2(n9117), .A3(n9110), .A4(n8883), .ZN(n9018)
         );
  AND2_X1 U10082 ( .A1(n8978), .A2(n8884), .ZN(n8885) );
  NAND2_X1 U10083 ( .A1(n8979), .A2(n8885), .ZN(n9021) );
  NAND2_X1 U10084 ( .A1(n8886), .A2(n9094), .ZN(n8888) );
  NAND2_X1 U10085 ( .A1(n8973), .A2(n8959), .ZN(n8887) );
  MUX2_X1 U10086 ( .A(n8888), .B(n8887), .S(n9011), .Z(n8889) );
  INV_X1 U10087 ( .A(n8889), .ZN(n8967) );
  INV_X1 U10088 ( .A(n8890), .ZN(n9093) );
  NOR2_X1 U10089 ( .A1(n8957), .A2(n9093), .ZN(n8956) );
  AND2_X1 U10090 ( .A1(n9078), .A2(n8895), .ZN(n8903) );
  INV_X1 U10091 ( .A(n8891), .ZN(n8892) );
  NAND2_X1 U10092 ( .A1(n8894), .A2(n8892), .ZN(n8893) );
  AND2_X1 U10093 ( .A1(n8893), .A2(n9077), .ZN(n8900) );
  NAND2_X1 U10094 ( .A1(n8895), .A2(n8894), .ZN(n9075) );
  INV_X1 U10095 ( .A(n8896), .ZN(n8897) );
  AND2_X1 U10096 ( .A1(n9077), .A2(n8897), .ZN(n8898) );
  NOR2_X1 U10097 ( .A1(n9075), .A2(n8898), .ZN(n8899) );
  INV_X1 U10098 ( .A(n9011), .ZN(n9002) );
  MUX2_X1 U10099 ( .A(n8900), .B(n8899), .S(n9002), .Z(n8932) );
  INV_X1 U10100 ( .A(n8901), .ZN(n8902) );
  NAND2_X1 U10101 ( .A1(n8940), .A2(n8931), .ZN(n9080) );
  NAND2_X1 U10102 ( .A1(n8904), .A2(n9058), .ZN(n8906) );
  NAND3_X1 U10103 ( .A1(n8906), .A2(n9061), .A3(n8905), .ZN(n8907) );
  NAND3_X1 U10104 ( .A1(n8907), .A2(n9057), .A3(n9063), .ZN(n8909) );
  MUX2_X1 U10105 ( .A(n8909), .B(n8908), .S(n9011), .Z(n8918) );
  INV_X1 U10106 ( .A(n9064), .ZN(n8913) );
  OR2_X1 U10107 ( .A1(n8913), .A2(n8910), .ZN(n8912) );
  NAND2_X1 U10108 ( .A1(n8912), .A2(n8911), .ZN(n9066) );
  MUX2_X1 U10109 ( .A(n9066), .B(n8913), .S(n9011), .Z(n8915) );
  NOR2_X1 U10110 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  OAI21_X1 U10111 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(n8920) );
  MUX2_X1 U10112 ( .A(n9070), .B(n9067), .S(n9011), .Z(n8919) );
  NAND3_X1 U10113 ( .A1(n8920), .A2(n5397), .A3(n8919), .ZN(n8925) );
  MUX2_X1 U10114 ( .A(n8922), .B(n8921), .S(n9002), .Z(n8923) );
  NAND3_X1 U10115 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n8930) );
  OR2_X1 U10116 ( .A1(n8926), .A2(n9002), .ZN(n8927) );
  NAND4_X1 U10117 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n8933)
         );
  NAND3_X1 U10118 ( .A1(n8933), .A2(n8932), .A3(n8931), .ZN(n8934) );
  NAND2_X1 U10119 ( .A1(n8935), .A2(n8934), .ZN(n8941) );
  NAND2_X1 U10120 ( .A1(n8941), .A2(n9078), .ZN(n8936) );
  NAND2_X1 U10121 ( .A1(n8936), .A2(n9083), .ZN(n8939) );
  NAND2_X1 U10122 ( .A1(n8948), .A2(n9084), .ZN(n8937) );
  AOI21_X1 U10123 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n8946) );
  NAND2_X1 U10124 ( .A1(n8947), .A2(n8942), .ZN(n9053) );
  AOI21_X1 U10125 ( .B1(n8944), .B2(n8943), .A(n9053), .ZN(n8945) );
  NAND2_X1 U10126 ( .A1(n9087), .A2(n8947), .ZN(n8949) );
  NAND2_X1 U10127 ( .A1(n8950), .A2(n8948), .ZN(n9052) );
  MUX2_X1 U10128 ( .A(n8949), .B(n9052), .S(n9011), .Z(n8953) );
  MUX2_X1 U10129 ( .A(n8950), .B(n9087), .S(n9011), .Z(n8951) );
  OAI211_X1 U10130 ( .C1(n8954), .C2(n8953), .A(n8952), .B(n8951), .ZN(n8962)
         );
  INV_X1 U10131 ( .A(n8961), .ZN(n8955) );
  AOI21_X1 U10132 ( .B1(n8956), .B2(n8962), .A(n8955), .ZN(n8964) );
  INV_X1 U10133 ( .A(n8957), .ZN(n8958) );
  NAND2_X1 U10134 ( .A1(n8959), .A2(n8958), .ZN(n9051) );
  AND2_X1 U10135 ( .A1(n8961), .A2(n8960), .ZN(n9091) );
  MUX2_X1 U10136 ( .A(n8964), .B(n8963), .S(n9002), .Z(n8965) );
  NAND2_X1 U10137 ( .A1(n8965), .A2(n9094), .ZN(n8966) );
  INV_X1 U10138 ( .A(n8974), .ZN(n8968) );
  NAND2_X1 U10139 ( .A1(n8982), .A2(n8969), .ZN(n8970) );
  NAND2_X1 U10140 ( .A1(n8970), .A2(n8979), .ZN(n9023) );
  OAI211_X1 U10141 ( .C1(n9021), .C2(n8971), .A(n9023), .B(n9011), .ZN(n8972)
         );
  INV_X1 U10142 ( .A(n8989), .ZN(n8985) );
  AND2_X1 U10143 ( .A1(n8974), .A2(n8973), .ZN(n9050) );
  INV_X1 U10144 ( .A(n8975), .ZN(n8976) );
  AOI21_X1 U10145 ( .B1(n8977), .B2(n9050), .A(n8976), .ZN(n8980) );
  OAI211_X1 U10146 ( .C1(n8981), .C2(n8980), .A(n8979), .B(n8978), .ZN(n8983)
         );
  NAND2_X1 U10147 ( .A1(n8983), .A2(n8982), .ZN(n8984) );
  OAI211_X1 U10148 ( .C1(n8985), .C2(n8984), .A(n9024), .B(n8991), .ZN(n8986)
         );
  NAND2_X1 U10149 ( .A1(n8987), .A2(n8992), .ZN(n8988) );
  NAND2_X1 U10150 ( .A1(n8992), .A2(n8991), .ZN(n9105) );
  NAND2_X1 U10151 ( .A1(n8993), .A2(n9028), .ZN(n8994) );
  NAND2_X1 U10152 ( .A1(n8994), .A2(n9011), .ZN(n8995) );
  NAND2_X1 U10153 ( .A1(n8996), .A2(n8995), .ZN(n8999) );
  MUX2_X1 U10154 ( .A(n9029), .B(n9019), .S(n9011), .Z(n8997) );
  OAI211_X1 U10155 ( .C1(n8999), .C2(n10508), .A(n8998), .B(n8997), .ZN(n9001)
         );
  MUX2_X1 U10156 ( .A(n9020), .B(n9031), .S(n9011), .Z(n9000) );
  AOI21_X1 U10157 ( .B1(n10475), .B2(n9937), .A(n10779), .ZN(n9007) );
  INV_X1 U10158 ( .A(n9111), .ZN(n9035) );
  NOR2_X1 U10159 ( .A1(n9007), .A2(n9035), .ZN(n9003) );
  MUX2_X1 U10160 ( .A(n9003), .B(n9032), .S(n9002), .Z(n9005) );
  NAND2_X1 U10161 ( .A1(n9004), .A2(n10475), .ZN(n9034) );
  INV_X1 U10162 ( .A(n9007), .ZN(n9037) );
  NAND2_X1 U10163 ( .A1(n9010), .A2(n9009), .ZN(n9013) );
  NAND2_X1 U10164 ( .A1(n9034), .A2(n9039), .ZN(n9012) );
  AOI211_X1 U10165 ( .C1(n9015), .C2(n9014), .A(n9018), .B(n9016), .ZN(n9046)
         );
  INV_X1 U10166 ( .A(n9018), .ZN(n9043) );
  AND2_X1 U10167 ( .A1(n9020), .A2(n9019), .ZN(n9047) );
  INV_X1 U10168 ( .A(n9021), .ZN(n9022) );
  AND2_X1 U10169 ( .A1(n9024), .A2(n9022), .ZN(n9049) );
  INV_X1 U10170 ( .A(n9023), .ZN(n9025) );
  NAND2_X1 U10171 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  NAND3_X1 U10172 ( .A1(n9027), .A2(n10532), .A3(n9026), .ZN(n9103) );
  AOI21_X1 U10173 ( .B1(n9049), .B2(n10613), .A(n9103), .ZN(n9030) );
  AND2_X1 U10174 ( .A1(n9029), .A2(n9028), .ZN(n9048) );
  OAI21_X1 U10175 ( .B1(n9030), .B2(n9105), .A(n9048), .ZN(n9033) );
  NAND2_X1 U10176 ( .A1(n9032), .A2(n9031), .ZN(n9113) );
  AOI21_X1 U10177 ( .B1(n9047), .B2(n9033), .A(n9113), .ZN(n9036) );
  OAI21_X1 U10178 ( .B1(n9036), .B2(n9035), .A(n9034), .ZN(n9038) );
  NAND3_X1 U10179 ( .A1(n9038), .A2(n9037), .A3(n9118), .ZN(n9041) );
  NAND3_X1 U10180 ( .A1(n9041), .A2(n9040), .A3(n9039), .ZN(n9042) );
  AOI21_X1 U10181 ( .B1(n9043), .B2(n9042), .A(n10464), .ZN(n9044) );
  NOR4_X1 U10182 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9120), .ZN(n9130)
         );
  INV_X1 U10183 ( .A(n9047), .ZN(n9109) );
  INV_X1 U10184 ( .A(n9048), .ZN(n9107) );
  INV_X1 U10185 ( .A(n9049), .ZN(n9101) );
  INV_X1 U10186 ( .A(n9050), .ZN(n9099) );
  INV_X1 U10187 ( .A(n9051), .ZN(n9097) );
  INV_X1 U10188 ( .A(n9052), .ZN(n9090) );
  INV_X1 U10189 ( .A(n9053), .ZN(n9086) );
  AOI21_X1 U10190 ( .B1(n6434), .B2(n5941), .A(n9054), .ZN(n9056) );
  AND2_X1 U10191 ( .A1(n9056), .A2(n9055), .ZN(n9059) );
  OAI211_X1 U10192 ( .C1(n9060), .C2(n9059), .A(n9058), .B(n9057), .ZN(n9062)
         );
  NAND2_X1 U10193 ( .A1(n9062), .A2(n9061), .ZN(n9065) );
  NAND3_X1 U10194 ( .A1(n9065), .A2(n9064), .A3(n9063), .ZN(n9069) );
  INV_X1 U10195 ( .A(n9066), .ZN(n9068) );
  NAND3_X1 U10196 ( .A1(n9069), .A2(n9068), .A3(n9067), .ZN(n9072) );
  NAND3_X1 U10197 ( .A1(n9072), .A2(n9071), .A3(n9070), .ZN(n9074) );
  NAND2_X1 U10198 ( .A1(n9074), .A2(n9073), .ZN(n9076) );
  AOI21_X1 U10199 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9081) );
  OAI211_X1 U10200 ( .C1(n9081), .C2(n9080), .A(n9079), .B(n9078), .ZN(n9082)
         );
  NAND3_X1 U10201 ( .A1(n9084), .A2(n9083), .A3(n9082), .ZN(n9085) );
  NAND2_X1 U10202 ( .A1(n9086), .A2(n9085), .ZN(n9089) );
  INV_X1 U10203 ( .A(n9087), .ZN(n9088) );
  AOI21_X1 U10204 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9092) );
  OAI21_X1 U10205 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9096) );
  INV_X1 U10206 ( .A(n9094), .ZN(n9095) );
  AOI21_X1 U10207 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9098) );
  NOR2_X1 U10208 ( .A1(n9099), .A2(n9098), .ZN(n9100) );
  NOR2_X1 U10209 ( .A1(n9101), .A2(n9100), .ZN(n9102) );
  NOR2_X1 U10210 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  NOR2_X1 U10211 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  NOR2_X1 U10212 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  NOR2_X1 U10213 ( .A1(n9109), .A2(n9108), .ZN(n9114) );
  INV_X1 U10214 ( .A(n9110), .ZN(n9112) );
  OAI211_X1 U10215 ( .C1(n9114), .C2(n9113), .A(n9112), .B(n9111), .ZN(n9115)
         );
  INV_X1 U10216 ( .A(n9115), .ZN(n9116) );
  OR2_X1 U10217 ( .A1(n9117), .A2(n9116), .ZN(n9119) );
  NAND2_X1 U10218 ( .A1(n9119), .A2(n9118), .ZN(n9123) );
  NAND3_X1 U10219 ( .A1(n9123), .A2(n10464), .A3(n9120), .ZN(n9122) );
  INV_X1 U10220 ( .A(n9126), .ZN(n9121) );
  OAI211_X1 U10221 ( .C1(n9123), .C2(n6420), .A(n9122), .B(n9121), .ZN(n9129)
         );
  NOR2_X1 U10222 ( .A1(n9125), .A2(n9124), .ZN(n9128) );
  OAI21_X1 U10223 ( .B1(n9126), .B2(n6419), .A(P1_B_REG_SCAN_IN), .ZN(n9127)
         );
  INV_X1 U10224 ( .A(n9131), .ZN(n9133) );
  XNOR2_X1 U10225 ( .A(n9190), .B(n7528), .ZN(n9320) );
  NAND2_X1 U10226 ( .A1(n9320), .A2(n9688), .ZN(n9136) );
  NOR2_X1 U10227 ( .A1(n9320), .A2(n9688), .ZN(n9135) );
  AOI21_X2 U10228 ( .B1(n9319), .B2(n9136), .A(n9135), .ZN(n9234) );
  XNOR2_X1 U10229 ( .A(n9232), .B(n7528), .ZN(n9137) );
  XNOR2_X1 U10230 ( .A(n9137), .B(n9669), .ZN(n9233) );
  XNOR2_X1 U10231 ( .A(n9768), .B(n7528), .ZN(n9138) );
  XNOR2_X1 U10232 ( .A(n9138), .B(n9774), .ZN(n9366) );
  NOR2_X1 U10233 ( .A1(n9137), .A2(n9382), .ZN(n9367) );
  NAND2_X1 U10234 ( .A1(n9235), .A2(n5754), .ZN(n9369) );
  INV_X1 U10235 ( .A(n9138), .ZN(n9139) );
  NAND2_X1 U10236 ( .A1(n9139), .A2(n9694), .ZN(n9140) );
  NAND2_X1 U10237 ( .A1(n9369), .A2(n9140), .ZN(n9282) );
  XNOR2_X1 U10238 ( .A(n9661), .B(n7528), .ZN(n9141) );
  XNOR2_X1 U10239 ( .A(n9141), .B(n9767), .ZN(n9283) );
  NAND2_X1 U10240 ( .A1(n9141), .A2(n9645), .ZN(n9142) );
  XNOR2_X1 U10241 ( .A(n9755), .B(n7528), .ZN(n9144) );
  XNOR2_X1 U10242 ( .A(n9144), .B(n9628), .ZN(n9293) );
  XNOR2_X1 U10243 ( .A(n9748), .B(n7528), .ZN(n9146) );
  XNOR2_X1 U10244 ( .A(n9146), .B(n9757), .ZN(n9342) );
  NOR2_X1 U10245 ( .A1(n9144), .A2(n9628), .ZN(n9343) );
  NOR2_X1 U10246 ( .A1(n9342), .A2(n9343), .ZN(n9145) );
  NAND2_X1 U10247 ( .A1(n9291), .A2(n9145), .ZN(n9345) );
  INV_X1 U10248 ( .A(n9146), .ZN(n9147) );
  NAND2_X1 U10249 ( .A1(n9345), .A2(n9148), .ZN(n9255) );
  XNOR2_X1 U10250 ( .A(n9616), .B(n7528), .ZN(n9254) );
  OR2_X1 U10251 ( .A1(n9254), .A2(n9347), .ZN(n9149) );
  XNOR2_X1 U10252 ( .A(n9740), .B(n9158), .ZN(n9150) );
  NAND2_X1 U10253 ( .A1(n9150), .A2(n9268), .ZN(n9152) );
  OAI21_X1 U10254 ( .B1(n9150), .B2(n9268), .A(n9152), .ZN(n9312) );
  NAND2_X1 U10255 ( .A1(n9310), .A2(n9152), .ZN(n9263) );
  XNOR2_X1 U10256 ( .A(n9736), .B(n7528), .ZN(n9153) );
  XNOR2_X1 U10257 ( .A(n9153), .B(n9337), .ZN(n9264) );
  NAND2_X1 U10258 ( .A1(n9263), .A2(n9264), .ZN(n9262) );
  XNOR2_X1 U10259 ( .A(n9732), .B(n7528), .ZN(n9155) );
  XNOR2_X1 U10260 ( .A(n9155), .B(n9593), .ZN(n9332) );
  NOR2_X1 U10261 ( .A1(n9153), .A2(n9602), .ZN(n9333) );
  NOR2_X1 U10262 ( .A1(n9332), .A2(n9333), .ZN(n9154) );
  XNOR2_X1 U10263 ( .A(n8637), .B(n7528), .ZN(n9243) );
  XNOR2_X1 U10264 ( .A(n9725), .B(n9158), .ZN(n9159) );
  NAND2_X1 U10265 ( .A1(n9159), .A2(n9277), .ZN(n9161) );
  OAI21_X1 U10266 ( .B1(n9159), .B2(n9277), .A(n9161), .ZN(n9301) );
  AOI21_X1 U10267 ( .B1(n9578), .B2(n9243), .A(n9301), .ZN(n9160) );
  NAND2_X1 U10268 ( .A1(n9303), .A2(n9161), .ZN(n9273) );
  XNOR2_X1 U10269 ( .A(n9721), .B(n7528), .ZN(n9163) );
  XNOR2_X1 U10270 ( .A(n9163), .B(n9362), .ZN(n9274) );
  NAND2_X1 U10271 ( .A1(n9273), .A2(n9274), .ZN(n9272) );
  XNOR2_X1 U10272 ( .A(n9717), .B(n7528), .ZN(n9165) );
  XNOR2_X1 U10273 ( .A(n9165), .B(n9538), .ZN(n9353) );
  NOR2_X1 U10274 ( .A1(n9163), .A2(n9549), .ZN(n9354) );
  NOR2_X1 U10275 ( .A1(n9353), .A2(n9354), .ZN(n9164) );
  NAND2_X1 U10276 ( .A1(n9272), .A2(n9164), .ZN(n9356) );
  NAND2_X1 U10277 ( .A1(n9165), .A2(n9538), .ZN(n9166) );
  XNOR2_X1 U10278 ( .A(n9713), .B(n7528), .ZN(n9167) );
  XNOR2_X1 U10279 ( .A(n9167), .B(n9531), .ZN(n9224) );
  XNOR2_X1 U10280 ( .A(n9506), .B(n7528), .ZN(n9168) );
  NOR2_X1 U10281 ( .A1(n9348), .A2(n9502), .ZN(n9171) );
  AOI22_X1 U10282 ( .A1(n9373), .A2(n9716), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n9169) );
  OAI21_X1 U10283 ( .B1(n9505), .B2(n9375), .A(n9169), .ZN(n9170) );
  AOI211_X1 U10284 ( .C1(n9708), .C2(n9327), .A(n9171), .B(n9170), .ZN(n9172)
         );
  INV_X1 U10285 ( .A(n9175), .ZN(n9176) );
  OAI21_X1 U10286 ( .B1(n9177), .B2(n9176), .A(n9926), .ZN(n9181) );
  AOI22_X1 U10287 ( .A1(n10502), .A2(n9917), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9178) );
  OAI21_X1 U10288 ( .B1(n10694), .B2(n9912), .A(n9178), .ZN(n9179) );
  AOI21_X1 U10289 ( .B1(n9938), .B2(n9932), .A(n9179), .ZN(n9180) );
  OAI211_X1 U10290 ( .C1(n5433), .C2(n9936), .A(n9181), .B(n9180), .ZN(
        P1_U3214) );
  INV_X1 U10291 ( .A(n9703), .ZN(n9217) );
  NAND2_X1 U10292 ( .A1(n9183), .A2(n9182), .ZN(n9514) );
  NAND2_X1 U10293 ( .A1(n9514), .A2(n5749), .ZN(n9186) );
  NAND2_X1 U10294 ( .A1(n9186), .A2(n9185), .ZN(n9507) );
  NAND2_X1 U10295 ( .A1(n9507), .A2(n9506), .ZN(n9509) );
  NAND2_X1 U10296 ( .A1(n9509), .A2(n9187), .ZN(n9189) );
  INV_X1 U10297 ( .A(n9204), .ZN(n9211) );
  NAND2_X1 U10298 ( .A1(n9328), .A2(n9383), .ZN(n9192) );
  NAND2_X1 U10299 ( .A1(n9193), .A2(n9192), .ZN(n9686) );
  NAND2_X1 U10300 ( .A1(n9661), .A2(n9645), .ZN(n9195) );
  INV_X1 U10301 ( .A(n9268), .ZN(n9612) );
  NOR2_X1 U10302 ( .A1(n9740), .A2(n9612), .ZN(n9590) );
  INV_X1 U10303 ( .A(n9582), .ZN(n9577) );
  INV_X1 U10304 ( .A(n8637), .ZN(n9572) );
  INV_X1 U10305 ( .A(n9532), .ZN(n9526) );
  XNOR2_X1 U10306 ( .A(n9202), .B(n9201), .ZN(n9209) );
  NAND2_X1 U10307 ( .A1(n9204), .A2(n9203), .ZN(n9207) );
  NAND2_X1 U10308 ( .A1(n7130), .A2(P2_B_REG_SCAN_IN), .ZN(n9205) );
  AND2_X1 U10309 ( .A1(n7160), .A2(n9205), .ZN(n9492) );
  AOI22_X1 U10310 ( .A1(n9381), .A2(n9492), .B1(n7162), .B2(n9517), .ZN(n9206)
         );
  NAND2_X1 U10311 ( .A1(n9207), .A2(n9206), .ZN(n9208) );
  AOI21_X2 U10312 ( .B1(n9209), .B2(n9643), .A(n9208), .ZN(n9706) );
  OAI21_X1 U10313 ( .B1(n9211), .B2(n9210), .A(n9706), .ZN(n9212) );
  NAND2_X1 U10314 ( .A1(n9212), .A2(n9692), .ZN(n9216) );
  OR2_X1 U10315 ( .A1(n11105), .A2(n9213), .ZN(n9214) );
  NAND2_X1 U10316 ( .A1(n9692), .A2(n9214), .ZN(n9494) );
  OAI21_X1 U10317 ( .B1(P2_REG2_REG_29__SCAN_IN), .B2(n11118), .A(n9494), .ZN(
        n9215) );
  OAI211_X1 U10318 ( .C1(n9217), .C2(n9662), .A(n9216), .B(n9215), .ZN(
        P2_U3204) );
  INV_X1 U10319 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10055) );
  OAI222_X1 U10320 ( .A1(n6421), .A2(P1_U3086), .B1(n9222), .B2(n9218), .C1(
        n10055), .C2(n9220), .ZN(P1_U3336) );
  INV_X1 U10321 ( .A(n9219), .ZN(n9805) );
  OAI222_X1 U10322 ( .A1(n9223), .A2(P1_U3086), .B1(n9222), .B2(n9805), .C1(
        n9221), .C2(n9220), .ZN(P1_U3325) );
  XNOR2_X1 U10323 ( .A(n9225), .B(n9224), .ZN(n9231) );
  NOR2_X1 U10324 ( .A1(n9348), .A2(n9521), .ZN(n9229) );
  AOI22_X1 U10325 ( .A1(n9373), .A2(n9538), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9226) );
  OAI21_X1 U10326 ( .B1(n9227), .B2(n9375), .A(n9226), .ZN(n9228) );
  AOI211_X1 U10327 ( .C1(n9713), .C2(n9327), .A(n9229), .B(n9228), .ZN(n9230)
         );
  OAI21_X1 U10328 ( .B1(n9231), .B2(n9330), .A(n9230), .ZN(P2_U3154) );
  INV_X1 U10329 ( .A(n9232), .ZN(n9776) );
  NOR2_X1 U10330 ( .A1(n9234), .A2(n9233), .ZN(n9236) );
  OAI21_X1 U10331 ( .B1(n9236), .B2(n9368), .A(n9370), .ZN(n9242) );
  INV_X1 U10332 ( .A(n9691), .ZN(n9240) );
  NOR2_X1 U10333 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9237), .ZN(n9400) );
  AOI21_X1 U10334 ( .B1(n9373), .B2(n9383), .A(n9400), .ZN(n9238) );
  OAI21_X1 U10335 ( .B1(n9774), .B2(n9375), .A(n9238), .ZN(n9239) );
  AOI21_X1 U10336 ( .B1(n9377), .B2(n9240), .A(n9239), .ZN(n9241) );
  OAI211_X1 U10337 ( .C1(n9776), .C2(n9380), .A(n9242), .B(n9241), .ZN(
        P2_U3155) );
  NOR2_X1 U10338 ( .A1(n9244), .A2(n9243), .ZN(n9299) );
  AOI21_X1 U10339 ( .B1(n9244), .B2(n9243), .A(n9299), .ZN(n9245) );
  NAND2_X1 U10340 ( .A1(n9245), .A2(n9246), .ZN(n9302) );
  OAI21_X1 U10341 ( .B1(n9246), .B2(n9245), .A(n9302), .ZN(n9247) );
  NAND2_X1 U10342 ( .A1(n9247), .A2(n9370), .ZN(n9253) );
  INV_X1 U10343 ( .A(n9248), .ZN(n9570) );
  AOI22_X1 U10344 ( .A1(n9359), .A2(n9561), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9249) );
  OAI21_X1 U10345 ( .B1(n9250), .B2(n9361), .A(n9249), .ZN(n9251) );
  AOI21_X1 U10346 ( .B1(n9377), .B2(n9570), .A(n9251), .ZN(n9252) );
  OAI211_X1 U10347 ( .C1(n9572), .C2(n9380), .A(n9253), .B(n9252), .ZN(
        P2_U3156) );
  XNOR2_X1 U10348 ( .A(n9255), .B(n9254), .ZN(n9261) );
  OAI21_X1 U10349 ( .B1(n9375), .B2(n9268), .A(n9256), .ZN(n9257) );
  AOI21_X1 U10350 ( .B1(n9373), .B2(n9613), .A(n9257), .ZN(n9258) );
  OAI21_X1 U10351 ( .B1(n9348), .B2(n9618), .A(n9258), .ZN(n9259) );
  AOI21_X1 U10352 ( .B1(n9744), .B2(n9327), .A(n9259), .ZN(n9260) );
  OAI21_X1 U10353 ( .B1(n9261), .B2(n9330), .A(n9260), .ZN(P2_U3159) );
  INV_X1 U10354 ( .A(n9736), .ZN(n9598) );
  OAI21_X1 U10355 ( .B1(n9264), .B2(n9263), .A(n9262), .ZN(n9265) );
  NAND2_X1 U10356 ( .A1(n9265), .A2(n9370), .ZN(n9271) );
  INV_X1 U10357 ( .A(n9266), .ZN(n9596) );
  AOI22_X1 U10358 ( .A1(n9359), .A2(n9593), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n9267) );
  OAI21_X1 U10359 ( .B1(n9268), .B2(n9361), .A(n9267), .ZN(n9269) );
  AOI21_X1 U10360 ( .B1(n9377), .B2(n9596), .A(n9269), .ZN(n9270) );
  OAI211_X1 U10361 ( .C1(n9598), .C2(n9380), .A(n9271), .B(n9270), .ZN(
        P2_U3163) );
  OAI21_X1 U10362 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9275) );
  NAND2_X1 U10363 ( .A1(n9275), .A2(n9370), .ZN(n9281) );
  INV_X1 U10364 ( .A(n9540), .ZN(n9279) );
  AOI22_X1 U10365 ( .A1(n9359), .A2(n9538), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9276) );
  OAI21_X1 U10366 ( .B1(n9277), .B2(n9361), .A(n9276), .ZN(n9278) );
  AOI21_X1 U10367 ( .B1(n9377), .B2(n9279), .A(n9278), .ZN(n9280) );
  OAI211_X1 U10368 ( .C1(n9541), .C2(n9380), .A(n9281), .B(n9280), .ZN(
        P2_U3165) );
  XNOR2_X1 U10369 ( .A(n9282), .B(n9283), .ZN(n9290) );
  NOR2_X1 U10370 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9284), .ZN(n9438) );
  NOR2_X1 U10371 ( .A1(n9375), .A2(n9761), .ZN(n9285) );
  AOI211_X1 U10372 ( .C1(n9373), .C2(n9694), .A(n9438), .B(n9285), .ZN(n9286)
         );
  OAI21_X1 U10373 ( .B1(n9348), .B2(n9287), .A(n9286), .ZN(n9288) );
  AOI21_X1 U10374 ( .B1(n9661), .B2(n9327), .A(n9288), .ZN(n9289) );
  OAI21_X1 U10375 ( .B1(n9290), .B2(n9330), .A(n9289), .ZN(P2_U3166) );
  INV_X1 U10376 ( .A(n9291), .ZN(n9344) );
  AOI21_X1 U10377 ( .B1(n9293), .B2(n9292), .A(n9344), .ZN(n9298) );
  NAND2_X1 U10378 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9459) );
  OAI21_X1 U10379 ( .B1(n9375), .B2(n9757), .A(n9459), .ZN(n9294) );
  AOI21_X1 U10380 ( .B1(n9373), .B2(n9645), .A(n9294), .ZN(n9295) );
  OAI21_X1 U10381 ( .B1(n9348), .B2(n9648), .A(n9295), .ZN(n9296) );
  AOI21_X1 U10382 ( .B1(n9755), .B2(n9327), .A(n9296), .ZN(n9297) );
  OAI21_X1 U10383 ( .B1(n9298), .B2(n9330), .A(n9297), .ZN(P2_U3168) );
  INV_X1 U10384 ( .A(n9299), .ZN(n9300) );
  NAND3_X1 U10385 ( .A1(n9302), .A2(n9301), .A3(n9300), .ZN(n9304) );
  AND2_X1 U10386 ( .A1(n9304), .A2(n9303), .ZN(n9309) );
  AOI22_X1 U10387 ( .A1(n9359), .A2(n9549), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9306) );
  NAND2_X1 U10388 ( .A1(n9373), .A2(n9578), .ZN(n9305) );
  OAI211_X1 U10389 ( .C1(n9348), .C2(n9555), .A(n9306), .B(n9305), .ZN(n9307)
         );
  AOI21_X1 U10390 ( .B1(n9725), .B2(n9327), .A(n9307), .ZN(n9308) );
  OAI21_X1 U10391 ( .B1(n9309), .B2(n9330), .A(n9308), .ZN(P2_U3169) );
  INV_X1 U10392 ( .A(n9310), .ZN(n9311) );
  AOI21_X1 U10393 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9318) );
  AOI22_X1 U10394 ( .A1(n9359), .A2(n9602), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9315) );
  NAND2_X1 U10395 ( .A1(n9373), .A2(n9629), .ZN(n9314) );
  OAI211_X1 U10396 ( .C1(n9348), .C2(n9604), .A(n9315), .B(n9314), .ZN(n9316)
         );
  AOI21_X1 U10397 ( .B1(n9740), .B2(n9327), .A(n9316), .ZN(n9317) );
  OAI21_X1 U10398 ( .B1(n9318), .B2(n9330), .A(n9317), .ZN(P2_U3173) );
  XNOR2_X1 U10399 ( .A(n9320), .B(n9383), .ZN(n9321) );
  XNOR2_X1 U10400 ( .A(n9319), .B(n9321), .ZN(n9331) );
  NAND2_X1 U10401 ( .A1(n9377), .A2(n9322), .ZN(n9325) );
  AOI21_X1 U10402 ( .B1(n9373), .B2(n9384), .A(n9323), .ZN(n9324) );
  OAI211_X1 U10403 ( .C1(n9669), .C2(n9375), .A(n9325), .B(n9324), .ZN(n9326)
         );
  AOI21_X1 U10404 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9329) );
  OAI21_X1 U10405 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(P2_U3174) );
  INV_X1 U10406 ( .A(n9262), .ZN(n9334) );
  OAI21_X1 U10407 ( .B1(n9334), .B2(n9333), .A(n9332), .ZN(n9336) );
  NAND3_X1 U10408 ( .A1(n9336), .A2(n9370), .A3(n9335), .ZN(n9341) );
  INV_X1 U10409 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10024) );
  OAI22_X1 U10410 ( .A1(n9361), .A2(n9337), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10024), .ZN(n9339) );
  NOR2_X1 U10411 ( .A1(n9348), .A2(n9584), .ZN(n9338) );
  AOI211_X1 U10412 ( .C1(n9359), .C2(n9578), .A(n9339), .B(n9338), .ZN(n9340)
         );
  OAI211_X1 U10413 ( .C1(n9587), .C2(n9380), .A(n9341), .B(n9340), .ZN(
        P2_U3175) );
  OAI21_X1 U10414 ( .B1(n9344), .B2(n9343), .A(n9342), .ZN(n9346) );
  NAND3_X1 U10415 ( .A1(n9346), .A2(n9370), .A3(n9345), .ZN(n9352) );
  NAND2_X1 U10416 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9478) );
  OAI21_X1 U10417 ( .B1(n9375), .B2(n9347), .A(n9478), .ZN(n9350) );
  NOR2_X1 U10418 ( .A1(n9348), .A2(n9632), .ZN(n9349) );
  AOI211_X1 U10419 ( .C1(n9373), .C2(n9628), .A(n9350), .B(n9349), .ZN(n9351)
         );
  OAI211_X1 U10420 ( .C1(n9748), .C2(n9380), .A(n9352), .B(n9351), .ZN(
        P2_U3178) );
  INV_X1 U10421 ( .A(n9272), .ZN(n9355) );
  OAI21_X1 U10422 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(n9357) );
  NAND3_X1 U10423 ( .A1(n9357), .A2(n9370), .A3(n9356), .ZN(n9365) );
  INV_X1 U10424 ( .A(n9358), .ZN(n9529) );
  AOI22_X1 U10425 ( .A1(n9359), .A2(n9716), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9360) );
  OAI21_X1 U10426 ( .B1(n9362), .B2(n9361), .A(n9360), .ZN(n9363) );
  AOI21_X1 U10427 ( .B1(n9377), .B2(n9529), .A(n9363), .ZN(n9364) );
  OAI211_X1 U10428 ( .C1(n5459), .C2(n9380), .A(n9365), .B(n9364), .ZN(
        P2_U3180) );
  OAI21_X1 U10429 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9371) );
  NAND3_X1 U10430 ( .A1(n9371), .A2(n9370), .A3(n9369), .ZN(n9379) );
  INV_X1 U10431 ( .A(n9372), .ZN(n9675) );
  INV_X1 U10432 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U10433 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10231), .ZN(n9419) );
  AOI21_X1 U10434 ( .B1(n9373), .B2(n9382), .A(n9419), .ZN(n9374) );
  OAI21_X1 U10435 ( .B1(n9767), .B2(n9375), .A(n9374), .ZN(n9376) );
  AOI21_X1 U10436 ( .B1(n9377), .B2(n9675), .A(n9376), .ZN(n9378) );
  OAI211_X1 U10437 ( .C1(n9768), .C2(n9380), .A(n9379), .B(n9378), .ZN(
        P2_U3181) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9493), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10439 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9381), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10440 ( .A(n9505), .ZN(n9707) );
  MUX2_X1 U10441 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9707), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10442 ( .A(n9517), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9483), .Z(
        P2_U3519) );
  MUX2_X1 U10443 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9716), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10444 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9538), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10445 ( .A(n9549), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9483), .Z(
        P2_U3516) );
  MUX2_X1 U10446 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9561), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10447 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9578), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10448 ( .A(n9593), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9483), .Z(
        P2_U3513) );
  MUX2_X1 U10449 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9602), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10450 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9612), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10451 ( .A(n9629), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9483), .Z(
        P2_U3510) );
  MUX2_X1 U10452 ( .A(n9613), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9483), .Z(
        P2_U3509) );
  MUX2_X1 U10453 ( .A(n9628), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9483), .Z(
        P2_U3508) );
  MUX2_X1 U10454 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9645), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10455 ( .A(n9694), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9483), .Z(
        P2_U3506) );
  MUX2_X1 U10456 ( .A(n9382), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9483), .Z(
        P2_U3505) );
  MUX2_X1 U10457 ( .A(n9383), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9483), .Z(
        P2_U3504) );
  MUX2_X1 U10458 ( .A(n9384), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9483), .Z(
        P2_U3503) );
  MUX2_X1 U10459 ( .A(n9385), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9483), .Z(
        P2_U3502) );
  MUX2_X1 U10460 ( .A(n9386), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9483), .Z(
        P2_U3501) );
  MUX2_X1 U10461 ( .A(n9387), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9483), .Z(
        P2_U3500) );
  MUX2_X1 U10462 ( .A(n9388), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9483), .Z(
        P2_U3499) );
  MUX2_X1 U10463 ( .A(n9389), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9483), .Z(
        P2_U3498) );
  MUX2_X1 U10464 ( .A(n9390), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9483), .Z(
        P2_U3497) );
  MUX2_X1 U10465 ( .A(n9391), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9483), .Z(
        P2_U3496) );
  MUX2_X1 U10466 ( .A(n9392), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9483), .Z(
        P2_U3495) );
  MUX2_X1 U10467 ( .A(n9393), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9483), .Z(
        P2_U3494) );
  MUX2_X1 U10468 ( .A(n7305), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9483), .Z(
        P2_U3492) );
  MUX2_X1 U10469 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7164), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U10470 ( .A(n9394), .ZN(n9395) );
  AOI21_X1 U10471 ( .B1(n5224), .B2(n9396), .A(n9395), .ZN(n9412) );
  OAI21_X1 U10472 ( .B1(n9399), .B2(n9398), .A(n9397), .ZN(n9410) );
  INV_X1 U10473 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9403) );
  AOI21_X1 U10474 ( .B1(n11033), .B2(n9401), .A(n9400), .ZN(n9402) );
  OAI21_X1 U10475 ( .B1(n11040), .B2(n9403), .A(n9402), .ZN(n9409) );
  NAND2_X1 U10476 ( .A1(n9405), .A2(n9404), .ZN(n9406) );
  AOI21_X1 U10477 ( .B1(n9407), .B2(n9406), .A(n11090), .ZN(n9408) );
  AOI211_X1 U10478 ( .C1(n11086), .C2(n9410), .A(n9409), .B(n9408), .ZN(n9411)
         );
  OAI21_X1 U10479 ( .B1(n9412), .B2(n11081), .A(n9411), .ZN(P2_U3196) );
  AOI21_X1 U10480 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(n9431) );
  OAI21_X1 U10481 ( .B1(n9418), .B2(n9417), .A(n9416), .ZN(n9429) );
  INV_X1 U10482 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9422) );
  AOI21_X1 U10483 ( .B1(n11033), .B2(n9420), .A(n9419), .ZN(n9421) );
  OAI21_X1 U10484 ( .B1(n11040), .B2(n9422), .A(n9421), .ZN(n9428) );
  AOI21_X1 U10485 ( .B1(n9425), .B2(n9424), .A(n9423), .ZN(n9426) );
  NOR2_X1 U10486 ( .A1(n9426), .A2(n11090), .ZN(n9427) );
  AOI211_X1 U10487 ( .C1(n11086), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9430)
         );
  OAI21_X1 U10488 ( .B1(n9431), .B2(n11081), .A(n9430), .ZN(P2_U3197) );
  AOI21_X1 U10489 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9450) );
  OAI21_X1 U10490 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9448) );
  INV_X1 U10491 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9441) );
  AOI21_X1 U10492 ( .B1(n11033), .B2(n9439), .A(n9438), .ZN(n9440) );
  OAI21_X1 U10493 ( .B1(n11040), .B2(n9441), .A(n9440), .ZN(n9447) );
  AOI21_X1 U10494 ( .B1(n9444), .B2(n9443), .A(n9442), .ZN(n9445) );
  NOR2_X1 U10495 ( .A1(n9445), .A2(n11090), .ZN(n9446) );
  AOI211_X1 U10496 ( .C1(n11086), .C2(n9448), .A(n9447), .B(n9446), .ZN(n9449)
         );
  OAI21_X1 U10497 ( .B1(n9450), .B2(n11081), .A(n9449), .ZN(P2_U3198) );
  AOI21_X1 U10498 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9469) );
  INV_X1 U10499 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9454) );
  NOR2_X1 U10500 ( .A1(n11040), .A2(n9454), .ZN(n9462) );
  AOI21_X1 U10501 ( .B1(n9456), .B2(n9455), .A(n9473), .ZN(n9460) );
  NAND2_X1 U10502 ( .A1(n11033), .A2(n9457), .ZN(n9458) );
  OAI211_X1 U10503 ( .C1(n11081), .C2(n9460), .A(n9459), .B(n9458), .ZN(n9461)
         );
  NOR2_X1 U10504 ( .A1(n9462), .A2(n9461), .ZN(n9468) );
  OAI21_X1 U10505 ( .B1(n9465), .B2(n9464), .A(n9463), .ZN(n9466) );
  NAND2_X1 U10506 ( .A1(n9466), .A2(n11086), .ZN(n9467) );
  OAI211_X1 U10507 ( .C1(n9469), .C2(n11090), .A(n9468), .B(n9467), .ZN(
        P2_U3199) );
  AOI21_X1 U10508 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9491) );
  NOR2_X1 U10509 ( .A1(n5510), .A2(n9473), .ZN(n9476) );
  INV_X1 U10510 ( .A(n9474), .ZN(n9475) );
  XNOR2_X1 U10511 ( .A(n9476), .B(n9475), .ZN(n9477) );
  NAND2_X1 U10512 ( .A1(n9477), .A2(n8377), .ZN(n9479) );
  NAND2_X1 U10513 ( .A1(n9479), .A2(n9478), .ZN(n9490) );
  INV_X1 U10514 ( .A(n9480), .ZN(n9481) );
  NOR2_X1 U10515 ( .A1(n9482), .A2(n9481), .ZN(n9485) );
  INV_X1 U10516 ( .A(n9485), .ZN(n9484) );
  OAI21_X1 U10517 ( .B1(n9484), .B2(n9483), .A(n11096), .ZN(n9488) );
  NOR2_X1 U10518 ( .A1(n9485), .A2(n11020), .ZN(n9487) );
  MUX2_X1 U10519 ( .A(n9488), .B(n9487), .S(n9486), .Z(n9489) );
  NAND2_X1 U10520 ( .A1(n9493), .A2(n9492), .ZN(n9701) );
  INV_X1 U10521 ( .A(n9701), .ZN(n9495) );
  NOR2_X1 U10522 ( .A1(n9495), .A2(n9494), .ZN(n9498) );
  NOR2_X1 U10523 ( .A1(n9692), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9496) );
  OAI22_X1 U10524 ( .A1(n9700), .A2(n9662), .B1(n9498), .B2(n9496), .ZN(
        P2_U3202) );
  NOR2_X1 U10525 ( .A1(n9692), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9497) );
  OAI22_X1 U10526 ( .A1(n9702), .A2(n9662), .B1(n9498), .B2(n9497), .ZN(
        P2_U3203) );
  XNOR2_X1 U10527 ( .A(n9500), .B(n9499), .ZN(n9501) );
  INV_X1 U10528 ( .A(n9502), .ZN(n9503) );
  AOI22_X1 U10529 ( .A1(n11124), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n11118), 
        .B2(n9503), .ZN(n9504) );
  OAI21_X1 U10530 ( .B1(n9505), .B2(n9678), .A(n9504), .ZN(n9511) );
  OR2_X1 U10531 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  NAND2_X1 U10532 ( .A1(n9509), .A2(n9508), .ZN(n9711) );
  NOR2_X1 U10533 ( .A1(n9711), .A2(n9698), .ZN(n9510) );
  AOI211_X1 U10534 ( .C1(n11116), .C2(n9708), .A(n9511), .B(n9510), .ZN(n9512)
         );
  OAI21_X1 U10535 ( .B1(n9710), .B2(n11124), .A(n9512), .ZN(P2_U3205) );
  NAND2_X1 U10536 ( .A1(n9514), .A2(n9513), .ZN(n9515) );
  XNOR2_X1 U10537 ( .A(n9515), .B(n9516), .ZN(n9715) );
  OAI21_X1 U10538 ( .B1(n5185), .B2(n9516), .A(n9643), .ZN(n9520) );
  AOI22_X1 U10539 ( .A1(n9538), .A2(n7162), .B1(n9517), .B2(n7160), .ZN(n9518)
         );
  OAI21_X1 U10540 ( .B1(n9520), .B2(n9519), .A(n9518), .ZN(n9712) );
  NAND2_X1 U10541 ( .A1(n9712), .A2(n9692), .ZN(n9525) );
  OAI22_X1 U10542 ( .A1(n9692), .A2(n9522), .B1(n9521), .B2(n11105), .ZN(n9523) );
  AOI21_X1 U10543 ( .B1(n9713), .B2(n11116), .A(n9523), .ZN(n9524) );
  OAI211_X1 U10544 ( .C1(n9698), .C2(n9715), .A(n9525), .B(n9524), .ZN(
        P2_U3206) );
  XNOR2_X1 U10545 ( .A(n9527), .B(n9526), .ZN(n9528) );
  AOI22_X1 U10546 ( .A1(n9528), .A2(n9643), .B1(n7162), .B2(n9549), .ZN(n9719)
         );
  AOI22_X1 U10547 ( .A1(n11124), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n11118), 
        .B2(n9529), .ZN(n9530) );
  OAI21_X1 U10548 ( .B1(n9531), .B2(n9678), .A(n9530), .ZN(n9534) );
  XNOR2_X1 U10549 ( .A(n9183), .B(n9532), .ZN(n9720) );
  NOR2_X1 U10550 ( .A1(n9720), .A2(n9698), .ZN(n9533) );
  AOI211_X1 U10551 ( .C1(n11116), .C2(n9717), .A(n9534), .B(n9533), .ZN(n9535)
         );
  OAI21_X1 U10552 ( .B1(n9719), .B2(n11124), .A(n9535), .ZN(P2_U3207) );
  XNOR2_X1 U10553 ( .A(n9537), .B(n9536), .ZN(n9539) );
  AOI222_X1 U10554 ( .A1(n9643), .A2(n9539), .B1(n9538), .B2(n7160), .C1(n9561), .C2(n7162), .ZN(n9724) );
  INV_X1 U10555 ( .A(n9724), .ZN(n9543) );
  OAI22_X1 U10556 ( .A1(n9541), .A2(n11103), .B1(n9540), .B2(n11105), .ZN(
        n9542) );
  OAI21_X1 U10557 ( .B1(n9543), .B2(n9542), .A(n9692), .ZN(n9547) );
  OAI21_X1 U10558 ( .B1(n5184), .B2(n9545), .A(n9544), .ZN(n9722) );
  AOI22_X1 U10559 ( .A1(n9722), .A2(n11120), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n11124), .ZN(n9546) );
  NAND2_X1 U10560 ( .A1(n9547), .A2(n9546), .ZN(P2_U3208) );
  INV_X1 U10561 ( .A(n11103), .ZN(n9552) );
  XNOR2_X1 U10562 ( .A(n9548), .B(n9553), .ZN(n9550) );
  AOI222_X1 U10563 ( .A1(n9643), .A2(n9550), .B1(n9549), .B2(n7160), .C1(n9578), .C2(n7162), .ZN(n9728) );
  INV_X1 U10564 ( .A(n9728), .ZN(n9551) );
  AOI21_X1 U10565 ( .B1(n9552), .B2(n9725), .A(n9551), .ZN(n9559) );
  XNOR2_X1 U10566 ( .A(n9554), .B(n9553), .ZN(n9726) );
  OAI22_X1 U10567 ( .A1(n9692), .A2(n9556), .B1(n9555), .B2(n11105), .ZN(n9557) );
  AOI21_X1 U10568 ( .B1(n9726), .B2(n11120), .A(n9557), .ZN(n9558) );
  OAI21_X1 U10569 ( .B1(n9559), .B2(n11124), .A(n9558), .ZN(P2_U3209) );
  XNOR2_X1 U10570 ( .A(n9560), .B(n9569), .ZN(n9562) );
  AOI222_X1 U10571 ( .A1(n9643), .A2(n9562), .B1(n9561), .B2(n7160), .C1(n9593), .C2(n7162), .ZN(n9731) );
  NAND2_X1 U10572 ( .A1(n9563), .A2(n9564), .ZN(n9566) );
  NAND2_X1 U10573 ( .A1(n9566), .A2(n9565), .ZN(n9580) );
  NAND2_X1 U10574 ( .A1(n9581), .A2(n9567), .ZN(n9568) );
  XOR2_X1 U10575 ( .A(n9569), .B(n9568), .Z(n9729) );
  AOI22_X1 U10576 ( .A1(n11124), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n11118), 
        .B2(n9570), .ZN(n9571) );
  OAI21_X1 U10577 ( .B1(n9572), .B2(n9662), .A(n9571), .ZN(n9573) );
  AOI21_X1 U10578 ( .B1(n9729), .B2(n11120), .A(n9573), .ZN(n9574) );
  OAI21_X1 U10579 ( .B1(n9731), .B2(n11124), .A(n9574), .ZN(P2_U3210) );
  OAI21_X1 U10580 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9579) );
  AOI222_X1 U10581 ( .A1(n9643), .A2(n9579), .B1(n9602), .B2(n7162), .C1(n9578), .C2(n7160), .ZN(n9735) );
  INV_X1 U10582 ( .A(n9580), .ZN(n9583) );
  OAI21_X1 U10583 ( .B1(n9583), .B2(n9582), .A(n9581), .ZN(n9733) );
  INV_X1 U10584 ( .A(n9584), .ZN(n9585) );
  AOI22_X1 U10585 ( .A1(n11124), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n11118), 
        .B2(n9585), .ZN(n9586) );
  OAI21_X1 U10586 ( .B1(n9587), .B2(n9662), .A(n9586), .ZN(n9588) );
  AOI21_X1 U10587 ( .B1(n9733), .B2(n11120), .A(n9588), .ZN(n9589) );
  OAI21_X1 U10588 ( .B1(n9735), .B2(n11124), .A(n9589), .ZN(P2_U3211) );
  OR3_X1 U10589 ( .A1(n5199), .A2(n9590), .A3(n9595), .ZN(n9591) );
  NAND2_X1 U10590 ( .A1(n9592), .A2(n9591), .ZN(n9594) );
  AOI222_X1 U10591 ( .A1(n9643), .A2(n9594), .B1(n9593), .B2(n7160), .C1(n9612), .C2(n7162), .ZN(n9739) );
  XNOR2_X1 U10592 ( .A(n9563), .B(n9595), .ZN(n9737) );
  AOI22_X1 U10593 ( .A1(n11124), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n11118), 
        .B2(n9596), .ZN(n9597) );
  OAI21_X1 U10594 ( .B1(n9598), .B2(n9662), .A(n9597), .ZN(n9599) );
  AOI21_X1 U10595 ( .B1(n9737), .B2(n11120), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10596 ( .B1(n9739), .B2(n11124), .A(n9600), .ZN(P2_U3212) );
  INV_X1 U10597 ( .A(n5199), .ZN(n9601) );
  OAI21_X1 U10598 ( .B1(n5178), .B2(n9607), .A(n9601), .ZN(n9603) );
  AOI222_X1 U10599 ( .A1(n9643), .A2(n9603), .B1(n9602), .B2(n7160), .C1(n9629), .C2(n7162), .ZN(n9743) );
  OAI22_X1 U10600 ( .A1(n9692), .A2(n9605), .B1(n9604), .B2(n11105), .ZN(n9606) );
  AOI21_X1 U10601 ( .B1(n9740), .B2(n11116), .A(n9606), .ZN(n9610) );
  XNOR2_X1 U10602 ( .A(n9608), .B(n9607), .ZN(n9741) );
  NAND2_X1 U10603 ( .A1(n9741), .A2(n11120), .ZN(n9609) );
  OAI211_X1 U10604 ( .C1(n9743), .C2(n11124), .A(n9610), .B(n9609), .ZN(
        P2_U3213) );
  XOR2_X1 U10605 ( .A(n9616), .B(n9611), .Z(n9614) );
  AOI222_X1 U10606 ( .A1(n9643), .A2(n9614), .B1(n9613), .B2(n7162), .C1(n9612), .C2(n7160), .ZN(n9747) );
  XNOR2_X1 U10607 ( .A(n9615), .B(n9616), .ZN(n9745) );
  NOR2_X1 U10608 ( .A1(n9617), .A2(n9662), .ZN(n9620) );
  OAI22_X1 U10609 ( .A1(n9692), .A2(n8376), .B1(n9618), .B2(n11105), .ZN(n9619) );
  AOI211_X1 U10610 ( .C1(n9745), .C2(n11120), .A(n9620), .B(n9619), .ZN(n9621)
         );
  OAI21_X1 U10611 ( .B1(n9747), .B2(n11124), .A(n9621), .ZN(P2_U3214) );
  OR2_X1 U10612 ( .A1(n9623), .A2(n9622), .ZN(n9624) );
  NAND2_X1 U10613 ( .A1(n9625), .A2(n9624), .ZN(n9749) );
  XNOR2_X1 U10614 ( .A(n5304), .B(n9626), .ZN(n9627) );
  NAND2_X1 U10615 ( .A1(n9627), .A2(n9643), .ZN(n9631) );
  AOI22_X1 U10616 ( .A1(n7160), .A2(n9629), .B1(n9628), .B2(n7162), .ZN(n9630)
         );
  NAND2_X1 U10617 ( .A1(n9631), .A2(n9630), .ZN(n9751) );
  NAND2_X1 U10618 ( .A1(n9751), .A2(n9692), .ZN(n9637) );
  OAI22_X1 U10619 ( .A1(n9692), .A2(n9633), .B1(n9632), .B2(n11105), .ZN(n9634) );
  AOI21_X1 U10620 ( .B1(n9635), .B2(n11116), .A(n9634), .ZN(n9636) );
  OAI211_X1 U10621 ( .C1(n9749), .C2(n9698), .A(n9637), .B(n9636), .ZN(
        P2_U3215) );
  OR2_X1 U10622 ( .A1(n9638), .A2(n9641), .ZN(n9639) );
  NAND2_X1 U10623 ( .A1(n9640), .A2(n9639), .ZN(n9753) );
  XNOR2_X1 U10624 ( .A(n9642), .B(n9641), .ZN(n9644) );
  NAND2_X1 U10625 ( .A1(n9644), .A2(n9643), .ZN(n9647) );
  NAND2_X1 U10626 ( .A1(n9645), .A2(n7162), .ZN(n9646) );
  NAND2_X1 U10627 ( .A1(n9647), .A2(n9646), .ZN(n9760) );
  NAND2_X1 U10628 ( .A1(n9760), .A2(n9692), .ZN(n9652) );
  NOR2_X1 U10629 ( .A1(n9678), .A2(n9757), .ZN(n9650) );
  OAI22_X1 U10630 ( .A1(n9692), .A2(n9455), .B1(n9648), .B2(n11105), .ZN(n9649) );
  AOI211_X1 U10631 ( .C1(n9755), .C2(n11116), .A(n9650), .B(n9649), .ZN(n9651)
         );
  OAI211_X1 U10632 ( .C1(n9753), .C2(n9698), .A(n9652), .B(n9651), .ZN(
        P2_U3216) );
  XNOR2_X1 U10633 ( .A(n9653), .B(n9660), .ZN(n9654) );
  OAI22_X1 U10634 ( .A1(n9654), .A2(n9689), .B1(n9774), .B2(n9687), .ZN(n9763)
         );
  AOI21_X1 U10635 ( .B1(n9655), .B2(n11118), .A(n9763), .ZN(n9666) );
  NAND2_X1 U10636 ( .A1(n9671), .A2(n9657), .ZN(n9659) );
  AOI21_X1 U10637 ( .B1(n9660), .B2(n9659), .A(n5755), .ZN(n9765) );
  INV_X1 U10638 ( .A(n9661), .ZN(n9762) );
  NOR2_X1 U10639 ( .A1(n9762), .A2(n9662), .ZN(n9664) );
  OAI22_X1 U10640 ( .A1(n9678), .A2(n9761), .B1(n8370), .B2(n9692), .ZN(n9663)
         );
  AOI211_X1 U10641 ( .C1(n9765), .C2(n11120), .A(n9664), .B(n9663), .ZN(n9665)
         );
  OAI21_X1 U10642 ( .B1(n9666), .B2(n11124), .A(n9665), .ZN(P2_U3217) );
  XNOR2_X1 U10643 ( .A(n9668), .B(n9667), .ZN(n9670) );
  OAI22_X1 U10644 ( .A1(n9670), .A2(n9689), .B1(n9669), .B2(n9687), .ZN(n9769)
         );
  INV_X1 U10645 ( .A(n9769), .ZN(n9681) );
  INV_X1 U10646 ( .A(n9656), .ZN(n9673) );
  OAI21_X1 U10647 ( .B1(n9673), .B2(n9672), .A(n9671), .ZN(n9771) );
  NAND2_X1 U10648 ( .A1(n9674), .A2(n11116), .ZN(n9677) );
  AOI22_X1 U10649 ( .A1(n11124), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11118), 
        .B2(n9675), .ZN(n9676) );
  OAI211_X1 U10650 ( .C1(n9767), .C2(n9678), .A(n9677), .B(n9676), .ZN(n9679)
         );
  AOI21_X1 U10651 ( .B1(n9771), .B2(n11120), .A(n9679), .ZN(n9680) );
  OAI21_X1 U10652 ( .B1(n9681), .B2(n11124), .A(n9680), .ZN(P2_U3218) );
  INV_X1 U10653 ( .A(n9682), .ZN(n9683) );
  AOI21_X1 U10654 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9780) );
  INV_X1 U10655 ( .A(n9780), .ZN(n9699) );
  XNOR2_X1 U10656 ( .A(n9686), .B(n9685), .ZN(n9690) );
  OAI22_X1 U10657 ( .A1(n9690), .A2(n9689), .B1(n9688), .B2(n9687), .ZN(n9777)
         );
  OAI22_X1 U10658 ( .A1(n9776), .A2(n11103), .B1(n9691), .B2(n11105), .ZN(
        n9693) );
  OAI21_X1 U10659 ( .B1(n9777), .B2(n9693), .A(n9692), .ZN(n9697) );
  AOI22_X1 U10660 ( .A1(n9695), .A2(n9694), .B1(n11124), .B2(
        P2_REG2_REG_14__SCAN_IN), .ZN(n9696) );
  OAI211_X1 U10661 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(
        P2_U3219) );
  OAI21_X1 U10662 ( .B1(n9700), .B2(n9775), .A(n9701), .ZN(n9782) );
  MUX2_X1 U10663 ( .A(n9782), .B(P2_REG1_REG_31__SCAN_IN), .S(n5132), .Z(
        P2_U3490) );
  OAI21_X1 U10664 ( .B1(n9702), .B2(n9775), .A(n9701), .ZN(n9783) );
  MUX2_X1 U10665 ( .A(n9783), .B(P2_REG1_REG_30__SCAN_IN), .S(n5132), .Z(
        P2_U3489) );
  AOI22_X1 U10666 ( .A1(n9204), .A2(n9704), .B1(n9754), .B2(n9703), .ZN(n9705)
         );
  NAND2_X1 U10667 ( .A1(n9706), .A2(n9705), .ZN(n9784) );
  MUX2_X1 U10668 ( .A(n9784), .B(P2_REG1_REG_29__SCAN_IN), .S(n5132), .Z(
        P2_U3488) );
  AOI22_X1 U10669 ( .A1(n9708), .A2(n9754), .B1(n7160), .B2(n9707), .ZN(n9709)
         );
  OAI211_X1 U10670 ( .C1(n9752), .C2(n9711), .A(n9710), .B(n9709), .ZN(n9785)
         );
  MUX2_X1 U10671 ( .A(n9785), .B(P2_REG1_REG_28__SCAN_IN), .S(n5132), .Z(
        P2_U3487) );
  AOI21_X1 U10672 ( .B1(n9754), .B2(n9713), .A(n9712), .ZN(n9714) );
  OAI21_X1 U10673 ( .B1(n9752), .B2(n9715), .A(n9714), .ZN(n9786) );
  MUX2_X1 U10674 ( .A(n9786), .B(P2_REG1_REG_27__SCAN_IN), .S(n5132), .Z(
        P2_U3486) );
  AOI22_X1 U10675 ( .A1(n9717), .A2(n9754), .B1(n7160), .B2(n9716), .ZN(n9718)
         );
  OAI211_X1 U10676 ( .C1(n9752), .C2(n9720), .A(n9719), .B(n9718), .ZN(n9787)
         );
  MUX2_X1 U10677 ( .A(n9787), .B(P2_REG1_REG_26__SCAN_IN), .S(n5132), .Z(
        P2_U3485) );
  AOI22_X1 U10678 ( .A1(n9722), .A2(n9779), .B1(n9754), .B2(n9721), .ZN(n9723)
         );
  NAND2_X1 U10679 ( .A1(n9724), .A2(n9723), .ZN(n9788) );
  MUX2_X1 U10680 ( .A(n9788), .B(P2_REG1_REG_25__SCAN_IN), .S(n5132), .Z(
        P2_U3484) );
  AOI22_X1 U10681 ( .A1(n9726), .A2(n9779), .B1(n9754), .B2(n9725), .ZN(n9727)
         );
  NAND2_X1 U10682 ( .A1(n9728), .A2(n9727), .ZN(n9789) );
  MUX2_X1 U10683 ( .A(n9789), .B(P2_REG1_REG_24__SCAN_IN), .S(n5132), .Z(
        P2_U3483) );
  AOI22_X1 U10684 ( .A1(n9729), .A2(n9779), .B1(n9754), .B2(n8637), .ZN(n9730)
         );
  NAND2_X1 U10685 ( .A1(n9731), .A2(n9730), .ZN(n9790) );
  MUX2_X1 U10686 ( .A(n9790), .B(P2_REG1_REG_23__SCAN_IN), .S(n5132), .Z(
        P2_U3482) );
  AOI22_X1 U10687 ( .A1(n9733), .A2(n9779), .B1(n9754), .B2(n9732), .ZN(n9734)
         );
  NAND2_X1 U10688 ( .A1(n9735), .A2(n9734), .ZN(n9791) );
  MUX2_X1 U10689 ( .A(n9791), .B(P2_REG1_REG_22__SCAN_IN), .S(n5132), .Z(
        P2_U3481) );
  AOI22_X1 U10690 ( .A1(n9737), .A2(n9779), .B1(n9754), .B2(n9736), .ZN(n9738)
         );
  NAND2_X1 U10691 ( .A1(n9739), .A2(n9738), .ZN(n9792) );
  MUX2_X1 U10692 ( .A(n9792), .B(P2_REG1_REG_21__SCAN_IN), .S(n5132), .Z(
        P2_U3480) );
  AOI22_X1 U10693 ( .A1(n9741), .A2(n9779), .B1(n9754), .B2(n9740), .ZN(n9742)
         );
  NAND2_X1 U10694 ( .A1(n9743), .A2(n9742), .ZN(n9793) );
  MUX2_X1 U10695 ( .A(n9793), .B(P2_REG1_REG_20__SCAN_IN), .S(n5132), .Z(
        P2_U3479) );
  AOI22_X1 U10696 ( .A1(n9745), .A2(n9779), .B1(n9754), .B2(n9744), .ZN(n9746)
         );
  NAND2_X1 U10697 ( .A1(n9747), .A2(n9746), .ZN(n9794) );
  MUX2_X1 U10698 ( .A(n9794), .B(P2_REG1_REG_19__SCAN_IN), .S(n5132), .Z(
        P2_U3478) );
  OAI22_X1 U10699 ( .A1(n9749), .A2(n9752), .B1(n9748), .B2(n9775), .ZN(n9750)
         );
  MUX2_X1 U10700 ( .A(n9795), .B(P2_REG1_REG_18__SCAN_IN), .S(n5132), .Z(
        P2_U3477) );
  NOR2_X1 U10701 ( .A1(n9753), .A2(n9752), .ZN(n9759) );
  NAND2_X1 U10702 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  OAI21_X1 U10703 ( .B1(n9757), .B2(n9773), .A(n9756), .ZN(n9758) );
  MUX2_X1 U10704 ( .A(n9796), .B(P2_REG1_REG_17__SCAN_IN), .S(n5132), .Z(
        P2_U3476) );
  OAI22_X1 U10705 ( .A1(n9762), .A2(n9775), .B1(n9761), .B2(n9773), .ZN(n9764)
         );
  AOI211_X1 U10706 ( .C1(n9765), .C2(n9779), .A(n9764), .B(n9763), .ZN(n11194)
         );
  NAND2_X1 U10707 ( .A1(n5132), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9766) );
  OAI21_X1 U10708 ( .B1(n11194), .B2(n5132), .A(n9766), .ZN(P2_U3475) );
  OAI22_X1 U10709 ( .A1(n9768), .A2(n9775), .B1(n9767), .B2(n9773), .ZN(n9770)
         );
  AOI211_X1 U10710 ( .C1(n9779), .C2(n9771), .A(n9770), .B(n9769), .ZN(n11191)
         );
  NAND2_X1 U10711 ( .A1(n5132), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9772) );
  OAI21_X1 U10712 ( .B1(n11191), .B2(n5132), .A(n9772), .ZN(P2_U3474) );
  OAI22_X1 U10713 ( .A1(n9776), .A2(n9775), .B1(n9774), .B2(n9773), .ZN(n9778)
         );
  AOI211_X1 U10714 ( .C1(n9780), .C2(n9779), .A(n9778), .B(n9777), .ZN(n11189)
         );
  NAND2_X1 U10715 ( .A1(n5132), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9781) );
  OAI21_X1 U10716 ( .B1(n11189), .B2(n5132), .A(n9781), .ZN(P2_U3473) );
  MUX2_X1 U10717 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9782), .S(n11195), .Z(
        P2_U3458) );
  MUX2_X1 U10718 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9783), .S(n11195), .Z(
        P2_U3457) );
  MUX2_X1 U10719 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9784), .S(n11195), .Z(
        P2_U3456) );
  MUX2_X1 U10720 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9785), .S(n11195), .Z(
        P2_U3455) );
  MUX2_X1 U10721 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9786), .S(n11195), .Z(
        P2_U3454) );
  MUX2_X1 U10722 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9787), .S(n11195), .Z(
        P2_U3453) );
  MUX2_X1 U10723 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9788), .S(n11195), .Z(
        P2_U3452) );
  MUX2_X1 U10724 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9789), .S(n11195), .Z(
        P2_U3451) );
  MUX2_X1 U10725 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9790), .S(n11195), .Z(
        P2_U3450) );
  MUX2_X1 U10726 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9791), .S(n11195), .Z(
        P2_U3449) );
  MUX2_X1 U10727 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9792), .S(n11195), .Z(
        P2_U3448) );
  MUX2_X1 U10728 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9793), .S(n11195), .Z(
        P2_U3447) );
  MUX2_X1 U10729 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9794), .S(n11195), .Z(
        P2_U3446) );
  MUX2_X1 U10730 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9795), .S(n11195), .Z(
        P2_U3444) );
  MUX2_X1 U10731 ( .A(n9796), .B(P2_REG0_REG_17__SCAN_IN), .S(n11192), .Z(
        P2_U3441) );
  INV_X1 U10732 ( .A(n10821), .ZN(n9801) );
  NOR4_X1 U10733 ( .A1(n9797), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n7131), .ZN(n9798) );
  AOI21_X1 U10734 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9802), .A(n9798), .ZN(
        n9799) );
  OAI21_X1 U10735 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(P2_U3264) );
  AOI22_X1 U10736 ( .A1(n7097), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9802), .ZN(n9803) );
  OAI21_X1 U10737 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(P2_U3265) );
  INV_X1 U10738 ( .A(n9806), .ZN(n9807) );
  MUX2_X1 U10739 ( .A(n9807), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10740 ( .B1(n9809), .B2(n9900), .A(n9808), .ZN(n9810) );
  NAND2_X1 U10741 ( .A1(n9810), .A2(n9926), .ZN(n9816) );
  NOR2_X1 U10742 ( .A1(n10567), .A2(n9930), .ZN(n9814) );
  OAI22_X1 U10743 ( .A1(n9812), .A2(n9912), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9811), .ZN(n9813) );
  AOI211_X1 U10744 ( .C1(n9932), .C2(n10710), .A(n9814), .B(n9813), .ZN(n9815)
         );
  OAI211_X1 U10745 ( .C1(n10793), .C2(n9936), .A(n9816), .B(n9815), .ZN(
        P1_U3216) );
  XOR2_X1 U10746 ( .A(n9817), .B(n9884), .Z(n9822) );
  NAND2_X1 U10747 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10465)
         );
  OAI21_X1 U10748 ( .B1(n10645), .B2(n9878), .A(n10465), .ZN(n9818) );
  AOI21_X1 U10749 ( .B1(n9928), .B2(n10344), .A(n9818), .ZN(n9819) );
  OAI21_X1 U10750 ( .B1(n10660), .B2(n9930), .A(n9819), .ZN(n9820) );
  AOI21_X1 U10751 ( .B1(n10657), .B2(n9904), .A(n9820), .ZN(n9821) );
  OAI21_X1 U10752 ( .B1(n9822), .B2(n9919), .A(n9821), .ZN(P1_U3219) );
  NAND2_X1 U10753 ( .A1(n10709), .A2(n9932), .ZN(n9824) );
  AOI22_X1 U10754 ( .A1(n10616), .A2(n9928), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9823) );
  OAI211_X1 U10755 ( .C1(n9930), .C2(n10609), .A(n9824), .B(n9823), .ZN(n9832)
         );
  NAND2_X1 U10756 ( .A1(n9826), .A2(n9825), .ZN(n9830) );
  INV_X1 U10757 ( .A(n9827), .ZN(n9828) );
  AOI211_X1 U10758 ( .C1(n9830), .C2(n9829), .A(n9919), .B(n9828), .ZN(n9831)
         );
  AOI211_X1 U10759 ( .C1(n10725), .C2(n9904), .A(n9832), .B(n9831), .ZN(n9833)
         );
  INV_X1 U10760 ( .A(n9833), .ZN(P1_U3223) );
  AOI21_X1 U10761 ( .B1(n9835), .B2(n9834), .A(n9924), .ZN(n9840) );
  NAND2_X1 U10762 ( .A1(n10503), .A2(n9932), .ZN(n9837) );
  AOI22_X1 U10763 ( .A1(n10710), .A2(n9928), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9836) );
  OAI211_X1 U10764 ( .C1(n9930), .C2(n10540), .A(n9837), .B(n9836), .ZN(n9838)
         );
  AOI21_X1 U10765 ( .B1(n10538), .B2(n9904), .A(n9838), .ZN(n9839) );
  OAI21_X1 U10766 ( .B1(n9840), .B2(n9919), .A(n9839), .ZN(P1_U3225) );
  INV_X1 U10767 ( .A(n9841), .ZN(n9842) );
  AOI21_X1 U10768 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(n9851) );
  NAND2_X1 U10769 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10409)
         );
  NAND2_X1 U10770 ( .A1(n9928), .A2(n10346), .ZN(n9845) );
  OAI211_X1 U10771 ( .C1(n9878), .C2(n10740), .A(n10409), .B(n9845), .ZN(n9848) );
  NOR2_X1 U10772 ( .A1(n9846), .A2(n9936), .ZN(n9847) );
  AOI211_X1 U10773 ( .C1(n9917), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9850)
         );
  OAI21_X1 U10774 ( .B1(n9851), .B2(n9919), .A(n9850), .ZN(P1_U3226) );
  OAI21_X1 U10775 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  NAND2_X1 U10776 ( .A1(n9855), .A2(n9926), .ZN(n9861) );
  NAND2_X1 U10777 ( .A1(n10344), .A2(n9932), .ZN(n9856) );
  NAND2_X1 U10778 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10446)
         );
  OAI211_X1 U10779 ( .C1(n9857), .C2(n9912), .A(n9856), .B(n10446), .ZN(n9858)
         );
  AOI21_X1 U10780 ( .B1(n9859), .B2(n9917), .A(n9858), .ZN(n9860) );
  OAI211_X1 U10781 ( .C1(n9862), .C2(n9936), .A(n9861), .B(n9860), .ZN(
        P1_U3228) );
  NAND2_X1 U10782 ( .A1(n5221), .A2(n9863), .ZN(n9864) );
  XNOR2_X1 U10783 ( .A(n9865), .B(n9864), .ZN(n9873) );
  INV_X1 U10784 ( .A(n10555), .ZN(n9870) );
  NAND2_X1 U10785 ( .A1(n10520), .A2(n9932), .ZN(n9869) );
  NOR2_X1 U10786 ( .A1(n9866), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9867) );
  AOI21_X1 U10787 ( .B1(n10590), .B2(n9928), .A(n9867), .ZN(n9868) );
  OAI211_X1 U10788 ( .C1(n9930), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9871)
         );
  AOI21_X1 U10789 ( .B1(n10556), .B2(n9904), .A(n9871), .ZN(n9872) );
  OAI21_X1 U10790 ( .B1(n9873), .B2(n9919), .A(n9872), .ZN(P1_U3229) );
  OAI211_X1 U10791 ( .C1(n9876), .C2(n9875), .A(n9874), .B(n9926), .ZN(n9883)
         );
  AOI22_X1 U10792 ( .A1(n9904), .A2(n5979), .B1(n10356), .B2(n9928), .ZN(n9882) );
  AND2_X1 U10793 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10376) );
  NOR2_X1 U10794 ( .A1(n9878), .A2(n9877), .ZN(n9879) );
  AOI211_X1 U10795 ( .C1(n9917), .C2(n9880), .A(n10376), .B(n9879), .ZN(n9881)
         );
  NAND3_X1 U10796 ( .A1(n9883), .A2(n9882), .A3(n9881), .ZN(P1_U3230) );
  NAND2_X1 U10797 ( .A1(n9817), .A2(n9884), .ZN(n9886) );
  NAND2_X1 U10798 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  XOR2_X1 U10799 ( .A(n9888), .B(n9887), .Z(n9893) );
  AOI22_X1 U10800 ( .A1(n10589), .A2(n9932), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9890) );
  NAND2_X1 U10801 ( .A1(n9917), .A2(n10633), .ZN(n9889) );
  OAI211_X1 U10802 ( .C1(n10742), .C2(n9912), .A(n9890), .B(n9889), .ZN(n9891)
         );
  AOI21_X1 U10803 ( .B1(n10631), .B2(n9904), .A(n9891), .ZN(n9892) );
  OAI21_X1 U10804 ( .B1(n9893), .B2(n9919), .A(n9892), .ZN(P1_U3233) );
  INV_X1 U10805 ( .A(n9894), .ZN(n9899) );
  AOI21_X1 U10806 ( .B1(n9897), .B2(n5332), .A(n9896), .ZN(n9898) );
  AOI21_X1 U10807 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9906) );
  AOI22_X1 U10808 ( .A1(n10589), .A2(n9928), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9902) );
  NAND2_X1 U10809 ( .A1(n10590), .A2(n9932), .ZN(n9901) );
  OAI211_X1 U10810 ( .C1(n9930), .C2(n10596), .A(n9902), .B(n9901), .ZN(n9903)
         );
  AOI21_X1 U10811 ( .B1(n10595), .B2(n9904), .A(n9903), .ZN(n9905) );
  OAI21_X1 U10812 ( .B1(n9906), .B2(n9919), .A(n9905), .ZN(P1_U3235) );
  XNOR2_X1 U10813 ( .A(n9908), .B(n9907), .ZN(n9909) );
  XNOR2_X1 U10814 ( .A(n9910), .B(n9909), .ZN(n9920) );
  NAND2_X1 U10815 ( .A1(n10343), .A2(n9932), .ZN(n9911) );
  NAND2_X1 U10816 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10935)
         );
  OAI211_X1 U10817 ( .C1(n10740), .C2(n9912), .A(n9911), .B(n10935), .ZN(n9915) );
  NOR2_X1 U10818 ( .A1(n9913), .A2(n9936), .ZN(n9914) );
  AOI211_X1 U10819 ( .C1(n9917), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9918)
         );
  OAI21_X1 U10820 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(P1_U3238) );
  OAI21_X1 U10821 ( .B1(n9924), .B2(n9923), .A(n9922), .ZN(n9925) );
  NAND3_X1 U10822 ( .A1(n5337), .A2(n9926), .A3(n9925), .ZN(n9935) );
  AOI22_X1 U10823 ( .A1(n10520), .A2(n9928), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9929) );
  OAI21_X1 U10824 ( .B1(n10518), .B2(n9930), .A(n9929), .ZN(n9931) );
  AOI21_X1 U10825 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(n9934) );
  OAI211_X1 U10826 ( .C1(n10517), .C2(n9936), .A(n9935), .B(n9934), .ZN(
        P1_U3240) );
  MUX2_X1 U10827 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10475), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10828 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9937), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10829 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9938), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10830 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10503), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10831 ( .A(n10520), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10357), .Z(
        P1_U3579) );
  MUX2_X1 U10832 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10710), .S(P1_U3973), .Z(
        n10342) );
  XNOR2_X1 U10833 ( .A(n9939), .B(keyinput_129), .ZN(n9943) );
  XOR2_X1 U10834 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n9942) );
  XNOR2_X1 U10835 ( .A(SI_29_), .B(keyinput_131), .ZN(n9941) );
  XOR2_X1 U10836 ( .A(SI_30_), .B(keyinput_130), .Z(n9940) );
  AOI211_X1 U10837 ( .C1(n9943), .C2(n9942), .A(n9941), .B(n9940), .ZN(n9946)
         );
  XNOR2_X1 U10838 ( .A(SI_28_), .B(keyinput_132), .ZN(n9945) );
  XNOR2_X1 U10839 ( .A(SI_27_), .B(keyinput_133), .ZN(n9944) );
  NOR3_X1 U10840 ( .A1(n9946), .A2(n9945), .A3(n9944), .ZN(n9952) );
  XNOR2_X1 U10841 ( .A(n10141), .B(keyinput_134), .ZN(n9951) );
  XNOR2_X1 U10842 ( .A(SI_25_), .B(keyinput_135), .ZN(n9949) );
  XNOR2_X1 U10843 ( .A(SI_24_), .B(keyinput_136), .ZN(n9948) );
  XNOR2_X1 U10844 ( .A(SI_23_), .B(keyinput_137), .ZN(n9947) );
  NOR3_X1 U10845 ( .A1(n9949), .A2(n9948), .A3(n9947), .ZN(n9950) );
  OAI21_X1 U10846 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(n9955) );
  XNOR2_X1 U10847 ( .A(SI_22_), .B(keyinput_138), .ZN(n9954) );
  XNOR2_X1 U10848 ( .A(SI_21_), .B(keyinput_139), .ZN(n9953) );
  AOI21_X1 U10849 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9960) );
  XNOR2_X1 U10850 ( .A(n9956), .B(keyinput_140), .ZN(n9959) );
  XOR2_X1 U10851 ( .A(SI_18_), .B(keyinput_142), .Z(n9958) );
  XNOR2_X1 U10852 ( .A(SI_19_), .B(keyinput_141), .ZN(n9957) );
  OAI211_X1 U10853 ( .C1(n9960), .C2(n9959), .A(n9958), .B(n9957), .ZN(n9963)
         );
  XNOR2_X1 U10854 ( .A(n10159), .B(keyinput_143), .ZN(n9962) );
  XNOR2_X1 U10855 ( .A(SI_16_), .B(keyinput_144), .ZN(n9961) );
  AOI21_X1 U10856 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n9970) );
  XNOR2_X1 U10857 ( .A(SI_15_), .B(keyinput_145), .ZN(n9969) );
  XOR2_X1 U10858 ( .A(SI_13_), .B(keyinput_147), .Z(n9967) );
  XNOR2_X1 U10859 ( .A(SI_11_), .B(keyinput_149), .ZN(n9966) );
  XNOR2_X1 U10860 ( .A(SI_14_), .B(keyinput_146), .ZN(n9965) );
  XNOR2_X1 U10861 ( .A(SI_12_), .B(keyinput_148), .ZN(n9964) );
  NOR4_X1 U10862 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(n9968)
         );
  OAI21_X1 U10863 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9974) );
  XOR2_X1 U10864 ( .A(SI_10_), .B(keyinput_150), .Z(n9973) );
  XNOR2_X1 U10865 ( .A(n10170), .B(keyinput_151), .ZN(n9972) );
  XNOR2_X1 U10866 ( .A(SI_8_), .B(keyinput_152), .ZN(n9971) );
  AOI211_X1 U10867 ( .C1(n9974), .C2(n9973), .A(n9972), .B(n9971), .ZN(n9978)
         );
  XNOR2_X1 U10868 ( .A(SI_7_), .B(keyinput_153), .ZN(n9977) );
  XNOR2_X1 U10869 ( .A(SI_6_), .B(keyinput_154), .ZN(n9976) );
  XNOR2_X1 U10870 ( .A(SI_5_), .B(keyinput_155), .ZN(n9975) );
  OAI211_X1 U10871 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9982)
         );
  XNOR2_X1 U10872 ( .A(SI_4_), .B(keyinput_156), .ZN(n9981) );
  XOR2_X1 U10873 ( .A(SI_3_), .B(keyinput_157), .Z(n9980) );
  XNOR2_X1 U10874 ( .A(SI_2_), .B(keyinput_158), .ZN(n9979) );
  AOI211_X1 U10875 ( .C1(n9982), .C2(n9981), .A(n9980), .B(n9979), .ZN(n9986)
         );
  XNOR2_X1 U10876 ( .A(SI_1_), .B(keyinput_159), .ZN(n9985) );
  XNOR2_X1 U10877 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n9984) );
  XNOR2_X1 U10878 ( .A(SI_0_), .B(keyinput_160), .ZN(n9983) );
  OAI211_X1 U10879 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n9983), .ZN(n9989)
         );
  XNOR2_X1 U10880 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n9988) );
  XNOR2_X1 U10881 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n9987)
         );
  AOI21_X1 U10882 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(n9993) );
  XNOR2_X1 U10883 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n9992)
         );
  XOR2_X1 U10884 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n9991) );
  XNOR2_X1 U10885 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n9990)
         );
  OAI211_X1 U10886 ( .C1(n9993), .C2(n9992), .A(n9991), .B(n9990), .ZN(n9996)
         );
  XOR2_X1 U10887 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n9995) );
  XOR2_X1 U10888 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .Z(n9994) );
  AOI21_X1 U10889 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n10000) );
  XNOR2_X1 U10890 ( .A(n10195), .B(keyinput_169), .ZN(n9999) );
  XNOR2_X1 U10891 ( .A(n10196), .B(keyinput_171), .ZN(n9998) );
  XNOR2_X1 U10892 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n9997)
         );
  NOR4_X1 U10893 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(n10009) );
  XOR2_X1 U10894 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .Z(n10006)
         );
  XOR2_X1 U10895 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n10005) );
  XNOR2_X1 U10896 ( .A(n10001), .B(keyinput_175), .ZN(n10004) );
  XNOR2_X1 U10897 ( .A(n10002), .B(keyinput_173), .ZN(n10003) );
  NAND4_X1 U10898 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        n10008) );
  XNOR2_X1 U10899 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n10007)
         );
  OAI21_X1 U10900 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10021) );
  XOR2_X1 U10901 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n10014) );
  XNOR2_X1 U10902 ( .A(n10210), .B(keyinput_177), .ZN(n10013) );
  XNOR2_X1 U10903 ( .A(n10010), .B(keyinput_179), .ZN(n10012) );
  XNOR2_X1 U10904 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n10011)
         );
  NOR4_X1 U10905 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10020) );
  XOR2_X1 U10906 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n10018) );
  XOR2_X1 U10907 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .Z(n10017)
         );
  XNOR2_X1 U10908 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n10016)
         );
  XNOR2_X1 U10909 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n10015)
         );
  NAND4_X1 U10910 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n10019) );
  AOI21_X1 U10911 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10029) );
  AOI22_X1 U10912 ( .A1(n10223), .A2(keyinput_186), .B1(keyinput_187), .B2(
        n11106), .ZN(n10022) );
  OAI221_X1 U10913 ( .B1(n10223), .B2(keyinput_186), .C1(n11106), .C2(
        keyinput_187), .A(n10022), .ZN(n10028) );
  INV_X1 U10914 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10025) );
  AOI22_X1 U10915 ( .A1(n10025), .A2(keyinput_188), .B1(n10024), .B2(
        keyinput_185), .ZN(n10023) );
  OAI221_X1 U10916 ( .B1(n10025), .B2(keyinput_188), .C1(n10024), .C2(
        keyinput_185), .A(n10023), .ZN(n10027) );
  XNOR2_X1 U10917 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n10026)
         );
  NOR4_X1 U10918 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10033) );
  XNOR2_X1 U10919 ( .A(n10231), .B(keyinput_191), .ZN(n10032) );
  XNOR2_X1 U10920 ( .A(n10232), .B(keyinput_190), .ZN(n10031) );
  XNOR2_X1 U10921 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n10030) );
  NOR4_X1 U10922 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n10037) );
  XNOR2_X1 U10923 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n10036) );
  XOR2_X1 U10924 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n10035)
         );
  XOR2_X1 U10925 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .Z(n10034)
         );
  OAI211_X1 U10926 ( .C1(n10037), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10047) );
  XOR2_X1 U10927 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .Z(n10046)
         );
  XOR2_X1 U10928 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n10041)
         );
  XOR2_X1 U10929 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .Z(n10040)
         );
  XNOR2_X1 U10930 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n10039) );
  XNOR2_X1 U10931 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n10038) );
  NOR4_X1 U10932 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10044) );
  XOR2_X1 U10933 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .Z(n10043)
         );
  XOR2_X1 U10934 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .Z(n10042)
         );
  NAND3_X1 U10935 ( .A1(n10044), .A2(n10043), .A3(n10042), .ZN(n10045) );
  AOI21_X1 U10936 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(n10049) );
  XOR2_X1 U10937 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n10048)
         );
  NOR2_X1 U10938 ( .A1(n10049), .A2(n10048), .ZN(n10059) );
  AOI22_X1 U10939 ( .A1(n10052), .A2(keyinput_207), .B1(n10051), .B2(
        keyinput_206), .ZN(n10050) );
  OAI221_X1 U10940 ( .B1(n10052), .B2(keyinput_207), .C1(n10051), .C2(
        keyinput_206), .A(n10050), .ZN(n10058) );
  AOI22_X1 U10941 ( .A1(n10055), .A2(keyinput_205), .B1(n10054), .B2(
        keyinput_204), .ZN(n10053) );
  OAI221_X1 U10942 ( .B1(n10055), .B2(keyinput_205), .C1(n10054), .C2(
        keyinput_204), .A(n10053), .ZN(n10057) );
  XNOR2_X1 U10943 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n10056) );
  NOR4_X1 U10944 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10066) );
  XNOR2_X1 U10945 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n10065) );
  XOR2_X1 U10946 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n10063)
         );
  XOR2_X1 U10947 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .Z(n10062)
         );
  XOR2_X1 U10948 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n10061)
         );
  XOR2_X1 U10949 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .Z(n10060)
         );
  NOR4_X1 U10950 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10064) );
  OAI21_X1 U10951 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(n10069) );
  XOR2_X1 U10952 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .Z(n10068)
         );
  XNOR2_X1 U10953 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n10067)
         );
  AOI21_X1 U10954 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10072) );
  XOR2_X1 U10955 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .Z(n10071)
         );
  XNOR2_X1 U10956 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n10070)
         );
  NOR3_X1 U10957 ( .A1(n10072), .A2(n10071), .A3(n10070), .ZN(n10075) );
  XNOR2_X1 U10958 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_218), .ZN(n10074) );
  XNOR2_X1 U10959 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .ZN(n10073) );
  NOR3_X1 U10960 ( .A1(n10075), .A2(n10074), .A3(n10073), .ZN(n10078) );
  XNOR2_X1 U10961 ( .A(n10276), .B(keyinput_220), .ZN(n10077) );
  XNOR2_X1 U10962 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n10076) );
  OAI21_X1 U10963 ( .B1(n10078), .B2(n10077), .A(n10076), .ZN(n10082) );
  XNOR2_X1 U10964 ( .A(n10079), .B(keyinput_223), .ZN(n10081) );
  XNOR2_X1 U10965 ( .A(n5971), .B(keyinput_222), .ZN(n10080) );
  NAND3_X1 U10966 ( .A1(n10082), .A2(n10081), .A3(n10080), .ZN(n10085) );
  XNOR2_X1 U10967 ( .A(n10284), .B(keyinput_225), .ZN(n10084) );
  XNOR2_X1 U10968 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .ZN(n10083) );
  NAND3_X1 U10969 ( .A1(n10085), .A2(n10084), .A3(n10083), .ZN(n10089) );
  XNOR2_X1 U10970 ( .A(n6058), .B(keyinput_227), .ZN(n10088) );
  XNOR2_X1 U10971 ( .A(n10288), .B(keyinput_226), .ZN(n10087) );
  XNOR2_X1 U10972 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_228), .ZN(n10086)
         );
  NAND4_X1 U10973 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10092) );
  XNOR2_X1 U10974 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .ZN(n10091)
         );
  XNOR2_X1 U10975 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_229), .ZN(n10090)
         );
  NAND3_X1 U10976 ( .A1(n10092), .A2(n10091), .A3(n10090), .ZN(n10095) );
  XNOR2_X1 U10977 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n10094)
         );
  XNOR2_X1 U10978 ( .A(n10296), .B(keyinput_232), .ZN(n10093) );
  AOI21_X1 U10979 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(n10099) );
  XNOR2_X1 U10980 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_233), .ZN(n10098)
         );
  XNOR2_X1 U10981 ( .A(n10096), .B(keyinput_234), .ZN(n10097) );
  OAI21_X1 U10982 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(n10103) );
  XOR2_X1 U10983 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_236), .Z(n10102) );
  XNOR2_X1 U10984 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_235), .ZN(n10101)
         );
  XNOR2_X1 U10985 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_237), .ZN(n10100)
         );
  NAND4_X1 U10986 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10106) );
  XNOR2_X1 U10987 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_238), .ZN(n10105)
         );
  XNOR2_X1 U10988 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_239), .ZN(n10104)
         );
  AOI21_X1 U10989 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(n10109) );
  XNOR2_X1 U10990 ( .A(n10312), .B(keyinput_240), .ZN(n10108) );
  XNOR2_X1 U10991 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_241), .ZN(n10107)
         );
  NOR3_X1 U10992 ( .A1(n10109), .A2(n10108), .A3(n10107), .ZN(n10116) );
  XNOR2_X1 U10993 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_243), .ZN(n10113)
         );
  XNOR2_X1 U10994 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_242), .ZN(n10112)
         );
  XNOR2_X1 U10995 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .ZN(n10111)
         );
  XNOR2_X1 U10996 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_245), .ZN(n10110)
         );
  NAND4_X1 U10997 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10115) );
  XNOR2_X1 U10998 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_246), .ZN(n10114)
         );
  OAI21_X1 U10999 ( .B1(n10116), .B2(n10115), .A(n10114), .ZN(n10119) );
  XNOR2_X1 U11000 ( .A(n10325), .B(keyinput_247), .ZN(n10118) );
  XNOR2_X1 U11001 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .ZN(n10117)
         );
  AOI21_X1 U11002 ( .B1(n10119), .B2(n10118), .A(n10117), .ZN(n10122) );
  XNOR2_X1 U11003 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .ZN(n10121)
         );
  XNOR2_X1 U11004 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .ZN(n10120) );
  OAI21_X1 U11005 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n10125) );
  INV_X1 U11006 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10824) );
  XNOR2_X1 U11007 ( .A(n10824), .B(keyinput_252), .ZN(n10124) );
  XNOR2_X1 U11008 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .ZN(n10123) );
  NAND3_X1 U11009 ( .A1(n10125), .A2(n10124), .A3(n10123), .ZN(n10129) );
  XOR2_X1 U11010 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_253), .Z(n10128) );
  XNOR2_X1 U11011 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_255), .ZN(n10127) );
  XNOR2_X1 U11012 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_254), .ZN(n10126) );
  AOI211_X1 U11013 ( .C1(n10129), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10340) );
  INV_X1 U11014 ( .A(keyinput_38), .ZN(n10130) );
  XNOR2_X1 U11015 ( .A(n10130), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n10132) );
  XNOR2_X1 U11016 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n10131)
         );
  AND2_X1 U11017 ( .A1(n10132), .A2(n10131), .ZN(n10188) );
  INV_X1 U11018 ( .A(n10188), .ZN(n10194) );
  XNOR2_X1 U11019 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n10193)
         );
  XNOR2_X1 U11020 ( .A(SI_31_), .B(keyinput_1), .ZN(n10136) );
  XNOR2_X1 U11021 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n10135) );
  XOR2_X1 U11022 ( .A(SI_30_), .B(keyinput_2), .Z(n10134) );
  XNOR2_X1 U11023 ( .A(SI_29_), .B(keyinput_3), .ZN(n10133) );
  OAI211_X1 U11024 ( .C1(n10136), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10140) );
  XNOR2_X1 U11025 ( .A(n10137), .B(keyinput_4), .ZN(n10139) );
  XNOR2_X1 U11026 ( .A(SI_27_), .B(keyinput_5), .ZN(n10138) );
  NAND3_X1 U11027 ( .A1(n10140), .A2(n10139), .A3(n10138), .ZN(n10149) );
  XNOR2_X1 U11028 ( .A(n10141), .B(keyinput_6), .ZN(n10148) );
  XNOR2_X1 U11029 ( .A(n10142), .B(keyinput_9), .ZN(n10146) );
  XNOR2_X1 U11030 ( .A(n10143), .B(keyinput_8), .ZN(n10145) );
  XNOR2_X1 U11031 ( .A(SI_25_), .B(keyinput_7), .ZN(n10144) );
  NAND3_X1 U11032 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n10147) );
  AOI21_X1 U11033 ( .B1(n10149), .B2(n10148), .A(n10147), .ZN(n10153) );
  XNOR2_X1 U11034 ( .A(n10150), .B(keyinput_10), .ZN(n10152) );
  XOR2_X1 U11035 ( .A(SI_21_), .B(keyinput_11), .Z(n10151) );
  OAI21_X1 U11036 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10158) );
  XNOR2_X1 U11037 ( .A(SI_20_), .B(keyinput_12), .ZN(n10157) );
  XNOR2_X1 U11038 ( .A(n10154), .B(keyinput_13), .ZN(n10156) );
  XNOR2_X1 U11039 ( .A(SI_18_), .B(keyinput_14), .ZN(n10155) );
  AOI211_X1 U11040 ( .C1(n10158), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        n10162) );
  XNOR2_X1 U11041 ( .A(n10159), .B(keyinput_15), .ZN(n10161) );
  XNOR2_X1 U11042 ( .A(SI_16_), .B(keyinput_16), .ZN(n10160) );
  OAI21_X1 U11043 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(n10169) );
  XOR2_X1 U11044 ( .A(SI_15_), .B(keyinput_17), .Z(n10168) );
  XOR2_X1 U11045 ( .A(SI_14_), .B(keyinput_18), .Z(n10166) );
  XOR2_X1 U11046 ( .A(SI_12_), .B(keyinput_20), .Z(n10165) );
  XNOR2_X1 U11047 ( .A(SI_11_), .B(keyinput_21), .ZN(n10164) );
  XNOR2_X1 U11048 ( .A(SI_13_), .B(keyinput_19), .ZN(n10163) );
  NAND4_X1 U11049 ( .A1(n10166), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10167) );
  AOI21_X1 U11050 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(n10174) );
  XOR2_X1 U11051 ( .A(SI_10_), .B(keyinput_22), .Z(n10173) );
  XNOR2_X1 U11052 ( .A(n10170), .B(keyinput_23), .ZN(n10172) );
  XNOR2_X1 U11053 ( .A(SI_8_), .B(keyinput_24), .ZN(n10171) );
  OAI211_X1 U11054 ( .C1(n10174), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10178) );
  XNOR2_X1 U11055 ( .A(SI_7_), .B(keyinput_25), .ZN(n10177) );
  XOR2_X1 U11056 ( .A(SI_5_), .B(keyinput_27), .Z(n10176) );
  XNOR2_X1 U11057 ( .A(SI_6_), .B(keyinput_26), .ZN(n10175) );
  AOI211_X1 U11058 ( .C1(n10178), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10182) );
  XNOR2_X1 U11059 ( .A(SI_4_), .B(keyinput_28), .ZN(n10181) );
  XNOR2_X1 U11060 ( .A(SI_3_), .B(keyinput_29), .ZN(n10180) );
  XNOR2_X1 U11061 ( .A(SI_2_), .B(keyinput_30), .ZN(n10179) );
  OAI211_X1 U11062 ( .C1(n10182), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10186) );
  XOR2_X1 U11063 ( .A(SI_1_), .B(keyinput_31), .Z(n10185) );
  XOR2_X1 U11064 ( .A(SI_0_), .B(keyinput_32), .Z(n10184) );
  XNOR2_X1 U11065 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n10183) );
  AOI211_X1 U11066 ( .C1(n10186), .C2(n10185), .A(n10184), .B(n10183), .ZN(
        n10190) );
  XNOR2_X1 U11067 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n10189) );
  XNOR2_X1 U11068 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n10187)
         );
  OAI211_X1 U11069 ( .C1(n10190), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10192) );
  XNOR2_X1 U11070 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n10191)
         );
  OAI211_X1 U11071 ( .C1(n10194), .C2(n10193), .A(n10192), .B(n10191), .ZN(
        n10202) );
  XNOR2_X1 U11072 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n10201)
         );
  XNOR2_X1 U11073 ( .A(n10195), .B(keyinput_41), .ZN(n10199) );
  XNOR2_X1 U11074 ( .A(n10196), .B(keyinput_43), .ZN(n10198) );
  XNOR2_X1 U11075 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n10197)
         );
  NAND3_X1 U11076 ( .A1(n10199), .A2(n10198), .A3(n10197), .ZN(n10200) );
  AOI21_X1 U11077 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(n10209) );
  XNOR2_X1 U11078 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n10206)
         );
  XNOR2_X1 U11079 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n10205)
         );
  XNOR2_X1 U11080 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n10204)
         );
  XNOR2_X1 U11081 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n10203)
         );
  NAND4_X1 U11082 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10208) );
  XOR2_X1 U11083 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .Z(n10207) );
  OAI21_X1 U11084 ( .B1(n10209), .B2(n10208), .A(n10207), .ZN(n10221) );
  XNOR2_X1 U11085 ( .A(n10210), .B(keyinput_49), .ZN(n10214) );
  XNOR2_X1 U11086 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n10213)
         );
  XNOR2_X1 U11087 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n10212)
         );
  XNOR2_X1 U11088 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n10211)
         );
  NOR4_X1 U11089 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10220) );
  XOR2_X1 U11090 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n10218) );
  XOR2_X1 U11091 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .Z(n10217) );
  XNOR2_X1 U11092 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n10216)
         );
  XNOR2_X1 U11093 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n10215)
         );
  NAND4_X1 U11094 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10219) );
  AOI21_X1 U11095 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(n10230) );
  OAI22_X1 U11096 ( .A1(n10223), .A2(keyinput_58), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(keyinput_61), .ZN(n10222) );
  AOI21_X1 U11097 ( .B1(n10223), .B2(keyinput_58), .A(n10222), .ZN(n10226) );
  XNOR2_X1 U11098 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n10225)
         );
  NAND2_X1 U11099 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_61), .ZN(n10224)
         );
  NAND3_X1 U11100 ( .A1(n10226), .A2(n10225), .A3(n10224), .ZN(n10229) );
  XNOR2_X1 U11101 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n10228)
         );
  XNOR2_X1 U11102 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n10227)
         );
  NOR4_X1 U11103 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10236) );
  XOR2_X1 U11104 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .Z(n10235) );
  XNOR2_X1 U11105 ( .A(n10231), .B(keyinput_63), .ZN(n10234) );
  XNOR2_X1 U11106 ( .A(n10232), .B(keyinput_62), .ZN(n10233) );
  NOR4_X1 U11107 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10240) );
  XOR2_X1 U11108 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n10239)
         );
  XNOR2_X1 U11109 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n10238)
         );
  XNOR2_X1 U11110 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n10237)
         );
  OAI211_X1 U11111 ( .C1(n10240), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10250) );
  XNOR2_X1 U11112 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n10249)
         );
  XOR2_X1 U11113 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n10244)
         );
  XOR2_X1 U11114 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n10243)
         );
  XOR2_X1 U11115 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .Z(n10242)
         );
  XOR2_X1 U11116 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .Z(n10241)
         );
  NOR4_X1 U11117 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10247) );
  XNOR2_X1 U11118 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n10246)
         );
  XNOR2_X1 U11119 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n10245)
         );
  NAND3_X1 U11120 ( .A1(n10247), .A2(n10246), .A3(n10245), .ZN(n10248) );
  AOI21_X1 U11121 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(n10259) );
  XOR2_X1 U11122 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n10258)
         );
  XOR2_X1 U11123 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .Z(n10253)
         );
  XNOR2_X1 U11124 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n10252)
         );
  XNOR2_X1 U11125 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n10251)
         );
  NAND3_X1 U11126 ( .A1(n10253), .A2(n10252), .A3(n10251), .ZN(n10256) );
  XOR2_X1 U11127 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n10255)
         );
  XOR2_X1 U11128 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n10254)
         );
  NOR3_X1 U11129 ( .A1(n10256), .A2(n10255), .A3(n10254), .ZN(n10257) );
  OAI21_X1 U11130 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10266) );
  XNOR2_X1 U11131 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n10265)
         );
  XOR2_X1 U11132 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n10263)
         );
  XOR2_X1 U11133 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n10262)
         );
  XNOR2_X1 U11134 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n10261)
         );
  XNOR2_X1 U11135 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n10260)
         );
  NAND4_X1 U11136 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10264) );
  AOI21_X1 U11137 ( .B1(n10266), .B2(n10265), .A(n10264), .ZN(n10269) );
  XOR2_X1 U11138 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n10268)
         );
  XOR2_X1 U11139 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n10267) );
  OAI21_X1 U11140 ( .B1(n10269), .B2(n10268), .A(n10267), .ZN(n10272) );
  XOR2_X1 U11141 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n10271) );
  XNOR2_X1 U11142 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n10270)
         );
  NAND3_X1 U11143 ( .A1(n10272), .A2(n10271), .A3(n10270), .ZN(n10275) );
  XOR2_X1 U11144 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_90), .Z(n10274) );
  XOR2_X1 U11145 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .Z(n10273) );
  NAND3_X1 U11146 ( .A1(n10275), .A2(n10274), .A3(n10273), .ZN(n10279) );
  XNOR2_X1 U11147 ( .A(n10276), .B(keyinput_92), .ZN(n10278) );
  XNOR2_X1 U11148 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n10277) );
  AOI21_X1 U11149 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(n10282) );
  XNOR2_X1 U11150 ( .A(n5971), .B(keyinput_94), .ZN(n10281) );
  XNOR2_X1 U11151 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n10280) );
  NOR3_X1 U11152 ( .A1(n10282), .A2(n10281), .A3(n10280), .ZN(n10287) );
  XNOR2_X1 U11153 ( .A(n10283), .B(keyinput_96), .ZN(n10286) );
  XNOR2_X1 U11154 ( .A(n10284), .B(keyinput_97), .ZN(n10285) );
  NOR3_X1 U11155 ( .A1(n10287), .A2(n10286), .A3(n10285), .ZN(n10292) );
  XNOR2_X1 U11156 ( .A(n10288), .B(keyinput_98), .ZN(n10291) );
  XNOR2_X1 U11157 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_99), .ZN(n10290) );
  XNOR2_X1 U11158 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_100), .ZN(n10289)
         );
  NOR4_X1 U11159 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10295) );
  XOR2_X1 U11160 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .Z(n10294) );
  XNOR2_X1 U11161 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_101), .ZN(n10293)
         );
  NOR3_X1 U11162 ( .A1(n10295), .A2(n10294), .A3(n10293), .ZN(n10299) );
  XOR2_X1 U11163 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .Z(n10298) );
  XNOR2_X1 U11164 ( .A(n10296), .B(keyinput_104), .ZN(n10297) );
  OAI21_X1 U11165 ( .B1(n10299), .B2(n10298), .A(n10297), .ZN(n10302) );
  XNOR2_X1 U11166 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_105), .ZN(n10301)
         );
  XNOR2_X1 U11167 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .ZN(n10300)
         );
  AOI21_X1 U11168 ( .B1(n10302), .B2(n10301), .A(n10300), .ZN(n10307) );
  XNOR2_X1 U11169 ( .A(n10303), .B(keyinput_109), .ZN(n10306) );
  XNOR2_X1 U11170 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n10305)
         );
  XNOR2_X1 U11171 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_108), .ZN(n10304)
         );
  NOR4_X1 U11172 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10310) );
  XOR2_X1 U11173 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_110), .Z(n10309) );
  XNOR2_X1 U11174 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_111), .ZN(n10308)
         );
  OAI21_X1 U11175 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(n10315) );
  XNOR2_X1 U11176 ( .A(n10311), .B(keyinput_113), .ZN(n10314) );
  XNOR2_X1 U11177 ( .A(n10312), .B(keyinput_112), .ZN(n10313) );
  NAND3_X1 U11178 ( .A1(n10315), .A2(n10314), .A3(n10313), .ZN(n10324) );
  XOR2_X1 U11179 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .Z(n10320) );
  XNOR2_X1 U11180 ( .A(n5838), .B(keyinput_114), .ZN(n10319) );
  XNOR2_X1 U11181 ( .A(n10316), .B(keyinput_117), .ZN(n10318) );
  XNOR2_X1 U11182 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_115), .ZN(n10317)
         );
  NOR4_X1 U11183 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10323) );
  XNOR2_X1 U11184 ( .A(n10321), .B(keyinput_118), .ZN(n10322) );
  AOI21_X1 U11185 ( .B1(n10324), .B2(n10323), .A(n10322), .ZN(n10328) );
  XNOR2_X1 U11186 ( .A(n10325), .B(keyinput_119), .ZN(n10327) );
  XNOR2_X1 U11187 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .ZN(n10326)
         );
  OAI21_X1 U11188 ( .B1(n10328), .B2(n10327), .A(n10326), .ZN(n10331) );
  XOR2_X1 U11189 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .Z(n10330) );
  XNOR2_X1 U11190 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .ZN(n10329) );
  AOI21_X1 U11191 ( .B1(n10331), .B2(n10330), .A(n10329), .ZN(n10334) );
  XNOR2_X1 U11192 ( .A(n10824), .B(keyinput_124), .ZN(n10333) );
  XNOR2_X1 U11193 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .ZN(n10332) );
  NOR3_X1 U11194 ( .A1(n10334), .A2(n10333), .A3(n10332), .ZN(n10338) );
  XNOR2_X1 U11195 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_125), .ZN(n10337) );
  XOR2_X1 U11196 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_127), .Z(n10336) );
  XNOR2_X1 U11197 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_126), .ZN(n10335) );
  OAI211_X1 U11198 ( .C1(n10338), .C2(n10337), .A(n10336), .B(n10335), .ZN(
        n10339) );
  NOR2_X1 U11199 ( .A1(n10340), .A2(n10339), .ZN(n10341) );
  XOR2_X1 U11200 ( .A(n10342), .B(n10341), .Z(P1_U3578) );
  MUX2_X1 U11201 ( .A(n10590), .B(P1_DATAO_REG_23__SCAN_IN), .S(n10357), .Z(
        P1_U3577) );
  MUX2_X1 U11202 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10709), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11203 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10589), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11204 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10616), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11205 ( .A(n10343), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10357), .Z(
        P1_U3573) );
  MUX2_X1 U11206 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10344), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11207 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10345), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11208 ( .A(n10346), .B(P1_DATAO_REG_15__SCAN_IN), .S(n10357), .Z(
        P1_U3569) );
  MUX2_X1 U11209 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10347), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11210 ( .A(n10348), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10357), .Z(
        P1_U3567) );
  MUX2_X1 U11211 ( .A(n11154), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10357), .Z(
        P1_U3566) );
  INV_X1 U11212 ( .A(n10349), .ZN(n10350) );
  MUX2_X1 U11213 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10350), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11214 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n11157), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11215 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10351), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11216 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10352), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11217 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10353), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U11218 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10354), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U11219 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10355), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U11220 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10356), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11221 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5320), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U11222 ( .A(n6434), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10357), .Z(
        P1_U3555) );
  INV_X1 U11223 ( .A(n10358), .ZN(n10362) );
  INV_X1 U11224 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10360) );
  OAI21_X1 U11225 ( .B1(n10967), .B2(n10360), .A(n10359), .ZN(n10361) );
  AOI21_X1 U11226 ( .B1(n10362), .B2(n10962), .A(n10361), .ZN(n10371) );
  OAI211_X1 U11227 ( .C1(n10365), .C2(n10364), .A(n10910), .B(n10363), .ZN(
        n10370) );
  OAI211_X1 U11228 ( .C1(n10368), .C2(n10367), .A(n10916), .B(n10366), .ZN(
        n10369) );
  NAND3_X1 U11229 ( .A1(n10371), .A2(n10370), .A3(n10369), .ZN(P1_U3246) );
  INV_X1 U11230 ( .A(n10372), .ZN(n10386) );
  NOR2_X1 U11231 ( .A1(n10374), .A2(n10373), .ZN(n10375) );
  AOI211_X1 U11232 ( .C1(n10396), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10376), .B(
        n10375), .ZN(n10385) );
  OAI211_X1 U11233 ( .C1(n10379), .C2(n10378), .A(n10916), .B(n10377), .ZN(
        n10384) );
  OAI211_X1 U11234 ( .C1(n10382), .C2(n10381), .A(n10910), .B(n10380), .ZN(
        n10383) );
  NAND4_X1 U11235 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        P1_U3247) );
  OAI21_X1 U11236 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(n10390) );
  NAND2_X1 U11237 ( .A1(n10390), .A2(n10916), .ZN(n10401) );
  OAI21_X1 U11238 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(n10394) );
  NAND2_X1 U11239 ( .A1(n10394), .A2(n10910), .ZN(n10400) );
  AOI21_X1 U11240 ( .B1(n10396), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10395), .ZN(
        n10399) );
  NAND2_X1 U11241 ( .A1(n10962), .A2(n10397), .ZN(n10398) );
  NAND4_X1 U11242 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        P1_U3252) );
  XOR2_X1 U11243 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10441), .Z(n10438) );
  OR2_X1 U11244 ( .A1(n10412), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U11245 ( .A1(n10403), .A2(n10402), .ZN(n10944) );
  XNOR2_X1 U11246 ( .A(n10948), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U11247 ( .A1(n10948), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U11248 ( .A1(n10942), .A2(n10404), .ZN(n10896) );
  XNOR2_X1 U11249 ( .A(n10422), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U11250 ( .A1(n10896), .A2(n10897), .ZN(n10895) );
  NAND2_X1 U11251 ( .A1(n10904), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U11252 ( .A1(n10895), .A2(n10405), .ZN(n10406) );
  NOR2_X1 U11253 ( .A1(n10406), .A2(n10917), .ZN(n10407) );
  INV_X1 U11254 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10908) );
  NOR2_X1 U11255 ( .A1(n10909), .A2(n10908), .ZN(n10920) );
  NOR2_X1 U11256 ( .A1(n10408), .A2(n10920), .ZN(n10437) );
  XNOR2_X1 U11257 ( .A(n10438), .B(n10437), .ZN(n10433) );
  INV_X1 U11258 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U11259 ( .A1(n10962), .A2(n10441), .ZN(n10410) );
  OAI211_X1 U11260 ( .C1(n10967), .C2(n10411), .A(n10410), .B(n10409), .ZN(
        n10432) );
  INV_X1 U11261 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10421) );
  INV_X1 U11262 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10414) );
  INV_X1 U11263 ( .A(n10412), .ZN(n10413) );
  AOI22_X1 U11264 ( .A1(n10416), .A2(n10415), .B1(n10414), .B2(n10413), .ZN(
        n10939) );
  INV_X1 U11265 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U11266 ( .A1(n10948), .A2(n10418), .ZN(n10417) );
  OAI21_X1 U11267 ( .B1(n10948), .B2(n10418), .A(n10417), .ZN(n10938) );
  NAND2_X1 U11268 ( .A1(n10904), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10419) );
  OAI21_X1 U11269 ( .B1(n10904), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10419), 
        .ZN(n10900) );
  NOR2_X1 U11270 ( .A1(n10901), .A2(n10900), .ZN(n10899) );
  INV_X1 U11271 ( .A(n10899), .ZN(n10420) );
  OAI21_X1 U11272 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(n10423) );
  AND2_X1 U11273 ( .A1(n10423), .A2(n10917), .ZN(n10428) );
  INV_X1 U11274 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10913) );
  INV_X1 U11275 ( .A(n10428), .ZN(n10427) );
  INV_X1 U11276 ( .A(n10423), .ZN(n10425) );
  INV_X1 U11277 ( .A(n10917), .ZN(n10424) );
  NAND2_X1 U11278 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NAND2_X1 U11279 ( .A1(n10427), .A2(n10426), .ZN(n10914) );
  NOR2_X1 U11280 ( .A1(n10428), .A2(n10912), .ZN(n10430) );
  XNOR2_X1 U11281 ( .A(n10441), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10429) );
  NOR2_X1 U11282 ( .A1(n10429), .A2(n10430), .ZN(n10440) );
  AOI211_X1 U11283 ( .C1(n10430), .C2(n10429), .A(n10440), .B(n10952), .ZN(
        n10431) );
  AOI211_X1 U11284 ( .C1(n10910), .C2(n10433), .A(n10432), .B(n10431), .ZN(
        n10434) );
  INV_X1 U11285 ( .A(n10434), .ZN(P1_U3259) );
  INV_X1 U11286 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10436) );
  INV_X1 U11287 ( .A(n10441), .ZN(n10435) );
  AOI22_X1 U11288 ( .A1(n10438), .A2(n10437), .B1(n10436), .B2(n10435), .ZN(
        n10459) );
  XNOR2_X1 U11289 ( .A(n10457), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10458) );
  XNOR2_X1 U11290 ( .A(n10459), .B(n10458), .ZN(n10445) );
  XNOR2_X1 U11291 ( .A(n10439), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n10443) );
  AOI21_X1 U11292 ( .B1(n10441), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10440), 
        .ZN(n10442) );
  NAND2_X1 U11293 ( .A1(n10442), .A2(n10443), .ZN(n10451) );
  OAI21_X1 U11294 ( .B1(n10443), .B2(n10442), .A(n10451), .ZN(n10444) );
  AOI22_X1 U11295 ( .A1(n10910), .A2(n10445), .B1(n10916), .B2(n10444), .ZN(
        n10450) );
  INV_X1 U11296 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10447) );
  OAI21_X1 U11297 ( .B1(n10967), .B2(n10447), .A(n10446), .ZN(n10448) );
  AOI21_X1 U11298 ( .B1(n10457), .B2(n10962), .A(n10448), .ZN(n10449) );
  NAND2_X1 U11299 ( .A1(n10450), .A2(n10449), .ZN(P1_U3260) );
  OAI21_X1 U11300 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10457), .A(n10451), 
        .ZN(n10930) );
  NAND2_X1 U11301 ( .A1(n10934), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10452) );
  OAI21_X1 U11302 ( .B1(n10934), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10452), 
        .ZN(n10931) );
  INV_X1 U11303 ( .A(n10452), .ZN(n10453) );
  NOR2_X1 U11304 ( .A1(n10929), .A2(n10453), .ZN(n10456) );
  INV_X1 U11305 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10454) );
  MUX2_X1 U11306 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10454), .S(n6421), .Z(
        n10455) );
  XNOR2_X1 U11307 ( .A(n10456), .B(n10455), .ZN(n10470) );
  OAI22_X1 U11308 ( .A1(n10459), .A2(n10458), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n10457), .ZN(n10927) );
  NAND2_X1 U11309 ( .A1(n10934), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10460) );
  OAI21_X1 U11310 ( .B1(n10934), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10460), 
        .ZN(n10928) );
  NOR2_X1 U11311 ( .A1(n10927), .A2(n10928), .ZN(n10926) );
  INV_X1 U11312 ( .A(n10460), .ZN(n10461) );
  NOR2_X1 U11313 ( .A1(n10926), .A2(n10461), .ZN(n10463) );
  XNOR2_X1 U11314 ( .A(n6421), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10462) );
  XNOR2_X1 U11315 ( .A(n10463), .B(n10462), .ZN(n10468) );
  NAND2_X1 U11316 ( .A1(n10962), .A2(n10464), .ZN(n10466) );
  OAI211_X1 U11317 ( .C1(n5757), .C2(n10967), .A(n10466), .B(n10465), .ZN(
        n10467) );
  AOI21_X1 U11318 ( .B1(n10468), .B2(n10910), .A(n10467), .ZN(n10469) );
  OAI21_X1 U11319 ( .B1(n10470), .B2(n10952), .A(n10469), .ZN(P1_U3262) );
  XNOR2_X1 U11320 ( .A(n10473), .B(n10472), .ZN(n10668) );
  NAND2_X1 U11321 ( .A1(n10668), .A2(n10480), .ZN(n10478) );
  INV_X1 U11322 ( .A(n10671), .ZN(n10476) );
  NOR2_X1 U11323 ( .A1(n10476), .A2(n7511), .ZN(n10481) );
  AOI21_X1 U11324 ( .B1(n7511), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10481), .ZN(
        n10477) );
  OAI211_X1 U11325 ( .C1(n10775), .C2(n10658), .A(n10478), .B(n10477), .ZN(
        P1_U3263) );
  XNOR2_X1 U11326 ( .A(n10779), .B(n10479), .ZN(n10673) );
  NAND2_X1 U11327 ( .A1(n10673), .A2(n10480), .ZN(n10483) );
  AOI21_X1 U11328 ( .B1(n7511), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10481), .ZN(
        n10482) );
  OAI211_X1 U11329 ( .C1(n10779), .C2(n10658), .A(n10483), .B(n10482), .ZN(
        P1_U3264) );
  INV_X1 U11330 ( .A(n10484), .ZN(n10498) );
  NAND2_X1 U11331 ( .A1(n10485), .A2(n10651), .ZN(n10497) );
  INV_X1 U11332 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10486) );
  OAI22_X1 U11333 ( .A1(n10487), .A2(n10572), .B1(n10601), .B2(n10486), .ZN(
        n10490) );
  NOR2_X1 U11334 ( .A1(n10685), .A2(n10488), .ZN(n10489) );
  AOI211_X1 U11335 ( .C1(n10632), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        n10492) );
  OAI21_X1 U11336 ( .B1(n10493), .B2(n10658), .A(n10492), .ZN(n10494) );
  AOI21_X1 U11337 ( .B1(n10495), .B2(n10664), .A(n10494), .ZN(n10496) );
  OAI211_X1 U11338 ( .C1(n10498), .C2(n10583), .A(n10497), .B(n10496), .ZN(
        P1_U3265) );
  AOI21_X1 U11339 ( .B1(n10500), .B2(n10499), .A(n5210), .ZN(n10683) );
  AOI211_X1 U11340 ( .C1(n10679), .C2(n10515), .A(n10655), .B(n10501), .ZN(
        n10677) );
  NOR2_X1 U11341 ( .A1(n5433), .A2(n10658), .ZN(n10507) );
  AOI22_X1 U11342 ( .A1(n10502), .A2(n10632), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n7511), .ZN(n10505) );
  NAND2_X1 U11343 ( .A1(n10503), .A2(n10569), .ZN(n10504) );
  OAI211_X1 U11344 ( .C1(n10676), .C2(n10572), .A(n10505), .B(n10504), .ZN(
        n10506) );
  AOI211_X1 U11345 ( .C1(n10677), .C2(n10664), .A(n10507), .B(n10506), .ZN(
        n10511) );
  XNOR2_X1 U11346 ( .A(n10509), .B(n10508), .ZN(n10680) );
  NAND2_X1 U11347 ( .A1(n10680), .A2(n10529), .ZN(n10510) );
  OAI211_X1 U11348 ( .C1(n10683), .C2(n10638), .A(n10511), .B(n10510), .ZN(
        P1_U3266) );
  OAI21_X1 U11349 ( .B1(n10513), .B2(n10526), .A(n10512), .ZN(n10692) );
  INV_X1 U11350 ( .A(n10515), .ZN(n10516) );
  AOI211_X1 U11351 ( .C1(n10688), .C2(n10537), .A(n10655), .B(n10516), .ZN(
        n10686) );
  NOR2_X1 U11352 ( .A1(n10517), .A2(n10658), .ZN(n10524) );
  INV_X1 U11353 ( .A(n10518), .ZN(n10519) );
  AOI22_X1 U11354 ( .A1(n10519), .A2(n10632), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n7511), .ZN(n10522) );
  NAND2_X1 U11355 ( .A1(n10520), .A2(n10569), .ZN(n10521) );
  OAI211_X1 U11356 ( .C1(n10685), .C2(n10572), .A(n10522), .B(n10521), .ZN(
        n10523) );
  AOI211_X1 U11357 ( .C1(n10686), .C2(n10664), .A(n10524), .B(n10523), .ZN(
        n10531) );
  AOI21_X1 U11358 ( .B1(n10527), .B2(n10526), .A(n10525), .ZN(n10528) );
  INV_X1 U11359 ( .A(n10528), .ZN(n10689) );
  NAND2_X1 U11360 ( .A1(n10689), .A2(n10529), .ZN(n10530) );
  OAI211_X1 U11361 ( .C1(n10692), .C2(n10638), .A(n10531), .B(n10530), .ZN(
        P1_U3267) );
  NAND2_X1 U11362 ( .A1(n5583), .A2(n10532), .ZN(n10534) );
  AOI21_X1 U11363 ( .B1(n10536), .B2(n10534), .A(n10533), .ZN(n10698) );
  XOR2_X1 U11364 ( .A(n10535), .B(n10536), .Z(n10700) );
  NAND2_X1 U11365 ( .A1(n10700), .A2(n10651), .ZN(n10546) );
  AOI211_X1 U11366 ( .C1(n10538), .C2(n10554), .A(n10655), .B(n10514), .ZN(
        n10696) );
  INV_X1 U11367 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10539) );
  OAI22_X1 U11368 ( .A1(n10540), .A2(n10659), .B1(n10539), .B2(n10601), .ZN(
        n10542) );
  NOR2_X1 U11369 ( .A1(n10694), .A2(n10572), .ZN(n10541) );
  AOI211_X1 U11370 ( .C1(n10569), .C2(n10710), .A(n10542), .B(n10541), .ZN(
        n10543) );
  OAI21_X1 U11371 ( .B1(n10785), .B2(n10658), .A(n10543), .ZN(n10544) );
  AOI21_X1 U11372 ( .B1(n10696), .B2(n10664), .A(n10544), .ZN(n10545) );
  OAI211_X1 U11373 ( .C1(n10698), .C2(n10583), .A(n10546), .B(n10545), .ZN(
        P1_U3268) );
  XNOR2_X1 U11374 ( .A(n10547), .B(n10550), .ZN(n10705) );
  AOI211_X1 U11375 ( .C1(n10550), .C2(n10549), .A(n10713), .B(n10548), .ZN(
        n10553) );
  OAI22_X1 U11376 ( .A1(n10684), .A2(n10741), .B1(n10551), .B2(n10763), .ZN(
        n10552) );
  NOR2_X1 U11377 ( .A1(n10553), .A2(n10552), .ZN(n10704) );
  INV_X1 U11378 ( .A(n10704), .ZN(n10560) );
  OAI211_X1 U11379 ( .C1(n10789), .C2(n10574), .A(n10672), .B(n10554), .ZN(
        n10703) );
  AOI22_X1 U11380 ( .A1(n10555), .A2(n10632), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n7511), .ZN(n10558) );
  NAND2_X1 U11381 ( .A1(n10556), .A2(n10580), .ZN(n10557) );
  OAI211_X1 U11382 ( .C1(n10703), .C2(n10576), .A(n10558), .B(n10557), .ZN(
        n10559) );
  AOI21_X1 U11383 ( .B1(n10560), .B2(n10601), .A(n10559), .ZN(n10561) );
  OAI21_X1 U11384 ( .B1(n10705), .B2(n10638), .A(n10561), .ZN(P1_U3269) );
  OAI21_X1 U11385 ( .B1(n10563), .B2(n10566), .A(n10562), .ZN(n10564) );
  INV_X1 U11386 ( .A(n10564), .ZN(n10714) );
  XOR2_X1 U11387 ( .A(n10566), .B(n10565), .Z(n10716) );
  NAND2_X1 U11388 ( .A1(n10716), .A2(n10651), .ZN(n10582) );
  INV_X1 U11389 ( .A(n10567), .ZN(n10568) );
  AOI22_X1 U11390 ( .A1(n10568), .A2(n10632), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n7511), .ZN(n10571) );
  NAND2_X1 U11391 ( .A1(n10709), .A2(n10569), .ZN(n10570) );
  OAI211_X1 U11392 ( .C1(n10693), .C2(n10572), .A(n10571), .B(n10570), .ZN(
        n10578) );
  INV_X1 U11393 ( .A(n10573), .ZN(n10594) );
  INV_X1 U11394 ( .A(n10574), .ZN(n10575) );
  OAI211_X1 U11395 ( .C1(n10793), .C2(n10594), .A(n10575), .B(n10672), .ZN(
        n10711) );
  NOR2_X1 U11396 ( .A1(n10711), .A2(n10576), .ZN(n10577) );
  AOI211_X1 U11397 ( .C1(n10580), .C2(n10579), .A(n10578), .B(n10577), .ZN(
        n10581) );
  OAI211_X1 U11398 ( .C1(n10714), .C2(n10583), .A(n10582), .B(n10581), .ZN(
        P1_U3270) );
  OAI21_X1 U11399 ( .B1(n10585), .B2(n10586), .A(n10584), .ZN(n10721) );
  INV_X1 U11400 ( .A(n10721), .ZN(n10603) );
  XNOR2_X1 U11401 ( .A(n10587), .B(n10586), .ZN(n10588) );
  NAND2_X1 U11402 ( .A1(n10588), .A2(n10746), .ZN(n10592) );
  AOI22_X1 U11403 ( .A1(n11155), .A2(n10590), .B1(n10589), .B2(n11156), .ZN(
        n10591) );
  NAND2_X1 U11404 ( .A1(n10592), .A2(n10591), .ZN(n10719) );
  INV_X1 U11405 ( .A(n10595), .ZN(n10797) );
  AOI211_X1 U11406 ( .C1(n10595), .C2(n10608), .A(n10655), .B(n10594), .ZN(
        n10720) );
  NAND2_X1 U11407 ( .A1(n10720), .A2(n10664), .ZN(n10599) );
  INV_X1 U11408 ( .A(n10596), .ZN(n10597) );
  AOI22_X1 U11409 ( .A1(n10597), .A2(n10632), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n7511), .ZN(n10598) );
  OAI211_X1 U11410 ( .C1(n10797), .C2(n10658), .A(n10599), .B(n10598), .ZN(
        n10600) );
  AOI21_X1 U11411 ( .B1(n10601), .B2(n10719), .A(n10600), .ZN(n10602) );
  OAI21_X1 U11412 ( .B1(n10603), .B2(n10638), .A(n10602), .ZN(P1_U3271) );
  OAI21_X1 U11413 ( .B1(n10606), .B2(n10605), .A(n10604), .ZN(n10607) );
  INV_X1 U11414 ( .A(n10607), .ZN(n10728) );
  AOI211_X1 U11415 ( .C1(n10725), .C2(n10630), .A(n10655), .B(n10593), .ZN(
        n10724) );
  INV_X1 U11416 ( .A(n10725), .ZN(n10612) );
  INV_X1 U11417 ( .A(n10609), .ZN(n10610) );
  AOI22_X1 U11418 ( .A1(n10610), .A2(n10632), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n7511), .ZN(n10611) );
  OAI21_X1 U11419 ( .B1(n10612), .B2(n10658), .A(n10611), .ZN(n10619) );
  OAI21_X1 U11420 ( .B1(n10615), .B2(n10614), .A(n10613), .ZN(n10617) );
  AOI222_X1 U11421 ( .A1(n10746), .A2(n10617), .B1(n10616), .B2(n11156), .C1(
        n10709), .C2(n11155), .ZN(n10727) );
  NOR2_X1 U11422 ( .A1(n10727), .A2(n7511), .ZN(n10618) );
  AOI211_X1 U11423 ( .C1(n10724), .C2(n10664), .A(n10619), .B(n10618), .ZN(
        n10620) );
  OAI21_X1 U11424 ( .B1(n10728), .B2(n10638), .A(n10620), .ZN(P1_U3272) );
  XNOR2_X1 U11425 ( .A(n10621), .B(n10624), .ZN(n10731) );
  INV_X1 U11426 ( .A(n10731), .ZN(n10639) );
  OAI21_X1 U11427 ( .B1(n10624), .B2(n10623), .A(n10622), .ZN(n10625) );
  NAND2_X1 U11428 ( .A1(n10625), .A2(n10746), .ZN(n10629) );
  OAI22_X1 U11429 ( .A1(n10626), .A2(n10741), .B1(n10742), .B2(n10763), .ZN(
        n10627) );
  INV_X1 U11430 ( .A(n10627), .ZN(n10628) );
  NAND2_X1 U11431 ( .A1(n10629), .A2(n10628), .ZN(n10729) );
  INV_X1 U11432 ( .A(n10631), .ZN(n10802) );
  AOI211_X1 U11433 ( .C1(n10631), .C2(n10653), .A(n10655), .B(n5439), .ZN(
        n10730) );
  NAND2_X1 U11434 ( .A1(n10730), .A2(n10664), .ZN(n10635) );
  AOI22_X1 U11435 ( .A1(n10633), .A2(n10632), .B1(n7511), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n10634) );
  OAI211_X1 U11436 ( .C1(n10802), .C2(n10658), .A(n10635), .B(n10634), .ZN(
        n10636) );
  AOI21_X1 U11437 ( .B1(n10729), .B2(n10601), .A(n10636), .ZN(n10637) );
  OAI21_X1 U11438 ( .B1(n10639), .B2(n10638), .A(n10637), .ZN(P1_U3273) );
  OAI21_X1 U11439 ( .B1(n10642), .B2(n10641), .A(n10640), .ZN(n10643) );
  NAND2_X1 U11440 ( .A1(n10643), .A2(n10746), .ZN(n10648) );
  OAI22_X1 U11441 ( .A1(n10645), .A2(n10741), .B1(n10644), .B2(n10763), .ZN(
        n10646) );
  INV_X1 U11442 ( .A(n10646), .ZN(n10647) );
  NAND2_X1 U11443 ( .A1(n10648), .A2(n10647), .ZN(n10734) );
  INV_X1 U11444 ( .A(n10734), .ZN(n10667) );
  XNOR2_X1 U11445 ( .A(n10650), .B(n10649), .ZN(n10736) );
  NAND2_X1 U11446 ( .A1(n10736), .A2(n10651), .ZN(n10666) );
  INV_X1 U11447 ( .A(n10652), .ZN(n10656) );
  INV_X1 U11448 ( .A(n10653), .ZN(n10654) );
  AOI211_X1 U11449 ( .C1(n10657), .C2(n10656), .A(n10655), .B(n10654), .ZN(
        n10735) );
  NOR2_X1 U11450 ( .A1(n10807), .A2(n10658), .ZN(n10663) );
  OAI22_X1 U11451 ( .A1(n10661), .A2(n10454), .B1(n10660), .B2(n10659), .ZN(
        n10662) );
  AOI211_X1 U11452 ( .C1(n10735), .C2(n10664), .A(n10663), .B(n10662), .ZN(
        n10665) );
  OAI211_X1 U11453 ( .C1(n7511), .C2(n10667), .A(n10666), .B(n10665), .ZN(
        P1_U3274) );
  INV_X1 U11454 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10669) );
  AOI21_X1 U11455 ( .B1(n10668), .B2(n10672), .A(n10671), .ZN(n10772) );
  MUX2_X1 U11456 ( .A(n10669), .B(n10772), .S(n11181), .Z(n10670) );
  OAI21_X1 U11457 ( .B1(n10775), .B2(n10739), .A(n10670), .ZN(P1_U3553) );
  AOI21_X1 U11458 ( .B1(n10673), .B2(n10672), .A(n10671), .ZN(n10776) );
  MUX2_X1 U11459 ( .A(n10674), .B(n10776), .S(n11181), .Z(n10675) );
  OAI21_X1 U11460 ( .B1(n10779), .B2(n10739), .A(n10675), .ZN(P1_U3552) );
  OAI22_X1 U11461 ( .A1(n10676), .A2(n10741), .B1(n10694), .B2(n10763), .ZN(
        n10678) );
  AOI211_X1 U11462 ( .C1(n11127), .C2(n10679), .A(n10678), .B(n10677), .ZN(
        n10682) );
  NAND2_X1 U11463 ( .A1(n10680), .A2(n10746), .ZN(n10681) );
  OAI211_X1 U11464 ( .C1(n10683), .C2(n10770), .A(n10682), .B(n10681), .ZN(
        n10780) );
  MUX2_X1 U11465 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10780), .S(n11181), .Z(
        P1_U3549) );
  OAI22_X1 U11466 ( .A1(n10685), .A2(n10741), .B1(n10684), .B2(n10763), .ZN(
        n10687) );
  AOI211_X1 U11467 ( .C1(n11127), .C2(n10688), .A(n10687), .B(n10686), .ZN(
        n10691) );
  NAND2_X1 U11468 ( .A1(n10689), .A2(n10746), .ZN(n10690) );
  OAI211_X1 U11469 ( .C1(n10692), .C2(n10770), .A(n10691), .B(n10690), .ZN(
        n10781) );
  MUX2_X1 U11470 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10781), .S(n11181), .Z(
        P1_U3548) );
  OAI22_X1 U11471 ( .A1(n10694), .A2(n10741), .B1(n10693), .B2(n10763), .ZN(
        n10695) );
  NOR2_X1 U11472 ( .A1(n10696), .A2(n10695), .ZN(n10697) );
  OAI21_X1 U11473 ( .B1(n10698), .B2(n10713), .A(n10697), .ZN(n10699) );
  AOI21_X1 U11474 ( .B1(n10700), .B2(n11178), .A(n10699), .ZN(n10782) );
  MUX2_X1 U11475 ( .A(n10701), .B(n10782), .S(n11181), .Z(n10702) );
  OAI21_X1 U11476 ( .B1(n10785), .B2(n10739), .A(n10702), .ZN(P1_U3547) );
  OAI211_X1 U11477 ( .C1(n10705), .C2(n10770), .A(n10704), .B(n10703), .ZN(
        n10706) );
  INV_X1 U11478 ( .A(n10706), .ZN(n10786) );
  MUX2_X1 U11479 ( .A(n10707), .B(n10786), .S(n11181), .Z(n10708) );
  OAI21_X1 U11480 ( .B1(n10789), .B2(n10739), .A(n10708), .ZN(P1_U3546) );
  AOI22_X1 U11481 ( .A1(n10710), .A2(n11155), .B1(n11156), .B2(n10709), .ZN(
        n10712) );
  OAI211_X1 U11482 ( .C1(n10714), .C2(n10713), .A(n10712), .B(n10711), .ZN(
        n10715) );
  AOI21_X1 U11483 ( .B1(n10716), .B2(n11178), .A(n10715), .ZN(n10790) );
  MUX2_X1 U11484 ( .A(n10717), .B(n10790), .S(n11181), .Z(n10718) );
  OAI21_X1 U11485 ( .B1(n10793), .B2(n10739), .A(n10718), .ZN(P1_U3545) );
  AOI211_X1 U11486 ( .C1(n10721), .C2(n11178), .A(n10720), .B(n10719), .ZN(
        n10794) );
  MUX2_X1 U11487 ( .A(n10722), .B(n10794), .S(n11181), .Z(n10723) );
  OAI21_X1 U11488 ( .B1(n10797), .B2(n10739), .A(n10723), .ZN(P1_U3544) );
  AOI21_X1 U11489 ( .B1(n11127), .B2(n10725), .A(n10724), .ZN(n10726) );
  OAI211_X1 U11490 ( .C1(n10728), .C2(n10770), .A(n10727), .B(n10726), .ZN(
        n10798) );
  MUX2_X1 U11491 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10798), .S(n11181), .Z(
        P1_U3543) );
  INV_X1 U11492 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10732) );
  AOI211_X1 U11493 ( .C1(n10731), .C2(n11178), .A(n10730), .B(n10729), .ZN(
        n10799) );
  MUX2_X1 U11494 ( .A(n10732), .B(n10799), .S(n11181), .Z(n10733) );
  OAI21_X1 U11495 ( .B1(n10802), .B2(n10739), .A(n10733), .ZN(P1_U3542) );
  INV_X1 U11496 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10737) );
  AOI211_X1 U11497 ( .C1(n10736), .C2(n11178), .A(n10735), .B(n10734), .ZN(
        n10803) );
  MUX2_X1 U11498 ( .A(n10737), .B(n10803), .S(n11181), .Z(n10738) );
  OAI21_X1 U11499 ( .B1(n10807), .B2(n10739), .A(n10738), .ZN(P1_U3541) );
  OAI22_X1 U11500 ( .A1(n10742), .A2(n10741), .B1(n10740), .B2(n10763), .ZN(
        n10744) );
  AOI211_X1 U11501 ( .C1(n11127), .C2(n10745), .A(n10744), .B(n10743), .ZN(
        n10749) );
  NAND2_X1 U11502 ( .A1(n10747), .A2(n10746), .ZN(n10748) );
  OAI211_X1 U11503 ( .C1(n10750), .C2(n10770), .A(n10749), .B(n10748), .ZN(
        n10808) );
  MUX2_X1 U11504 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10808), .S(n11181), .Z(
        P1_U3540) );
  AOI211_X1 U11505 ( .C1(n11127), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        n10754) );
  OAI21_X1 U11506 ( .B1(n10755), .B2(n10770), .A(n10754), .ZN(n10809) );
  MUX2_X1 U11507 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10809), .S(n11181), .Z(
        P1_U3539) );
  NOR2_X1 U11508 ( .A1(n10756), .A2(n10763), .ZN(n10758) );
  AOI211_X1 U11509 ( .C1(n11127), .C2(n10759), .A(n10758), .B(n10757), .ZN(
        n10760) );
  OAI211_X1 U11510 ( .C1(n10762), .C2(n10770), .A(n10761), .B(n10760), .ZN(
        n10810) );
  MUX2_X1 U11511 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10810), .S(n11181), .Z(
        P1_U3538) );
  NOR2_X1 U11512 ( .A1(n10764), .A2(n10763), .ZN(n10766) );
  AOI211_X1 U11513 ( .C1(n11127), .C2(n10767), .A(n10766), .B(n10765), .ZN(
        n10768) );
  OAI211_X1 U11514 ( .C1(n10771), .C2(n10770), .A(n10769), .B(n10768), .ZN(
        n10811) );
  MUX2_X1 U11515 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10811), .S(n11181), .Z(
        P1_U3537) );
  INV_X1 U11516 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10773) );
  MUX2_X1 U11517 ( .A(n10773), .B(n10772), .S(n11185), .Z(n10774) );
  OAI21_X1 U11518 ( .B1(n10775), .B2(n10806), .A(n10774), .ZN(P1_U3521) );
  INV_X1 U11519 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10777) );
  MUX2_X1 U11520 ( .A(n10777), .B(n10776), .S(n11185), .Z(n10778) );
  OAI21_X1 U11521 ( .B1(n10779), .B2(n10806), .A(n10778), .ZN(P1_U3520) );
  MUX2_X1 U11522 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10780), .S(n11185), .Z(
        P1_U3517) );
  MUX2_X1 U11523 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10781), .S(n11185), .Z(
        P1_U3516) );
  INV_X1 U11524 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10783) );
  MUX2_X1 U11525 ( .A(n10783), .B(n10782), .S(n11185), .Z(n10784) );
  OAI21_X1 U11526 ( .B1(n10785), .B2(n10806), .A(n10784), .ZN(P1_U3515) );
  INV_X1 U11527 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10787) );
  MUX2_X1 U11528 ( .A(n10787), .B(n10786), .S(n11185), .Z(n10788) );
  OAI21_X1 U11529 ( .B1(n10789), .B2(n10806), .A(n10788), .ZN(P1_U3514) );
  INV_X1 U11530 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10791) );
  MUX2_X1 U11531 ( .A(n10791), .B(n10790), .S(n11185), .Z(n10792) );
  OAI21_X1 U11532 ( .B1(n10793), .B2(n10806), .A(n10792), .ZN(P1_U3513) );
  INV_X1 U11533 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10795) );
  MUX2_X1 U11534 ( .A(n10795), .B(n10794), .S(n11185), .Z(n10796) );
  OAI21_X1 U11535 ( .B1(n10797), .B2(n10806), .A(n10796), .ZN(P1_U3512) );
  MUX2_X1 U11536 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10798), .S(n11185), .Z(
        P1_U3511) );
  INV_X1 U11537 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10800) );
  MUX2_X1 U11538 ( .A(n10800), .B(n10799), .S(n11185), .Z(n10801) );
  OAI21_X1 U11539 ( .B1(n10802), .B2(n10806), .A(n10801), .ZN(P1_U3510) );
  INV_X1 U11540 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10804) );
  MUX2_X1 U11541 ( .A(n10804), .B(n10803), .S(n11185), .Z(n10805) );
  OAI21_X1 U11542 ( .B1(n10807), .B2(n10806), .A(n10805), .ZN(P1_U3509) );
  MUX2_X1 U11543 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10808), .S(n11185), .Z(
        P1_U3507) );
  MUX2_X1 U11544 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10809), .S(n11185), .Z(
        P1_U3504) );
  MUX2_X1 U11545 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10810), .S(n11185), .Z(
        P1_U3501) );
  MUX2_X1 U11546 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10811), .S(n11185), .Z(
        P1_U3498) );
  AND2_X1 U11547 ( .A1(n10813), .A2(n10812), .ZN(n10826) );
  MUX2_X1 U11548 ( .A(P1_D_REG_1__SCAN_IN), .B(n10814), .S(n10826), .Z(
        P1_U3440) );
  MUX2_X1 U11549 ( .A(P1_D_REG_0__SCAN_IN), .B(n10815), .S(n10826), .Z(
        P1_U3439) );
  INV_X1 U11550 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10816) );
  NAND3_X1 U11551 ( .A1(n10816), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10818) );
  OAI22_X1 U11552 ( .A1(n5868), .A2(n10818), .B1(n10817), .B2(n9220), .ZN(
        n10819) );
  AOI21_X1 U11553 ( .B1(n10821), .B2(n10820), .A(n10819), .ZN(n10822) );
  INV_X1 U11554 ( .A(n10822), .ZN(P1_U3324) );
  MUX2_X1 U11555 ( .A(n10823), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11556 ( .A1(n10826), .A2(n10824), .ZN(P1_U3323) );
  AND2_X1 U11557 ( .A1(n10827), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  INV_X1 U11558 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10825) );
  NOR2_X1 U11559 ( .A1(n10826), .A2(n10825), .ZN(P1_U3321) );
  AND2_X1 U11560 ( .A1(n10827), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11561 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10827), .ZN(P1_U3319) );
  AND2_X1 U11562 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10827), .ZN(P1_U3318) );
  AND2_X1 U11563 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10827), .ZN(P1_U3317) );
  AND2_X1 U11564 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10827), .ZN(P1_U3316) );
  AND2_X1 U11565 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10827), .ZN(P1_U3315) );
  AND2_X1 U11566 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10827), .ZN(P1_U3314) );
  AND2_X1 U11567 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10827), .ZN(P1_U3313) );
  AND2_X1 U11568 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10827), .ZN(P1_U3312) );
  AND2_X1 U11569 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10827), .ZN(P1_U3311) );
  AND2_X1 U11570 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10827), .ZN(P1_U3310) );
  AND2_X1 U11571 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10827), .ZN(P1_U3309) );
  AND2_X1 U11572 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10827), .ZN(P1_U3308) );
  AND2_X1 U11573 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10827), .ZN(P1_U3307) );
  AND2_X1 U11574 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10827), .ZN(P1_U3306) );
  AND2_X1 U11575 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10827), .ZN(P1_U3305) );
  AND2_X1 U11576 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10827), .ZN(P1_U3304) );
  AND2_X1 U11577 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10827), .ZN(P1_U3303) );
  AND2_X1 U11578 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10827), .ZN(P1_U3302) );
  AND2_X1 U11579 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10827), .ZN(P1_U3301) );
  AND2_X1 U11580 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10827), .ZN(P1_U3300) );
  AND2_X1 U11581 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10827), .ZN(P1_U3299) );
  AND2_X1 U11582 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10827), .ZN(P1_U3298) );
  AND2_X1 U11583 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10827), .ZN(P1_U3297) );
  AND2_X1 U11584 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10827), .ZN(P1_U3296) );
  AND2_X1 U11585 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10827), .ZN(P1_U3295) );
  AND2_X1 U11586 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10827), .ZN(P1_U3294) );
  XOR2_X1 U11587 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11588 ( .A1(n10992), .A2(n10831), .B1(n10992), .B2(n10830), .C1(
        n10829), .C2(n10828), .ZN(ADD_1068_U5) );
  AOI21_X1 U11589 ( .B1(n10834), .B2(n10833), .A(n10832), .ZN(ADD_1068_U54) );
  AOI21_X1 U11590 ( .B1(n10837), .B2(n10836), .A(n10835), .ZN(ADD_1068_U53) );
  OAI21_X1 U11591 ( .B1(n10840), .B2(n10839), .A(n10838), .ZN(ADD_1068_U52) );
  OAI21_X1 U11592 ( .B1(n10843), .B2(n10842), .A(n10841), .ZN(ADD_1068_U51) );
  OAI21_X1 U11593 ( .B1(n10846), .B2(n10845), .A(n10844), .ZN(ADD_1068_U50) );
  OAI21_X1 U11594 ( .B1(n10849), .B2(n10848), .A(n10847), .ZN(ADD_1068_U49) );
  OAI21_X1 U11595 ( .B1(n10852), .B2(n10851), .A(n10850), .ZN(ADD_1068_U48) );
  OAI21_X1 U11596 ( .B1(n10855), .B2(n10854), .A(n10853), .ZN(ADD_1068_U47) );
  OAI21_X1 U11597 ( .B1(n10858), .B2(n10857), .A(n10856), .ZN(ADD_1068_U63) );
  OAI21_X1 U11598 ( .B1(n10861), .B2(n10860), .A(n10859), .ZN(ADD_1068_U62) );
  OAI21_X1 U11599 ( .B1(n10864), .B2(n10863), .A(n10862), .ZN(ADD_1068_U61) );
  OAI21_X1 U11600 ( .B1(n10867), .B2(n10866), .A(n10865), .ZN(ADD_1068_U60) );
  OAI21_X1 U11601 ( .B1(n10870), .B2(n10869), .A(n10868), .ZN(ADD_1068_U59) );
  OAI21_X1 U11602 ( .B1(n10873), .B2(n10872), .A(n10871), .ZN(ADD_1068_U58) );
  OAI21_X1 U11603 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(ADD_1068_U57) );
  OAI21_X1 U11604 ( .B1(n10879), .B2(n10878), .A(n10877), .ZN(ADD_1068_U56) );
  OAI21_X1 U11605 ( .B1(n10882), .B2(n10881), .A(n10880), .ZN(ADD_1068_U55) );
  INV_X1 U11606 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10894) );
  AOI211_X1 U11607 ( .C1(n10885), .C2(n10884), .A(n10883), .B(n10952), .ZN(
        n10890) );
  AOI211_X1 U11608 ( .C1(n10888), .C2(n10887), .A(n10886), .B(n10956), .ZN(
        n10889) );
  AOI211_X1 U11609 ( .C1(n10962), .C2(n10891), .A(n10890), .B(n10889), .ZN(
        n10893) );
  OAI211_X1 U11610 ( .C1(n10967), .C2(n10894), .A(n10893), .B(n10892), .ZN(
        P1_U3254) );
  INV_X1 U11611 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10907) );
  OAI211_X1 U11612 ( .C1(n10897), .C2(n10896), .A(n10910), .B(n10895), .ZN(
        n10898) );
  INV_X1 U11613 ( .A(n10898), .ZN(n10903) );
  AOI211_X1 U11614 ( .C1(n10901), .C2(n10900), .A(n10899), .B(n10952), .ZN(
        n10902) );
  AOI211_X1 U11615 ( .C1(n10962), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10906) );
  NAND2_X1 U11616 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10905)
         );
  OAI211_X1 U11617 ( .C1(n10967), .C2(n10907), .A(n10906), .B(n10905), .ZN(
        P1_U3257) );
  INV_X1 U11618 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10925) );
  NAND2_X1 U11619 ( .A1(n10909), .A2(n10908), .ZN(n10911) );
  NAND2_X1 U11620 ( .A1(n10911), .A2(n10910), .ZN(n10919) );
  AOI21_X1 U11621 ( .B1(n10914), .B2(n10913), .A(n10912), .ZN(n10915) );
  AOI22_X1 U11622 ( .A1(n10917), .A2(n10962), .B1(n10916), .B2(n10915), .ZN(
        n10918) );
  OAI21_X1 U11623 ( .B1(n10920), .B2(n10919), .A(n10918), .ZN(n10921) );
  INV_X1 U11624 ( .A(n10921), .ZN(n10924) );
  INV_X1 U11625 ( .A(n10922), .ZN(n10923) );
  OAI211_X1 U11626 ( .C1(n10967), .C2(n10925), .A(n10924), .B(n10923), .ZN(
        P1_U3258) );
  INV_X1 U11627 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10937) );
  AOI211_X1 U11628 ( .C1(n10928), .C2(n10927), .A(n10956), .B(n10926), .ZN(
        n10933) );
  AOI211_X1 U11629 ( .C1(n10931), .C2(n10930), .A(n10952), .B(n10929), .ZN(
        n10932) );
  AOI211_X1 U11630 ( .C1(n10962), .C2(n10934), .A(n10933), .B(n10932), .ZN(
        n10936) );
  OAI211_X1 U11631 ( .C1(n10967), .C2(n10937), .A(n10936), .B(n10935), .ZN(
        P1_U3261) );
  INV_X1 U11632 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10951) );
  NOR2_X1 U11633 ( .A1(n10939), .A2(n10938), .ZN(n10940) );
  NOR3_X1 U11634 ( .A1(n10952), .A2(n10941), .A3(n10940), .ZN(n10947) );
  INV_X1 U11635 ( .A(n10942), .ZN(n10943) );
  AOI211_X1 U11636 ( .C1(n10945), .C2(n10944), .A(n10943), .B(n10956), .ZN(
        n10946) );
  AOI211_X1 U11637 ( .C1(n10962), .C2(n10948), .A(n10947), .B(n10946), .ZN(
        n10950) );
  OAI211_X1 U11638 ( .C1(n10967), .C2(n10951), .A(n10950), .B(n10949), .ZN(
        P1_U3256) );
  INV_X1 U11639 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10966) );
  AOI211_X1 U11640 ( .C1(n10955), .C2(n10954), .A(n10953), .B(n10952), .ZN(
        n10961) );
  AOI211_X1 U11641 ( .C1(n10959), .C2(n10958), .A(n10957), .B(n10956), .ZN(
        n10960) );
  AOI211_X1 U11642 ( .C1(n10963), .C2(n10962), .A(n10961), .B(n10960), .ZN(
        n10965) );
  OAI211_X1 U11643 ( .C1(n10967), .C2(n10966), .A(n10965), .B(n10964), .ZN(
        P1_U3253) );
  AOI22_X1 U11644 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n11076), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10973) );
  INV_X1 U11645 ( .A(n10968), .ZN(n10971) );
  OAI21_X1 U11646 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10969), .A(n10988), .ZN(
        n10970) );
  OAI21_X1 U11647 ( .B1(n10971), .B2(n11086), .A(n10970), .ZN(n10972) );
  OAI211_X1 U11648 ( .C1(n11096), .C2(n10974), .A(n10973), .B(n10972), .ZN(
        P2_U3182) );
  INV_X1 U11649 ( .A(n10975), .ZN(n10979) );
  NAND2_X1 U11650 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  AOI21_X1 U11651 ( .B1(n10979), .B2(n10978), .A(n11081), .ZN(n10986) );
  AND2_X1 U11652 ( .A1(n10981), .A2(n10980), .ZN(n10982) );
  NOR2_X1 U11653 ( .A1(n10983), .A2(n10982), .ZN(n10984) );
  OAI22_X1 U11654 ( .A1(n11096), .A2(n7234), .B1(n11090), .B2(n10984), .ZN(
        n10985) );
  AOI211_X1 U11655 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3151), .A(n10986), 
        .B(n10985), .ZN(n10991) );
  XOR2_X1 U11656 ( .A(n10988), .B(n10987), .Z(n10989) );
  NAND2_X1 U11657 ( .A1(n10989), .A2(n11086), .ZN(n10990) );
  OAI211_X1 U11658 ( .C1(n10992), .C2(n11040), .A(n10991), .B(n10990), .ZN(
        P2_U3183) );
  AOI21_X1 U11659 ( .B1(n10995), .B2(n10994), .A(n10993), .ZN(n10996) );
  OAI22_X1 U11660 ( .A1(n11081), .A2(n10996), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11106), .ZN(n11002) );
  AOI21_X1 U11661 ( .B1(n10999), .B2(n10998), .A(n10997), .ZN(n11000) );
  OAI22_X1 U11662 ( .A1(n11096), .A2(n7237), .B1(n11090), .B2(n11000), .ZN(
        n11001) );
  AOI211_X1 U11663 ( .C1(n11076), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n11002), .B(
        n11001), .ZN(n11007) );
  XOR2_X1 U11664 ( .A(n11003), .B(n11004), .Z(n11005) );
  NAND2_X1 U11665 ( .A1(n11005), .A2(n11086), .ZN(n11006) );
  NAND2_X1 U11666 ( .A1(n11007), .A2(n11006), .ZN(P2_U3184) );
  INV_X1 U11667 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n11024) );
  AOI21_X1 U11668 ( .B1(n7697), .B2(n11009), .A(n11008), .ZN(n11013) );
  AOI21_X1 U11669 ( .B1(n7212), .B2(n11011), .A(n11010), .ZN(n11012) );
  OAI22_X1 U11670 ( .A1(n11013), .A2(n11081), .B1(n11090), .B2(n11012), .ZN(
        n11014) );
  AOI211_X1 U11671 ( .C1(n11016), .C2(n11033), .A(n11015), .B(n11014), .ZN(
        n11023) );
  AOI21_X1 U11672 ( .B1(n11019), .B2(n11018), .A(n11017), .ZN(n11021) );
  OR2_X1 U11673 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  OAI211_X1 U11674 ( .C1(n11024), .C2(n11040), .A(n11023), .B(n11022), .ZN(
        P2_U3185) );
  INV_X1 U11675 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n11041) );
  AOI21_X1 U11676 ( .B1(n11026), .B2(n11025), .A(n5239), .ZN(n11030) );
  AOI21_X1 U11677 ( .B1(n5241), .B2(n11028), .A(n11027), .ZN(n11029) );
  OAI22_X1 U11678 ( .A1(n11030), .A2(n11081), .B1(n11090), .B2(n11029), .ZN(
        n11031) );
  AOI211_X1 U11679 ( .C1(n11034), .C2(n11033), .A(n11032), .B(n11031), .ZN(
        n11039) );
  OAI211_X1 U11680 ( .C1(n11037), .C2(n11036), .A(n11035), .B(n11086), .ZN(
        n11038) );
  OAI211_X1 U11681 ( .C1(n11041), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        P2_U3186) );
  AOI21_X1 U11682 ( .B1(n11044), .B2(n11043), .A(n11042), .ZN(n11045) );
  OAI22_X1 U11683 ( .A1(n11096), .A2(n11046), .B1(n11090), .B2(n11045), .ZN(
        n11047) );
  AOI21_X1 U11684 ( .B1(n11076), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n11047), .ZN(
        n11058) );
  XOR2_X1 U11685 ( .A(n11049), .B(n11048), .Z(n11050) );
  NAND2_X1 U11686 ( .A1(n11050), .A2(n11086), .ZN(n11056) );
  AOI21_X1 U11687 ( .B1(n11053), .B2(n11052), .A(n11051), .ZN(n11054) );
  OR2_X1 U11688 ( .A1(n11081), .A2(n11054), .ZN(n11055) );
  NAND4_X1 U11689 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(
        P2_U3187) );
  AOI21_X1 U11690 ( .B1(n5240), .B2(n11060), .A(n11059), .ZN(n11062) );
  OAI22_X1 U11691 ( .A1(n11062), .A2(n11090), .B1(n11096), .B2(n11061), .ZN(
        n11063) );
  AOI21_X1 U11692 ( .B1(n11076), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n11063), .ZN(
        n11075) );
  OAI21_X1 U11693 ( .B1(n11066), .B2(n11065), .A(n11064), .ZN(n11067) );
  NAND2_X1 U11694 ( .A1(n11067), .A2(n11086), .ZN(n11073) );
  AOI21_X1 U11695 ( .B1(n11070), .B2(n11069), .A(n11068), .ZN(n11071) );
  OR2_X1 U11696 ( .A1(n11081), .A2(n11071), .ZN(n11072) );
  NAND4_X1 U11697 ( .A1(n11075), .A2(n11074), .A3(n11073), .A4(n11072), .ZN(
        P2_U3188) );
  AOI22_X1 U11698 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n11076), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(P2_U3151), .ZN(n11094) );
  AOI21_X1 U11699 ( .B1(n8014), .B2(n11078), .A(n11077), .ZN(n11091) );
  AOI21_X1 U11700 ( .B1(n8017), .B2(n11080), .A(n11079), .ZN(n11082) );
  OR2_X1 U11701 ( .A1(n11082), .A2(n11081), .ZN(n11089) );
  OAI21_X1 U11702 ( .B1(n11085), .B2(n11084), .A(n11083), .ZN(n11087) );
  NAND2_X1 U11703 ( .A1(n11087), .A2(n11086), .ZN(n11088) );
  OAI211_X1 U11704 ( .C1(n11091), .C2(n11090), .A(n11089), .B(n11088), .ZN(
        n11092) );
  INV_X1 U11705 ( .A(n11092), .ZN(n11093) );
  OAI211_X1 U11706 ( .C1(n11096), .C2(n11095), .A(n11094), .B(n11093), .ZN(
        P2_U3193) );
  XOR2_X1 U11707 ( .A(P1_RD_REG_SCAN_IN), .B(n11097), .Z(U126) );
  INV_X1 U11708 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U11709 ( .A1(n11195), .A2(n11099), .B1(n11098), .B2(n11192), .ZN(
        P2_U3393) );
  INV_X1 U11710 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U11711 ( .A1(n11195), .A2(n11101), .B1(n11100), .B2(n11192), .ZN(
        P2_U3396) );
  INV_X1 U11712 ( .A(n11102), .ZN(n11109) );
  OAI22_X1 U11713 ( .A1(n11106), .A2(n11105), .B1(n11104), .B2(n11103), .ZN(
        n11108) );
  AOI211_X1 U11714 ( .C1(n11110), .C2(n11109), .A(n11108), .B(n11107), .ZN(
        n11111) );
  AOI22_X1 U11715 ( .A1(n11124), .A2(n7125), .B1(n11111), .B2(n9692), .ZN(
        P2_U3231) );
  INV_X1 U11716 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U11717 ( .A1(n11195), .A2(n11113), .B1(n11112), .B2(n11192), .ZN(
        P2_U3399) );
  INV_X1 U11718 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U11719 ( .A1(n11195), .A2(n11115), .B1(n11114), .B2(n11192), .ZN(
        P2_U3402) );
  AOI222_X1 U11720 ( .A1(n11121), .A2(n11120), .B1(n11119), .B2(n11118), .C1(
        n11117), .C2(n11116), .ZN(n11122) );
  OAI221_X1 U11721 ( .B1(n11124), .B2(n11123), .C1(n9692), .C2(n7331), .A(
        n11122), .ZN(P2_U3229) );
  INV_X1 U11722 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U11723 ( .A1(n11195), .A2(n11126), .B1(n11125), .B2(n11192), .ZN(
        P2_U3405) );
  INV_X1 U11724 ( .A(n11127), .ZN(n11174) );
  OAI21_X1 U11725 ( .B1(n11129), .B2(n11174), .A(n11128), .ZN(n11131) );
  AOI211_X1 U11726 ( .C1(n11178), .C2(n11132), .A(n11131), .B(n11130), .ZN(
        n11135) );
  INV_X1 U11727 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U11728 ( .A1(n11181), .A2(n11135), .B1(n11133), .B2(n11180), .ZN(
        P1_U3527) );
  INV_X1 U11729 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U11730 ( .A1(n11185), .A2(n11135), .B1(n11134), .B2(n11182), .ZN(
        P1_U3468) );
  INV_X1 U11731 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11136) );
  AOI22_X1 U11732 ( .A1(n11195), .A2(n11137), .B1(n11136), .B2(n11192), .ZN(
        P2_U3408) );
  OAI21_X1 U11733 ( .B1(n11139), .B2(n11174), .A(n11138), .ZN(n11141) );
  AOI211_X1 U11734 ( .C1(n11178), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        n11145) );
  INV_X1 U11735 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U11736 ( .A1(n11181), .A2(n11145), .B1(n11143), .B2(n11180), .ZN(
        P1_U3529) );
  INV_X1 U11737 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U11738 ( .A1(n11185), .A2(n11145), .B1(n11144), .B2(n11182), .ZN(
        P1_U3474) );
  INV_X1 U11739 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U11740 ( .A1(n11195), .A2(n11147), .B1(n11146), .B2(n11192), .ZN(
        P2_U3411) );
  INV_X1 U11741 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U11742 ( .A1(n11195), .A2(n11149), .B1(n11148), .B2(n11192), .ZN(
        P2_U3417) );
  INV_X1 U11743 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11150) );
  AOI22_X1 U11744 ( .A1(n11195), .A2(n11151), .B1(n11150), .B2(n11192), .ZN(
        P2_U3420) );
  INV_X1 U11745 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U11746 ( .A1(n11195), .A2(n11153), .B1(n11152), .B2(n11192), .ZN(
        P2_U3423) );
  AOI22_X1 U11747 ( .A1(n11157), .A2(n11156), .B1(n11155), .B2(n11154), .ZN(
        n11158) );
  OAI211_X1 U11748 ( .C1(n11160), .C2(n11174), .A(n11159), .B(n11158), .ZN(
        n11162) );
  AOI211_X1 U11749 ( .C1(n11164), .C2(n11163), .A(n11162), .B(n11161), .ZN(
        n11165) );
  OAI21_X1 U11750 ( .B1(n11167), .B2(n11166), .A(n11165), .ZN(n11168) );
  INV_X1 U11751 ( .A(n11168), .ZN(n11170) );
  AOI22_X1 U11752 ( .A1(n11181), .A2(n11170), .B1(n7633), .B2(n11180), .ZN(
        P1_U3533) );
  INV_X1 U11753 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U11754 ( .A1(n11185), .A2(n11170), .B1(n11169), .B2(n11182), .ZN(
        P1_U3486) );
  INV_X1 U11755 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U11756 ( .A1(n11195), .A2(n11172), .B1(n11171), .B2(n11192), .ZN(
        P2_U3426) );
  OAI21_X1 U11757 ( .B1(n11175), .B2(n11174), .A(n11173), .ZN(n11176) );
  AOI211_X1 U11758 ( .C1(n11179), .C2(n11178), .A(n11177), .B(n11176), .ZN(
        n11184) );
  AOI22_X1 U11759 ( .A1(n11181), .A2(n11184), .B1(n7634), .B2(n11180), .ZN(
        P1_U3534) );
  INV_X1 U11760 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U11761 ( .A1(n11185), .A2(n11184), .B1(n11183), .B2(n11182), .ZN(
        P1_U3489) );
  INV_X1 U11762 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U11763 ( .A1(n11195), .A2(n11187), .B1(n11186), .B2(n11192), .ZN(
        P2_U3429) );
  INV_X1 U11764 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U11765 ( .A1(n11195), .A2(n11189), .B1(n11188), .B2(n11192), .ZN(
        P2_U3432) );
  INV_X1 U11766 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U11767 ( .A1(n11195), .A2(n11191), .B1(n11190), .B2(n11192), .ZN(
        P2_U3435) );
  INV_X1 U11768 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U11769 ( .A1(n11195), .A2(n11194), .B1(n11193), .B2(n11192), .ZN(
        P2_U3438) );
  XNOR2_X1 U11770 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U5202 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7131) );
  INV_X1 U5198 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10288) );
  CLKBUF_X1 U5209 ( .A(n7532), .Z(n5140) );
  INV_X1 U5357 ( .A(n7539), .ZN(n8711) );
endmodule

