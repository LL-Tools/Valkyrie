

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4399, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372;

  INV_X4 U4904 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4906 ( .A(n5147), .ZN(n6648) );
  NAND2_X1 U4908 ( .A1(n5595), .A2(n5578), .ZN(n6792) );
  CLKBUF_X2 U4909 ( .A(n5135), .Z(n5508) );
  NAND3_X1 U4910 ( .A1(n5764), .A2(n5763), .A3(n5762), .ZN(n10246) );
  AND2_X1 U4911 ( .A1(n5105), .A2(n7994), .ZN(n5107) );
  CLKBUF_X3 U4912 ( .A(n6214), .Z(n6387) );
  OR2_X1 U4913 ( .A1(n6432), .A2(n8318), .ZN(n8604) );
  AND2_X1 U4914 ( .A1(n4409), .A2(n8320), .ZN(n4410) );
  INV_X1 U4915 ( .A(n6687), .ZN(n6982) );
  INV_X1 U4916 ( .A(n5745), .ZN(n6051) );
  NAND2_X1 U4917 ( .A1(n5697), .A2(n5696), .ZN(n5746) );
  INV_X1 U4918 ( .A(n5200), .ZN(n5234) );
  AND2_X1 U4919 ( .A1(n5401), .A2(n8088), .ZN(n9125) );
  INV_X1 U4920 ( .A(n6763), .ZN(n4401) );
  INV_X1 U4921 ( .A(n5723), .ZN(n8142) );
  INV_X1 U4922 ( .A(n9989), .ZN(n10019) );
  XNOR2_X1 U4923 ( .A(n5565), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5653) );
  INV_X1 U4924 ( .A(n5696), .ZN(n5698) );
  NAND2_X1 U4925 ( .A1(n6497), .A2(n5043), .ZN(n4399) );
  NAND2_X1 U4926 ( .A1(n6497), .A2(n5043), .ZN(n5753) );
  NAND2_X2 U4927 ( .A1(n9453), .A2(n5467), .ZN(n9456) );
  NAND2_X2 U4928 ( .A1(n9474), .A2(n9471), .ZN(n9453) );
  OAI21_X2 U4929 ( .B1(n7060), .B2(n4736), .A(n4734), .ZN(n7288) );
  OAI21_X2 U4930 ( .B1(n7951), .B2(n7947), .A(n7948), .ZN(n8034) );
  XNOR2_X2 U4931 ( .A(n5692), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5697) );
  NAND2_X2 U4932 ( .A1(n7989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5692) );
  XNOR2_X2 U4933 ( .A(n4944), .B(n4943), .ZN(n5156) );
  XNOR2_X2 U4934 ( .A(n5123), .B(n9211), .ZN(n5607) );
  NAND4_X2 U4935 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n9211)
         );
  NAND2_X1 U4936 ( .A1(n5654), .A2(n5653), .ZN(n6191) );
  NAND2_X1 U4937 ( .A1(n5655), .A2(n6415), .ZN(n6192) );
  XNOR2_X2 U4938 ( .A(n5705), .B(n5704), .ZN(n6073) );
  NAND2_X1 U4939 ( .A1(n6344), .A2(n6343), .ZN(n8369) );
  AND2_X1 U4940 ( .A1(n8315), .A2(n4802), .ZN(n4409) );
  NAND2_X1 U4941 ( .A1(n5485), .A2(n5484), .ZN(n9430) );
  OR2_X1 U4942 ( .A1(n6132), .A2(n8632), .ZN(n6133) );
  BUF_X1 U4943 ( .A(n10297), .Z(n4403) );
  INV_X1 U4944 ( .A(n7436), .ZN(n10023) );
  AND2_X1 U4945 ( .A1(n8203), .A2(n8217), .ZN(n8150) );
  INV_X2 U4946 ( .A(n6196), .ZN(n6395) );
  INV_X1 U4947 ( .A(n10246), .ZN(n6695) );
  INV_X1 U4948 ( .A(n7645), .ZN(n7186) );
  AND4_X1 U4949 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n6949)
         );
  AND2_X2 U4950 ( .A1(n8094), .A2(n5698), .ZN(n5744) );
  INV_X1 U4951 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5549) );
  AND2_X1 U4952 ( .A1(n4589), .A2(n4588), .ZN(n4587) );
  AND2_X1 U4953 ( .A1(n8406), .A2(n8405), .ZN(n9566) );
  AND2_X1 U4954 ( .A1(n9560), .A2(n9561), .ZN(n4760) );
  AOI21_X1 U4955 ( .B1(n4824), .B2(n8184), .A(n4822), .ZN(n4911) );
  NAND2_X1 U4956 ( .A1(n6466), .A2(n6465), .ZN(n8383) );
  OAI21_X1 U4957 ( .B1(n9128), .B2(n4469), .A(n4528), .ZN(n4524) );
  AND2_X1 U4958 ( .A1(n8399), .A2(n8398), .ZN(n9425) );
  AND2_X1 U4959 ( .A1(n4637), .A2(n4457), .ZN(n8425) );
  INV_X1 U4960 ( .A(n9036), .ZN(n8931) );
  NAND2_X1 U4961 ( .A1(n8146), .A2(n8145), .ZN(n8598) );
  NAND2_X1 U4962 ( .A1(n8342), .A2(n8181), .ZN(n8335) );
  OR2_X1 U4963 ( .A1(n8099), .A2(n6167), .ZN(n8342) );
  NAND2_X1 U4964 ( .A1(n5529), .A2(n5528), .ZN(n9558) );
  AOI21_X1 U4965 ( .B1(n8091), .B2(n8142), .A(n7999), .ZN(n8180) );
  XNOR2_X1 U4966 ( .A(n6658), .B(n6657), .ZN(n8143) );
  OAI22_X1 U4967 ( .A1(n6654), .A2(n6653), .B1(SI_30_), .B2(n6652), .ZN(n6658)
         );
  AOI22_X1 U4968 ( .A1(n8694), .A2(n8693), .B1(n8681), .B2(n8760), .ZN(n8680)
         );
  AND2_X1 U4969 ( .A1(n6133), .A2(n8311), .ZN(n8315) );
  NAND2_X1 U4970 ( .A1(n7689), .A2(n7688), .ZN(n7763) );
  AND2_X1 U4971 ( .A1(n8117), .A2(n8643), .ZN(n8118) );
  NAND2_X1 U4972 ( .A1(n6001), .A2(n6000), .ZN(n8469) );
  NAND2_X1 U4973 ( .A1(n7733), .A2(n6127), .ZN(n7806) );
  AND2_X1 U4974 ( .A1(n4901), .A2(n5892), .ZN(n4900) );
  OR2_X1 U4975 ( .A1(n4902), .A2(n5881), .ZN(n4901) );
  XNOR2_X1 U4976 ( .A(n5443), .B(n5442), .ZN(n7394) );
  OAI21_X1 U4977 ( .B1(n5434), .B2(n5433), .A(n5037), .ZN(n5443) );
  OR2_X1 U4978 ( .A1(n7890), .A2(n8512), .ZN(n5919) );
  NAND2_X1 U4979 ( .A1(n5032), .A2(n5031), .ZN(n5434) );
  AOI21_X1 U4980 ( .B1(n6714), .B2(n7193), .A(n4670), .ZN(n4668) );
  OR2_X1 U4981 ( .A1(n7476), .A2(n7827), .ZN(n8253) );
  AND2_X1 U4982 ( .A1(n5849), .A2(n5848), .ZN(n10291) );
  NAND2_X1 U4983 ( .A1(n5274), .A2(n5273), .ZN(n10008) );
  AOI21_X1 U4984 ( .B1(n5395), .B2(n5023), .A(n4909), .ZN(n5027) );
  NAND2_X1 U4985 ( .A1(n5261), .A2(n5260), .ZN(n7759) );
  NAND2_X1 U4986 ( .A1(n5195), .A2(n5194), .ZN(n6810) );
  AND3_X1 U4987 ( .A1(n5833), .A2(n5832), .A3(n5831), .ZN(n10286) );
  XOR2_X1 U4988 ( .A(n6218), .B(n6220), .Z(n7146) );
  INV_X1 U4989 ( .A(n7639), .ZN(n10073) );
  OAI21_X1 U4990 ( .B1(n5253), .B2(n4765), .A(n4763), .ZN(n5349) );
  OR2_X1 U4991 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  NAND2_X1 U4992 ( .A1(n4614), .A2(n4617), .ZN(n5195) );
  OAI211_X1 U4993 ( .C1(n6794), .C2(n9240), .A(n5248), .B(n5247), .ZN(n7436)
         );
  AND2_X1 U4994 ( .A1(n5394), .A2(n5017), .ZN(n5023) );
  INV_X2 U4995 ( .A(n6252), .ZN(n6392) );
  INV_X1 U4996 ( .A(n6199), .ZN(n7609) );
  NAND2_X1 U4997 ( .A1(n4577), .A2(n4953), .ZN(n5246) );
  AND2_X1 U4998 ( .A1(n5379), .A2(n5018), .ZN(n5394) );
  AND2_X1 U4999 ( .A1(n5366), .A2(n5007), .ZN(n5379) );
  NAND2_X1 U5000 ( .A1(n4950), .A2(n4949), .ZN(n5189) );
  AND2_X1 U5001 ( .A1(n5001), .A2(n5000), .ZN(n5366) );
  OR2_X1 U5002 ( .A1(n5352), .A2(n5350), .ZN(n5001) );
  AND3_X1 U5003 ( .A1(n4828), .A2(n4449), .A3(n5737), .ZN(n6948) );
  NAND4_X1 U5004 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(n9209)
         );
  OAI211_X1 U5005 ( .C1(n6497), .C2(n6762), .A(n5769), .B(n5768), .ZN(n10265)
         );
  AND4_X1 U5006 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n7160)
         );
  AND2_X1 U5007 ( .A1(n4998), .A2(n4997), .ZN(n5350) );
  OR2_X1 U5008 ( .A1(n5340), .A2(n5118), .ZN(n5120) );
  OR2_X1 U5009 ( .A1(n4994), .A2(n5332), .ZN(n4998) );
  NAND2_X2 U5010 ( .A1(n6794), .A2(n6763), .ZN(n6649) );
  INV_X1 U5011 ( .A(n8184), .ZN(n8196) );
  OR2_X1 U5012 ( .A1(n4993), .A2(n4992), .ZN(n5332) );
  AND2_X2 U5013 ( .A1(n5106), .A2(n5107), .ZN(n5489) );
  AND2_X1 U5014 ( .A1(n5316), .A2(n4991), .ZN(n4992) );
  INV_X1 U5015 ( .A(n6531), .ZN(n6074) );
  XNOR2_X1 U5016 ( .A(n6061), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8184) );
  XNOR2_X1 U5017 ( .A(n5550), .B(n5549), .ZN(n6415) );
  XNOR2_X1 U5018 ( .A(n4503), .B(P2_IR_REG_27__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U5019 ( .A1(n5548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U5020 ( .A1(n4504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U5021 ( .A1(n5703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5705) );
  NOR2_X1 U5022 ( .A1(n5544), .A2(n5543), .ZN(n5547) );
  NAND2_X1 U5023 ( .A1(n5083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U5024 ( .A(n4939), .B(SI_2_), .ZN(n5145) );
  AND2_X1 U5025 ( .A1(n5702), .A2(n5704), .ZN(n5693) );
  INV_X2 U5026 ( .A(n6763), .ZN(n4402) );
  AND2_X1 U5027 ( .A1(n5707), .A2(n5706), .ZN(n5702) );
  NOR2_X1 U5028 ( .A1(n4641), .A2(n4640), .ZN(n4639) );
  AND2_X1 U5029 ( .A1(n6087), .A2(n5688), .ZN(n5706) );
  AND3_X1 U5030 ( .A1(n5680), .A2(n5679), .A3(n5678), .ZN(n5682) );
  AND3_X1 U5031 ( .A1(n4712), .A2(n5140), .A3(n5070), .ZN(n4708) );
  NOR2_X1 U5032 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n4424), .ZN(n5081) );
  AND3_X1 U5033 ( .A1(n5675), .A2(n5674), .A3(n5673), .ZN(n5679) );
  NAND4_X1 U5034 ( .A1(n5257), .A2(n5228), .A3(n4506), .A4(n4505), .ZN(n4710)
         );
  NOR2_X1 U5035 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4712) );
  INV_X1 U5036 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5228) );
  INV_X1 U5037 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5196) );
  NOR2_X1 U5038 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4643) );
  INV_X1 U5039 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5257) );
  INV_X1 U5040 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4505) );
  INV_X1 U5041 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4506) );
  INV_X1 U5042 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5069) );
  INV_X4 U5043 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5044 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4645) );
  INV_X1 U5045 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5399) );
  INV_X1 U5046 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5751) );
  INV_X1 U5047 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5542) );
  AOI211_X2 U5048 ( .C1(n9570), .C2(n6629), .A(n9569), .B(n9568), .ZN(n9635)
         );
  INV_X2 U5049 ( .A(n7133), .ZN(n5123) );
  NOR2_X2 U5050 ( .A1(n5927), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5929) );
  OR2_X2 U5051 ( .A1(n5911), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5927) );
  INV_X2 U5052 ( .A(n8508), .ZN(n8643) );
  NAND2_X4 U5053 ( .A1(n6683), .A2(n6682), .ZN(n6685) );
  NAND2_X1 U5054 ( .A1(n4966), .A2(n4965), .ZN(n4969) );
  NOR2_X1 U5055 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5685) );
  NOR2_X1 U5056 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5684) );
  NOR2_X1 U5057 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5683) );
  NOR2_X1 U5058 ( .A1(n4912), .A2(n4725), .ZN(n4724) );
  INV_X1 U5059 ( .A(n4726), .ZN(n4725) );
  NAND2_X1 U5060 ( .A1(n5349), .A2(n4985), .ZN(n5395) );
  XNOR2_X1 U5061 ( .A(n4999), .B(SI_16_), .ZN(n5352) );
  NAND2_X1 U5062 ( .A1(n4990), .A2(n4989), .ZN(n5318) );
  OR2_X1 U5063 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  AND2_X1 U5064 ( .A1(n8391), .A2(n4573), .ZN(n9401) );
  NOR2_X1 U5065 ( .A1(n9558), .A2(n4574), .ZN(n4573) );
  INV_X1 U5066 ( .A(n4575), .ZN(n4574) );
  NAND2_X1 U5067 ( .A1(n6794), .A2(n5043), .ZN(n5147) );
  NAND2_X2 U5068 ( .A1(n5554), .A2(n5558), .ZN(n6794) );
  NAND2_X1 U5069 ( .A1(n8947), .A2(n9141), .ZN(n4543) );
  OAI21_X1 U5070 ( .B1(n4537), .B2(n4539), .A(n9044), .ZN(n4534) );
  INV_X1 U5071 ( .A(n4543), .ZN(n4539) );
  OAI21_X1 U5072 ( .B1(n9141), .B2(n4541), .A(n8947), .ZN(n4535) );
  NAND2_X1 U5073 ( .A1(n4440), .A2(n8354), .ZN(n4599) );
  NAND2_X1 U5074 ( .A1(n4602), .A2(n8349), .ZN(n4601) );
  NAND2_X1 U5075 ( .A1(n8339), .A2(n4603), .ZN(n4602) );
  NOR2_X1 U5076 ( .A1(n7961), .A2(n7965), .ZN(n8272) );
  NAND2_X1 U5077 ( .A1(n4621), .A2(n4960), .ZN(n4620) );
  INV_X1 U5078 ( .A(n5214), .ZN(n4621) );
  AOI21_X1 U5079 ( .B1(n4663), .B2(n4664), .A(n8449), .ZN(n4661) );
  OAI21_X1 U5080 ( .B1(n8178), .B2(n8177), .A(n8183), .ZN(n4825) );
  OR2_X1 U5081 ( .A1(n8185), .A2(n8184), .ZN(n4823) );
  NOR2_X1 U5082 ( .A1(n4808), .A2(n4809), .ZN(n4807) );
  INV_X1 U5083 ( .A(n8202), .ZN(n4809) );
  OR2_X1 U5084 ( .A1(n6431), .A2(n6045), .ZN(n6039) );
  AND2_X1 U5085 ( .A1(n6042), .A2(n6041), .ZN(n6433) );
  OR2_X1 U5086 ( .A1(n8803), .A2(n8642), .ZN(n8309) );
  OR2_X1 U5087 ( .A1(n7961), .A2(n8511), .ZN(n7948) );
  NOR2_X1 U5088 ( .A1(n6272), .A2(n6271), .ZN(n6273) );
  OR2_X1 U5089 ( .A1(n6369), .A2(n8134), .ZN(n6382) );
  NAND2_X1 U5090 ( .A1(n4421), .A2(n4513), .ZN(n4512) );
  NOR2_X1 U5091 ( .A1(n4519), .A2(n4516), .ZN(n4513) );
  NOR2_X1 U5092 ( .A1(n9020), .A2(n9092), .ZN(n4516) );
  NAND2_X1 U5093 ( .A1(n4421), .A2(n4515), .ZN(n4514) );
  NOR2_X1 U5094 ( .A1(n9101), .A2(n9125), .ZN(n4515) );
  NAND2_X1 U5095 ( .A1(n6647), .A2(n6646), .ZN(n6654) );
  NAND2_X1 U5096 ( .A1(n5483), .A2(n5059), .ZN(n5501) );
  NAND2_X1 U5097 ( .A1(n5027), .A2(n5026), .ZN(n5426) );
  NOR2_X1 U5098 ( .A1(n4908), .A2(n5025), .ZN(n5026) );
  INV_X1 U5099 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5071) );
  INV_X1 U5100 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4859) );
  INV_X1 U5101 ( .A(n4710), .ZN(n4707) );
  INV_X1 U5102 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5070) );
  AND2_X1 U5103 ( .A1(n4969), .A2(n4968), .ZN(n5192) );
  AND2_X1 U5104 ( .A1(n5140), .A2(n5069), .ZN(n5183) );
  INV_X1 U5105 ( .A(n4663), .ZN(n4662) );
  NOR2_X1 U5106 ( .A1(n6875), .A2(n6876), .ZN(n6874) );
  NOR2_X1 U5107 ( .A1(n8592), .A2(n8591), .ZN(n8590) );
  OAI22_X1 U5108 ( .A1(n8706), .A2(n5957), .B1(n8696), .B2(n5956), .ZN(n8694)
         );
  AND2_X1 U5109 ( .A1(n8330), .A2(n8331), .ZN(n8327) );
  NAND2_X1 U5110 ( .A1(n4800), .A2(n4798), .ZN(n8602) );
  INV_X1 U5111 ( .A(n8321), .ZN(n4799) );
  AND2_X1 U5112 ( .A1(n8276), .A2(n8283), .ZN(n8705) );
  NOR2_X1 U5113 ( .A1(n4797), .A2(n4796), .ZN(n4795) );
  INV_X1 U5114 ( .A(n8281), .ZN(n4796) );
  INV_X1 U5115 ( .A(n8287), .ZN(n4797) );
  INV_X1 U5116 ( .A(n5753), .ZN(n5962) );
  AND2_X1 U5117 ( .A1(n6076), .A2(n8354), .ZN(n10248) );
  NAND2_X1 U5118 ( .A1(n5694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5695) );
  CLKBUF_X1 U5119 ( .A(n5719), .Z(n5941) );
  AND2_X1 U5120 ( .A1(n6265), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U5121 ( .A1(n4724), .A2(n4722), .ZN(n4721) );
  INV_X1 U5122 ( .A(n4724), .ZN(n4723) );
  NAND2_X1 U5123 ( .A1(n8369), .A2(n6355), .ZN(n6466) );
  NAND2_X1 U5124 ( .A1(n6963), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4477) );
  AND2_X1 U5125 ( .A1(n4488), .A2(n4487), .ZN(n9306) );
  NAND2_X1 U5126 ( .A1(n9302), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4487) );
  INV_X1 U5127 ( .A(n9632), .ZN(n9405) );
  NAND2_X1 U5128 ( .A1(n8391), .A2(n4575), .ZN(n6627) );
  NOR2_X1 U5129 ( .A1(n9444), .A2(n9430), .ZN(n8391) );
  NAND2_X1 U5130 ( .A1(n4775), .A2(n4779), .ZN(n9419) );
  NAND2_X1 U5131 ( .A1(n7940), .A2(n5365), .ZN(n7901) );
  INV_X1 U5132 ( .A(n10002), .ZN(n9980) );
  INV_X1 U5133 ( .A(n10010), .ZN(n9968) );
  OR2_X1 U5134 ( .A1(n6619), .A2(n6622), .ZN(n6620) );
  OR2_X1 U5135 ( .A1(n7927), .A2(n5147), .ZN(n5529) );
  NAND2_X1 U5136 ( .A1(n5356), .A2(n5355), .ZN(n7908) );
  NAND2_X1 U5137 ( .A1(n5323), .A2(n5322), .ZN(n7794) );
  NAND2_X1 U5138 ( .A1(n5524), .A2(SI_29_), .ZN(n6647) );
  XNOR2_X1 U5139 ( .A(n5569), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U5140 ( .A1(n5573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U5141 ( .A1(n5545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5546) );
  AND2_X1 U5142 ( .A1(n5397), .A2(n5396), .ZN(n5411) );
  INV_X1 U5143 ( .A(n8507), .ZN(n8459) );
  NOR2_X1 U5144 ( .A1(n7069), .A2(n7070), .ZN(n7068) );
  NAND2_X1 U5145 ( .A1(n10222), .A2(n10223), .ZN(n10221) );
  NAND2_X1 U5146 ( .A1(n4694), .A2(n4693), .ZN(n8578) );
  OR2_X1 U5147 ( .A1(n10230), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U5148 ( .A1(n4696), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5149 ( .A1(n5089), .A2(n5088), .ZN(n9026) );
  NAND2_X1 U5150 ( .A1(n4480), .A2(n5654), .ZN(n4479) );
  NAND2_X1 U5151 ( .A1(n4482), .A2(n4481), .ZN(n4480) );
  NAND2_X1 U5152 ( .A1(n9398), .A2(n9961), .ZN(n4481) );
  NAND2_X1 U5153 ( .A1(n9396), .A2(n9397), .ZN(n4482) );
  AOI21_X1 U5154 ( .B1(n9193), .B2(n9985), .A(n5560), .ZN(n5561) );
  INV_X1 U5155 ( .A(n4532), .ZN(n4531) );
  OAI21_X1 U5156 ( .B1(n4535), .B2(n4536), .A(n8944), .ZN(n4532) );
  INV_X1 U5157 ( .A(n4541), .ZN(n4536) );
  OAI21_X1 U5158 ( .B1(n4543), .B2(n4538), .A(n8949), .ZN(n4537) );
  NOR2_X1 U5159 ( .A1(n4896), .A2(n6007), .ZN(n4895) );
  INV_X1 U5160 ( .A(n4899), .ZN(n4896) );
  INV_X1 U5161 ( .A(n9427), .ZN(n9029) );
  NAND2_X1 U5162 ( .A1(n4792), .A2(n5498), .ZN(n4791) );
  NAND2_X1 U5163 ( .A1(n4782), .A2(n5647), .ZN(n4781) );
  INV_X1 U5164 ( .A(n9421), .ZN(n5499) );
  AOI21_X1 U5165 ( .B1(n8473), .B2(n4667), .A(n4918), .ZN(n4663) );
  XNOR2_X1 U5166 ( .A(n6685), .B(n10265), .ZN(n6698) );
  INV_X1 U5167 ( .A(n7839), .ZN(n4648) );
  OAI21_X1 U5168 ( .B1(n4652), .B2(n8021), .A(n8020), .ZN(n4651) );
  OR3_X1 U5169 ( .A1(n8335), .A2(n8334), .A3(n8333), .ZN(n8344) );
  NAND2_X1 U5170 ( .A1(n4601), .A2(n4599), .ZN(n4598) );
  INV_X1 U5171 ( .A(n4596), .ZN(n4595) );
  OAI22_X1 U5172 ( .A1(n4601), .A2(n4415), .B1(n4599), .B2(n4437), .ZN(n4596)
         );
  AND2_X1 U5173 ( .A1(n6508), .A2(n4681), .ZN(n4676) );
  INV_X1 U5174 ( .A(n6510), .ZN(n4681) );
  AND2_X1 U5175 ( .A1(n4678), .A2(n4677), .ZN(n6513) );
  NOR2_X1 U5176 ( .A1(n4680), .A2(n6511), .ZN(n4677) );
  AOI21_X1 U5177 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6800), .A(n7335), .ZN(
        n6514) );
  NAND2_X1 U5178 ( .A1(n4853), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4852) );
  AND2_X1 U5179 ( .A1(n10140), .A2(n4427), .ZN(n4850) );
  AND2_X1 U5180 ( .A1(n8572), .A2(n6551), .ZN(n6552) );
  NAND2_X1 U5181 ( .A1(n5850), .A2(n4875), .ZN(n4874) );
  INV_X1 U5182 ( .A(n5835), .ZN(n4875) );
  AND2_X1 U5183 ( .A1(n4403), .A2(n8516), .ZN(n8235) );
  INV_X1 U5184 ( .A(n5796), .ZN(n4880) );
  INV_X1 U5185 ( .A(n5808), .ZN(n4877) );
  NAND2_X1 U5186 ( .A1(n8204), .A2(n8202), .ZN(n6120) );
  AND2_X1 U5187 ( .A1(n8786), .A2(n8459), .ZN(n8147) );
  NAND2_X1 U5188 ( .A1(n4893), .A2(n4892), .ZN(n4891) );
  INV_X1 U5189 ( .A(n4895), .ZN(n4892) );
  OR2_X1 U5190 ( .A1(n8786), .A2(n8459), .ZN(n8324) );
  OR2_X1 U5191 ( .A1(n8809), .A2(n8111), .ZN(n8300) );
  OR2_X1 U5192 ( .A1(n7815), .A2(n8513), .ZN(n7805) );
  AND2_X1 U5193 ( .A1(n5686), .A2(n5942), .ZN(n6058) );
  INV_X1 U5194 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5944) );
  NAND3_X1 U5195 ( .A1(n4645), .A2(n5717), .A3(n5751), .ZN(n4640) );
  OR2_X1 U5196 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  INV_X1 U5197 ( .A(n6225), .ZN(n4740) );
  OAI21_X1 U5198 ( .B1(n9070), .B2(n4788), .A(n5651), .ZN(n4787) );
  NAND2_X1 U5199 ( .A1(n5650), .A2(n5649), .ZN(n4788) );
  AND2_X1 U5200 ( .A1(n4789), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U5201 ( .A1(n4779), .A2(n4778), .ZN(n4777) );
  NOR2_X1 U5202 ( .A1(n9070), .A2(n4790), .ZN(n4789) );
  INV_X1 U5203 ( .A(n4782), .ZN(n4778) );
  NAND2_X1 U5204 ( .A1(n4776), .A2(n4780), .ZN(n4773) );
  OR2_X1 U5205 ( .A1(n9564), .A2(n9029), .ZN(n9079) );
  OR2_X1 U5206 ( .A1(n9430), .A2(n9443), .ZN(n9078) );
  NOR2_X1 U5207 ( .A1(n5497), .A2(n4869), .ZN(n4868) );
  INV_X1 U5208 ( .A(n9081), .ZN(n4869) );
  OR2_X1 U5209 ( .A1(n9420), .A2(n5499), .ZN(n5497) );
  NOR2_X1 U5210 ( .A1(n9575), .A2(n5498), .ZN(n9420) );
  NOR2_X1 U5211 ( .A1(n9530), .A2(n9597), .ZN(n4572) );
  OAI21_X1 U5212 ( .B1(n8011), .B2(n4839), .A(n9546), .ZN(n4838) );
  OAI21_X1 U5213 ( .B1(n9054), .B2(n4833), .A(n9046), .ZN(n4831) );
  NAND2_X1 U5214 ( .A1(n4562), .A2(n10079), .ZN(n4565) );
  INV_X1 U5215 ( .A(n4567), .ZN(n4562) );
  AND2_X1 U5216 ( .A1(n7637), .A2(n10073), .ZN(n7583) );
  AND2_X1 U5217 ( .A1(n5523), .A2(n5522), .ZN(n6645) );
  NAND2_X1 U5218 ( .A1(n5501), .A2(n5500), .ZN(n5521) );
  NAND2_X1 U5219 ( .A1(n5481), .A2(n5480), .ZN(n5483) );
  NAND2_X1 U5220 ( .A1(n5049), .A2(n5048), .ZN(n5469) );
  NAND2_X1 U5221 ( .A1(n5028), .A2(n5425), .ZN(n5032) );
  OR2_X1 U5222 ( .A1(n5021), .A2(n5020), .ZN(n5396) );
  AOI21_X1 U5223 ( .B1(n4771), .B2(n4769), .A(n4768), .ZN(n4767) );
  INV_X1 U5224 ( .A(n4977), .ZN(n4768) );
  NOR2_X1 U5225 ( .A1(n5269), .A2(n4770), .ZN(n4769) );
  INV_X1 U5226 ( .A(n4972), .ZN(n4770) );
  INV_X1 U5227 ( .A(n5252), .ZN(n4771) );
  AOI21_X1 U5228 ( .B1(n4620), .B2(n4964), .A(n4618), .ZN(n4617) );
  INV_X1 U5229 ( .A(n5192), .ZN(n4618) );
  INV_X1 U5230 ( .A(n4620), .ZN(n4616) );
  NAND2_X1 U5231 ( .A1(n4964), .A2(n4963), .ZN(n5214) );
  NAND2_X1 U5232 ( .A1(n6088), .A2(n5706), .ZN(n4504) );
  NAND2_X1 U5233 ( .A1(n6948), .A2(n6979), .ZN(n8195) );
  NAND2_X1 U5234 ( .A1(n8473), .A2(n4665), .ZN(n4664) );
  INV_X1 U5235 ( .A(n8440), .ZN(n4665) );
  NOR2_X1 U5236 ( .A1(n7970), .A2(n4653), .ZN(n4652) );
  INV_X1 U5237 ( .A(n7967), .ZN(n4653) );
  NOR2_X1 U5238 ( .A1(n4659), .A2(n4656), .ZN(n4655) );
  OAI21_X1 U5239 ( .B1(n4658), .B2(n4656), .A(n4460), .ZN(n4654) );
  NAND2_X1 U5240 ( .A1(n4823), .A2(n8347), .ZN(n4822) );
  NAND2_X1 U5241 ( .A1(n4825), .A2(n4435), .ZN(n4824) );
  INV_X1 U5242 ( .A(n5914), .ZN(n6174) );
  NAND2_X1 U5243 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  NAND2_X1 U5244 ( .A1(n8361), .A2(n5736), .ZN(n4496) );
  OR2_X1 U5245 ( .A1(n8361), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4497) );
  OR2_X1 U5246 ( .A1(n6874), .A2(n4426), .ZN(n4829) );
  NAND2_X1 U5247 ( .A1(n6509), .A2(n6508), .ZN(n7076) );
  AOI21_X1 U5248 ( .B1(n7338), .B2(n7336), .A(n7337), .ZN(n7335) );
  OAI22_X1 U5249 ( .A1(n7276), .A2(n7277), .B1(n6589), .B2(n7283), .ZN(n7331)
         );
  NOR2_X1 U5250 ( .A1(n7327), .A2(n6543), .ZN(n6544) );
  AND2_X1 U5251 ( .A1(n6800), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U5252 ( .A1(n6544), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U5253 ( .A1(n4851), .A2(n4850), .ZN(n10139) );
  OR2_X1 U5254 ( .A1(n5893), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5894) );
  OR2_X1 U5255 ( .A1(n10195), .A2(n4691), .ZN(n4689) );
  OR2_X1 U5256 ( .A1(n10212), .A2(n10194), .ZN(n4691) );
  OR2_X1 U5257 ( .A1(n4422), .A2(n10212), .ZN(n4690) );
  OR2_X1 U5258 ( .A1(n10195), .A2(n10194), .ZN(n4692) );
  NAND2_X1 U5259 ( .A1(n10186), .A2(n6548), .ZN(n10204) );
  AOI21_X1 U5260 ( .B1(n10204), .B2(n10201), .A(n4840), .ZN(n6549) );
  NOR2_X1 U5261 ( .A1(n10202), .A2(n5913), .ZN(n4840) );
  OR2_X1 U5262 ( .A1(n8570), .A2(n8569), .ZN(n8572) );
  XNOR2_X1 U5263 ( .A(n6552), .B(n10218), .ZN(n10225) );
  XNOR2_X1 U5264 ( .A(n6525), .B(n7192), .ZN(n10230) );
  AND2_X1 U5265 ( .A1(n6011), .A2(n6010), .ZN(n6020) );
  AND2_X1 U5266 ( .A1(n6020), .A2(n8494), .ZN(n6032) );
  OR2_X1 U5267 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  AOI21_X1 U5268 ( .B1(n4886), .B2(n4889), .A(n4444), .ZN(n4884) );
  OR2_X1 U5269 ( .A1(n7714), .A2(n8516), .ZN(n5862) );
  NOR2_X1 U5270 ( .A1(n8235), .A2(n4820), .ZN(n4819) );
  INV_X1 U5271 ( .A(n8236), .ZN(n4820) );
  OR2_X1 U5272 ( .A1(n7418), .A2(n7421), .ZN(n4821) );
  AND4_X1 U5273 ( .A1(n5842), .A2(n5841), .A3(n5840), .A4(n5839), .ZN(n7451)
         );
  AND4_X1 U5274 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(n7827)
         );
  NAND2_X1 U5275 ( .A1(n7214), .A2(n5821), .ZN(n7320) );
  AND4_X1 U5276 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n7199)
         );
  NAND2_X1 U5277 ( .A1(n10242), .A2(n4807), .ZN(n4804) );
  NAND2_X1 U5278 ( .A1(n6919), .A2(n6979), .ZN(n6946) );
  NAND2_X1 U5279 ( .A1(n6030), .A2(n6029), .ZN(n8122) );
  NAND2_X1 U5280 ( .A1(n6173), .A2(n6184), .ZN(n6185) );
  NAND2_X1 U5281 ( .A1(n8325), .A2(n8324), .ZN(n8605) );
  NAND2_X1 U5282 ( .A1(n8312), .A2(n4803), .ZN(n4802) );
  INV_X1 U5283 ( .A(n8309), .ZN(n4803) );
  OR2_X1 U5284 ( .A1(n8803), .A2(n8671), .ZN(n5998) );
  NAND2_X1 U5285 ( .A1(n8815), .A2(n8697), .ZN(n8663) );
  AND2_X1 U5286 ( .A1(n5972), .A2(n5971), .ZN(n8108) );
  NAND2_X1 U5287 ( .A1(n8187), .A2(n8663), .ZN(n8679) );
  AND2_X1 U5288 ( .A1(n8286), .A2(n8705), .ZN(n4793) );
  NOR2_X1 U5289 ( .A1(n8034), .A2(n8033), .ZN(n8037) );
  AND2_X1 U5290 ( .A1(n8266), .A2(n8273), .ZN(n4814) );
  NAND2_X1 U5291 ( .A1(n7881), .A2(n8269), .ZN(n4815) );
  INV_X1 U5292 ( .A(n8710), .ZN(n10247) );
  AND3_X1 U5293 ( .A1(n5794), .A2(n5793), .A3(n5792), .ZN(n10277) );
  XNOR2_X1 U5294 ( .A(n6090), .B(P2_B_REG_SCAN_IN), .ZN(n6089) );
  AND2_X1 U5295 ( .A1(n5681), .A2(n9796), .ZN(n4882) );
  OR2_X1 U5296 ( .A1(n5804), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5817) );
  AND2_X1 U5297 ( .A1(n4644), .A2(n5751), .ZN(n5777) );
  AND2_X1 U5298 ( .A1(n4642), .A2(n4645), .ZN(n4644) );
  NOR2_X1 U5299 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4642) );
  INV_X1 U5300 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9796) );
  INV_X1 U5301 ( .A(n5725), .ZN(n4843) );
  NAND2_X1 U5302 ( .A1(n6310), .A2(n4744), .ZN(n4743) );
  OAI21_X1 U5303 ( .B1(n7288), .B2(n7291), .A(n7289), .ZN(n7383) );
  NOR2_X1 U5304 ( .A1(n5147), .A2(n6764), .ZN(n4507) );
  OAI22_X1 U5305 ( .A1(n6649), .A2(n4929), .B1(n6794), .B2(n9219), .ZN(n4508)
         );
  OAI22_X1 U5306 ( .A1(n7135), .A2(n6253), .B1(n6213), .B2(n8082), .ZN(n6206)
         );
  NAND2_X1 U5307 ( .A1(n5093), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5429) );
  INV_X1 U5308 ( .A(n5420), .ZN(n5093) );
  NAND2_X1 U5309 ( .A1(n4719), .A2(n4717), .ZN(n7777) );
  AOI21_X1 U5310 ( .B1(n4720), .B2(n4723), .A(n4718), .ZN(n4717) );
  INV_X1 U5311 ( .A(n7779), .ZN(n4718) );
  NAND2_X1 U5312 ( .A1(n5096), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U5313 ( .A1(n6214), .A2(n7645), .ZN(n6216) );
  OR2_X1 U5314 ( .A1(n6383), .A2(n6467), .ZN(n6482) );
  NAND2_X1 U5315 ( .A1(n6466), .A2(n6378), .ZN(n6484) );
  AND2_X1 U5316 ( .A1(n8382), .A2(n6382), .ZN(n6467) );
  NAND2_X1 U5317 ( .A1(n4728), .A2(n6290), .ZN(n4729) );
  INV_X1 U5318 ( .A(n5489), .ZN(n5530) );
  AOI21_X1 U5319 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6848), .A(n9951), .ZN(
        n9232) );
  AOI21_X1 U5320 ( .B1(n6842), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6907), .ZN(
        n6845) );
  NAND2_X1 U5321 ( .A1(n4474), .A2(n4472), .ZN(n4476) );
  NOR2_X1 U5322 ( .A1(n9244), .A2(n4473), .ZN(n4472) );
  NAND2_X1 U5323 ( .A1(n6845), .A2(n4477), .ZN(n4474) );
  AND2_X1 U5324 ( .A1(n6844), .A2(n4477), .ZN(n4473) );
  OR2_X1 U5325 ( .A1(n6845), .A2(n6844), .ZN(n4478) );
  NAND2_X1 U5326 ( .A1(n7490), .A2(n7491), .ZN(n7492) );
  OR2_X1 U5327 ( .A1(n7494), .A2(n7495), .ZN(n4488) );
  OR2_X1 U5328 ( .A1(n9306), .A2(n9305), .ZN(n9314) );
  AND2_X1 U5329 ( .A1(n9079), .A2(n9092), .ZN(n9070) );
  NOR2_X1 U5330 ( .A1(n9492), .A2(n9588), .ZN(n9477) );
  NAND2_X1 U5331 ( .A1(n5645), .A2(n5644), .ZN(n9451) );
  AOI21_X1 U5332 ( .B1(n5642), .B2(n4748), .A(n4747), .ZN(n4746) );
  AND2_X1 U5333 ( .A1(n9538), .A2(n9541), .ZN(n9539) );
  AND2_X1 U5334 ( .A1(n9171), .A2(n9175), .ZN(n9546) );
  NAND2_X1 U5335 ( .A1(n8010), .A2(n8011), .ZN(n8009) );
  AND2_X1 U5336 ( .A1(n5632), .A2(n9165), .ZN(n4854) );
  OR2_X1 U5337 ( .A1(n7908), .A2(n8877), .ZN(n9165) );
  OR2_X1 U5338 ( .A1(n9970), .A2(n9969), .ZN(n9971) );
  NAND2_X1 U5339 ( .A1(n7459), .A2(n9054), .ZN(n7458) );
  AOI22_X1 U5340 ( .A1(n5612), .A2(n7245), .B1(n5611), .B2(n9052), .ZN(n7432)
         );
  INV_X1 U5341 ( .A(n6625), .ZN(n4846) );
  AND2_X1 U5342 ( .A1(n6628), .A2(n6627), .ZN(n9410) );
  NAND2_X1 U5343 ( .A1(n5339), .A2(n5338), .ZN(n9623) );
  AND2_X1 U5344 ( .A1(n5551), .A2(n8930), .ZN(n10002) );
  NOR2_X1 U5345 ( .A1(n5287), .A2(n4857), .ZN(n4855) );
  NAND2_X1 U5346 ( .A1(n4858), .A2(n5101), .ZN(n4857) );
  XNOR2_X1 U5347 ( .A(n6654), .B(n6653), .ZN(n8091) );
  XNOR2_X1 U5348 ( .A(n6645), .B(n6643), .ZN(n5524) );
  NAND2_X1 U5349 ( .A1(n4445), .A2(n4559), .ZN(n5083) );
  NOR2_X1 U5350 ( .A1(n5287), .A2(n4856), .ZN(n4559) );
  INV_X1 U5351 ( .A(n5083), .ZN(n5085) );
  NOR2_X1 U5352 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5084) );
  NOR2_X1 U5353 ( .A1(n5287), .A2(n4553), .ZN(n4551) );
  NAND2_X1 U5354 ( .A1(n5081), .A2(n4858), .ZN(n4553) );
  NAND2_X1 U5355 ( .A1(n5568), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5571) );
  XNOR2_X1 U5356 ( .A(n5469), .B(n5468), .ZN(n7515) );
  XNOR2_X1 U5357 ( .A(n5383), .B(n5382), .ZN(n7116) );
  NAND2_X1 U5358 ( .A1(n5381), .A2(n5380), .ZN(n5383) );
  XNOR2_X1 U5359 ( .A(n4927), .B(n5367), .ZN(n7153) );
  XNOR2_X1 U5360 ( .A(n5353), .B(n5352), .ZN(n7053) );
  XNOR2_X1 U5361 ( .A(n5336), .B(n5335), .ZN(n7055) );
  AOI21_X1 U5362 ( .B1(n5349), .B2(n5334), .A(n5333), .ZN(n5336) );
  INV_X1 U5363 ( .A(n5332), .ZN(n5333) );
  XNOR2_X1 U5364 ( .A(n5319), .B(n5318), .ZN(n7111) );
  AOI21_X1 U5365 ( .B1(n4763), .B2(n4765), .A(n5301), .ZN(n4762) );
  CLKBUF_X1 U5366 ( .A(n5287), .Z(n5288) );
  NAND2_X1 U5367 ( .A1(n4952), .A2(SI_5_), .ZN(n4953) );
  AND2_X1 U5368 ( .A1(n5187), .A2(n5186), .ZN(n6963) );
  OAI21_X1 U5369 ( .B1(n8490), .B2(n4635), .A(n4633), .ZN(n4638) );
  AOI21_X1 U5370 ( .B1(n4636), .B2(n4634), .A(n8124), .ZN(n4633) );
  INV_X1 U5371 ( .A(n4636), .ZN(n4635) );
  INV_X1 U5372 ( .A(n8491), .ZN(n4634) );
  AND4_X1 U5373 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n8709)
         );
  NAND2_X1 U5374 ( .A1(n4495), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6826) );
  XNOR2_X1 U5375 ( .A(n4829), .B(n6770), .ZN(n6992) );
  NAND2_X1 U5376 ( .A1(n6993), .A2(n4499), .ZN(n7069) );
  OR2_X1 U5377 ( .A1(n6585), .A2(n6997), .ZN(n4499) );
  NOR2_X1 U5378 ( .A1(n7328), .A2(n7329), .ZN(n7327) );
  NAND2_X1 U5379 ( .A1(n8563), .A2(n6602), .ZN(n10222) );
  OAI21_X1 U5380 ( .B1(n8590), .B2(n4433), .A(n10209), .ZN(n4864) );
  NOR2_X1 U5381 ( .A1(n8593), .A2(n4862), .ZN(n4861) );
  NOR2_X1 U5382 ( .A1(n4863), .A2(n8585), .ZN(n4862) );
  NOR2_X1 U5383 ( .A1(n8578), .A2(n6528), .ZN(n6529) );
  OAI211_X1 U5384 ( .C1(n6608), .C2(n10127), .A(n4502), .B(n4501), .ZN(n4500)
         );
  INV_X1 U5385 ( .A(n6609), .ZN(n4501) );
  NAND2_X1 U5386 ( .A1(n10219), .A2(n6610), .ZN(n4502) );
  OAI21_X1 U5387 ( .B1(n7927), .B2(n5723), .A(n6166), .ZN(n8099) );
  NAND2_X1 U5388 ( .A1(n5964), .A2(n5963), .ZN(n8760) );
  NAND2_X1 U5389 ( .A1(n5884), .A2(n5883), .ZN(n10313) );
  INV_X1 U5390 ( .A(n8747), .ZN(n8767) );
  XNOR2_X1 U5391 ( .A(n6170), .B(n8171), .ZN(n8784) );
  NAND2_X1 U5392 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  NAND2_X1 U5393 ( .A1(n8607), .A2(n10248), .ZN(n6077) );
  OAI21_X1 U5394 ( .B1(n6439), .B2(n10252), .A(n6438), .ZN(n6613) );
  NOR2_X1 U5395 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NOR2_X1 U5396 ( .A1(n8459), .A2(n8719), .ZN(n6436) );
  NAND2_X1 U5397 ( .A1(n6091), .A2(n6090), .ZN(n6786) );
  NAND2_X1 U5398 ( .A1(n5458), .A2(n5457), .ZN(n9464) );
  INV_X1 U5399 ( .A(n9208), .ZN(n7063) );
  NAND2_X1 U5400 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  NAND2_X1 U5401 ( .A1(n9186), .A2(n4525), .ZN(n4522) );
  INV_X1 U5402 ( .A(n4524), .ZN(n4523) );
  NOR2_X1 U5403 ( .A1(n9191), .A2(n5601), .ZN(n4525) );
  AND2_X1 U5404 ( .A1(n9188), .A2(n4530), .ZN(n4526) );
  NAND2_X1 U5405 ( .A1(n4530), .A2(n5601), .ZN(n4527) );
  OAI21_X1 U5406 ( .B1(n4509), .B2(n4510), .A(n4511), .ZN(n9043) );
  OAI21_X1 U5407 ( .B1(n9396), .B2(n9958), .A(n4485), .ZN(n4484) );
  AND2_X1 U5408 ( .A1(n9395), .A2(n9956), .ZN(n4485) );
  NOR2_X1 U5409 ( .A1(n6660), .A2(n9968), .ZN(n8410) );
  NAND2_X1 U5410 ( .A1(n4925), .A2(n6620), .ZN(n9418) );
  OR2_X1 U5411 ( .A1(n5604), .A2(n9988), .ZN(n10022) );
  OR2_X1 U5412 ( .A1(n9975), .A2(n5604), .ZN(n9554) );
  NAND2_X1 U5413 ( .A1(n6659), .A2(n6794), .ZN(n9036) );
  MUX2_X1 U5414 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8143), .S(n5043), .Z(n6659) );
  OAI211_X1 U5415 ( .C1(n9034), .C2(n5652), .A(n4756), .B(n4755), .ZN(n9562)
         );
  OR2_X1 U5416 ( .A1(n6620), .A2(n9034), .ZN(n4756) );
  NOR2_X1 U5417 ( .A1(n9073), .A2(n4759), .ZN(n4758) );
  OAI21_X1 U5418 ( .B1(n9561), .B2(n10099), .A(n4464), .ZN(n4754) );
  AOI22_X1 U5419 ( .A1(n9559), .A2(n10010), .B1(n9624), .B2(n9558), .ZN(n9560)
         );
  AND2_X1 U5420 ( .A1(n5597), .A2(n5596), .ZN(n9941) );
  NAND2_X1 U5421 ( .A1(n4714), .A2(n4713), .ZN(n5400) );
  AOI21_X1 U5422 ( .B1(n4716), .B2(n7993), .A(n7993), .ZN(n4713) );
  NAND2_X1 U5423 ( .A1(n8245), .A2(n8354), .ZN(n4628) );
  NAND2_X1 U5424 ( .A1(n4630), .A2(n8349), .ZN(n4629) );
  INV_X1 U5425 ( .A(n4534), .ZN(n4533) );
  INV_X1 U5426 ( .A(n4605), .ZN(n4607) );
  AND2_X1 U5427 ( .A1(n8263), .A2(n8264), .ZN(n4606) );
  NAND2_X1 U5428 ( .A1(n4612), .A2(n8258), .ZN(n4609) );
  NAND2_X1 U5429 ( .A1(n4611), .A2(n4610), .ZN(n8280) );
  AND2_X1 U5430 ( .A1(n8271), .A2(n8270), .ZN(n4610) );
  OAI211_X1 U5431 ( .C1(n8251), .C2(n4609), .A(n4608), .B(n4607), .ZN(n4611)
         );
  MUX2_X1 U5432 ( .A(n8269), .B(n8268), .S(n8349), .Z(n8271) );
  AOI21_X1 U5433 ( .B1(n4556), .B2(n4555), .A(n4554), .ZN(n8982) );
  AND2_X1 U5434 ( .A1(n9163), .A2(n9125), .ZN(n4554) );
  NOR2_X1 U5435 ( .A1(n8976), .A2(n9060), .ZN(n4555) );
  AND3_X1 U5436 ( .A1(n8305), .A2(n8663), .A3(n8304), .ZN(n8307) );
  NOR2_X1 U5437 ( .A1(n8354), .A2(n4626), .ZN(n4625) );
  INV_X1 U5438 ( .A(n8302), .ZN(n4626) );
  NAND2_X1 U5439 ( .A1(n8341), .A2(n8342), .ZN(n4604) );
  NAND2_X1 U5440 ( .A1(n4623), .A2(n8317), .ZN(n8319) );
  NAND2_X1 U5441 ( .A1(n10221), .A2(n4468), .ZN(n6605) );
  NAND2_X1 U5442 ( .A1(n6684), .A2(n6687), .ZN(n8198) );
  NAND2_X1 U5443 ( .A1(n6982), .A2(n6950), .ZN(n8197) );
  AOI21_X1 U5444 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n4550) );
  INV_X1 U5445 ( .A(n9013), .ZN(n4547) );
  NAND2_X1 U5446 ( .A1(n4549), .A2(n4750), .ZN(n4548) );
  NAND2_X1 U5447 ( .A1(n9085), .A2(n9125), .ZN(n4549) );
  INV_X1 U5448 ( .A(n5649), .ZN(n4790) );
  INV_X1 U5449 ( .A(n8481), .ZN(n4656) );
  NAND2_X1 U5450 ( .A1(n6818), .A2(n6502), .ZN(n8532) );
  OR2_X1 U5451 ( .A1(n10116), .A2(n10319), .ZN(n6878) );
  AOI21_X1 U5452 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6833), .A(n10145), .ZN(
        n6517) );
  AOI21_X1 U5453 ( .B1(n4850), .B2(n4848), .A(n4436), .ZN(n4847) );
  INV_X1 U5454 ( .A(n4850), .ZN(n4849) );
  INV_X1 U5455 ( .A(n4852), .ZN(n4848) );
  AND3_X1 U5456 ( .A1(n4690), .A2(n4689), .A3(n4466), .ZN(n6521) );
  NOR2_X1 U5457 ( .A1(n6605), .A2(n6604), .ZN(n8580) );
  OR2_X1 U5458 ( .A1(n8781), .A2(n8337), .ZN(n6171) );
  INV_X1 U5459 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5783) );
  OR2_X1 U5460 ( .A1(n8318), .A2(n6040), .ZN(n6431) );
  NAND2_X1 U5461 ( .A1(n4894), .A2(n4897), .ZN(n6432) );
  OR2_X1 U5462 ( .A1(n8122), .A2(n8497), .ZN(n8330) );
  AOI21_X1 U5463 ( .B1(n8033), .B2(n4887), .A(n8722), .ZN(n4886) );
  NAND2_X1 U5464 ( .A1(n4903), .A2(n5891), .ZN(n4902) );
  INV_X1 U5465 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4646) );
  INV_X1 U5466 ( .A(n7482), .ZN(n4722) );
  NOR2_X1 U5467 ( .A1(n5238), .A2(n9253), .ZN(n5206) );
  NAND2_X1 U5468 ( .A1(n6247), .A2(n4727), .ZN(n4726) );
  AND2_X1 U5469 ( .A1(n6377), .A2(n6468), .ZN(n6379) );
  AOI21_X1 U5470 ( .B1(n4546), .B2(n4545), .A(n4544), .ZN(n9023) );
  INV_X1 U5471 ( .A(n9014), .ZN(n4544) );
  AND2_X1 U5472 ( .A1(n9012), .A2(n9011), .ZN(n4545) );
  OAI21_X1 U5473 ( .B1(n4550), .B2(n4548), .A(n4547), .ZN(n4546) );
  NOR2_X1 U5474 ( .A1(n9564), .A2(n9026), .ZN(n4575) );
  INV_X1 U5475 ( .A(n4868), .ZN(n4867) );
  AOI21_X1 U5476 ( .B1(n4868), .B2(n4866), .A(n4442), .ZN(n4865) );
  INV_X1 U5477 ( .A(n5467), .ZN(n4866) );
  NAND2_X1 U5478 ( .A1(n9430), .A2(n9443), .ZN(n9094) );
  NOR2_X1 U5479 ( .A1(n5648), .A2(n4783), .ZN(n4782) );
  INV_X1 U5480 ( .A(n5646), .ZN(n4783) );
  AND2_X1 U5481 ( .A1(n9575), .A2(n9458), .ZN(n5648) );
  OAI21_X1 U5482 ( .B1(n4749), .B2(n9484), .A(n9473), .ZN(n4747) );
  OR2_X1 U5483 ( .A1(n9464), .A2(n9442), .ZN(n9081) );
  NOR2_X1 U5484 ( .A1(n7790), .A2(n9060), .ZN(n5331) );
  OR2_X1 U5485 ( .A1(n7794), .A2(n8922), .ZN(n9160) );
  NAND2_X1 U5486 ( .A1(n7794), .A2(n8922), .ZN(n8934) );
  NOR2_X1 U5487 ( .A1(n5263), .A2(n7755), .ZN(n5262) );
  AND2_X1 U5488 ( .A1(n5161), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5175) );
  AND2_X1 U5489 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5161) );
  NAND2_X1 U5490 ( .A1(n7063), .A2(n7682), .ZN(n9139) );
  OR2_X1 U5491 ( .A1(n9558), .A2(n5537), .ZN(n9101) );
  NAND2_X1 U5492 ( .A1(n9539), .A2(n4413), .ZN(n9492) );
  NAND2_X1 U5493 ( .A1(n5055), .A2(n5054), .ZN(n5481) );
  NAND2_X1 U5494 ( .A1(n5469), .A2(n5468), .ZN(n5055) );
  NAND2_X1 U5495 ( .A1(n5042), .A2(n5041), .ZN(n5456) );
  AND2_X1 U5496 ( .A1(n5334), .A2(n5335), .ZN(n5348) );
  INV_X1 U5497 ( .A(n5318), .ZN(n4991) );
  INV_X1 U5498 ( .A(n4407), .ZN(n4765) );
  AOI21_X1 U5499 ( .B1(n4407), .B2(n4764), .A(n4441), .ZN(n4763) );
  INV_X1 U5500 ( .A(n4769), .ZN(n4764) );
  OR3_X1 U5501 ( .A1(n5216), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n5254) );
  OAI21_X1 U5502 ( .B1(n4401), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4938), .ZN(
        n4939) );
  NAND2_X1 U5503 ( .A1(n4402), .A2(n9797), .ZN(n4938) );
  NAND2_X1 U5504 ( .A1(n6763), .A2(n6758), .ZN(n4932) );
  INV_X1 U5505 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4582) );
  AND2_X1 U5506 ( .A1(n4457), .A2(n8424), .ZN(n4636) );
  NOR2_X1 U5507 ( .A1(n5810), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5822) );
  INV_X1 U5508 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9838) );
  XNOR2_X1 U5509 ( .A(n6685), .B(n6684), .ZN(n6688) );
  XNOR2_X1 U5510 ( .A(n8116), .B(n8115), .ZN(n8433) );
  AOI21_X1 U5511 ( .B1(n4661), .B2(n4662), .A(n4461), .ZN(n4658) );
  INV_X1 U5512 ( .A(n4661), .ZN(n4659) );
  INV_X1 U5513 ( .A(n4651), .ZN(n4650) );
  OR2_X1 U5514 ( .A1(n4648), .A2(n8021), .ZN(n4647) );
  AND2_X1 U5515 ( .A1(n8180), .A2(n8505), .ZN(n8353) );
  NAND2_X1 U5516 ( .A1(n4597), .A2(n4595), .ZN(n8346) );
  AND2_X1 U5517 ( .A1(n7212), .A2(n6072), .ZN(n6167) );
  AND4_X1 U5518 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n8111)
         );
  NAND2_X1 U5519 ( .A1(n4678), .A2(n4679), .ZN(n6512) );
  NAND2_X1 U5520 ( .A1(n7071), .A2(n4432), .ZN(n4842) );
  AOI22_X1 U5521 ( .A1(n7411), .A2(P2_REG1_REG_9__SCAN_IN), .B1(n4853), .B2(
        n6515), .ZN(n10147) );
  XNOR2_X1 U5522 ( .A(n6517), .B(n10153), .ZN(n10162) );
  OAI21_X1 U5523 ( .B1(n10162), .B2(n4698), .A(n4697), .ZN(n10178) );
  NAND2_X1 U5524 ( .A1(n4699), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5525 ( .A1(n6518), .A2(n4699), .ZN(n4697) );
  INV_X1 U5526 ( .A(n10179), .ZN(n4699) );
  NOR2_X1 U5527 ( .A1(n10162), .A2(n5873), .ZN(n10161) );
  XNOR2_X1 U5528 ( .A(n6547), .B(n10185), .ZN(n10187) );
  NAND2_X1 U5529 ( .A1(n10187), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U5530 ( .A1(n8545), .A2(n6550), .ZN(n8570) );
  OAI211_X1 U5531 ( .C1(n8551), .C2(n4685), .A(n4684), .B(n6523), .ZN(n6525)
         );
  OR2_X1 U5532 ( .A1(n8562), .A2(n9899), .ZN(n4685) );
  NAND2_X1 U5533 ( .A1(n6522), .A2(n4686), .ZN(n4684) );
  NOR2_X1 U5534 ( .A1(n6553), .A2(n10224), .ZN(n8592) );
  INV_X1 U5535 ( .A(n8594), .ZN(n4863) );
  INV_X1 U5536 ( .A(n8579), .ZN(n4696) );
  OR2_X1 U5537 ( .A1(n8647), .A2(n8627), .ZN(n8632) );
  NAND2_X1 U5538 ( .A1(n5982), .A2(n5981), .ZN(n5992) );
  NAND2_X1 U5539 ( .A1(n8292), .A2(n8304), .ZN(n8693) );
  NAND2_X1 U5540 ( .A1(n5949), .A2(n5669), .ZN(n5965) );
  AND2_X1 U5541 ( .A1(n5929), .A2(n5710), .ZN(n5949) );
  NAND2_X1 U5542 ( .A1(n5899), .A2(n5898), .ZN(n5911) );
  OR2_X1 U5543 ( .A1(n5875), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5885) );
  NOR2_X2 U5544 ( .A1(n5885), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U5545 ( .A1(n4818), .A2(n4816), .ZN(n7731) );
  INV_X1 U5546 ( .A(n8255), .ZN(n4817) );
  OR2_X1 U5547 ( .A1(n5856), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U5548 ( .A1(n4873), .A2(n4434), .ZN(n7449) );
  NAND2_X1 U5549 ( .A1(n7320), .A2(n4411), .ZN(n4873) );
  AND2_X1 U5550 ( .A1(n5822), .A2(n9838), .ZN(n5837) );
  NAND2_X1 U5551 ( .A1(n5837), .A2(n5836), .ZN(n5856) );
  NAND2_X1 U5552 ( .A1(n7320), .A2(n8157), .ZN(n7319) );
  NOR2_X1 U5553 ( .A1(n7119), .A2(n4812), .ZN(n4811) );
  INV_X1 U5554 ( .A(n8221), .ZN(n4812) );
  NAND2_X1 U5555 ( .A1(n4878), .A2(n4876), .ZN(n7215) );
  OR2_X1 U5556 ( .A1(n4877), .A2(n4879), .ZN(n4876) );
  NOR2_X1 U5557 ( .A1(n5809), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U5558 ( .A1(n5784), .A2(n5783), .ZN(n5797) );
  OR2_X1 U5559 ( .A1(n5797), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U5560 ( .A1(n10242), .A2(n8202), .ZN(n7018) );
  NAND2_X1 U5561 ( .A1(n6051), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4828) );
  AND2_X1 U5562 ( .A1(n6093), .A2(n8349), .ZN(n6448) );
  AOI21_X1 U5563 ( .B1(n4890), .B2(n4893), .A(n4443), .ZN(n6165) );
  INV_X1 U5564 ( .A(n5999), .ZN(n4890) );
  NOR2_X1 U5565 ( .A1(n8337), .A2(n8710), .ZN(n6437) );
  NAND2_X1 U5566 ( .A1(n8797), .A2(n8627), .ZN(n4899) );
  NOR2_X1 U5567 ( .A1(n4827), .A2(n8298), .ZN(n4826) );
  INV_X1 U5568 ( .A(n8187), .ZN(n4827) );
  AND2_X1 U5569 ( .A1(n8300), .A2(n8306), .ZN(n8668) );
  AND4_X1 U5570 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n8720)
         );
  INV_X1 U5571 ( .A(n4886), .ZN(n4885) );
  NOR2_X1 U5572 ( .A1(n8037), .A2(n4889), .ZN(n8721) );
  AND2_X1 U5573 ( .A1(n8287), .A2(n8286), .ZN(n8722) );
  INV_X1 U5574 ( .A(n8164), .ZN(n8264) );
  AOI21_X1 U5575 ( .B1(n6814), .B2(n8142), .A(n4631), .ZN(n10297) );
  INV_X1 U5576 ( .A(n5854), .ZN(n4631) );
  INV_X1 U5577 ( .A(n10314), .ZN(n10303) );
  XNOR2_X1 U5578 ( .A(n4674), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U5579 ( .A1(n4675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4674) );
  AND2_X1 U5580 ( .A1(n4423), .A2(n6087), .ZN(n4673) );
  NAND2_X1 U5581 ( .A1(n6065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6061) );
  AND2_X1 U5582 ( .A1(n6058), .A2(n6057), .ZN(n6062) );
  OR2_X1 U5583 ( .A1(n5817), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5843) );
  OR2_X1 U5584 ( .A1(n5790), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U5585 ( .A1(n5175), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U5586 ( .A(n6350), .B(n6196), .ZN(n8370) );
  AND2_X1 U5587 ( .A1(n6258), .A2(n6257), .ZN(n7752) );
  INV_X1 U5588 ( .A(n9209), .ZN(n7044) );
  OR2_X1 U5589 ( .A1(n5406), .A2(n8842), .ZN(n5420) );
  NOR2_X1 U5590 ( .A1(n8838), .A2(n4742), .ZN(n4741) );
  INV_X1 U5591 ( .A(n4913), .ZN(n4742) );
  NAND2_X1 U5592 ( .A1(n4730), .A2(n4739), .ZN(n4733) );
  INV_X1 U5593 ( .A(n5448), .ZN(n5095) );
  XNOR2_X1 U5594 ( .A(n8369), .B(n8370), .ZN(n8891) );
  NAND2_X1 U5595 ( .A1(n8891), .A2(n8892), .ZN(n8890) );
  OR2_X1 U5596 ( .A1(n5372), .A2(n8873), .ZN(n5388) );
  NAND2_X1 U5597 ( .A1(n4467), .A2(n4529), .ZN(n4528) );
  INV_X1 U5598 ( .A(n9190), .ZN(n4529) );
  NOR2_X2 U5599 ( .A1(n8931), .A2(n9035), .ZN(n9182) );
  NOR2_X1 U5600 ( .A1(n9020), .A2(n4518), .ZN(n4517) );
  INV_X1 U5601 ( .A(n9078), .ZN(n4518) );
  AND2_X1 U5602 ( .A1(n8931), .A2(n9035), .ZN(n9039) );
  AND4_X1 U5603 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n7135)
         );
  AND2_X1 U5604 ( .A1(n9954), .A2(n9953), .ZN(n9951) );
  AND2_X1 U5605 ( .A1(n4476), .A2(n4475), .ZN(n9259) );
  NAND2_X1 U5606 ( .A1(n6965), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4475) );
  NOR2_X1 U5607 ( .A1(n9257), .A2(n4494), .ZN(n9272) );
  AND2_X1 U5608 ( .A1(n6966), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4494) );
  NOR2_X1 U5609 ( .A1(n9272), .A2(n9271), .ZN(n9270) );
  NOR2_X1 U5610 ( .A1(n9270), .A2(n4493), .ZN(n6969) );
  AND2_X1 U5611 ( .A1(n6968), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U5612 ( .A1(n6969), .A2(n6970), .ZN(n7086) );
  NOR2_X1 U5613 ( .A1(n7350), .A2(n4459), .ZN(n9289) );
  NOR2_X1 U5614 ( .A1(n9289), .A2(n9288), .ZN(n9287) );
  NAND2_X1 U5615 ( .A1(n9352), .A2(n4489), .ZN(n9376) );
  AND2_X1 U5616 ( .A1(n9353), .A2(n9351), .ZN(n4489) );
  NAND2_X1 U5617 ( .A1(n9352), .A2(n9351), .ZN(n4492) );
  AND2_X1 U5618 ( .A1(n9376), .A2(n9375), .ZN(n9381) );
  NAND2_X1 U5619 ( .A1(n4774), .A2(n4772), .ZN(n6619) );
  AND2_X1 U5620 ( .A1(n4773), .A2(n4786), .ZN(n4772) );
  INV_X1 U5621 ( .A(n4787), .ZN(n4786) );
  AND2_X1 U5622 ( .A1(n9100), .A2(n9091), .ZN(n6622) );
  NAND2_X1 U5623 ( .A1(n8391), .A2(n9025), .ZN(n8392) );
  AND2_X1 U5624 ( .A1(n5505), .A2(n5488), .ZN(n9431) );
  AND2_X1 U5625 ( .A1(n9078), .A2(n9094), .ZN(n9421) );
  NAND2_X1 U5626 ( .A1(n9456), .A2(n4868), .ZN(n8399) );
  NAND2_X1 U5627 ( .A1(n9456), .A2(n9081), .ZN(n9440) );
  NAND2_X1 U5628 ( .A1(n9539), .A2(n9931), .ZN(n9527) );
  NAND2_X1 U5629 ( .A1(n9539), .A2(n4572), .ZN(n9502) );
  NAND2_X1 U5630 ( .A1(n4836), .A2(n4834), .ZN(n9520) );
  AOI21_X1 U5631 ( .B1(n4837), .B2(n4839), .A(n4835), .ZN(n4834) );
  INV_X1 U5632 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U5633 ( .A1(n8004), .A2(n5634), .ZN(n9537) );
  OAI21_X1 U5634 ( .B1(n7977), .B2(n5632), .A(n5633), .ZN(n8005) );
  NAND2_X1 U5635 ( .A1(n8005), .A2(n9066), .ZN(n8004) );
  AND2_X1 U5636 ( .A1(n7936), .A2(n4418), .ZN(n9538) );
  NAND2_X1 U5637 ( .A1(n7936), .A2(n4408), .ZN(n8006) );
  NAND2_X1 U5638 ( .A1(n7936), .A2(n4406), .ZN(n7983) );
  AND2_X1 U5639 ( .A1(n7936), .A2(n8929), .ZN(n7937) );
  AND2_X1 U5640 ( .A1(n9162), .A2(n8977), .ZN(n9062) );
  NAND2_X1 U5641 ( .A1(n5622), .A2(n5621), .ZN(n9974) );
  NOR2_X1 U5642 ( .A1(n4428), .A2(n4405), .ZN(n5622) );
  NOR2_X1 U5643 ( .A1(n9971), .A2(n7794), .ZN(n7936) );
  NAND2_X1 U5644 ( .A1(n9160), .A2(n8934), .ZN(n9060) );
  NAND2_X1 U5645 ( .A1(n5275), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5307) );
  OR2_X1 U5646 ( .A1(n5307), .A2(n5306), .ZN(n5325) );
  NAND2_X1 U5647 ( .A1(n5305), .A2(n5304), .ZN(n9969) );
  OR2_X1 U5648 ( .A1(n7562), .A2(n4563), .ZN(n9970) );
  INV_X1 U5649 ( .A(n4565), .ZN(n4561) );
  NAND2_X1 U5650 ( .A1(n9154), .A2(n9976), .ZN(n9059) );
  INV_X1 U5651 ( .A(n4831), .ZN(n4830) );
  NOR2_X1 U5652 ( .A1(n7435), .A2(n7436), .ZN(n7637) );
  NAND2_X1 U5653 ( .A1(n7232), .A2(n8945), .ZN(n7566) );
  NAND2_X1 U5654 ( .A1(n7678), .A2(n4560), .ZN(n7435) );
  AND2_X1 U5655 ( .A1(n7264), .A2(n7609), .ZN(n4560) );
  NAND2_X1 U5656 ( .A1(n7675), .A2(n5610), .ZN(n7245) );
  NAND2_X1 U5657 ( .A1(n7678), .A2(n7609), .ZN(n7251) );
  NOR2_X1 U5658 ( .A1(n7677), .A2(n7682), .ZN(n7678) );
  NAND2_X1 U5659 ( .A1(n9139), .A2(n9134), .ZN(n8936) );
  NAND2_X1 U5660 ( .A1(n8935), .A2(n9135), .ZN(n9047) );
  INV_X1 U5661 ( .A(n5652), .ZN(n4759) );
  NAND2_X1 U5662 ( .A1(n5405), .A2(n5404), .ZN(n9608) );
  INV_X1 U5663 ( .A(n6649), .ZN(n5403) );
  INV_X1 U5664 ( .A(n6794), .ZN(n5402) );
  CLKBUF_X1 U5665 ( .A(n5123), .Z(n10062) );
  XNOR2_X1 U5666 ( .A(n5068), .B(n5067), .ZN(n7741) );
  XNOR2_X1 U5667 ( .A(n5501), .B(n5500), .ZN(n7727) );
  AND2_X1 U5668 ( .A1(n4860), .A2(n4552), .ZN(n5574) );
  NOR2_X1 U5669 ( .A1(n5080), .A2(n4856), .ZN(n4552) );
  AOI21_X1 U5670 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_18__SCAN_IN), .ZN(n4716) );
  XNOR2_X1 U5671 ( .A(n5411), .B(n5410), .ZN(n7183) );
  INV_X1 U5672 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5673 ( .A1(n4710), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U5674 ( .A1(n4712), .A2(n5140), .ZN(n4706) );
  NAND2_X1 U5675 ( .A1(n4766), .A2(n4767), .ZN(n5284) );
  INV_X1 U5676 ( .A(n4615), .ZN(n5193) );
  AOI21_X1 U5677 ( .B1(n4622), .B2(n4616), .A(n4619), .ZN(n4615) );
  NAND2_X1 U5678 ( .A1(n4622), .A2(n4960), .ZN(n5215) );
  XNOR2_X1 U5679 ( .A(n4958), .B(SI_7_), .ZN(n5226) );
  NAND2_X1 U5680 ( .A1(n4948), .A2(SI_4_), .ZN(n4949) );
  XNOR2_X1 U5681 ( .A(n4951), .B(SI_5_), .ZN(n5188) );
  XNOR2_X1 U5682 ( .A(n4947), .B(SI_4_), .ZN(n5171) );
  INV_X1 U5683 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9795) );
  AND2_X1 U5684 ( .A1(n5144), .A2(n5143), .ZN(n6848) );
  OR2_X1 U5685 ( .A1(n6763), .A2(n4751), .ZN(n4934) );
  NAND2_X1 U5686 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4751) );
  AND2_X1 U5687 ( .A1(n6750), .A2(n6749), .ZN(n8474) );
  AOI21_X1 U5688 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n7838) );
  AND3_X1 U5689 ( .A1(n5997), .A2(n5996), .A3(n5995), .ZN(n8642) );
  INV_X1 U5690 ( .A(n8672), .ZN(n8697) );
  NOR2_X1 U5691 ( .A1(n4660), .A2(n4662), .ZN(n8448) );
  NOR2_X1 U5692 ( .A1(n8441), .A2(n4664), .ZN(n4660) );
  NAND2_X1 U5693 ( .A1(n6009), .A2(n6008), .ZN(n8461) );
  AND2_X1 U5694 ( .A1(n7968), .A2(n4652), .ZN(n8022) );
  AND2_X1 U5695 ( .A1(n6932), .A2(n6700), .ZN(n7027) );
  OAI21_X1 U5696 ( .B1(n8441), .B2(n8440), .A(n4666), .ZN(n8472) );
  OAI21_X1 U5697 ( .B1(n8441), .B2(n4659), .A(n4658), .ZN(n8480) );
  NAND2_X1 U5698 ( .A1(n4671), .A2(n6708), .ZN(n7303) );
  NOR2_X1 U5699 ( .A1(n8360), .A2(n6678), .ZN(n4585) );
  OR2_X1 U5700 ( .A1(n8366), .A2(n8365), .ZN(n4591) );
  NAND2_X1 U5701 ( .A1(n4587), .A2(n4592), .ZN(n4586) );
  INV_X1 U5702 ( .A(n8642), .ZN(n8671) );
  INV_X1 U5703 ( .A(n6948), .ZN(n6919) );
  OAI21_X1 U5704 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n4495), .A(n6826), .ZN(n6802) );
  OR2_X1 U5705 ( .A1(n6816), .A2(n5729), .ZN(n6818) );
  INV_X1 U5706 ( .A(n4829), .ZN(n6540) );
  NAND2_X1 U5707 ( .A1(n7072), .A2(n7073), .ZN(n7071) );
  AND2_X1 U5708 ( .A1(n7076), .A2(n7075), .ZN(n7078) );
  XNOR2_X1 U5709 ( .A(n4842), .B(n6511), .ZN(n7278) );
  NOR2_X1 U5710 ( .A1(n7068), .A2(n4498), .ZN(n7276) );
  AND2_X1 U5711 ( .A1(n6587), .A2(n6588), .ZN(n4498) );
  AOI21_X1 U5712 ( .B1(n7278), .B2(P2_REG2_REG_7__SCAN_IN), .A(n4841), .ZN(
        n7328) );
  AND2_X1 U5713 ( .A1(n4842), .A2(n7283), .ZN(n4841) );
  XNOR2_X1 U5714 ( .A(n6544), .B(n6593), .ZN(n7408) );
  AND2_X1 U5715 ( .A1(n4851), .A2(n4427), .ZN(n10141) );
  NAND2_X1 U5716 ( .A1(n4690), .A2(n4689), .ZN(n10211) );
  OR2_X1 U5717 ( .A1(n8551), .A2(n9899), .ZN(n4688) );
  OR2_X1 U5718 ( .A1(n6049), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8097) );
  OR2_X1 U5719 ( .A1(n6032), .A2(n6021), .ZN(n8614) );
  NAND2_X1 U5720 ( .A1(n6151), .A2(n6150), .ZN(n8621) );
  NAND2_X1 U5721 ( .A1(n6148), .A2(n8684), .ZN(n6151) );
  NAND2_X1 U5722 ( .A1(n5948), .A2(n5947), .ZN(n8764) );
  NAND2_X1 U5723 ( .A1(n4455), .A2(n5881), .ZN(n7734) );
  NAND2_X1 U5724 ( .A1(n4821), .A2(n4819), .ZN(n7474) );
  NAND2_X1 U5725 ( .A1(n4821), .A2(n8236), .ZN(n7448) );
  INV_X1 U5726 ( .A(n4403), .ZN(n7714) );
  NAND2_X1 U5727 ( .A1(n6124), .A2(n8221), .ZN(n7118) );
  NAND2_X1 U5728 ( .A1(n4881), .A2(n5796), .ZN(n7120) );
  NAND2_X1 U5729 ( .A1(n7105), .A2(n5795), .ZN(n4881) );
  OR2_X1 U5730 ( .A1(n4399), .A2(n6761), .ZN(n5768) );
  AND2_X1 U5731 ( .A1(n6185), .A2(n10333), .ZN(n4872) );
  NAND2_X1 U5732 ( .A1(n6019), .A2(n6018), .ZN(n8786) );
  NAND2_X1 U5733 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U5734 ( .A1(n4801), .A2(n4409), .ZN(n6159) );
  OR2_X1 U5735 ( .A1(n6131), .A2(n6132), .ZN(n4801) );
  NAND2_X1 U5736 ( .A1(n5989), .A2(n5988), .ZN(n8803) );
  NAND2_X1 U5737 ( .A1(n5980), .A2(n5979), .ZN(n8809) );
  INV_X1 U5738 ( .A(n8108), .ZN(n8815) );
  NAND2_X1 U5739 ( .A1(n8692), .A2(n8292), .ZN(n8678) );
  AND2_X1 U5740 ( .A1(n4794), .A2(n8286), .ZN(n8704) );
  NAND2_X1 U5741 ( .A1(n5936), .A2(n5935), .ZN(n8829) );
  NAND2_X1 U5742 ( .A1(n5722), .A2(n5721), .ZN(n8048) );
  AND2_X1 U5743 ( .A1(n8039), .A2(n8038), .ZN(n8047) );
  NAND2_X1 U5744 ( .A1(n5926), .A2(n5925), .ZN(n7961) );
  NAND2_X1 U5745 ( .A1(n7055), .A2(n8142), .ZN(n5926) );
  NAND2_X1 U5746 ( .A1(n5910), .A2(n5909), .ZN(n7890) );
  NAND2_X1 U5747 ( .A1(n5896), .A2(n5895), .ZN(n7815) );
  NAND2_X1 U5748 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  NAND2_X1 U5749 ( .A1(n6081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6082) );
  AND3_X1 U5750 ( .A1(n5682), .A2(n5777), .A3(n4882), .ZN(n5716) );
  NAND2_X1 U5751 ( .A1(n4843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U5752 ( .A1(n5726), .A2(n4843), .ZN(n6830) );
  MUX2_X1 U5753 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5724), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5726) );
  NAND2_X1 U5754 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5724) );
  NAND2_X1 U5755 ( .A1(n8052), .A2(n4702), .ZN(n8054) );
  NAND2_X1 U5756 ( .A1(n6287), .A2(n6288), .ZN(n4704) );
  OAI21_X1 U5757 ( .B1(n7145), .B2(n7146), .A(n6221), .ZN(n7042) );
  OR2_X1 U5758 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  NAND2_X1 U5759 ( .A1(n6472), .A2(n6391), .ZN(n6488) );
  INV_X1 U5760 ( .A(n5606), .ZN(n10087) );
  OAI21_X1 U5761 ( .B1(n7483), .B2(n4723), .A(n4720), .ZN(n7778) );
  NAND2_X1 U5762 ( .A1(n7483), .A2(n7482), .ZN(n7481) );
  AOI21_X1 U5763 ( .B1(n4731), .B2(n4737), .A(n4412), .ZN(n4734) );
  AOI21_X1 U5764 ( .B1(n6471), .B2(n6470), .A(n8912), .ZN(n6473) );
  INV_X1 U5765 ( .A(n8909), .ZN(n8928) );
  AND2_X1 U5766 ( .A1(n6422), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8924) );
  AND2_X1 U5767 ( .A1(n4729), .A2(n6293), .ZN(n8914) );
  AND3_X1 U5768 ( .A1(n6413), .A2(n7037), .A3(n6414), .ZN(n8917) );
  NAND2_X1 U5769 ( .A1(n5513), .A2(n5512), .ZN(n9427) );
  OR2_X1 U5770 ( .A1(n8395), .A2(n5530), .ZN(n5513) );
  NAND4_X1 U5771 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n9208)
         );
  NAND2_X1 U5772 ( .A1(n5174), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5122) );
  AND2_X1 U5773 ( .A1(n4478), .A2(n4477), .ZN(n9245) );
  NOR2_X1 U5774 ( .A1(n9287), .A2(n4486), .ZN(n7490) );
  AND2_X1 U5775 ( .A1(n7357), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4486) );
  INV_X1 U5776 ( .A(n4488), .ZN(n9301) );
  INV_X1 U5777 ( .A(n9314), .ZN(n9313) );
  AOI211_X1 U5778 ( .C1(n9405), .C2(n9404), .A(n9968), .B(n9403), .ZN(n9556)
         );
  AOI21_X1 U5779 ( .B1(n9193), .B2(n9982), .A(n8404), .ZN(n8405) );
  NOR2_X1 U5780 ( .A1(n9443), .A2(n9549), .ZN(n8404) );
  NAND2_X1 U5781 ( .A1(n4785), .A2(n5649), .ZN(n8390) );
  OR2_X1 U5782 ( .A1(n9419), .A2(n5650), .ZN(n4785) );
  NAND2_X1 U5783 ( .A1(n4784), .A2(n5646), .ZN(n9438) );
  OR2_X1 U5784 ( .A1(n9451), .A2(n5647), .ZN(n4784) );
  NAND2_X1 U5785 ( .A1(n5445), .A2(n5444), .ZN(n9588) );
  OAI21_X1 U5786 ( .B1(n5642), .B2(n4750), .A(n4748), .ZN(n9472) );
  NAND2_X1 U5787 ( .A1(n5642), .A2(n5641), .ZN(n9485) );
  NAND2_X1 U5788 ( .A1(n8009), .A2(n8995), .ZN(n9545) );
  NAND2_X1 U5789 ( .A1(n7901), .A2(n9165), .ZN(n7980) );
  NAND2_X1 U5790 ( .A1(n7458), .A2(n9151), .ZN(n10000) );
  OR2_X1 U5791 ( .A1(n6639), .A2(n6636), .ZN(n10110) );
  AND2_X1 U5792 ( .A1(n6651), .A2(n6650), .ZN(n9632) );
  INV_X1 U5793 ( .A(n9418), .ZN(n6630) );
  NOR2_X1 U5794 ( .A1(n9410), .A2(n4846), .ZN(n4845) );
  CLKBUF_X1 U5795 ( .A(n10044), .Z(n10060) );
  OR2_X1 U5796 ( .A1(n7395), .A2(n5579), .ZN(n9940) );
  NAND2_X1 U5797 ( .A1(n6647), .A2(n5527), .ZN(n7927) );
  NAND2_X1 U5798 ( .A1(n5082), .A2(n4919), .ZN(n5087) );
  XNOR2_X1 U5799 ( .A(n5416), .B(n5415), .ZN(n7227) );
  NAND2_X1 U5800 ( .A1(n5413), .A2(n5412), .ZN(n5416) );
  OR2_X1 U5801 ( .A1(n5411), .A2(n5410), .ZN(n5413) );
  NAND2_X1 U5802 ( .A1(n5384), .A2(n5542), .ZN(n4715) );
  XNOR2_X1 U5803 ( .A(n5115), .B(n5114), .ZN(n9219) );
  XNOR2_X1 U5804 ( .A(n4638), .B(n8125), .ZN(n8131) );
  NAND2_X1 U5805 ( .A1(n10219), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6804) );
  AOI211_X1 U5806 ( .C1(n10237), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n10238) );
  AND2_X1 U5807 ( .A1(n4864), .A2(n4861), .ZN(n8596) );
  AOI21_X1 U5808 ( .B1(n4416), .B2(n10209), .A(n4500), .ZN(n6611) );
  OAI21_X1 U5809 ( .B1(n8784), .B2(n8731), .A(n6141), .ZN(n6142) );
  INV_X1 U5810 ( .A(n6462), .ZN(n6463) );
  OAI21_X1 U5811 ( .B1(n6616), .B2(n8731), .A(n6461), .ZN(n6462) );
  NAND2_X1 U5812 ( .A1(n8736), .A2(n8735), .ZN(n8738) );
  NOR2_X1 U5813 ( .A1(n4917), .A2(n6186), .ZN(n6187) );
  MUX2_X1 U5814 ( .A(n8780), .B(n8779), .S(n10315), .Z(n8783) );
  AND2_X1 U5815 ( .A1(n6443), .A2(n6442), .ZN(n6444) );
  AOI21_X1 U5816 ( .B1(n9187), .B2(n4526), .A(n4521), .ZN(n4520) );
  NAND2_X1 U5817 ( .A1(n4484), .A2(n5401), .ZN(n4483) );
  OAI21_X1 U5818 ( .B1(n9562), .B2(n9554), .A(n5666), .ZN(n5667) );
  AOI21_X1 U5819 ( .B1(n9559), .B2(n7512), .A(n5665), .ZN(n5666) );
  NAND2_X1 U5820 ( .A1(n6626), .A2(n6625), .ZN(n9416) );
  OR2_X1 U5821 ( .A1(n9036), .A2(n9616), .ZN(n6670) );
  NAND2_X1 U5822 ( .A1(n10101), .A2(n6629), .ZN(n4757) );
  OR2_X1 U5823 ( .A1(n9560), .A2(n10099), .ZN(n4752) );
  INV_X1 U5824 ( .A(n4754), .ZN(n4753) );
  INV_X1 U5825 ( .A(n10008), .ZN(n10079) );
  NAND2_X2 U5826 ( .A1(n8094), .A2(n5696), .ZN(n5745) );
  OR2_X1 U5827 ( .A1(n7928), .A2(n9062), .ZN(n4404) );
  NOR2_X1 U5828 ( .A1(n5606), .A2(n9984), .ZN(n4405) );
  AND2_X1 U5829 ( .A1(n8868), .A2(n8929), .ZN(n4406) );
  AND2_X1 U5830 ( .A1(n4767), .A2(n5283), .ZN(n4407) );
  AND2_X1 U5831 ( .A1(n4406), .A2(n4570), .ZN(n4408) );
  AND2_X1 U5832 ( .A1(n8157), .A2(n5850), .ZN(n4411) );
  AND2_X1 U5833 ( .A1(n4735), .A2(n6227), .ZN(n4412) );
  AND2_X1 U5834 ( .A1(n4572), .A2(n4571), .ZN(n4413) );
  NOR2_X1 U5835 ( .A1(n6039), .A2(n4898), .ZN(n4893) );
  AND3_X1 U5836 ( .A1(n4683), .A2(n4686), .A3(n4682), .ZN(n4414) );
  AOI21_X1 U5837 ( .B1(n8034), .B2(n4887), .A(n4885), .ZN(n4883) );
  AND2_X1 U5838 ( .A1(n8339), .A2(n8336), .ZN(n4415) );
  XOR2_X1 U5839 ( .A(n6556), .B(n6565), .Z(n4416) );
  AND2_X1 U5840 ( .A1(n7026), .A2(n6700), .ZN(n4417) );
  AND2_X1 U5841 ( .A1(n4408), .A2(n4569), .ZN(n4418) );
  OR2_X1 U5842 ( .A1(n4590), .A2(n8367), .ZN(n4419) );
  INV_X1 U5843 ( .A(n8995), .ZN(n4839) );
  INV_X1 U5844 ( .A(n6593), .ZN(n4853) );
  AND3_X1 U5845 ( .A1(n5701), .A2(n5700), .A3(n5699), .ZN(n8627) );
  OR2_X1 U5846 ( .A1(n6639), .A2(n9941), .ZN(n10099) );
  INV_X1 U5847 ( .A(n7577), .ZN(n4568) );
  NAND2_X1 U5848 ( .A1(n4813), .A2(n8230), .ZN(n7219) );
  NOR2_X1 U5849 ( .A1(n7562), .A2(n4567), .ZN(n4420) );
  INV_X1 U5850 ( .A(n6685), .ZN(n7690) );
  OR2_X1 U5851 ( .A1(n9037), .A2(n9041), .ZN(n4421) );
  OR2_X1 U5852 ( .A1(n10185), .A2(n6520), .ZN(n4422) );
  NAND2_X1 U5853 ( .A1(n6131), .A2(n8309), .ZN(n8631) );
  AND2_X1 U5854 ( .A1(n4645), .A2(n4646), .ZN(n5725) );
  NAND2_X1 U5855 ( .A1(n5777), .A2(n9796), .ZN(n5790) );
  NAND2_X1 U5856 ( .A1(n6085), .A2(n6084), .ZN(n6090) );
  AND4_X1 U5857 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5944), .ZN(n4423)
         );
  NAND2_X1 U5858 ( .A1(n5291), .A2(n5290), .ZN(n5606) );
  OR2_X1 U5859 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4424) );
  NAND2_X1 U5860 ( .A1(n6695), .A2(n10265), .ZN(n8203) );
  INV_X1 U5861 ( .A(n8203), .ZN(n4808) );
  AND2_X1 U5862 ( .A1(n6252), .A2(n6196), .ZN(n6213) );
  INV_X1 U5863 ( .A(n6950), .ZN(n6684) );
  AND4_X1 U5864 ( .A1(n4711), .A2(n5196), .A3(n5069), .A4(n4709), .ZN(n4425)
         );
  NAND2_X1 U5865 ( .A1(n9101), .A2(n9110), .ZN(n9073) );
  AND2_X1 U5866 ( .A1(n6889), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4426) );
  OR2_X1 U5867 ( .A1(n4508), .A2(n4507), .ZN(n7133) );
  AOI21_X1 U5868 ( .B1(n6182), .B2(n8684), .A(n6181), .ZN(n8096) );
  NAND2_X1 U5869 ( .A1(n5503), .A2(n5502), .ZN(n9564) );
  NAND2_X1 U5870 ( .A1(n4743), .A2(n4913), .ZN(n8837) );
  NAND2_X1 U5871 ( .A1(n6593), .A2(n7426), .ZN(n4427) );
  AND2_X1 U5872 ( .A1(n8316), .A2(n8633), .ZN(n8312) );
  AND2_X1 U5873 ( .A1(n9165), .A2(n9169), .ZN(n9063) );
  NAND2_X1 U5874 ( .A1(n5725), .A2(n5751), .ZN(n5765) );
  NOR2_X1 U5875 ( .A1(n5619), .A2(n7869), .ZN(n4428) );
  OR2_X1 U5876 ( .A1(n6649), .A2(n9797), .ZN(n4429) );
  NOR2_X1 U5877 ( .A1(n6526), .A2(n10229), .ZN(n4430) );
  AND2_X1 U5878 ( .A1(n5071), .A2(n4859), .ZN(n4858) );
  INV_X1 U5879 ( .A(n4858), .ZN(n4856) );
  INV_X1 U5880 ( .A(n4667), .ZN(n4666) );
  NOR2_X1 U5881 ( .A1(n8107), .A2(n8681), .ZN(n4667) );
  XNOR2_X1 U5882 ( .A(n4979), .B(SI_12_), .ZN(n5283) );
  OR2_X1 U5883 ( .A1(n6045), .A2(n6044), .ZN(n4431) );
  OR2_X1 U5884 ( .A1(n6588), .A2(n6541), .ZN(n4432) );
  AND2_X1 U5885 ( .A1(n8592), .A2(n8591), .ZN(n4433) );
  INV_X1 U5886 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7993) );
  INV_X1 U5887 ( .A(n7260), .ZN(n4737) );
  AND2_X1 U5888 ( .A1(n5851), .A2(n4874), .ZN(n4434) );
  INV_X1 U5889 ( .A(n8258), .ZN(n4613) );
  INV_X1 U5890 ( .A(n4680), .ZN(n4679) );
  NOR2_X1 U5891 ( .A1(n7075), .A2(n6510), .ZN(n4680) );
  NAND2_X1 U5892 ( .A1(n8353), .A2(n8598), .ZN(n4435) );
  INV_X1 U5893 ( .A(n4780), .ZN(n4779) );
  NAND2_X1 U5894 ( .A1(n4781), .A2(n4791), .ZN(n4780) );
  AND2_X1 U5895 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6833), .ZN(n4436) );
  OR2_X1 U5896 ( .A1(n8461), .A2(n8628), .ZN(n8320) );
  AND2_X1 U5897 ( .A1(n4600), .A2(n8336), .ZN(n4437) );
  OR2_X1 U5898 ( .A1(n8829), .A2(n8708), .ZN(n8287) );
  AND2_X1 U5899 ( .A1(n4586), .A2(n4591), .ZN(n4438) );
  OR2_X1 U5900 ( .A1(n4613), .A2(n8250), .ZN(n4439) );
  OR2_X1 U5901 ( .A1(n9026), .A2(n5517), .ZN(n9100) );
  OR2_X1 U5902 ( .A1(n4604), .A2(n8340), .ZN(n4440) );
  INV_X1 U5903 ( .A(n4749), .ZN(n4748) );
  OAI21_X1 U5904 ( .B1(n4750), .B2(n5641), .A(n5643), .ZN(n4749) );
  AND2_X1 U5905 ( .A1(n4980), .A2(SI_12_), .ZN(n4441) );
  NAND2_X1 U5906 ( .A1(n8398), .A2(n5514), .ZN(n4442) );
  NAND2_X1 U5907 ( .A1(n4431), .A2(n4891), .ZN(n4443) );
  INV_X1 U5908 ( .A(n4964), .ZN(n4619) );
  NAND2_X1 U5909 ( .A1(n4961), .A2(n9745), .ZN(n4964) );
  INV_X1 U5910 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5540) );
  AND2_X1 U5911 ( .A1(n8829), .A2(n8509), .ZN(n4444) );
  AND2_X1 U5912 ( .A1(n5077), .A2(n5079), .ZN(n4445) );
  INV_X1 U5913 ( .A(n9151), .ZN(n4833) );
  AND2_X1 U5914 ( .A1(n4858), .A2(n5073), .ZN(n4446) );
  AND2_X1 U5915 ( .A1(n5808), .A2(n5795), .ZN(n4447) );
  AND2_X1 U5916 ( .A1(n4964), .A2(n5226), .ZN(n4448) );
  AND2_X1 U5917 ( .A1(n5734), .A2(n5735), .ZN(n4449) );
  AND2_X1 U5918 ( .A1(n6484), .A2(n6482), .ZN(n6472) );
  AND2_X1 U5919 ( .A1(n4688), .A2(n4687), .ZN(n4450) );
  OR2_X1 U5920 ( .A1(n9128), .A2(n4527), .ZN(n4451) );
  AND2_X1 U5921 ( .A1(n5364), .A2(n5629), .ZN(n4452) );
  AND2_X1 U5922 ( .A1(n5106), .A2(n7868), .ZN(n5135) );
  INV_X1 U5923 ( .A(n5135), .ZN(n5125) );
  XNOR2_X1 U5924 ( .A(n5400), .B(n5399), .ZN(n5654) );
  INV_X1 U5925 ( .A(n7664), .ZN(n7264) );
  INV_X1 U5926 ( .A(n9484), .ZN(n4750) );
  AND2_X1 U5927 ( .A1(n7481), .A2(n4726), .ZN(n4453) );
  NAND2_X1 U5928 ( .A1(n4860), .A2(n4858), .ZN(n5354) );
  OR2_X1 U5929 ( .A1(n5287), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U5930 ( .A1(n5369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U5931 ( .A1(n5544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U5932 ( .A1(n6129), .A2(n8281), .ZN(n8718) );
  NAND2_X1 U5933 ( .A1(n4815), .A2(n8266), .ZN(n7946) );
  NAND2_X1 U5934 ( .A1(n4715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5398) );
  OR2_X1 U5935 ( .A1(n7471), .A2(n8162), .ZN(n4455) );
  INV_X1 U5936 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4711) );
  AND4_X1 U5937 ( .A1(n9091), .A2(n9125), .A3(n9094), .A4(n9092), .ZN(n4456)
         );
  INV_X1 U5938 ( .A(n9175), .ZN(n4835) );
  NAND2_X1 U5939 ( .A1(n4794), .A2(n4793), .ZN(n8703) );
  AND2_X1 U5940 ( .A1(n4425), .A2(n4705), .ZN(n5285) );
  NAND2_X1 U5941 ( .A1(n4700), .A2(n6792), .ZN(n6252) );
  NAND2_X1 U5942 ( .A1(n8121), .A2(n8459), .ZN(n4457) );
  INV_X1 U5943 ( .A(n5174), .ZN(n5200) );
  AND2_X1 U5944 ( .A1(n6056), .A2(n6055), .ZN(n8337) );
  INV_X1 U5945 ( .A(n8337), .ZN(n4603) );
  OR2_X1 U5946 ( .A1(n8760), .A2(n8709), .ZN(n8292) );
  NOR2_X1 U5947 ( .A1(n9461), .A2(n9575), .ZN(n5659) );
  NOR2_X1 U5948 ( .A1(n10161), .A2(n6518), .ZN(n4458) );
  AND2_X1 U5949 ( .A1(n7351), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4459) );
  INV_X1 U5950 ( .A(n5287), .ZN(n4860) );
  INV_X1 U5951 ( .A(n4898), .ZN(n4897) );
  NAND2_X1 U5952 ( .A1(n8114), .A2(n8642), .ZN(n4460) );
  INV_X1 U5953 ( .A(n8797), .ZN(n8647) );
  AND2_X1 U5954 ( .A1(n5709), .A2(n5708), .ZN(n8797) );
  NOR2_X1 U5955 ( .A1(n8113), .A2(n8682), .ZN(n4461) );
  XNOR2_X1 U5956 ( .A(n8340), .B(n8337), .ZN(n8171) );
  NAND2_X1 U5957 ( .A1(n9997), .A2(n7869), .ZN(n4462) );
  AND2_X1 U5958 ( .A1(n4692), .A2(n4422), .ZN(n4463) );
  AOI21_X1 U5960 ( .B1(n6109), .B2(n6789), .A(n6092), .ZN(n6677) );
  NAND2_X1 U5961 ( .A1(n5436), .A2(n5435), .ZN(n9494) );
  INV_X1 U5962 ( .A(n9494), .ZN(n4571) );
  NAND2_X1 U5963 ( .A1(n5386), .A2(n5385), .ZN(n8910) );
  INV_X1 U5964 ( .A(n8910), .ZN(n4569) );
  AOI21_X1 U5965 ( .B1(n6089), .B2(n7518), .A(n6091), .ZN(n6109) );
  NAND2_X1 U5966 ( .A1(n7018), .A2(n8150), .ZN(n7008) );
  NAND2_X1 U5967 ( .A1(n7303), .A2(n6714), .ZN(n7304) );
  OR2_X1 U5968 ( .A1(n7562), .A2(n7577), .ZN(n4566) );
  NAND2_X1 U5969 ( .A1(n6224), .A2(n4740), .ZN(n4739) );
  OR2_X1 U5970 ( .A1(n10101), .A2(n5533), .ZN(n4464) );
  NAND2_X1 U5971 ( .A1(n7319), .A2(n5835), .ZN(n7420) );
  INV_X1 U5972 ( .A(n4889), .ZN(n4887) );
  NAND2_X1 U5973 ( .A1(n5371), .A2(n5370), .ZN(n9619) );
  INV_X1 U5974 ( .A(n9619), .ZN(n4570) );
  NAND2_X1 U5975 ( .A1(n5471), .A2(n5470), .ZN(n9575) );
  INV_X1 U5976 ( .A(n9575), .ZN(n4792) );
  INV_X1 U5977 ( .A(n4564), .ZN(n10009) );
  OR2_X1 U5978 ( .A1(n7562), .A2(n4565), .ZN(n4564) );
  NAND2_X1 U5979 ( .A1(n4730), .A2(n4738), .ZN(n4465) );
  OR2_X1 U5980 ( .A1(n10202), .A2(n9853), .ZN(n4466) );
  AND2_X1 U5981 ( .A1(n5598), .A2(n6899), .ZN(n9985) );
  NAND2_X1 U5982 ( .A1(n5087), .A2(n5086), .ZN(n5558) );
  OR3_X1 U5983 ( .A1(n9337), .A2(n6190), .A3(n9189), .ZN(n4467) );
  INV_X1 U5984 ( .A(n8562), .ZN(n4686) );
  INV_X1 U5985 ( .A(n7366), .ZN(n4670) );
  OR2_X1 U5986 ( .A1(n6603), .A2(n7192), .ZN(n4468) );
  OR2_X1 U5987 ( .A1(n4527), .A2(n5401), .ZN(n4469) );
  INV_X1 U5988 ( .A(n8367), .ZN(n4592) );
  AND2_X1 U5989 ( .A1(n4592), .A2(n4585), .ZN(n4470) );
  INV_X1 U5990 ( .A(n5697), .ZN(n8094) );
  INV_X1 U5991 ( .A(n5654), .ZN(n5401) );
  XNOR2_X1 U5992 ( .A(n5960), .B(n5959), .ZN(n8360) );
  OR2_X1 U5993 ( .A1(n6610), .A2(n8359), .ZN(n4471) );
  INV_X2 U5994 ( .A(P2_U3893), .ZN(n8584) );
  INV_X1 U5995 ( .A(n4478), .ZN(n6962) );
  INV_X1 U5996 ( .A(n4476), .ZN(n9243) );
  NAND4_X1 U5997 ( .A1(n4483), .A2(n9399), .A3(n4479), .A4(n9400), .ZN(
        P1_U3262) );
  NAND2_X1 U5998 ( .A1(n9376), .A2(n4490), .ZN(n9354) );
  NAND2_X1 U5999 ( .A1(n4492), .A2(n4491), .ZN(n4490) );
  INV_X1 U6000 ( .A(n9353), .ZN(n4491) );
  NOR2_X1 U6001 ( .A1(n5140), .A2(n7993), .ZN(n5141) );
  NOR2_X2 U6002 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5140) );
  NOR2_X1 U6003 ( .A1(n9016), .A2(n4512), .ZN(n4509) );
  OAI21_X1 U6004 ( .B1(n4512), .B2(n4517), .A(n4514), .ZN(n4510) );
  NAND3_X1 U6005 ( .A1(n9024), .A2(n4456), .A3(n4514), .ZN(n4511) );
  NAND2_X1 U6006 ( .A1(n9034), .A2(n9033), .ZN(n4519) );
  OAI21_X1 U6007 ( .B1(n9129), .B2(n4451), .A(n4520), .ZN(P1_U3242) );
  INV_X1 U6008 ( .A(n9191), .ZN(n4530) );
  OAI21_X1 U6009 ( .B1(n8948), .B2(n4535), .A(n4531), .ZN(n4540) );
  OAI21_X1 U6010 ( .B1(n8948), .B2(n4537), .A(n4533), .ZN(n4542) );
  INV_X1 U6011 ( .A(n9142), .ZN(n4538) );
  NAND2_X1 U6012 ( .A1(n4542), .A2(n4540), .ZN(n8956) );
  NAND2_X1 U6013 ( .A1(n8949), .A2(n8945), .ZN(n4541) );
  NAND2_X1 U6014 ( .A1(n5079), .A2(n4551), .ZN(n5082) );
  NAND3_X1 U6015 ( .A1(n4558), .A2(n4557), .A3(n9978), .ZN(n4556) );
  NAND3_X1 U6016 ( .A1(n8973), .A2(n9125), .A3(n9154), .ZN(n4557) );
  NAND3_X1 U6017 ( .A1(n8967), .A2(n9976), .A3(n9044), .ZN(n4558) );
  NAND2_X1 U6018 ( .A1(n5658), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U6019 ( .A1(n4561), .A2(n10087), .ZN(n4563) );
  NAND2_X1 U6020 ( .A1(n4576), .A2(n4937), .ZN(n5146) );
  NAND2_X1 U6021 ( .A1(n5117), .A2(n5116), .ZN(n4576) );
  XNOR2_X1 U6022 ( .A(n4935), .B(SI_1_), .ZN(n5117) );
  NAND2_X1 U6023 ( .A1(n4931), .A2(n4932), .ZN(n4935) );
  NAND2_X1 U6024 ( .A1(n5246), .A2(n5245), .ZN(n4957) );
  NAND2_X1 U6025 ( .A1(n5189), .A2(n5188), .ZN(n4577) );
  INV_X1 U6026 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4583) );
  INV_X1 U6027 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4581) );
  INV_X1 U6028 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4580) );
  AND2_X4 U6029 ( .A1(n4579), .A2(n4578), .ZN(n6763) );
  NAND3_X1 U6030 ( .A1(n4583), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4578) );
  NAND3_X1 U6031 ( .A1(n4582), .A2(n4581), .A3(n4580), .ZN(n4579) );
  NAND2_X1 U6032 ( .A1(n4593), .A2(n8360), .ZN(n4590) );
  OR2_X2 U6033 ( .A1(n4911), .A2(n8359), .ZN(n4593) );
  NAND2_X1 U6034 ( .A1(n8358), .A2(n4470), .ZN(n4584) );
  OAI211_X1 U6035 ( .C1(n8358), .C2(n4419), .A(n4438), .B(n4584), .ZN(P2_U3296) );
  NAND2_X1 U6036 ( .A1(n4593), .A2(n4471), .ZN(n4588) );
  OR2_X1 U6037 ( .A1(n4593), .A2(n6610), .ZN(n4589) );
  INV_X1 U6038 ( .A(n8344), .ZN(n4594) );
  NAND2_X1 U6039 ( .A1(n4594), .A2(n4598), .ZN(n4597) );
  INV_X1 U6040 ( .A(n4604), .ZN(n4600) );
  INV_X1 U6041 ( .A(n8265), .ZN(n4612) );
  OAI21_X1 U6042 ( .B1(n8265), .B2(n4439), .A(n4606), .ZN(n4605) );
  NAND2_X1 U6043 ( .A1(n8257), .A2(n4612), .ZN(n4608) );
  NAND2_X1 U6044 ( .A1(n5227), .A2(n5226), .ZN(n4622) );
  NAND2_X1 U6045 ( .A1(n5227), .A2(n4448), .ZN(n4614) );
  NAND3_X1 U6046 ( .A1(n4627), .A2(n8314), .A3(n4624), .ZN(n4623) );
  NAND3_X1 U6047 ( .A1(n8303), .A2(n8633), .A3(n4625), .ZN(n4624) );
  NAND3_X1 U6048 ( .A1(n8310), .A2(n8354), .A3(n8309), .ZN(n4627) );
  NAND3_X1 U6049 ( .A1(n4629), .A2(n4628), .A3(n8246), .ZN(n8256) );
  NAND3_X1 U6050 ( .A1(n8247), .A2(n8237), .A3(n8236), .ZN(n4630) );
  OAI21_X1 U6051 ( .B1(n6916), .B2(n4632), .A(n6915), .ZN(n6917) );
  NAND2_X1 U6052 ( .A1(n4632), .A2(n6916), .ZN(n6915) );
  AND2_X1 U6053 ( .A1(n6691), .A2(n6689), .ZN(n4632) );
  NAND2_X1 U6054 ( .A1(n8490), .A2(n8491), .ZN(n4637) );
  NAND2_X1 U6055 ( .A1(n4637), .A2(n4636), .ZN(n8423) );
  NAND2_X1 U6056 ( .A1(n5682), .A2(n4639), .ZN(n5719) );
  NAND3_X1 U6057 ( .A1(n4643), .A2(n4646), .A3(n5681), .ZN(n4641) );
  NAND2_X1 U6058 ( .A1(n7840), .A2(n7839), .ZN(n7968) );
  OAI21_X2 U6059 ( .B1(n4649), .B2(n4647), .A(n4650), .ZN(n8064) );
  INV_X1 U6060 ( .A(n7840), .ZN(n4649) );
  NAND2_X1 U6061 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  INV_X1 U6062 ( .A(n8441), .ZN(n4657) );
  AOI21_X2 U6063 ( .B1(n4657), .B2(n4655), .A(n4654), .ZN(n8116) );
  INV_X1 U6064 ( .A(n7194), .ZN(n4671) );
  NAND2_X1 U6065 ( .A1(n4669), .A2(n4668), .ZN(n6715) );
  NAND2_X1 U6066 ( .A1(n7194), .A2(n6714), .ZN(n4669) );
  NAND2_X1 U6067 ( .A1(n7025), .A2(n7162), .ZN(n4672) );
  NAND2_X1 U6068 ( .A1(n4417), .A2(n6932), .ZN(n7025) );
  NAND2_X1 U6069 ( .A1(n4672), .A2(n7161), .ZN(n7165) );
  AND2_X2 U6070 ( .A1(n5686), .A2(n4423), .ZN(n6088) );
  NAND2_X1 U6071 ( .A1(n5686), .A2(n4673), .ZN(n4675) );
  INV_X1 U6072 ( .A(n6930), .ZN(n6696) );
  NAND2_X1 U6073 ( .A1(n5657), .A2(n7186), .ZN(n7677) );
  OAI21_X1 U6074 ( .B1(n9562), .B2(n9627), .A(n4760), .ZN(n9633) );
  NOR2_X1 U6075 ( .A1(n8346), .A2(n8345), .ZN(n8350) );
  NAND2_X1 U6076 ( .A1(n6509), .A2(n4676), .ZN(n4678) );
  NAND2_X1 U6077 ( .A1(n4687), .A2(n9899), .ZN(n4682) );
  NAND2_X1 U6078 ( .A1(n8551), .A2(n4687), .ZN(n4683) );
  INV_X1 U6079 ( .A(n4688), .ZN(n8550) );
  INV_X1 U6080 ( .A(n6522), .ZN(n4687) );
  INV_X1 U6081 ( .A(n4692), .ZN(n10193) );
  NAND2_X1 U6082 ( .A1(n6526), .A2(n4696), .ZN(n4693) );
  NOR2_X1 U6083 ( .A1(n10230), .A2(n10231), .ZN(n10229) );
  MUX2_X1 U6084 ( .A(n8834), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6085 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8834), .S(n6497), .Z(n6979) );
  NAND2_X1 U6086 ( .A1(n4701), .A2(n6191), .ZN(n4700) );
  NAND2_X1 U6087 ( .A1(n6190), .A2(n6192), .ZN(n4701) );
  NAND2_X1 U6088 ( .A1(n5654), .A2(n6415), .ZN(n6190) );
  NAND3_X1 U6089 ( .A1(n6287), .A2(n6288), .A3(n8053), .ZN(n8052) );
  NAND2_X1 U6090 ( .A1(n4704), .A2(n4703), .ZN(n4702) );
  INV_X1 U6091 ( .A(n8053), .ZN(n4703) );
  NAND3_X2 U6092 ( .A1(n4425), .A2(n4708), .A3(n4707), .ZN(n5287) );
  NAND2_X1 U6093 ( .A1(n5384), .A2(n4716), .ZN(n4714) );
  NAND2_X1 U6094 ( .A1(n7483), .A2(n4720), .ZN(n4719) );
  INV_X1 U6095 ( .A(n6248), .ZN(n4727) );
  NAND3_X1 U6096 ( .A1(n4729), .A2(n8916), .A3(n6293), .ZN(n8915) );
  NAND2_X1 U6097 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  INV_X1 U6098 ( .A(n6292), .ZN(n4728) );
  CLKBUF_X1 U6099 ( .A(n7060), .Z(n4730) );
  INV_X1 U6100 ( .A(n4731), .ZN(n4738) );
  NAND2_X1 U6101 ( .A1(n4739), .A2(n4732), .ZN(n4731) );
  INV_X1 U6102 ( .A(n6227), .ZN(n4732) );
  NAND2_X1 U6103 ( .A1(n4733), .A2(n6227), .ZN(n7259) );
  INV_X1 U6104 ( .A(n4739), .ZN(n4735) );
  NOR2_X1 U6105 ( .A1(n6227), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U6106 ( .A1(n7062), .A2(n7061), .ZN(n7060) );
  NAND2_X1 U6107 ( .A1(n4743), .A2(n4741), .ZN(n8835) );
  NAND2_X1 U6108 ( .A1(n6310), .A2(n8870), .ZN(n8899) );
  NOR2_X1 U6109 ( .A1(n4745), .A2(n6318), .ZN(n4744) );
  INV_X1 U6110 ( .A(n8870), .ZN(n4745) );
  NAND2_X1 U6111 ( .A1(n4860), .A2(n4446), .ZN(n5544) );
  INV_X1 U6112 ( .A(n4746), .ZN(n5645) );
  NAND3_X1 U6113 ( .A1(n4404), .A2(n5630), .A3(n5629), .ZN(n7900) );
  NAND3_X1 U6114 ( .A1(n4404), .A2(n5630), .A3(n4452), .ZN(n7898) );
  INV_X4 U6115 ( .A(n6763), .ZN(n5043) );
  NAND2_X1 U6116 ( .A1(n6620), .A2(n4758), .ZN(n4755) );
  OAI211_X1 U6117 ( .C1(n9562), .C2(n4757), .A(n4753), .B(n4752), .ZN(P1_U3519) );
  NAND2_X1 U6118 ( .A1(n4761), .A2(n4762), .ZN(n5317) );
  NAND2_X1 U6119 ( .A1(n5253), .A2(n4763), .ZN(n4761) );
  NAND2_X1 U6120 ( .A1(n5253), .A2(n4769), .ZN(n4766) );
  OAI21_X1 U6121 ( .B1(n5253), .B2(n4771), .A(n4972), .ZN(n5270) );
  NAND2_X1 U6122 ( .A1(n9451), .A2(n4776), .ZN(n4774) );
  NAND2_X1 U6123 ( .A1(n9451), .A2(n4782), .ZN(n4775) );
  NAND2_X1 U6124 ( .A1(n6129), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U6125 ( .A1(n6131), .A2(n4410), .ZN(n4800) );
  AOI21_X2 U6126 ( .B1(n4410), .B2(n6132), .A(n4799), .ZN(n4798) );
  NAND2_X1 U6127 ( .A1(n4805), .A2(n4804), .ZN(n7009) );
  INV_X1 U6128 ( .A(n4806), .ZN(n4805) );
  OAI21_X1 U6129 ( .B1(n8150), .B2(n4808), .A(n8210), .ZN(n4806) );
  NAND2_X1 U6130 ( .A1(n6124), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U6131 ( .A1(n4810), .A2(n8223), .ZN(n7218) );
  INV_X1 U6132 ( .A(n7218), .ZN(n4813) );
  NAND2_X1 U6133 ( .A1(n4815), .A2(n4814), .ZN(n8031) );
  NAND2_X1 U6134 ( .A1(n7418), .A2(n4819), .ZN(n4818) );
  AOI21_X1 U6135 ( .B1(n4819), .B2(n7421), .A(n4817), .ZN(n4816) );
  NAND2_X1 U6136 ( .A1(n7731), .A2(n8253), .ZN(n6126) );
  NAND2_X1 U6137 ( .A1(n8692), .A2(n4826), .ZN(n8664) );
  NAND2_X1 U6138 ( .A1(n8664), .A2(n8188), .ZN(n6130) );
  INV_X1 U6139 ( .A(n5251), .ZN(n7459) );
  NAND2_X1 U6140 ( .A1(n4832), .A2(n4830), .ZN(n5282) );
  NAND2_X1 U6141 ( .A1(n5251), .A2(n9151), .ZN(n4832) );
  NAND2_X1 U6142 ( .A1(n8010), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U6143 ( .A1(n6626), .A2(n4845), .ZN(n4844) );
  AOI21_X1 U6144 ( .B1(n6630), .B2(n6629), .A(n4844), .ZN(n6640) );
  OAI21_X1 U6145 ( .B1(n6544), .B2(n4849), .A(n4847), .ZN(n6545) );
  NAND2_X1 U6146 ( .A1(n7901), .A2(n4854), .ZN(n7978) );
  NAND2_X1 U6147 ( .A1(n4445), .A2(n4855), .ZN(n5103) );
  OAI21_X1 U6148 ( .B1(n9453), .B2(n4867), .A(n4865), .ZN(n5516) );
  NAND2_X1 U6149 ( .A1(n4870), .A2(n10315), .ZN(n6188) );
  NAND2_X1 U6150 ( .A1(n8096), .A2(n6185), .ZN(n4870) );
  NAND2_X1 U6151 ( .A1(n4871), .A2(n6672), .ZN(n6675) );
  NAND2_X1 U6152 ( .A1(n8096), .A2(n4872), .ZN(n4871) );
  INV_X2 U6153 ( .A(n5746), .ZN(n5824) );
  XNOR2_X2 U6154 ( .A(n5695), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6155 ( .A1(n7105), .A2(n4447), .ZN(n4878) );
  INV_X1 U6156 ( .A(n5719), .ZN(n5686) );
  OAI21_X1 U6157 ( .B1(n8034), .B2(n4885), .A(n4884), .ZN(n4888) );
  INV_X1 U6158 ( .A(n4888), .ZN(n8706) );
  AND2_X1 U6159 ( .A1(n8048), .A2(n8510), .ZN(n4889) );
  NAND2_X1 U6160 ( .A1(n5999), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U6161 ( .A1(n5999), .A2(n4899), .ZN(n8625) );
  NOR2_X1 U6162 ( .A1(n8791), .A2(n8643), .ZN(n4898) );
  OAI21_X1 U6163 ( .B1(n7471), .B2(n4902), .A(n4900), .ZN(n7807) );
  NAND2_X1 U6164 ( .A1(n8162), .A2(n5881), .ZN(n4903) );
  XNOR2_X1 U6165 ( .A(n5284), .B(n5283), .ZN(n6986) );
  MUX2_X1 U6166 ( .A(n6118), .B(n8779), .S(n8714), .Z(n6144) );
  AOI21_X1 U6167 ( .B1(n6080), .B2(n8684), .A(n6079), .ZN(n8779) );
  NAND2_X1 U6168 ( .A1(n6613), .A2(n10315), .ZN(n6445) );
  AOI21_X1 U6169 ( .B1(n5553), .B2(n5552), .A(n10002), .ZN(n5563) );
  INV_X1 U6170 ( .A(n5106), .ZN(n8092) );
  NAND2_X1 U6171 ( .A1(n5607), .A2(n8070), .ZN(n8071) );
  XNOR2_X1 U6172 ( .A(n6217), .B(n6388), .ZN(n6220) );
  NAND2_X1 U6173 ( .A1(n8604), .A2(n6147), .ZN(n6148) );
  NAND2_X1 U6174 ( .A1(n8779), .A2(n10333), .ZN(n8736) );
  NAND2_X1 U6175 ( .A1(n8785), .A2(n10333), .ZN(n8741) );
  INV_X1 U6176 ( .A(n8195), .ZN(n6945) );
  NAND4_X2 U6177 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n6687)
         );
  XNOR2_X1 U6178 ( .A(n6165), .B(n8171), .ZN(n6080) );
  OAI21_X1 U6179 ( .B1(n6760), .B2(n10259), .A(n6533), .ZN(n8529) );
  NAND2_X1 U6180 ( .A1(n6760), .A2(n10259), .ZN(n6533) );
  NAND2_X1 U6181 ( .A1(n6760), .A2(n6500), .ZN(n6499) );
  AND2_X1 U6182 ( .A1(n7712), .A2(n8516), .ZN(n4904) );
  INV_X1 U6183 ( .A(n8708), .ZN(n8509) );
  OR2_X1 U6184 ( .A1(n6497), .A2(n6830), .ZN(n4905) );
  OR2_X1 U6185 ( .A1(n9414), .A2(n9936), .ZN(n4906) );
  OR2_X1 U6186 ( .A1(n6246), .A2(n6245), .ZN(n4907) );
  NOR2_X1 U6187 ( .A1(n5414), .A2(n5412), .ZN(n4908) );
  NOR2_X1 U6188 ( .A1(n5022), .A2(n5396), .ZN(n4909) );
  OR2_X1 U6189 ( .A1(n9340), .A2(n9339), .ZN(n4910) );
  OR2_X1 U6190 ( .A1(n6260), .A2(n6259), .ZN(n4912) );
  OR2_X1 U6191 ( .A1(n6317), .A2(n6316), .ZN(n4913) );
  OR2_X1 U6192 ( .A1(n9414), .A2(n9616), .ZN(n4914) );
  OR2_X1 U6193 ( .A1(n6674), .A2(n8747), .ZN(n4915) );
  OR2_X1 U6194 ( .A1(n8714), .A2(n6459), .ZN(n4916) );
  AND2_X1 U6195 ( .A1(n10317), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4917) );
  AND2_X1 U6196 ( .A1(n8110), .A2(n8697), .ZN(n4918) );
  AND2_X1 U6197 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4919) );
  AND2_X1 U6198 ( .A1(n7175), .A2(n6621), .ZN(n9627) );
  OR2_X1 U6199 ( .A1(n8116), .A2(n8115), .ZN(n4920) );
  NAND2_X1 U6200 ( .A1(n8064), .A2(n8063), .ZN(n8105) );
  INV_X1 U6201 ( .A(n5632), .ZN(n9065) );
  AND2_X1 U6202 ( .A1(n8987), .A2(n8994), .ZN(n5632) );
  INV_X1 U6203 ( .A(n5335), .ZN(n4994) );
  XNOR2_X1 U6204 ( .A(n4995), .B(SI_15_), .ZN(n5335) );
  NOR2_X1 U6205 ( .A1(n5614), .A2(n7437), .ZN(n4921) );
  AND2_X1 U6206 ( .A1(n9153), .A2(n9976), .ZN(n4922) );
  AND2_X1 U6207 ( .A1(n9154), .A2(n9149), .ZN(n4923) );
  AND2_X1 U6208 ( .A1(n6424), .A2(n8917), .ZN(n4924) );
  NAND2_X1 U6209 ( .A1(n6619), .A2(n6622), .ZN(n4925) );
  AND2_X1 U6210 ( .A1(n8273), .A2(n8281), .ZN(n4926) );
  NAND2_X1 U6211 ( .A1(n5395), .A2(n5366), .ZN(n4927) );
  AND2_X1 U6212 ( .A1(n6223), .A2(n6222), .ZN(n4928) );
  NAND2_X1 U6213 ( .A1(n5496), .A2(n5495), .ZN(n8403) );
  AOI21_X1 U6214 ( .B1(n7247), .B2(n8940), .A(n8939), .ZN(n8941) );
  OR2_X1 U6215 ( .A1(n8293), .A2(n8298), .ZN(n8294) );
  NAND2_X1 U6216 ( .A1(n8297), .A2(n8304), .ZN(n8305) );
  NAND2_X1 U6217 ( .A1(n9096), .A2(n9044), .ZN(n9005) );
  OAI211_X1 U6218 ( .C1(n9023), .C2(n9022), .A(n9078), .B(n9021), .ZN(n9024)
         );
  INV_X1 U6219 ( .A(n8359), .ZN(n6678) );
  INV_X1 U6220 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6221 ( .A1(n9100), .A2(n9019), .ZN(n9020) );
  NAND2_X1 U6222 ( .A1(n8196), .A2(n8359), .ZN(n6680) );
  AND2_X1 U6223 ( .A1(n7081), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U6224 ( .A1(n8523), .A2(n5757), .ZN(n8204) );
  OR2_X1 U6225 ( .A1(n6334), .A2(n8851), .ZN(n6336) );
  OR2_X1 U6226 ( .A1(n5410), .A2(n5414), .ZN(n5022) );
  INV_X1 U6227 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6500) );
  INV_X1 U6228 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6459) );
  NOR2_X1 U6229 ( .A1(n7850), .A2(n7752), .ZN(n6259) );
  AND2_X1 U6230 ( .A1(n8882), .A2(n6336), .ZN(n6335) );
  OR2_X1 U6231 ( .A1(n9015), .A2(n9070), .ZN(n5515) );
  OR2_X1 U6232 ( .A1(n5499), .A2(n9045), .ZN(n8398) );
  AND2_X1 U6233 ( .A1(n5348), .A2(n4984), .ZN(n4985) );
  INV_X1 U6234 ( .A(n8335), .ZN(n8173) );
  OR2_X1 U6235 ( .A1(n6261), .A2(n7848), .ZN(n6264) );
  OAI21_X1 U6236 ( .B1(n8374), .B2(n8373), .A(n6353), .ZN(n6354) );
  NAND2_X1 U6237 ( .A1(n9125), .A2(n5655), .ZN(n9126) );
  INV_X1 U6238 ( .A(n5459), .ZN(n5096) );
  OR2_X1 U6239 ( .A1(n5487), .A2(n5486), .ZN(n5505) );
  INV_X1 U6240 ( .A(n5388), .ZN(n5092) );
  INV_X1 U6241 ( .A(n7929), .ZN(n5623) );
  INV_X1 U6242 ( .A(n7759), .ZN(n5658) );
  INV_X1 U6243 ( .A(n8081), .ZN(n5657) );
  INV_X1 U6244 ( .A(n5024), .ZN(n5025) );
  AND2_X1 U6245 ( .A1(n5380), .A2(n5382), .ZN(n5020) );
  OAI21_X1 U6246 ( .B1(n10168), .B2(n7737), .A(n10169), .ZN(n6547) );
  NAND2_X1 U6247 ( .A1(n8608), .A2(n10248), .ZN(n8609) );
  OR2_X1 U6248 ( .A1(n8048), .A2(n8720), .ZN(n8281) );
  INV_X1 U6249 ( .A(n6497), .ZN(n5961) );
  AND2_X1 U6250 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  INV_X1 U6251 ( .A(n5357), .ZN(n5091) );
  INV_X1 U6252 ( .A(n6354), .ZN(n6355) );
  OR2_X1 U6253 ( .A1(n6376), .A2(n6375), .ZN(n6468) );
  INV_X1 U6254 ( .A(n5341), .ZN(n5090) );
  OR2_X1 U6255 ( .A1(n5472), .A2(n9904), .ZN(n5487) );
  NAND2_X1 U6256 ( .A1(n5095), .A2(n5094), .ZN(n5459) );
  INV_X1 U6257 ( .A(n9464), .ZN(n9579) );
  NAND2_X1 U6258 ( .A1(n5092), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5406) );
  AND2_X1 U6259 ( .A1(n5262), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5275) );
  OR2_X1 U6260 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  INV_X1 U6261 ( .A(n8607), .ZN(n8497) );
  OR2_X1 U6262 ( .A1(n6020), .A2(n6012), .ZN(n8617) );
  AND2_X1 U6263 ( .A1(n6460), .A2(n4916), .ZN(n6461) );
  INV_X1 U6264 ( .A(n8725), .ZN(n8696) );
  AND2_X1 U6265 ( .A1(n6048), .A2(n6047), .ZN(n8340) );
  OR2_X1 U6266 ( .A1(n8764), .A2(n8696), .ZN(n8276) );
  AND2_X1 U6267 ( .A1(n8281), .A2(n8274), .ZN(n8033) );
  INV_X1 U6268 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7988) );
  OR2_X1 U6269 ( .A1(n5325), .A2(n5324), .ZN(n5341) );
  NAND2_X1 U6270 ( .A1(n8369), .A2(n8371), .ZN(n8372) );
  OR2_X1 U6271 ( .A1(n6206), .A2(n6388), .ZN(n6207) );
  NAND2_X1 U6272 ( .A1(n5091), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5372) );
  OR2_X1 U6273 ( .A1(n5209), .A2(n6972), .ZN(n5263) );
  NAND2_X1 U6274 ( .A1(n7858), .A2(n7859), .ZN(n7857) );
  NAND2_X1 U6275 ( .A1(n5090), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5357) );
  INV_X1 U6276 ( .A(n9039), .ZN(n9183) );
  OR2_X1 U6277 ( .A1(n5429), .A2(n8852), .ZN(n5448) );
  INV_X1 U6278 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9253) );
  OR2_X1 U6279 ( .A1(n9334), .A2(n9335), .ZN(n9359) );
  XNOR2_X1 U6280 ( .A(n9402), .B(n8931), .ZN(n6660) );
  INV_X1 U6281 ( .A(n9564), .ZN(n9025) );
  AOI21_X1 U6282 ( .B1(n5150), .B2(n8935), .A(n5149), .ZN(n7673) );
  INV_X1 U6283 ( .A(n9627), .ZN(n6629) );
  XNOR2_X1 U6284 ( .A(n4970), .B(SI_10_), .ZN(n5252) );
  NAND2_X1 U6285 ( .A1(n4955), .A2(SI_6_), .ZN(n4956) );
  AOI21_X1 U6286 ( .B1(n8617), .B2(n5824), .A(n6016), .ZN(n8628) );
  AND4_X1 U6287 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n8708)
         );
  AND2_X1 U6288 ( .A1(n8320), .A2(n8321), .ZN(n8318) );
  INV_X1 U6289 ( .A(n8601), .ZN(n8728) );
  NAND2_X1 U6290 ( .A1(n6673), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6614) );
  INV_X1 U6291 ( .A(n8340), .ZN(n8781) );
  INV_X1 U6292 ( .A(n8469), .ZN(n8791) );
  AND2_X1 U6293 ( .A1(n7349), .A2(n8196), .ZN(n10314) );
  OAI21_X1 U6294 ( .B1(n9025), .B2(n8928), .A(n6492), .ZN(n6493) );
  AND2_X1 U6295 ( .A1(n6425), .A2(n4924), .ZN(n6406) );
  NAND2_X1 U6296 ( .A1(n5428), .A2(n5427), .ZN(n9597) );
  AOI21_X1 U6297 ( .B1(n7043), .B2(n7042), .A(n4928), .ZN(n7062) );
  OR2_X1 U6298 ( .A1(n6412), .A2(n5530), .ZN(n5113) );
  OR2_X1 U6299 ( .A1(n5340), .A2(n5151), .ZN(n5153) );
  INV_X1 U6300 ( .A(n5640), .ZN(n9510) );
  INV_X1 U6301 ( .A(n9467), .ZN(n10015) );
  AND2_X1 U6302 ( .A1(n5598), .A2(n5554), .ZN(n9982) );
  AND2_X1 U6303 ( .A1(n5603), .A2(n9994), .ZN(n5604) );
  NAND2_X1 U6304 ( .A1(n5418), .A2(n5417), .ZN(n9530) );
  AND2_X1 U6305 ( .A1(n9125), .A2(n6415), .ZN(n10084) );
  XNOR2_X1 U6306 ( .A(n4954), .B(SI_6_), .ZN(n5245) );
  AND2_X1 U6307 ( .A1(n6723), .A2(n6722), .ZN(n8488) );
  INV_X1 U6308 ( .A(n8627), .ZN(n8657) );
  INV_X1 U6309 ( .A(n8111), .ZN(n8682) );
  AND2_X1 U6310 ( .A1(n6140), .A2(n8711), .ZN(n10260) );
  NAND2_X1 U6311 ( .A1(n8741), .A2(n8740), .ZN(n8743) );
  INV_X1 U6312 ( .A(n8598), .ZN(n8773) );
  OR2_X1 U6313 ( .A1(n10317), .A2(n10309), .ZN(n8832) );
  AND2_X1 U6314 ( .A1(n6157), .A2(n6156), .ZN(n10317) );
  AND2_X1 U6315 ( .A1(n6101), .A2(n6787), .ZN(n6785) );
  INV_X1 U6316 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U6317 ( .A1(n6488), .A2(n6406), .ZN(n6429) );
  INV_X1 U6318 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U6319 ( .A1(n5113), .A2(n5112), .ZN(n9193) );
  OR2_X1 U6320 ( .A1(n5604), .A2(n5401), .ZN(n9467) );
  INV_X2 U6321 ( .A(n5604), .ZN(n9989) );
  OR2_X1 U6322 ( .A1(n9036), .A2(n9936), .ZN(n6666) );
  INV_X1 U6323 ( .A(n9530), .ZN(n9931) );
  INV_X1 U6324 ( .A(n7908), .ZN(n8868) );
  INV_X1 U6325 ( .A(n5107), .ZN(n7868) );
  INV_X1 U6326 ( .A(n5653), .ZN(n8088) );
  NAND2_X1 U6327 ( .A1(n6144), .A2(n6143), .ZN(P2_U3205) );
  NAND2_X1 U6328 ( .A1(n6445), .A2(n6444), .ZN(P2_U3454) );
  OAI21_X1 U6329 ( .B1(n9561), .B2(n5604), .A(n5668), .ZN(P1_U3356) );
  INV_X1 U6330 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6758) );
  INV_X1 U6331 ( .A(n6763), .ZN(n4930) );
  INV_X1 U6332 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6333 ( .A1(n4930), .A2(n4929), .ZN(n4931) );
  AND2_X1 U6334 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6335 ( .A1(n6763), .A2(n4933), .ZN(n5740) );
  NAND2_X1 U6336 ( .A1(n4934), .A2(n5740), .ZN(n5116) );
  INV_X1 U6337 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6338 ( .A1(n4936), .A2(SI_1_), .ZN(n4937) );
  INV_X1 U6339 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6759) );
  INV_X1 U6340 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U6341 ( .A1(n5146), .A2(n5145), .ZN(n4942) );
  INV_X1 U6342 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U6343 ( .A1(n4940), .A2(SI_2_), .ZN(n4941) );
  NAND2_X1 U6344 ( .A1(n4942), .A2(n4941), .ZN(n5157) );
  MUX2_X1 U6345 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5043), .Z(n4944) );
  INV_X1 U6346 ( .A(SI_3_), .ZN(n4943) );
  NAND2_X1 U6347 ( .A1(n5157), .A2(n5156), .ZN(n4946) );
  NAND2_X1 U6348 ( .A1(n4944), .A2(SI_3_), .ZN(n4945) );
  NAND2_X1 U6349 ( .A1(n4946), .A2(n4945), .ZN(n5170) );
  INV_X1 U6350 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6768) );
  INV_X1 U6351 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6767) );
  MUX2_X1 U6352 ( .A(n6768), .B(n6767), .S(n5043), .Z(n4947) );
  NAND2_X1 U6353 ( .A1(n5170), .A2(n5171), .ZN(n4950) );
  INV_X1 U6354 ( .A(n4947), .ZN(n4948) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6773) );
  MUX2_X1 U6356 ( .A(n9803), .B(n6773), .S(n5043), .Z(n4951) );
  INV_X1 U6357 ( .A(n4951), .ZN(n4952) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6776) );
  INV_X1 U6359 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6778) );
  MUX2_X1 U6360 ( .A(n6776), .B(n6778), .S(n5043), .Z(n4954) );
  INV_X1 U6361 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6362 ( .A1(n4957), .A2(n4956), .ZN(n5227) );
  INV_X1 U6363 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6781) );
  INV_X1 U6364 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6783) );
  MUX2_X1 U6365 ( .A(n6781), .B(n6783), .S(n5043), .Z(n4958) );
  INV_X1 U6366 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U6367 ( .A1(n4959), .A2(SI_7_), .ZN(n4960) );
  INV_X1 U6368 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6798) );
  INV_X1 U6369 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6797) );
  MUX2_X1 U6370 ( .A(n6798), .B(n6797), .S(n5043), .Z(n4961) );
  INV_X1 U6371 ( .A(SI_8_), .ZN(n9745) );
  INV_X1 U6372 ( .A(n4961), .ZN(n4962) );
  NAND2_X1 U6373 ( .A1(n4962), .A2(SI_8_), .ZN(n4963) );
  INV_X1 U6374 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6811) );
  INV_X1 U6375 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6813) );
  MUX2_X1 U6376 ( .A(n6811), .B(n6813), .S(n5043), .Z(n4966) );
  INV_X1 U6377 ( .A(SI_9_), .ZN(n4965) );
  INV_X1 U6378 ( .A(n4966), .ZN(n4967) );
  NAND2_X1 U6379 ( .A1(n4967), .A2(SI_9_), .ZN(n4968) );
  NAND2_X1 U6380 ( .A1(n5195), .A2(n4969), .ZN(n5253) );
  INV_X1 U6381 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6831) );
  INV_X1 U6382 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6815) );
  MUX2_X1 U6383 ( .A(n6831), .B(n6815), .S(n5043), .Z(n4970) );
  INV_X1 U6384 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6385 ( .A1(n4971), .A2(SI_10_), .ZN(n4972) );
  INV_X1 U6386 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6867) );
  INV_X1 U6387 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6870) );
  MUX2_X1 U6388 ( .A(n6867), .B(n6870), .S(n5043), .Z(n4974) );
  INV_X1 U6389 ( .A(SI_11_), .ZN(n4973) );
  NAND2_X1 U6390 ( .A1(n4974), .A2(n4973), .ZN(n4977) );
  INV_X1 U6391 ( .A(n4974), .ZN(n4975) );
  NAND2_X1 U6392 ( .A1(n4975), .A2(SI_11_), .ZN(n4976) );
  NAND2_X1 U6393 ( .A1(n4977), .A2(n4976), .ZN(n5269) );
  INV_X1 U6394 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7005) );
  INV_X1 U6395 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4978) );
  MUX2_X1 U6396 ( .A(n7005), .B(n4978), .S(n5043), .Z(n4979) );
  INV_X1 U6397 ( .A(n4979), .ZN(n4980) );
  MUX2_X1 U6398 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5043), .Z(n4986) );
  XNOR2_X1 U6399 ( .A(n4986), .B(SI_13_), .ZN(n5301) );
  INV_X1 U6400 ( .A(n5301), .ZN(n5315) );
  INV_X1 U6401 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7113) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7112) );
  MUX2_X1 U6403 ( .A(n7113), .B(n7112), .S(n5043), .Z(n4987) );
  INV_X1 U6404 ( .A(SI_14_), .ZN(n4981) );
  NAND2_X1 U6405 ( .A1(n4987), .A2(n4981), .ZN(n4990) );
  AND2_X1 U6406 ( .A1(n5315), .A2(n4990), .ZN(n5334) );
  INV_X1 U6407 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n4983) );
  INV_X1 U6408 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4982) );
  MUX2_X1 U6409 ( .A(n4983), .B(n4982), .S(n5043), .Z(n4995) );
  MUX2_X1 U6410 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4401), .Z(n4999) );
  INV_X1 U6411 ( .A(n5352), .ZN(n4984) );
  INV_X1 U6412 ( .A(n4990), .ZN(n4993) );
  NAND2_X1 U6413 ( .A1(n4986), .A2(SI_13_), .ZN(n5316) );
  INV_X1 U6414 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6415 ( .A1(n4988), .A2(SI_14_), .ZN(n4989) );
  INV_X1 U6416 ( .A(n4995), .ZN(n4996) );
  NAND2_X1 U6417 ( .A1(n4996), .A2(SI_15_), .ZN(n4997) );
  NAND2_X1 U6418 ( .A1(n4999), .A2(SI_16_), .ZN(n5000) );
  INV_X1 U6419 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7190) );
  INV_X1 U6420 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5002) );
  MUX2_X1 U6421 ( .A(n7190), .B(n5002), .S(n5043), .Z(n5004) );
  INV_X1 U6422 ( .A(SI_17_), .ZN(n5003) );
  NAND2_X1 U6423 ( .A1(n5004), .A2(n5003), .ZN(n5380) );
  INV_X1 U6424 ( .A(n5004), .ZN(n5005) );
  NAND2_X1 U6425 ( .A1(n5005), .A2(SI_17_), .ZN(n5006) );
  NAND2_X1 U6426 ( .A1(n5380), .A2(n5006), .ZN(n5367) );
  INV_X1 U6427 ( .A(n5367), .ZN(n5007) );
  INV_X1 U6428 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7156) );
  INV_X1 U6429 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5008) );
  MUX2_X1 U6430 ( .A(n7156), .B(n5008), .S(n4402), .Z(n5019) );
  INV_X1 U6431 ( .A(n5019), .ZN(n5009) );
  NAND2_X1 U6432 ( .A1(n5009), .A2(SI_18_), .ZN(n5018) );
  INV_X1 U6433 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7184) );
  INV_X1 U6434 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8421) );
  MUX2_X1 U6435 ( .A(n7184), .B(n8421), .S(n4401), .Z(n5010) );
  INV_X1 U6436 ( .A(SI_19_), .ZN(n9878) );
  NAND2_X1 U6437 ( .A1(n5010), .A2(n9878), .ZN(n5412) );
  INV_X1 U6438 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6439 ( .A1(n5011), .A2(SI_19_), .ZN(n5012) );
  NAND2_X1 U6440 ( .A1(n5412), .A2(n5012), .ZN(n5410) );
  INV_X1 U6441 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7228) );
  INV_X1 U6442 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7206) );
  MUX2_X1 U6443 ( .A(n7228), .B(n7206), .S(n4402), .Z(n5014) );
  INV_X1 U6444 ( .A(SI_20_), .ZN(n5013) );
  NAND2_X1 U6445 ( .A1(n5014), .A2(n5013), .ZN(n5024) );
  INV_X1 U6446 ( .A(n5014), .ZN(n5015) );
  NAND2_X1 U6447 ( .A1(n5015), .A2(SI_20_), .ZN(n5016) );
  NAND2_X1 U6448 ( .A1(n5024), .A2(n5016), .ZN(n5414) );
  INV_X1 U6449 ( .A(n5022), .ZN(n5017) );
  INV_X1 U6450 ( .A(n5018), .ZN(n5021) );
  XNOR2_X1 U6451 ( .A(n5019), .B(SI_18_), .ZN(n5382) );
  INV_X1 U6452 ( .A(n5426), .ZN(n5028) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7300) );
  INV_X1 U6454 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9902) );
  MUX2_X1 U6455 ( .A(n7300), .B(n9902), .S(n5043), .Z(n5029) );
  XNOR2_X1 U6456 ( .A(n5029), .B(SI_21_), .ZN(n5425) );
  INV_X1 U6457 ( .A(n5029), .ZN(n5030) );
  NAND2_X1 U6458 ( .A1(n5030), .A2(SI_21_), .ZN(n5031) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7348) );
  INV_X1 U6460 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8090) );
  MUX2_X1 U6461 ( .A(n7348), .B(n8090), .S(n4401), .Z(n5034) );
  INV_X1 U6462 ( .A(SI_22_), .ZN(n5033) );
  NAND2_X1 U6463 ( .A1(n5034), .A2(n5033), .ZN(n5037) );
  INV_X1 U6464 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6465 ( .A1(n5035), .A2(SI_22_), .ZN(n5036) );
  NAND2_X1 U6466 ( .A1(n5037), .A2(n5036), .ZN(n5433) );
  INV_X1 U6467 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7392) );
  INV_X1 U6468 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9710) );
  MUX2_X1 U6469 ( .A(n7392), .B(n9710), .S(n4402), .Z(n5038) );
  INV_X1 U6470 ( .A(SI_23_), .ZN(n9835) );
  NAND2_X1 U6471 ( .A1(n5038), .A2(n9835), .ZN(n5041) );
  INV_X1 U6472 ( .A(n5038), .ZN(n5039) );
  NAND2_X1 U6473 ( .A1(n5039), .A2(SI_23_), .ZN(n5040) );
  AND2_X1 U6474 ( .A1(n5041), .A2(n5040), .ZN(n5442) );
  NAND2_X1 U6475 ( .A1(n5443), .A2(n5442), .ZN(n5042) );
  INV_X1 U6476 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8416) );
  INV_X1 U6477 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7469) );
  MUX2_X1 U6478 ( .A(n8416), .B(n7469), .S(n5043), .Z(n5045) );
  INV_X1 U6479 ( .A(SI_24_), .ZN(n5044) );
  NAND2_X1 U6480 ( .A1(n5045), .A2(n5044), .ZN(n5048) );
  INV_X1 U6481 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6482 ( .A1(n5046), .A2(SI_24_), .ZN(n5047) );
  AND2_X1 U6483 ( .A1(n5048), .A2(n5047), .ZN(n5455) );
  NAND2_X1 U6484 ( .A1(n5456), .A2(n5455), .ZN(n5049) );
  INV_X1 U6485 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9822) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9794) );
  MUX2_X1 U6487 ( .A(n9822), .B(n9794), .S(n4401), .Z(n5051) );
  INV_X1 U6488 ( .A(SI_25_), .ZN(n5050) );
  NAND2_X1 U6489 ( .A1(n5051), .A2(n5050), .ZN(n5054) );
  INV_X1 U6490 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6491 ( .A1(n5052), .A2(SI_25_), .ZN(n5053) );
  AND2_X1 U6492 ( .A1(n5054), .A2(n5053), .ZN(n5468) );
  INV_X1 U6493 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6017) );
  INV_X1 U6494 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7726) );
  MUX2_X1 U6495 ( .A(n6017), .B(n7726), .S(n4402), .Z(n5056) );
  INV_X1 U6496 ( .A(SI_26_), .ZN(n9834) );
  NAND2_X1 U6497 ( .A1(n5056), .A2(n9834), .ZN(n5059) );
  INV_X1 U6498 ( .A(n5056), .ZN(n5057) );
  NAND2_X1 U6499 ( .A1(n5057), .A2(SI_26_), .ZN(n5058) );
  AND2_X1 U6500 ( .A1(n5059), .A2(n5058), .ZN(n5480) );
  INV_X1 U6501 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6028) );
  INV_X1 U6502 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7775) );
  MUX2_X1 U6503 ( .A(n6028), .B(n7775), .S(n5043), .Z(n5061) );
  INV_X1 U6504 ( .A(SI_27_), .ZN(n5060) );
  NAND2_X1 U6505 ( .A1(n5061), .A2(n5060), .ZN(n5519) );
  INV_X1 U6506 ( .A(n5061), .ZN(n5062) );
  NAND2_X1 U6507 ( .A1(n5062), .A2(SI_27_), .ZN(n5063) );
  AND2_X1 U6508 ( .A1(n5519), .A2(n5063), .ZN(n5500) );
  NAND2_X1 U6509 ( .A1(n5521), .A2(n5519), .ZN(n5068) );
  INV_X1 U6510 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6046) );
  INV_X1 U6511 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7802) );
  MUX2_X1 U6512 ( .A(n6046), .B(n7802), .S(n4401), .Z(n5065) );
  INV_X1 U6513 ( .A(SI_28_), .ZN(n5064) );
  NAND2_X1 U6514 ( .A1(n5065), .A2(n5064), .ZN(n5518) );
  INV_X1 U6515 ( .A(n5065), .ZN(n5066) );
  NAND2_X1 U6516 ( .A1(n5066), .A2(SI_28_), .ZN(n5522) );
  AND2_X1 U6517 ( .A1(n5518), .A2(n5522), .ZN(n5067) );
  INV_X1 U6518 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5072) );
  AND2_X1 U6519 ( .A1(n5072), .A2(n5081), .ZN(n5077) );
  NOR2_X1 U6520 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5074) );
  INV_X1 U6521 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5564) );
  INV_X1 U6522 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5073) );
  NAND4_X1 U6523 ( .A1(n5074), .A2(n5564), .A3(n5540), .A4(n5073), .ZN(n5076)
         );
  INV_X1 U6524 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9802) );
  NAND4_X1 U6525 ( .A1(n5542), .A2(n9802), .A3(n5549), .A4(n5399), .ZN(n5075)
         );
  NOR2_X1 U6526 ( .A1(n5076), .A2(n5075), .ZN(n5079) );
  INV_X1 U6527 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5101) );
  XNOR2_X2 U6528 ( .A(n5078), .B(n5101), .ZN(n5554) );
  INV_X1 U6529 ( .A(n5079), .ZN(n5080) );
  NOR2_X1 U6530 ( .A1(n5085), .A2(n5084), .ZN(n5086) );
  NAND2_X1 U6531 ( .A1(n7741), .A2(n6648), .ZN(n5089) );
  OR2_X1 U6532 ( .A1(n6649), .A2(n7802), .ZN(n5088) );
  NAND2_X1 U6533 ( .A1(n5206), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5209) );
  INV_X1 U6534 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6972) );
  INV_X1 U6535 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7755) );
  INV_X1 U6536 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5306) );
  INV_X1 U6537 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5324) );
  INV_X1 U6538 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8873) );
  INV_X1 U6539 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8842) );
  INV_X1 U6540 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8852) );
  AND2_X1 U6541 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5094) );
  INV_X1 U6542 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9904) );
  INV_X1 U6543 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5486) );
  INV_X1 U6544 ( .A(n5505), .ZN(n5097) );
  NAND2_X1 U6545 ( .A1(n5097), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5507) );
  INV_X1 U6546 ( .A(n5507), .ZN(n5098) );
  NAND2_X1 U6547 ( .A1(n5098), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5661) );
  INV_X1 U6548 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6549 ( .A1(n5507), .A2(n5099), .ZN(n5100) );
  NAND2_X1 U6550 ( .A1(n5661), .A2(n5100), .ZN(n6412) );
  OR2_X2 U6551 ( .A1(n5103), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n7994) );
  NAND2_X2 U6552 ( .A1(n7994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5102) );
  XNOR2_X2 U6553 ( .A(n5102), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6554 ( .A1(n5103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5104) );
  MUX2_X1 U6555 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5104), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5105) );
  INV_X1 U6556 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5110) );
  NAND2_X2 U6557 ( .A1(n8092), .A2(n7868), .ZN(n5340) );
  INV_X2 U6558 ( .A(n5340), .ZN(n5490) );
  NAND2_X1 U6559 ( .A1(n5490), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5109) );
  AND2_X2 U6560 ( .A1(n8092), .A2(n5107), .ZN(n5174) );
  NAND2_X1 U6561 ( .A1(n5174), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5108) );
  OAI211_X1 U6562 ( .C1(n5110), .C2(n5125), .A(n5109), .B(n5108), .ZN(n5111)
         );
  INV_X1 U6563 ( .A(n5111), .ZN(n5112) );
  INV_X1 U6564 ( .A(n9193), .ZN(n5517) );
  NAND2_X1 U6565 ( .A1(n9026), .A2(n5517), .ZN(n9091) );
  INV_X1 U6566 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6567 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5114) );
  XNOR2_X1 U6568 ( .A(n5117), .B(n5116), .ZN(n6764) );
  NAND2_X1 U6569 ( .A1(n5135), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5121) );
  INV_X1 U6570 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6571 ( .A1(n5489), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5119) );
  INV_X1 U6572 ( .A(n5607), .ZN(n5133) );
  NAND2_X1 U6573 ( .A1(n5489), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6574 ( .A1(n5174), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5129) );
  INV_X1 U6575 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5124) );
  OR2_X1 U6576 ( .A1(n5125), .A2(n5124), .ZN(n5128) );
  INV_X1 U6577 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5126) );
  OR2_X1 U6578 ( .A1(n5340), .A2(n5126), .ZN(n5127) );
  INV_X1 U6579 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9218) );
  INV_X1 U6580 ( .A(SI_0_), .ZN(n5131) );
  NOR2_X1 U6581 ( .A1(n6763), .A2(n5131), .ZN(n5132) );
  XNOR2_X1 U6582 ( .A(n5132), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U6583 ( .A(n9218), .B(n9942), .S(n6794), .Z(n8082) );
  INV_X1 U6584 ( .A(n8082), .ZN(n7511) );
  AND2_X1 U6585 ( .A1(n7135), .A2(n7511), .ZN(n6937) );
  NAND2_X1 U6586 ( .A1(n5133), .A2(n6937), .ZN(n8075) );
  INV_X1 U6587 ( .A(n9211), .ZN(n7148) );
  NAND2_X1 U6588 ( .A1(n7148), .A2(n7133), .ZN(n5134) );
  NAND2_X1 U6589 ( .A1(n8075), .A2(n5134), .ZN(n7174) );
  INV_X1 U6590 ( .A(n7174), .ZN(n5150) );
  NAND2_X1 U6591 ( .A1(n5489), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6592 ( .A1(n5174), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6593 ( .A1(n5508), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6594 ( .A1(n5490), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5136) );
  MUX2_X1 U6595 ( .A(n7993), .B(n5141), .S(P1_IR_REG_2__SCAN_IN), .Z(n5142) );
  INV_X1 U6596 ( .A(n5142), .ZN(n5144) );
  INV_X1 U6597 ( .A(n5183), .ZN(n5143) );
  INV_X1 U6598 ( .A(n6848), .ZN(n9955) );
  XNOR2_X1 U6599 ( .A(n5146), .B(n5145), .ZN(n6771) );
  OR2_X1 U6600 ( .A1(n5147), .A2(n6771), .ZN(n5148) );
  OAI211_X1 U6601 ( .C1(n6794), .C2(n9955), .A(n5148), .B(n4429), .ZN(n7645)
         );
  NAND2_X1 U6602 ( .A1(n7044), .A2(n7645), .ZN(n8935) );
  NAND2_X1 U6603 ( .A1(n9209), .A2(n7186), .ZN(n9135) );
  INV_X1 U6604 ( .A(n9135), .ZN(n5149) );
  NAND2_X1 U6605 ( .A1(n5174), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6606 ( .A1(n5508), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5154) );
  INV_X1 U6607 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5151) );
  INV_X1 U6608 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U6609 ( .A1(n5489), .A2(n7681), .ZN(n5152) );
  OR2_X1 U6610 ( .A1(n5183), .A2(n7993), .ZN(n5167) );
  XNOR2_X1 U6611 ( .A(n5167), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6847) );
  INV_X1 U6612 ( .A(n6847), .ZN(n9227) );
  XNOR2_X1 U6613 ( .A(n5157), .B(n5156), .ZN(n6765) );
  OR2_X1 U6614 ( .A1(n5147), .A2(n6765), .ZN(n5159) );
  INV_X1 U6615 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6766) );
  OR2_X1 U6616 ( .A1(n6649), .A2(n6766), .ZN(n5158) );
  OAI211_X1 U6617 ( .C1(n6794), .C2(n9227), .A(n5159), .B(n5158), .ZN(n7682)
         );
  INV_X1 U6618 ( .A(n7682), .ZN(n10067) );
  NAND2_X1 U6619 ( .A1(n9208), .A2(n10067), .ZN(n9134) );
  INV_X1 U6620 ( .A(n8936), .ZN(n9049) );
  NAND2_X1 U6621 ( .A1(n7673), .A2(n9049), .ZN(n7672) );
  NAND2_X1 U6622 ( .A1(n7672), .A2(n9139), .ZN(n7247) );
  NAND2_X1 U6623 ( .A1(n5490), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6624 ( .A1(n5174), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5165) );
  INV_X1 U6625 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6626 ( .A1(n7681), .A2(n5160), .ZN(n5162) );
  INV_X1 U6627 ( .A(n5161), .ZN(n5176) );
  AND2_X1 U6628 ( .A1(n5162), .A2(n5176), .ZN(n7059) );
  NAND2_X1 U6629 ( .A1(n5489), .A2(n7059), .ZN(n5164) );
  NAND2_X1 U6630 ( .A1(n5508), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5163) );
  NAND4_X1 U6631 ( .A1(n5166), .A2(n5165), .A3(n5164), .A4(n5163), .ZN(n9207)
         );
  INV_X1 U6632 ( .A(n9207), .ZN(n7235) );
  NAND2_X1 U6633 ( .A1(n5167), .A2(n9795), .ZN(n5168) );
  NAND2_X1 U6634 ( .A1(n5168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6635 ( .A(n5169), .B(n4711), .ZN(n6914) );
  XNOR2_X1 U6636 ( .A(n5170), .B(n5171), .ZN(n6769) );
  OR2_X1 U6637 ( .A1(n5147), .A2(n6769), .ZN(n5173) );
  OR2_X1 U6638 ( .A1(n6649), .A2(n6767), .ZN(n5172) );
  OAI211_X1 U6639 ( .C1(n6794), .C2(n6914), .A(n5173), .B(n5172), .ZN(n6199)
         );
  NAND2_X1 U6640 ( .A1(n7235), .A2(n6199), .ZN(n8946) );
  NAND2_X1 U6641 ( .A1(n9207), .A2(n7609), .ZN(n8940) );
  NAND2_X1 U6642 ( .A1(n8946), .A2(n8940), .ZN(n9051) );
  INV_X1 U6643 ( .A(n9051), .ZN(n7249) );
  NAND2_X1 U6644 ( .A1(n7247), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U6645 ( .A1(n7248), .A2(n8946), .ZN(n7233) );
  NAND2_X1 U6646 ( .A1(n5490), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6647 ( .A1(n5174), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5180) );
  INV_X1 U6648 ( .A(n5175), .ZN(n5236) );
  INV_X1 U6649 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9739) );
  NAND2_X1 U6650 ( .A1(n5176), .A2(n9739), .ZN(n5177) );
  AND2_X1 U6651 ( .A1(n5236), .A2(n5177), .ZN(n7663) );
  NAND2_X1 U6652 ( .A1(n5489), .A2(n7663), .ZN(n5179) );
  NAND2_X1 U6653 ( .A1(n5508), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5178) );
  NAND4_X1 U6654 ( .A1(n5181), .A2(n5180), .A3(n5179), .A4(n5178), .ZN(n9206)
         );
  INV_X1 U6655 ( .A(n9206), .ZN(n7293) );
  NOR2_X1 U6656 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5182) );
  NAND2_X1 U6657 ( .A1(n5183), .A2(n5182), .ZN(n5184) );
  NOR2_X1 U6658 ( .A1(n5184), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5243) );
  INV_X1 U6659 ( .A(n5243), .ZN(n5187) );
  NAND2_X1 U6660 ( .A1(n5184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5185) );
  MUX2_X1 U6661 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5185), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5186) );
  INV_X1 U6662 ( .A(n6963), .ZN(n6958) );
  XNOR2_X1 U6663 ( .A(n5189), .B(n5188), .ZN(n6772) );
  OR2_X1 U6664 ( .A1(n5147), .A2(n6772), .ZN(n5191) );
  OR2_X1 U6665 ( .A1(n6649), .A2(n6773), .ZN(n5190) );
  OAI211_X1 U6666 ( .C1(n6794), .C2(n6958), .A(n5191), .B(n5190), .ZN(n7664)
         );
  NAND2_X1 U6667 ( .A1(n7293), .A2(n7664), .ZN(n8945) );
  NAND2_X1 U6668 ( .A1(n9206), .A2(n7264), .ZN(n9141) );
  NAND2_X1 U6669 ( .A1(n8945), .A2(n9141), .ZN(n9052) );
  INV_X1 U6670 ( .A(n9052), .ZN(n7234) );
  NAND2_X1 U6671 ( .A1(n7233), .A2(n7234), .ZN(n7232) );
  NAND2_X1 U6672 ( .A1(n6810), .A2(n6648), .ZN(n5199) );
  NAND2_X1 U6673 ( .A1(n5243), .A2(n5196), .ZN(n5216) );
  NAND2_X1 U6674 ( .A1(n5254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5197) );
  XNOR2_X1 U6675 ( .A(n5197), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7089) );
  AOI22_X1 U6676 ( .A1(n5403), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5402), .B2(
        n7089), .ZN(n5198) );
  NAND2_X2 U6677 ( .A1(n5199), .A2(n5198), .ZN(n7577) );
  NAND2_X1 U6678 ( .A1(n5490), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6679 ( .A1(n5234), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6680 ( .A1(n5209), .A2(n6972), .ZN(n5201) );
  AND2_X1 U6681 ( .A1(n5263), .A2(n5201), .ZN(n7617) );
  NAND2_X1 U6682 ( .A1(n5489), .A2(n7617), .ZN(n5203) );
  NAND2_X1 U6683 ( .A1(n5508), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5202) );
  NAND4_X1 U6684 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n9202)
         );
  INV_X1 U6685 ( .A(n9202), .ZN(n7590) );
  OR2_X2 U6686 ( .A1(n7577), .A2(n7590), .ZN(n8968) );
  NAND2_X1 U6687 ( .A1(n5490), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6688 ( .A1(n5234), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5212) );
  INV_X1 U6689 ( .A(n5206), .ZN(n5221) );
  INV_X1 U6690 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6691 ( .A1(n5221), .A2(n5207), .ZN(n5208) );
  AND2_X1 U6692 ( .A1(n5209), .A2(n5208), .ZN(n7598) );
  NAND2_X1 U6693 ( .A1(n5489), .A2(n7598), .ZN(n5211) );
  NAND2_X1 U6694 ( .A1(n5508), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5210) );
  NAND4_X1 U6695 ( .A1(n5213), .A2(n5212), .A3(n5211), .A4(n5210), .ZN(n9203)
         );
  INV_X1 U6696 ( .A(n9203), .ZN(n7572) );
  XNOR2_X1 U6697 ( .A(n5215), .B(n5214), .ZN(n6796) );
  NAND2_X1 U6698 ( .A1(n6796), .A2(n6648), .ZN(n5219) );
  NAND2_X1 U6699 ( .A1(n5216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6700 ( .A1(n5229), .A2(n5228), .ZN(n5231) );
  NAND2_X1 U6701 ( .A1(n5231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U6702 ( .A(n5217), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U6703 ( .A1(n5403), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5402), .B2(
        n6968), .ZN(n5218) );
  NAND2_X1 U6704 ( .A1(n5219), .A2(n5218), .ZN(n7585) );
  OR2_X1 U6705 ( .A1(n7572), .A2(n7585), .ZN(n8951) );
  NAND2_X1 U6706 ( .A1(n8968), .A2(n8951), .ZN(n8959) );
  NAND2_X1 U6707 ( .A1(n7585), .A2(n7572), .ZN(n8957) );
  NAND2_X1 U6708 ( .A1(n5490), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6709 ( .A1(n5234), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6710 ( .A1(n5238), .A2(n9253), .ZN(n5220) );
  AND2_X1 U6711 ( .A1(n5221), .A2(n5220), .ZN(n7638) );
  NAND2_X1 U6712 ( .A1(n5489), .A2(n7638), .ZN(n5223) );
  NAND2_X1 U6713 ( .A1(n5508), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5222) );
  NAND4_X1 U6714 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(n9204)
         );
  INV_X1 U6715 ( .A(n9204), .ZN(n7589) );
  XNOR2_X1 U6716 ( .A(n5227), .B(n5226), .ZN(n6782) );
  OR2_X1 U6717 ( .A1(n6782), .A2(n5147), .ZN(n5233) );
  OR2_X1 U6718 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  AND2_X1 U6719 ( .A1(n5231), .A2(n5230), .ZN(n6966) );
  AOI22_X1 U6720 ( .A1(n5403), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5402), .B2(
        n6966), .ZN(n5232) );
  NAND2_X1 U6721 ( .A1(n5233), .A2(n5232), .ZN(n7639) );
  NAND2_X1 U6722 ( .A1(n7589), .A2(n7639), .ZN(n7567) );
  AND2_X1 U6723 ( .A1(n8957), .A2(n7567), .ZN(n8950) );
  NAND2_X1 U6724 ( .A1(n7577), .A2(n7590), .ZN(n8962) );
  OAI21_X1 U6725 ( .B1(n8959), .B2(n8950), .A(n8962), .ZN(n5250) );
  NAND2_X1 U6726 ( .A1(n5490), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6727 ( .A1(n5234), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5241) );
  INV_X1 U6728 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6729 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  AND2_X1 U6730 ( .A1(n5238), .A2(n5237), .ZN(n10018) );
  NAND2_X1 U6731 ( .A1(n5489), .A2(n10018), .ZN(n5240) );
  NAND2_X1 U6732 ( .A1(n5508), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5239) );
  NAND4_X1 U6733 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), .ZN(n9205)
         );
  INV_X1 U6734 ( .A(n9205), .ZN(n7385) );
  OR2_X1 U6735 ( .A1(n5243), .A2(n7993), .ZN(n5244) );
  XNOR2_X1 U6736 ( .A(n5244), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6965) );
  INV_X1 U6737 ( .A(n6965), .ZN(n9240) );
  XNOR2_X1 U6738 ( .A(n5246), .B(n5245), .ZN(n6777) );
  OR2_X1 U6739 ( .A1(n6777), .A2(n5147), .ZN(n5248) );
  OR2_X1 U6740 ( .A1(n6649), .A2(n6778), .ZN(n5247) );
  NAND2_X1 U6741 ( .A1(n7385), .A2(n7436), .ZN(n8949) );
  INV_X1 U6742 ( .A(n8949), .ZN(n7565) );
  OR2_X1 U6743 ( .A1(n5250), .A2(n7565), .ZN(n9147) );
  NAND2_X1 U6744 ( .A1(n10073), .A2(n9204), .ZN(n8955) );
  NAND2_X1 U6745 ( .A1(n9205), .A2(n10023), .ZN(n8947) );
  AND2_X1 U6746 ( .A1(n8955), .A2(n8947), .ZN(n5249) );
  AND3_X1 U6747 ( .A1(n8968), .A2(n5249), .A3(n8951), .ZN(n9056) );
  OR2_X1 U6748 ( .A1(n5250), .A2(n9056), .ZN(n9145) );
  OAI21_X1 U6749 ( .B1(n7566), .B2(n9147), .A(n9145), .ZN(n5251) );
  XNOR2_X1 U6750 ( .A(n5253), .B(n5252), .ZN(n6814) );
  NAND2_X1 U6751 ( .A1(n6814), .A2(n6648), .ZN(n5261) );
  OR2_X1 U6752 ( .A1(n5254), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5255) );
  AND2_X1 U6753 ( .A1(n5255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6754 ( .A1(n5256), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5259) );
  INV_X1 U6755 ( .A(n5256), .ZN(n5258) );
  NAND2_X1 U6756 ( .A1(n5258), .A2(n5257), .ZN(n5271) );
  AND2_X1 U6757 ( .A1(n5259), .A2(n5271), .ZN(n7351) );
  AOI22_X1 U6758 ( .A1(n5403), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5402), .B2(
        n7351), .ZN(n5260) );
  NAND2_X1 U6759 ( .A1(n5490), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6760 ( .A1(n5234), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5267) );
  INV_X1 U6761 ( .A(n5262), .ZN(n5276) );
  NAND2_X1 U6762 ( .A1(n5263), .A2(n7755), .ZN(n5264) );
  AND2_X1 U6763 ( .A1(n5276), .A2(n5264), .ZN(n7758) );
  NAND2_X1 U6764 ( .A1(n5489), .A2(n7758), .ZN(n5266) );
  NAND2_X1 U6765 ( .A1(n5508), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5265) );
  NAND4_X1 U6766 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n9201)
         );
  INV_X1 U6767 ( .A(n9201), .ZN(n7564) );
  OR2_X1 U6768 ( .A1(n7759), .A2(n7564), .ZN(n9146) );
  NAND2_X1 U6769 ( .A1(n7759), .A2(n7564), .ZN(n9151) );
  NAND2_X1 U6770 ( .A1(n9146), .A2(n9151), .ZN(n7456) );
  INV_X1 U6771 ( .A(n7456), .ZN(n9054) );
  XNOR2_X1 U6772 ( .A(n5270), .B(n5269), .ZN(n6866) );
  NAND2_X1 U6773 ( .A1(n6866), .A2(n6648), .ZN(n5274) );
  NAND2_X1 U6774 ( .A1(n5271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5272) );
  XNOR2_X1 U6775 ( .A(n5272), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7357) );
  AOI22_X1 U6776 ( .A1(n5403), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5402), .B2(
        n7357), .ZN(n5273) );
  NAND2_X1 U6777 ( .A1(n5490), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6778 ( .A1(n5234), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5280) );
  INV_X1 U6779 ( .A(n5275), .ZN(n5293) );
  INV_X1 U6780 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U6781 ( .A1(n5276), .A2(n9280), .ZN(n5277) );
  AND2_X1 U6782 ( .A1(n5293), .A2(n5277), .ZN(n10006) );
  NAND2_X1 U6783 ( .A1(n5489), .A2(n10006), .ZN(n5279) );
  NAND2_X1 U6784 ( .A1(n5508), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5278) );
  NAND4_X1 U6785 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n9200)
         );
  XNOR2_X1 U6786 ( .A(n10008), .B(n9200), .ZN(n9046) );
  INV_X1 U6787 ( .A(n9200), .ZN(n8965) );
  NAND2_X1 U6788 ( .A1(n10008), .A2(n8965), .ZN(n9153) );
  NAND2_X1 U6789 ( .A1(n5282), .A2(n9153), .ZN(n7872) );
  NAND2_X1 U6790 ( .A1(n6986), .A2(n6648), .ZN(n5291) );
  NOR2_X1 U6791 ( .A1(n5285), .A2(n7993), .ZN(n5286) );
  MUX2_X1 U6792 ( .A(n7993), .B(n5286), .S(P1_IR_REG_12__SCAN_IN), .Z(n5289)
         );
  NOR2_X1 U6793 ( .A1(n5289), .A2(n4860), .ZN(n7493) );
  AOI22_X1 U6794 ( .A1(n5403), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5402), .B2(
        n7493), .ZN(n5290) );
  NAND2_X1 U6795 ( .A1(n5234), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6796 ( .A1(n5508), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5297) );
  INV_X1 U6797 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6798 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  AND2_X1 U6799 ( .A1(n5307), .A2(n5294), .ZN(n7875) );
  NAND2_X1 U6800 ( .A1(n5489), .A2(n7875), .ZN(n5296) );
  NAND2_X1 U6801 ( .A1(n5490), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5295) );
  NAND4_X1 U6802 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n9984)
         );
  INV_X1 U6803 ( .A(n9984), .ZN(n5299) );
  OR2_X1 U6804 ( .A1(n5606), .A2(n5299), .ZN(n9154) );
  NAND2_X1 U6805 ( .A1(n5606), .A2(n5299), .ZN(n9976) );
  INV_X1 U6806 ( .A(n9059), .ZN(n5300) );
  NAND2_X1 U6807 ( .A1(n7872), .A2(n5300), .ZN(n9977) );
  XNOR2_X1 U6808 ( .A(n5349), .B(n5301), .ZN(n7049) );
  NAND2_X1 U6809 ( .A1(n7049), .A2(n6648), .ZN(n5305) );
  NAND2_X1 U6810 ( .A1(n5288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5302) );
  MUX2_X1 U6811 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5302), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5303) );
  AND2_X1 U6812 ( .A1(n5303), .A2(n4454), .ZN(n9302) );
  AOI22_X1 U6813 ( .A1(n5403), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5402), .B2(
        n9302), .ZN(n5304) );
  NAND2_X1 U6814 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6815 ( .A1(n5325), .A2(n5308), .ZN(n9995) );
  INV_X1 U6816 ( .A(n9995), .ZN(n7864) );
  NAND2_X1 U6817 ( .A1(n5489), .A2(n7864), .ZN(n5312) );
  NAND2_X1 U6818 ( .A1(n5234), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6819 ( .A1(n5508), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6820 ( .A1(n5490), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5309) );
  NAND4_X1 U6821 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n9199)
         );
  INV_X1 U6822 ( .A(n9199), .ZN(n8056) );
  AND2_X1 U6823 ( .A1(n9969), .A2(n8056), .ZN(n8975) );
  INV_X1 U6824 ( .A(n8975), .ZN(n9157) );
  AND2_X1 U6825 ( .A1(n9976), .A2(n9157), .ZN(n5313) );
  NAND2_X1 U6826 ( .A1(n9977), .A2(n5313), .ZN(n5314) );
  OR2_X1 U6827 ( .A1(n9969), .A2(n8056), .ZN(n9159) );
  NAND2_X1 U6828 ( .A1(n5314), .A2(n9159), .ZN(n7790) );
  NAND2_X1 U6829 ( .A1(n5317), .A2(n5316), .ZN(n5319) );
  NAND2_X1 U6830 ( .A1(n7111), .A2(n6648), .ZN(n5323) );
  NAND2_X1 U6831 ( .A1(n4454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5320) );
  MUX2_X1 U6832 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5320), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5321) );
  NAND2_X1 U6833 ( .A1(n5321), .A2(n5354), .ZN(n9316) );
  INV_X1 U6834 ( .A(n9316), .ZN(n9304) );
  AOI22_X1 U6835 ( .A1(n5403), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5402), .B2(
        n9304), .ZN(n5322) );
  NAND2_X1 U6836 ( .A1(n5490), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6837 ( .A1(n5234), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6838 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  AND2_X1 U6839 ( .A1(n5341), .A2(n5326), .ZN(n8058) );
  NAND2_X1 U6840 ( .A1(n5489), .A2(n8058), .ZN(n5328) );
  NAND2_X1 U6841 ( .A1(n5508), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5327) );
  NAND4_X1 U6842 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n9983)
         );
  INV_X1 U6843 ( .A(n9983), .ZN(n8922) );
  INV_X1 U6844 ( .A(n5331), .ZN(n7788) );
  NAND2_X1 U6845 ( .A1(n7788), .A2(n8934), .ZN(n7941) );
  NAND2_X1 U6846 ( .A1(n7055), .A2(n6648), .ZN(n5339) );
  NAND2_X1 U6847 ( .A1(n5354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5337) );
  XNOR2_X1 U6848 ( .A(n5337), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9328) );
  AOI22_X1 U6849 ( .A1(n5403), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5402), .B2(
        n9328), .ZN(n5338) );
  INV_X1 U6850 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9708) );
  OR2_X1 U6851 ( .A1(n5340), .A2(n9708), .ZN(n5346) );
  NAND2_X1 U6852 ( .A1(n5234), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5345) );
  INV_X1 U6853 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U6854 ( .A1(n5341), .A2(n9733), .ZN(n5342) );
  AND2_X1 U6855 ( .A1(n5357), .A2(n5342), .ZN(n8925) );
  NAND2_X1 U6856 ( .A1(n5489), .A2(n8925), .ZN(n5344) );
  NAND2_X1 U6857 ( .A1(n5508), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5343) );
  NAND4_X1 U6858 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), .ZN(n9198)
         );
  INV_X1 U6859 ( .A(n9198), .ZN(n5347) );
  OR2_X1 U6860 ( .A1(n9623), .A2(n5347), .ZN(n9162) );
  NAND2_X1 U6861 ( .A1(n9623), .A2(n5347), .ZN(n8977) );
  NAND2_X1 U6862 ( .A1(n7941), .A2(n9062), .ZN(n7940) );
  NAND2_X1 U6863 ( .A1(n5349), .A2(n5348), .ZN(n5351) );
  NAND2_X1 U6864 ( .A1(n5351), .A2(n5350), .ZN(n5353) );
  NAND2_X1 U6865 ( .A1(n7053), .A2(n6648), .ZN(n5356) );
  XNOR2_X1 U6866 ( .A(n5368), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9350) );
  AOI22_X1 U6867 ( .A1(n5403), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5402), .B2(
        n9350), .ZN(n5355) );
  INV_X1 U6868 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9762) );
  OR2_X1 U6869 ( .A1(n5340), .A2(n9762), .ZN(n5362) );
  NAND2_X1 U6870 ( .A1(n5234), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5361) );
  INV_X1 U6871 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U6872 ( .A1(n5357), .A2(n9747), .ZN(n5358) );
  AND2_X1 U6873 ( .A1(n5372), .A2(n5358), .ZN(n8865) );
  NAND2_X1 U6874 ( .A1(n5489), .A2(n8865), .ZN(n5360) );
  NAND2_X1 U6875 ( .A1(n5508), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5359) );
  NAND4_X1 U6876 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n9197)
         );
  INV_X1 U6877 ( .A(n9197), .ZN(n8877) );
  NAND2_X1 U6878 ( .A1(n7908), .A2(n8877), .ZN(n9169) );
  INV_X1 U6879 ( .A(n9063), .ZN(n5364) );
  INV_X1 U6880 ( .A(n8977), .ZN(n5363) );
  NOR2_X1 U6881 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  NAND2_X1 U6882 ( .A1(n7153), .A2(n6648), .ZN(n5371) );
  INV_X1 U6883 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U6884 ( .A1(n5368), .A2(n5541), .ZN(n5369) );
  XNOR2_X1 U6885 ( .A(n5384), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9367) );
  AOI22_X1 U6886 ( .A1(n5403), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5402), .B2(
        n9367), .ZN(n5370) );
  INV_X1 U6887 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9744) );
  OR2_X1 U6888 ( .A1(n5340), .A2(n9744), .ZN(n5377) );
  NAND2_X1 U6889 ( .A1(n5234), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6890 ( .A1(n5372), .A2(n8873), .ZN(n5373) );
  AND2_X1 U6891 ( .A1(n5388), .A2(n5373), .ZN(n8874) );
  NAND2_X1 U6892 ( .A1(n5489), .A2(n8874), .ZN(n5375) );
  NAND2_X1 U6893 ( .A1(n5508), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5374) );
  NAND4_X1 U6894 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n9196)
         );
  INV_X1 U6895 ( .A(n9196), .ZN(n5378) );
  OR2_X1 U6896 ( .A1(n9619), .A2(n5378), .ZN(n8987) );
  NAND2_X1 U6897 ( .A1(n9619), .A2(n5378), .ZN(n8994) );
  NAND2_X1 U6898 ( .A1(n7978), .A2(n8994), .ZN(n8010) );
  NAND2_X1 U6899 ( .A1(n5395), .A2(n5379), .ZN(n5381) );
  NAND2_X1 U6900 ( .A1(n7116), .A2(n6648), .ZN(n5386) );
  XNOR2_X1 U6901 ( .A(n5398), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9389) );
  AOI22_X1 U6902 ( .A1(n5403), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5402), .B2(
        n9389), .ZN(n5385) );
  INV_X1 U6903 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6904 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  NAND2_X1 U6905 ( .A1(n5406), .A2(n5389), .ZN(n8906) );
  OR2_X1 U6906 ( .A1(n5530), .A2(n8906), .ZN(n5393) );
  INV_X1 U6907 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9934) );
  OR2_X1 U6908 ( .A1(n5340), .A2(n9934), .ZN(n5392) );
  NAND2_X1 U6909 ( .A1(n5234), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6910 ( .A1(n5508), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5390) );
  NAND4_X1 U6911 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n9195)
         );
  INV_X1 U6912 ( .A(n9195), .ZN(n9548) );
  OR2_X1 U6913 ( .A1(n8910), .A2(n9548), .ZN(n9170) );
  NAND2_X1 U6914 ( .A1(n8910), .A2(n9548), .ZN(n8995) );
  NAND2_X1 U6915 ( .A1(n9170), .A2(n8995), .ZN(n9066) );
  INV_X1 U6916 ( .A(n9066), .ZN(n8011) );
  NAND2_X1 U6917 ( .A1(n5395), .A2(n5394), .ZN(n5397) );
  NAND2_X1 U6918 ( .A1(n7183), .A2(n6648), .ZN(n5405) );
  AOI22_X1 U6919 ( .A1(n5403), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5402), .B2(
        n5401), .ZN(n5404) );
  NAND2_X1 U6920 ( .A1(n5406), .A2(n8842), .ZN(n5407) );
  NAND2_X1 U6921 ( .A1(n5420), .A2(n5407), .ZN(n9542) );
  AOI22_X1 U6922 ( .A1(n5490), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n5234), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n5409) );
  INV_X1 U6923 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9879) );
  OR2_X1 U6924 ( .A1(n5125), .A2(n9879), .ZN(n5408) );
  OAI211_X1 U6925 ( .C1(n9542), .C2(n5530), .A(n5409), .B(n5408), .ZN(n9523)
         );
  INV_X1 U6926 ( .A(n9523), .ZN(n8886) );
  OR2_X1 U6927 ( .A1(n9608), .A2(n8886), .ZN(n9171) );
  NAND2_X1 U6928 ( .A1(n9608), .A2(n8886), .ZN(n9175) );
  INV_X1 U6929 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6930 ( .A1(n7227), .A2(n6648), .ZN(n5418) );
  OR2_X1 U6931 ( .A1(n6649), .A2(n7206), .ZN(n5417) );
  INV_X1 U6932 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5424) );
  INV_X1 U6933 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6934 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  NAND2_X1 U6935 ( .A1(n5429), .A2(n5421), .ZN(n8884) );
  OR2_X1 U6936 ( .A1(n8884), .A2(n5530), .ZN(n5423) );
  AOI22_X1 U6937 ( .A1(n5490), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n5234), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n5422) );
  OAI211_X1 U6938 ( .C1(n5125), .C2(n5424), .A(n5423), .B(n5422), .ZN(n9511)
         );
  INV_X1 U6939 ( .A(n9511), .ZN(n9550) );
  OR2_X1 U6940 ( .A1(n9530), .A2(n9550), .ZN(n9001) );
  NAND2_X1 U6941 ( .A1(n9530), .A2(n9550), .ZN(n8932) );
  NAND2_X1 U6942 ( .A1(n9001), .A2(n8932), .ZN(n9517) );
  INV_X1 U6943 ( .A(n9517), .ZN(n9521) );
  NAND2_X1 U6944 ( .A1(n9520), .A2(n9521), .ZN(n9519) );
  NAND2_X1 U6945 ( .A1(n9519), .A2(n8932), .ZN(n9509) );
  XNOR2_X1 U6946 ( .A(n5426), .B(n5425), .ZN(n7275) );
  NAND2_X1 U6947 ( .A1(n7275), .A2(n6648), .ZN(n5428) );
  OR2_X1 U6948 ( .A1(n6649), .A2(n9902), .ZN(n5427) );
  NAND2_X1 U6949 ( .A1(n5429), .A2(n8852), .ZN(n5430) );
  NAND2_X1 U6950 ( .A1(n5448), .A2(n5430), .ZN(n9504) );
  AOI22_X1 U6951 ( .A1(n5174), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5508), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6952 ( .A1(n5490), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5431) );
  OAI211_X1 U6953 ( .C1(n9504), .C2(n5530), .A(n5432), .B(n5431), .ZN(n9524)
         );
  INV_X1 U6954 ( .A(n9524), .ZN(n8895) );
  OR2_X1 U6955 ( .A1(n9597), .A2(n8895), .ZN(n9002) );
  NAND2_X1 U6956 ( .A1(n9597), .A2(n8895), .ZN(n9003) );
  NAND2_X1 U6957 ( .A1(n9002), .A2(n9003), .ZN(n5640) );
  NAND2_X1 U6958 ( .A1(n9509), .A2(n9510), .ZN(n9508) );
  NAND2_X1 U6959 ( .A1(n9508), .A2(n9003), .ZN(n9487) );
  XNOR2_X1 U6960 ( .A(n5434), .B(n5433), .ZN(n7347) );
  NAND2_X1 U6961 ( .A1(n7347), .A2(n6648), .ZN(n5436) );
  OR2_X1 U6962 ( .A1(n6649), .A2(n8090), .ZN(n5435) );
  XNOR2_X1 U6963 ( .A(n5448), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U6964 ( .A1(n9495), .A2(n5489), .ZN(n5441) );
  INV_X1 U6965 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U6966 ( .A1(n5174), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6967 ( .A1(n5508), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5437) );
  OAI211_X1 U6968 ( .C1(n5340), .C2(n9925), .A(n5438), .B(n5437), .ZN(n5439)
         );
  INV_X1 U6969 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6970 ( .A1(n5441), .A2(n5440), .ZN(n9512) );
  INV_X1 U6971 ( .A(n9512), .ZN(n9008) );
  XNOR2_X1 U6972 ( .A(n9494), .B(n9008), .ZN(n9484) );
  NAND2_X1 U6973 ( .A1(n9487), .A2(n4750), .ZN(n9486) );
  NAND2_X1 U6974 ( .A1(n9494), .A2(n9008), .ZN(n9007) );
  NAND2_X1 U6975 ( .A1(n9486), .A2(n9007), .ZN(n9474) );
  NAND2_X1 U6976 ( .A1(n7394), .A2(n6648), .ZN(n5445) );
  OR2_X1 U6977 ( .A1(n6649), .A2(n9710), .ZN(n5444) );
  INV_X1 U6978 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5447) );
  INV_X1 U6979 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5446) );
  OAI21_X1 U6980 ( .B1(n5448), .B2(n5447), .A(n5446), .ZN(n5449) );
  NAND2_X1 U6981 ( .A1(n5459), .A2(n5449), .ZN(n8377) );
  OR2_X1 U6982 ( .A1(n8377), .A2(n5530), .ZN(n5454) );
  INV_X1 U6983 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9764) );
  NAND2_X1 U6984 ( .A1(n5490), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6985 ( .A1(n5508), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5450) );
  OAI211_X1 U6986 ( .C1(n5200), .C2(n9764), .A(n5451), .B(n5450), .ZN(n5452)
         );
  INV_X1 U6987 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U6988 ( .A1(n5454), .A2(n5453), .ZN(n9489) );
  INV_X1 U6989 ( .A(n9489), .ZN(n8384) );
  OR2_X1 U6990 ( .A1(n9588), .A2(n8384), .ZN(n9010) );
  NAND2_X1 U6991 ( .A1(n9588), .A2(n8384), .ZN(n9452) );
  NAND2_X1 U6992 ( .A1(n9010), .A2(n9452), .ZN(n9473) );
  INV_X1 U6993 ( .A(n9473), .ZN(n9471) );
  XNOR2_X1 U6994 ( .A(n5456), .B(n5455), .ZN(n7468) );
  NAND2_X1 U6995 ( .A1(n7468), .A2(n6648), .ZN(n5458) );
  OR2_X1 U6996 ( .A1(n6649), .A2(n7469), .ZN(n5457) );
  INV_X1 U6997 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U6998 ( .A1(n5459), .A2(n9862), .ZN(n5460) );
  NAND2_X1 U6999 ( .A1(n5472), .A2(n5460), .ZN(n9462) );
  OR2_X1 U7000 ( .A1(n9462), .A2(n5530), .ZN(n5465) );
  INV_X1 U7001 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U7002 ( .A1(n5508), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7003 ( .A1(n5174), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5461) );
  OAI211_X1 U7004 ( .C1(n5340), .C2(n9641), .A(n5462), .B(n5461), .ZN(n5463)
         );
  INV_X1 U7005 ( .A(n5463), .ZN(n5464) );
  NAND2_X1 U7006 ( .A1(n5465), .A2(n5464), .ZN(n9194) );
  INV_X1 U7007 ( .A(n9194), .ZN(n9442) );
  NAND2_X1 U7008 ( .A1(n9464), .A2(n9442), .ZN(n9088) );
  NAND2_X1 U7009 ( .A1(n9081), .A2(n9088), .ZN(n9454) );
  INV_X1 U7010 ( .A(n9452), .ZN(n5466) );
  NOR2_X1 U7011 ( .A1(n9454), .A2(n5466), .ZN(n5467) );
  NAND2_X1 U7012 ( .A1(n7515), .A2(n6648), .ZN(n5471) );
  OR2_X1 U7013 ( .A1(n6649), .A2(n9794), .ZN(n5470) );
  NAND2_X1 U7014 ( .A1(n5472), .A2(n9904), .ZN(n5473) );
  NAND2_X1 U7015 ( .A1(n5487), .A2(n5473), .ZN(n9445) );
  OR2_X1 U7016 ( .A1(n9445), .A2(n5530), .ZN(n5479) );
  INV_X1 U7017 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7018 ( .A1(n5508), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7019 ( .A1(n5174), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5474) );
  OAI211_X1 U7020 ( .C1(n5340), .C2(n5476), .A(n5475), .B(n5474), .ZN(n5477)
         );
  INV_X1 U7021 ( .A(n5477), .ZN(n5478) );
  NAND2_X1 U7022 ( .A1(n5479), .A2(n5478), .ZN(n9458) );
  INV_X1 U7023 ( .A(n9458), .ZN(n5498) );
  OR2_X1 U7024 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U7025 ( .A1(n5483), .A2(n5482), .ZN(n7723) );
  NAND2_X1 U7026 ( .A1(n7723), .A2(n6648), .ZN(n5485) );
  OR2_X1 U7027 ( .A1(n6649), .A2(n7726), .ZN(n5484) );
  NAND2_X1 U7028 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  NAND2_X1 U7029 ( .A1(n9431), .A2(n5489), .ZN(n5496) );
  INV_X1 U7030 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7031 ( .A1(n5490), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7032 ( .A1(n5174), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5491) );
  OAI211_X1 U7033 ( .C1(n5493), .C2(n5125), .A(n5492), .B(n5491), .ZN(n5494)
         );
  INV_X1 U7034 ( .A(n5494), .ZN(n5495) );
  INV_X1 U7035 ( .A(n8403), .ZN(n9443) );
  NAND2_X1 U7036 ( .A1(n9575), .A2(n5498), .ZN(n9045) );
  NAND2_X1 U7037 ( .A1(n7727), .A2(n6648), .ZN(n5503) );
  OR2_X1 U7038 ( .A1(n6649), .A2(n7775), .ZN(n5502) );
  INV_X1 U7039 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7040 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  NAND2_X1 U7041 ( .A1(n5507), .A2(n5506), .ZN(n8395) );
  INV_X1 U7042 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U7043 ( .A1(n5174), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7044 ( .A1(n5508), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U7045 ( .C1(n5340), .C2(n9874), .A(n5510), .B(n5509), .ZN(n5511)
         );
  INV_X1 U7046 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U7047 ( .A1(n9564), .A2(n9029), .ZN(n9092) );
  AND2_X1 U7048 ( .A1(n9094), .A2(n9092), .ZN(n5514) );
  INV_X1 U7049 ( .A(n9092), .ZN(n9015) );
  NAND2_X1 U7050 ( .A1(n5516), .A2(n5515), .ZN(n6623) );
  INV_X1 U7051 ( .A(n9100), .ZN(n9017) );
  AOI21_X1 U7052 ( .B1(n6623), .B2(n9091), .A(n9017), .ZN(n5538) );
  AND2_X1 U7053 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  NAND2_X1 U7054 ( .A1(n5521), .A2(n5520), .ZN(n5523) );
  MUX2_X1 U7055 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4402), .Z(n6643) );
  INV_X1 U7056 ( .A(n5524), .ZN(n5526) );
  INV_X1 U7057 ( .A(SI_29_), .ZN(n5525) );
  NAND2_X1 U7058 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  INV_X1 U7059 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7867) );
  OR2_X1 U7060 ( .A1(n6649), .A2(n7867), .ZN(n5528) );
  OR2_X1 U7061 ( .A1(n5661), .A2(n5530), .ZN(n5536) );
  INV_X1 U7062 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7063 ( .A1(n5508), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7064 ( .A1(n5174), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5531) );
  OAI211_X1 U7065 ( .C1(n5340), .C2(n5533), .A(n5532), .B(n5531), .ZN(n5534)
         );
  INV_X1 U7066 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7067 ( .A1(n5536), .A2(n5535), .ZN(n9192) );
  INV_X1 U7068 ( .A(n9192), .ZN(n5537) );
  NAND2_X1 U7069 ( .A1(n9558), .A2(n5537), .ZN(n9110) );
  MUX2_X1 U7070 ( .A(n9091), .B(n5538), .S(n9073), .Z(n5553) );
  INV_X1 U7071 ( .A(n6623), .ZN(n5539) );
  INV_X1 U7072 ( .A(n9073), .ZN(n9034) );
  NAND3_X1 U7073 ( .A1(n5539), .A2(n9034), .A3(n9100), .ZN(n5552) );
  NAND4_X1 U7074 ( .A1(n5542), .A2(n5541), .A3(n5540), .A4(n5399), .ZN(n5543)
         );
  NAND2_X1 U7075 ( .A1(n5547), .A2(n5549), .ZN(n5545) );
  OAI21_X2 U7076 ( .B1(n5545), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7077 ( .A1(n5653), .A2(n5401), .ZN(n5551) );
  XNOR2_X2 U7078 ( .A(n5546), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5655) );
  INV_X1 U7079 ( .A(n5547), .ZN(n5548) );
  INV_X1 U7080 ( .A(n6415), .ZN(n5601) );
  NAND2_X1 U7081 ( .A1(n5655), .A2(n5601), .ZN(n8930) );
  NAND2_X1 U7082 ( .A1(n5653), .A2(n5655), .ZN(n9115) );
  INV_X1 U7083 ( .A(n9115), .ZN(n5598) );
  INV_X1 U7084 ( .A(n5554), .ZN(n6899) );
  NAND2_X1 U7085 ( .A1(n5174), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5557) );
  INV_X1 U7086 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9630) );
  OR2_X1 U7087 ( .A1(n5340), .A2(n9630), .ZN(n5556) );
  INV_X1 U7088 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9694) );
  OR2_X1 U7089 ( .A1(n5125), .A2(n9694), .ZN(n5555) );
  AND3_X1 U7090 ( .A1(n5557), .A2(n5556), .A3(n5555), .ZN(n9075) );
  INV_X1 U7091 ( .A(n5558), .ZN(n6846) );
  NAND2_X1 U7092 ( .A1(n6846), .A2(P1_B_REG_SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7093 ( .A1(n9982), .A2(n5559), .ZN(n6664) );
  NOR2_X1 U7094 ( .A1(n9075), .A2(n6664), .ZN(n5560) );
  INV_X1 U7095 ( .A(n5561), .ZN(n5562) );
  NOR2_X2 U7096 ( .A1(n5563), .A2(n5562), .ZN(n9561) );
  NAND2_X1 U7097 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U7098 ( .A1(n5566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7099 ( .A(n5567), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7395) );
  INV_X1 U7100 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7101 ( .A1(n5574), .A2(n5576), .ZN(n5568) );
  INV_X1 U7102 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7103 ( .A1(n5571), .A2(n5570), .ZN(n5573) );
  OR2_X1 U7104 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  NAND2_X1 U7105 ( .A1(n5573), .A2(n5572), .ZN(n7516) );
  INV_X1 U7106 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U7107 ( .A1(n5575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5577) );
  XNOR2_X1 U7108 ( .A(n5577), .B(n5576), .ZN(n7470) );
  NOR2_X1 U7109 ( .A1(n7516), .A2(n7470), .ZN(n5578) );
  NAND2_X1 U7110 ( .A1(n6792), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7111 ( .A1(n7516), .A2(P1_B_REG_SCAN_IN), .ZN(n5581) );
  INV_X1 U7112 ( .A(n7470), .ZN(n5580) );
  MUX2_X1 U7113 ( .A(n5581), .B(P1_B_REG_SCAN_IN), .S(n5580), .Z(n5582) );
  NAND2_X1 U7114 ( .A1(n5582), .A2(n5595), .ZN(n6401) );
  INV_X1 U7115 ( .A(n6401), .ZN(n5594) );
  NOR2_X2 U7116 ( .A1(n9940), .A2(n5594), .ZN(n10044) );
  NOR4_X1 U7117 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5583) );
  INV_X1 U7118 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10036) );
  INV_X1 U7119 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10035) );
  NAND3_X1 U7120 ( .A1(n5583), .A2(n10036), .A3(n10035), .ZN(n5589) );
  NOR4_X1 U7121 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5587) );
  NOR4_X1 U7122 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5586) );
  NOR4_X1 U7123 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5585) );
  NOR4_X1 U7124 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5584) );
  NAND4_X1 U7125 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n5588)
         );
  NOR4_X1 U7126 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n5589), .A4(n5588), .ZN(n5591) );
  INV_X1 U7127 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10039) );
  INV_X1 U7128 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10045) );
  INV_X1 U7129 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10042) );
  INV_X1 U7130 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10053) );
  NAND4_X1 U7131 ( .A1(n10039), .A2(n10045), .A3(n10042), .A4(n10053), .ZN(
        n5590) );
  NOR3_X1 U7132 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        n5590), .ZN(n9660) );
  AND2_X1 U7133 ( .A1(n5591), .A2(n9660), .ZN(n6400) );
  INV_X1 U7134 ( .A(n6400), .ZN(n5592) );
  NOR2_X1 U7135 ( .A1(n9940), .A2(n5592), .ZN(n5600) );
  INV_X1 U7136 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7137 ( .A1(n5594), .A2(n5593), .ZN(n5597) );
  INV_X1 U7138 ( .A(n5595), .ZN(n7724) );
  NAND2_X1 U7139 ( .A1(n7724), .A2(n7470), .ZN(n5596) );
  NAND2_X1 U7140 ( .A1(n7724), .A2(n7516), .ZN(n9939) );
  OAI21_X1 U7141 ( .B1(n6401), .B2(P1_D_REG_1__SCAN_IN), .A(n9939), .ZN(n6632)
         );
  NOR2_X1 U7142 ( .A1(n9941), .A2(n6632), .ZN(n5599) );
  AND2_X1 U7143 ( .A1(n6190), .A2(n5598), .ZN(n6418) );
  INV_X1 U7144 ( .A(n6418), .ZN(n6634) );
  OAI211_X1 U7145 ( .C1(n10060), .C2(n5600), .A(n5599), .B(n6634), .ZN(n5603)
         );
  NOR2_X1 U7146 ( .A1(n9940), .A2(n5655), .ZN(n5602) );
  NAND2_X1 U7147 ( .A1(n5602), .A2(n10084), .ZN(n9994) );
  NAND2_X1 U7148 ( .A1(n10008), .A2(n9200), .ZN(n7870) );
  NAND2_X1 U7149 ( .A1(n9059), .A2(n7870), .ZN(n5619) );
  OR2_X1 U7150 ( .A1(n7759), .A2(n9201), .ZN(n9996) );
  OR2_X1 U7151 ( .A1(n10008), .A2(n9200), .ZN(n5605) );
  AND2_X1 U7152 ( .A1(n9996), .A2(n5605), .ZN(n7869) );
  AND2_X1 U7153 ( .A1(n9051), .A2(n9052), .ZN(n5612) );
  INV_X1 U7154 ( .A(n7135), .ZN(n8073) );
  NAND2_X1 U7155 ( .A1(n8073), .A2(n7511), .ZN(n8070) );
  NAND2_X1 U7156 ( .A1(n7148), .A2(n10062), .ZN(n5608) );
  NAND2_X1 U7157 ( .A1(n8071), .A2(n5608), .ZN(n7170) );
  NAND2_X1 U7158 ( .A1(n7170), .A2(n9047), .ZN(n7172) );
  NAND2_X1 U7159 ( .A1(n7044), .A2(n7186), .ZN(n5609) );
  NAND2_X1 U7160 ( .A1(n7172), .A2(n5609), .ZN(n7676) );
  NAND2_X1 U7161 ( .A1(n7676), .A2(n8936), .ZN(n7675) );
  NAND2_X1 U7162 ( .A1(n7063), .A2(n10067), .ZN(n5610) );
  NAND2_X1 U7163 ( .A1(n7235), .A2(n7609), .ZN(n7230) );
  INV_X1 U7164 ( .A(n7230), .ZN(n5611) );
  NAND2_X1 U7165 ( .A1(n7293), .A2(n7264), .ZN(n7431) );
  NAND2_X1 U7166 ( .A1(n7385), .A2(n10023), .ZN(n5613) );
  AND2_X1 U7167 ( .A1(n7431), .A2(n5613), .ZN(n5615) );
  INV_X1 U7168 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7169 ( .A1(n8949), .A2(n8947), .ZN(n7437) );
  AOI21_X1 U7170 ( .B1(n7432), .B2(n5615), .A(n4921), .ZN(n7629) );
  NAND2_X1 U7171 ( .A1(n7567), .A2(n8955), .ZN(n7628) );
  NAND2_X1 U7172 ( .A1(n7629), .A2(n7628), .ZN(n7631) );
  NAND2_X1 U7173 ( .A1(n7589), .A2(n10073), .ZN(n5616) );
  NAND2_X1 U7174 ( .A1(n7631), .A2(n5616), .ZN(n7582) );
  NAND2_X1 U7175 ( .A1(n8951), .A2(n8957), .ZN(n7587) );
  NAND2_X1 U7176 ( .A1(n7582), .A2(n7587), .ZN(n7581) );
  OR2_X1 U7177 ( .A1(n9203), .A2(n7585), .ZN(n5617) );
  NAND2_X1 U7178 ( .A1(n7581), .A2(n5617), .ZN(n7561) );
  NAND2_X1 U7179 ( .A1(n8968), .A2(n8962), .ZN(n7570) );
  NAND2_X1 U7180 ( .A1(n7561), .A2(n7570), .ZN(n7560) );
  OR2_X1 U7181 ( .A1(n7577), .A2(n9202), .ZN(n5618) );
  NAND2_X1 U7182 ( .A1(n7560), .A2(n5618), .ZN(n7457) );
  NOR2_X1 U7183 ( .A1(n9054), .A2(n5619), .ZN(n5620) );
  NAND2_X1 U7184 ( .A1(n7457), .A2(n5620), .ZN(n5621) );
  INV_X1 U7185 ( .A(n9974), .ZN(n5624) );
  NOR2_X1 U7186 ( .A1(n9969), .A2(n9199), .ZN(n7929) );
  NAND2_X1 U7187 ( .A1(n5624), .A2(n5623), .ZN(n7786) );
  NAND2_X1 U7188 ( .A1(n9969), .A2(n9199), .ZN(n7785) );
  NAND2_X1 U7189 ( .A1(n7794), .A2(n9983), .ZN(n5627) );
  AND2_X1 U7190 ( .A1(n7785), .A2(n5627), .ZN(n7931) );
  INV_X1 U7191 ( .A(n9062), .ZN(n5625) );
  AND2_X1 U7192 ( .A1(n7931), .A2(n5625), .ZN(n5626) );
  NAND2_X1 U7193 ( .A1(n7786), .A2(n5626), .ZN(n5630) );
  INV_X1 U7194 ( .A(n5627), .ZN(n5628) );
  OR2_X1 U7195 ( .A1(n5628), .A2(n9060), .ZN(n7928) );
  OR2_X1 U7196 ( .A1(n9623), .A2(n9198), .ZN(n5629) );
  NAND2_X1 U7197 ( .A1(n7908), .A2(n9197), .ZN(n5631) );
  NAND2_X1 U7198 ( .A1(n7898), .A2(n5631), .ZN(n7977) );
  OR2_X1 U7199 ( .A1(n9619), .A2(n9196), .ZN(n5633) );
  OR2_X1 U7200 ( .A1(n8910), .A2(n9195), .ZN(n5634) );
  NAND2_X1 U7201 ( .A1(n9608), .A2(n9523), .ZN(n5635) );
  NAND2_X1 U7202 ( .A1(n9537), .A2(n5635), .ZN(n5637) );
  OR2_X1 U7203 ( .A1(n9608), .A2(n9523), .ZN(n5636) );
  NAND2_X1 U7204 ( .A1(n5637), .A2(n5636), .ZN(n9518) );
  NAND2_X1 U7205 ( .A1(n9518), .A2(n9517), .ZN(n5639) );
  OR2_X1 U7206 ( .A1(n9530), .A2(n9511), .ZN(n5638) );
  NAND2_X1 U7207 ( .A1(n5639), .A2(n5638), .ZN(n9501) );
  NAND2_X1 U7208 ( .A1(n9501), .A2(n5640), .ZN(n5642) );
  OR2_X1 U7209 ( .A1(n9597), .A2(n9524), .ZN(n5641) );
  OR2_X1 U7210 ( .A1(n9494), .A2(n9512), .ZN(n5643) );
  OR2_X1 U7211 ( .A1(n9588), .A2(n9489), .ZN(n5644) );
  NOR2_X1 U7212 ( .A1(n9464), .A2(n9194), .ZN(n5647) );
  NAND2_X1 U7213 ( .A1(n9464), .A2(n9194), .ZN(n5646) );
  NOR2_X1 U7214 ( .A1(n9430), .A2(n8403), .ZN(n5650) );
  NAND2_X1 U7215 ( .A1(n9430), .A2(n8403), .ZN(n5649) );
  OR2_X1 U7216 ( .A1(n9564), .A2(n9427), .ZN(n5651) );
  NAND2_X1 U7217 ( .A1(n9026), .A2(n9193), .ZN(n5652) );
  OR2_X1 U7218 ( .A1(n6191), .A2(n6192), .ZN(n6416) );
  INV_X1 U7219 ( .A(n5655), .ZN(n9132) );
  AND2_X1 U7220 ( .A1(n8088), .A2(n9132), .ZN(n6939) );
  INV_X1 U7221 ( .A(n6939), .ZN(n5660) );
  NAND2_X1 U7222 ( .A1(n6416), .A2(n5660), .ZN(n7509) );
  AND2_X1 U7223 ( .A1(n6190), .A2(n6191), .ZN(n5656) );
  OR2_X1 U7224 ( .A1(n7509), .A2(n5656), .ZN(n7175) );
  INV_X1 U7225 ( .A(n6192), .ZN(n6189) );
  NAND2_X1 U7226 ( .A1(n5401), .A2(n6189), .ZN(n7635) );
  AND2_X1 U7227 ( .A1(n7175), .A2(n7635), .ZN(n9975) );
  NAND2_X1 U7228 ( .A1(n5123), .A2(n8082), .ZN(n8081) );
  INV_X1 U7229 ( .A(n7585), .ZN(n7600) );
  NAND2_X1 U7230 ( .A1(n7583), .A2(n7600), .ZN(n7562) );
  INV_X1 U7231 ( .A(n9623), .ZN(n8929) );
  INV_X1 U7232 ( .A(n9608), .ZN(n9541) );
  NAND2_X1 U7233 ( .A1(n9579), .A2(n9477), .ZN(n9461) );
  INV_X1 U7234 ( .A(n5659), .ZN(n9444) );
  AOI21_X1 U7235 ( .B1(n9558), .B2(n6627), .A(n9401), .ZN(n9559) );
  AND2_X1 U7236 ( .A1(n6939), .A2(n6415), .ZN(n10010) );
  NOR2_X1 U7237 ( .A1(n9467), .A2(n9968), .ZN(n7512) );
  INV_X1 U7238 ( .A(n9558), .ZN(n5664) );
  OR2_X1 U7239 ( .A1(n5660), .A2(n6415), .ZN(n9988) );
  INV_X1 U7240 ( .A(n5661), .ZN(n5662) );
  INV_X1 U7241 ( .A(n9994), .ZN(n10017) );
  AOI22_X1 U7242 ( .A1(n5662), .A2(n10017), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10019), .ZN(n5663) );
  OAI21_X1 U7243 ( .B1(n5664), .B2(n10022), .A(n5663), .ZN(n5665) );
  INV_X1 U7244 ( .A(n5667), .ZN(n5668) );
  INV_X1 U7245 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6118) );
  NOR2_X2 U7246 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5784) );
  INV_X1 U7247 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5836) );
  INV_X1 U7248 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5898) );
  INV_X1 U7249 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5710) );
  NOR2_X1 U7250 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5669) );
  OR2_X2 U7251 ( .A1(n5965), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5973) );
  NOR2_X2 U7252 ( .A1(n5973), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5982) );
  INV_X1 U7253 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5981) );
  OR2_X2 U7254 ( .A1(n5992), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5994) );
  OR2_X2 U7255 ( .A1(n5994), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7256 ( .A1(n5994), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7257 ( .A1(n6002), .A2(n5670), .ZN(n8646) );
  NOR2_X1 U7258 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5672) );
  AND2_X1 U7259 ( .A1(n5672), .A2(n5671), .ZN(n5680) );
  INV_X1 U7260 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5675) );
  INV_X1 U7261 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5674) );
  INV_X1 U7262 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5673) );
  NOR2_X1 U7263 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5677) );
  NOR2_X1 U7264 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5676) );
  AND2_X1 U7265 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  INV_X1 U7266 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5681) );
  INV_X1 U7267 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5717) );
  INV_X1 U7268 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5707) );
  INV_X1 U7269 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5687) );
  INV_X1 U7270 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6081) );
  AND2_X1 U7271 ( .A1(n5687), .A2(n6081), .ZN(n6087) );
  INV_X1 U7272 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5688) );
  INV_X1 U7273 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5704) );
  INV_X1 U7274 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5689) );
  AND2_X1 U7275 ( .A1(n5693), .A2(n5689), .ZN(n5690) );
  NAND2_X1 U7276 ( .A1(n6088), .A2(n5690), .ZN(n7989) );
  INV_X1 U7277 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7278 ( .A1(n6088), .A2(n5693), .ZN(n5694) );
  NAND2_X1 U7279 ( .A1(n8646), .A2(n5824), .ZN(n5701) );
  AOI22_X1 U7280 ( .A1(n5744), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n6051), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5700) );
  NAND2_X2 U7281 ( .A1(n5698), .A2(n5697), .ZN(n5914) );
  NAND2_X1 U7282 ( .A1(n6174), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7283 ( .A1(n6088), .A2(n5702), .ZN(n5703) );
  NAND2_X4 U7284 ( .A1(n6073), .A2(n6074), .ZN(n6497) );
  NAND2_X1 U7285 ( .A1(n6497), .A2(n6763), .ZN(n5723) );
  NAND2_X1 U7286 ( .A1(n7394), .A2(n8142), .ZN(n5709) );
  OR2_X1 U7287 ( .A1(n5753), .A2(n7392), .ZN(n5708) );
  NAND2_X1 U7288 ( .A1(n6174), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5715) );
  INV_X1 U7289 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9771) );
  OR2_X1 U7290 ( .A1(n5745), .A2(n9771), .ZN(n5714) );
  NOR2_X1 U7291 ( .A1(n5929), .A2(n5710), .ZN(n5711) );
  OR2_X1 U7292 ( .A1(n5949), .A2(n5711), .ZN(n8044) );
  INV_X1 U7293 ( .A(n8044), .ZN(n7973) );
  OR2_X1 U7294 ( .A1(n5746), .A2(n7973), .ZN(n5713) );
  INV_X1 U7295 ( .A(n5744), .ZN(n6022) );
  INV_X1 U7296 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8040) );
  OR2_X1 U7297 ( .A1(n6022), .A2(n8040), .ZN(n5712) );
  INV_X1 U7298 ( .A(n8720), .ZN(n8510) );
  NAND2_X1 U7299 ( .A1(n7053), .A2(n8142), .ZN(n5722) );
  OR2_X1 U7300 ( .A1(n5716), .A2(n7988), .ZN(n5718) );
  MUX2_X1 U7301 ( .A(n5718), .B(P2_IR_REG_31__SCAN_IN), .S(n5717), .Z(n5720)
         );
  NAND2_X1 U7302 ( .A1(n5720), .A2(n5941), .ZN(n7102) );
  INV_X1 U7303 ( .A(n7102), .ZN(n8566) );
  AOI22_X1 U7304 ( .A1(n5962), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5961), .B2(
        n8566), .ZN(n5721) );
  OR2_X1 U7305 ( .A1(n4399), .A2(n6758), .ZN(n5728) );
  OR2_X1 U7306 ( .A1(n5723), .A2(n6764), .ZN(n5727) );
  NAND3_X1 U7307 ( .A1(n5728), .A2(n5727), .A3(n4905), .ZN(n6950) );
  INV_X1 U7308 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6819) );
  OR2_X1 U7309 ( .A1(n5914), .A2(n6819), .ZN(n5733) );
  INV_X1 U7310 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5729) );
  OR2_X1 U7311 ( .A1(n5745), .A2(n5729), .ZN(n5732) );
  NAND2_X1 U7312 ( .A1(n5744), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5731) );
  INV_X1 U7313 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7139) );
  OR2_X1 U7314 ( .A1(n5746), .A2(n7139), .ZN(n5730) );
  NAND2_X1 U7315 ( .A1(n8198), .A2(n8197), .ZN(n6943) );
  NAND2_X1 U7316 ( .A1(n5744), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5737) );
  INV_X1 U7317 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6896) );
  OR2_X1 U7318 ( .A1(n5914), .A2(n6896), .ZN(n5735) );
  NAND2_X1 U7319 ( .A1(n5824), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5734) );
  INV_X1 U7320 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7321 ( .A1(n6763), .A2(SI_0_), .ZN(n5739) );
  INV_X1 U7322 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7323 ( .A1(n5739), .A2(n5738), .ZN(n5741) );
  AND2_X1 U7324 ( .A1(n5741), .A2(n5740), .ZN(n8834) );
  NAND2_X1 U7325 ( .A1(n6943), .A2(n6946), .ZN(n5743) );
  NAND2_X1 U7326 ( .A1(n6982), .A2(n6684), .ZN(n5742) );
  NAND2_X1 U7327 ( .A1(n5743), .A2(n5742), .ZN(n10241) );
  NAND2_X1 U7328 ( .A1(n5744), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5750) );
  OR2_X1 U7329 ( .A1(n5745), .A2(n6500), .ZN(n5749) );
  INV_X1 U7330 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8537) );
  OR2_X1 U7331 ( .A1(n5746), .A2(n8537), .ZN(n5748) );
  OR2_X1 U7332 ( .A1(n5914), .A2(n10259), .ZN(n5747) );
  INV_X1 U7333 ( .A(n6949), .ZN(n8523) );
  XNOR2_X2 U7334 ( .A(n5752), .B(n5751), .ZN(n6760) );
  OR2_X1 U7335 ( .A1(n5723), .A2(n6771), .ZN(n5755) );
  OR2_X1 U7336 ( .A1(n5753), .A2(n6759), .ZN(n5754) );
  OAI211_X1 U7337 ( .C1(n6497), .C2(n6760), .A(n5755), .B(n5754), .ZN(n5756)
         );
  INV_X1 U7338 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7339 ( .A1(n6949), .A2(n5756), .ZN(n8202) );
  NAND2_X1 U7340 ( .A1(n10241), .A2(n6120), .ZN(n5759) );
  NAND2_X1 U7341 ( .A1(n6949), .A2(n5757), .ZN(n5758) );
  NAND2_X1 U7342 ( .A1(n5759), .A2(n5758), .ZN(n7019) );
  NAND2_X1 U7343 ( .A1(n6174), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7344 ( .A1(n6051), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5763) );
  OR2_X1 U7345 ( .A1(n5746), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7346 ( .A1(n5744), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5760) );
  AND2_X1 U7347 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  NAND2_X1 U7348 ( .A1(n5765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5767) );
  INV_X1 U7349 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5766) );
  XNOR2_X1 U7350 ( .A(n5767), .B(n5766), .ZN(n6762) );
  OR2_X1 U7351 ( .A1(n5723), .A2(n6765), .ZN(n5769) );
  INV_X1 U7352 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U7353 ( .A1(n10246), .A2(n10265), .ZN(n5771) );
  NAND2_X1 U7354 ( .A1(n10246), .A2(n10265), .ZN(n5770) );
  OAI21_X1 U7355 ( .B1(n7019), .B2(n5771), .A(n5770), .ZN(n7012) );
  NAND2_X1 U7356 ( .A1(n6051), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5776) );
  INV_X1 U7357 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9677) );
  OR2_X1 U7358 ( .A1(n6022), .A2(n9677), .ZN(n5775) );
  AND2_X1 U7359 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5772) );
  NOR2_X1 U7360 ( .A1(n5784), .A2(n5772), .ZN(n7033) );
  OR2_X1 U7361 ( .A1(n5746), .A2(n7033), .ZN(n5774) );
  INV_X1 U7362 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7014) );
  OR2_X1 U7363 ( .A1(n5914), .A2(n7014), .ZN(n5773) );
  OR2_X1 U7364 ( .A1(n5723), .A2(n6769), .ZN(n5781) );
  OR2_X1 U7365 ( .A1(n5753), .A2(n6768), .ZN(n5780) );
  OR2_X1 U7366 ( .A1(n5777), .A2(n7988), .ZN(n5778) );
  XNOR2_X1 U7367 ( .A(n5778), .B(n9796), .ZN(n6889) );
  OR2_X1 U7368 ( .A1(n6497), .A2(n6889), .ZN(n5779) );
  AND3_X1 U7369 ( .A1(n5781), .A2(n5780), .A3(n5779), .ZN(n10271) );
  NAND2_X1 U7370 ( .A1(n7160), .A2(n10271), .ZN(n6123) );
  NAND2_X1 U7371 ( .A1(n7012), .A2(n6123), .ZN(n5782) );
  INV_X1 U7372 ( .A(n7160), .ZN(n8522) );
  INV_X1 U7373 ( .A(n10271), .ZN(n7030) );
  NAND2_X1 U7374 ( .A1(n8522), .A2(n7030), .ZN(n6122) );
  NAND2_X1 U7375 ( .A1(n5782), .A2(n6122), .ZN(n7105) );
  NAND2_X1 U7376 ( .A1(n5744), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5789) );
  OR2_X1 U7377 ( .A1(n5745), .A2(n10323), .ZN(n5788) );
  OR2_X1 U7378 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  AND2_X1 U7379 ( .A1(n5797), .A2(n5785), .ZN(n7108) );
  OR2_X1 U7380 ( .A1(n5746), .A2(n7108), .ZN(n5787) );
  INV_X1 U7381 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7107) );
  OR2_X1 U7382 ( .A1(n5914), .A2(n7107), .ZN(n5786) );
  OR2_X1 U7383 ( .A1(n5723), .A2(n6772), .ZN(n5794) );
  OR2_X1 U7384 ( .A1(n5753), .A2(n9803), .ZN(n5793) );
  NAND2_X1 U7385 ( .A1(n5790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U7386 ( .A(n5791), .B(n5681), .ZN(n6770) );
  OR2_X1 U7387 ( .A1(n6497), .A2(n6770), .ZN(n5792) );
  NAND2_X1 U7388 ( .A1(n7199), .A2(n10277), .ZN(n5795) );
  INV_X1 U7389 ( .A(n7199), .ZN(n8521) );
  INV_X1 U7390 ( .A(n10277), .ZN(n7157) );
  NAND2_X1 U7391 ( .A1(n8521), .A2(n7157), .ZN(n5796) );
  NAND2_X1 U7392 ( .A1(n5797), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5798) );
  AND2_X1 U7393 ( .A1(n5810), .A2(n5798), .ZN(n7196) );
  OR2_X1 U7394 ( .A1(n5746), .A2(n7196), .ZN(n5802) );
  INV_X1 U7395 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6541) );
  OR2_X1 U7396 ( .A1(n5914), .A2(n6541), .ZN(n5801) );
  NAND2_X1 U7397 ( .A1(n5744), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7398 ( .A1(n6051), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5799) );
  NAND4_X1 U7399 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n8520)
         );
  NAND2_X1 U7400 ( .A1(n5804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  MUX2_X1 U7401 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5803), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5805) );
  NAND2_X1 U7402 ( .A1(n5805), .A2(n5817), .ZN(n7081) );
  OR2_X1 U7403 ( .A1(n5723), .A2(n6777), .ZN(n5807) );
  OR2_X1 U7404 ( .A1(n5753), .A2(n6776), .ZN(n5806) );
  OAI211_X1 U7405 ( .C1(n6497), .C2(n7081), .A(n5807), .B(n5806), .ZN(n7123)
         );
  AND2_X1 U7406 ( .A1(n8520), .A2(n7123), .ZN(n5809) );
  INV_X1 U7407 ( .A(n8520), .ZN(n6707) );
  INV_X1 U7408 ( .A(n7123), .ZN(n10281) );
  NAND2_X1 U7409 ( .A1(n6707), .A2(n10281), .ZN(n5808) );
  NAND2_X1 U7410 ( .A1(n6051), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5815) );
  AND2_X1 U7411 ( .A1(n5810), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5811) );
  NOR2_X1 U7412 ( .A1(n5822), .A2(n5811), .ZN(n7221) );
  OR2_X1 U7413 ( .A1(n5746), .A2(n7221), .ZN(n5814) );
  NAND2_X1 U7414 ( .A1(n5744), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7415 ( .A1(n6174), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5812) );
  NAND4_X1 U7416 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n8519)
         );
  NAND2_X1 U7417 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  MUX2_X1 U7418 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5816), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5818) );
  NAND2_X1 U7419 ( .A1(n5818), .A2(n5843), .ZN(n7283) );
  OR2_X1 U7420 ( .A1(n5723), .A2(n6782), .ZN(n5820) );
  OR2_X1 U7421 ( .A1(n5753), .A2(n6781), .ZN(n5819) );
  OAI211_X1 U7422 ( .C1(n6497), .C2(n7283), .A(n5820), .B(n5819), .ZN(n7308)
         );
  XNOR2_X1 U7423 ( .A(n8519), .B(n7308), .ZN(n8230) );
  NAND2_X1 U7424 ( .A1(n7215), .A2(n8159), .ZN(n7214) );
  NAND2_X1 U7425 ( .A1(n8519), .A2(n7308), .ZN(n5821) );
  NAND2_X1 U7426 ( .A1(n6051), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U7427 ( .A1(n5744), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5827) );
  NOR2_X1 U7428 ( .A1(n5822), .A2(n9838), .ZN(n5823) );
  OR2_X1 U7429 ( .A1(n5837), .A2(n5823), .ZN(n7376) );
  NAND2_X1 U7430 ( .A1(n5824), .A2(n7376), .ZN(n5826) );
  NAND2_X1 U7431 ( .A1(n6174), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5825) );
  NAND4_X1 U7432 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n8518)
         );
  NAND2_X1 U7433 ( .A1(n6796), .A2(n8142), .ZN(n5833) );
  NAND2_X1 U7434 ( .A1(n5843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  INV_X1 U7435 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U7436 ( .A(n5830), .B(n5829), .ZN(n6800) );
  OR2_X1 U7437 ( .A1(n6497), .A2(n6800), .ZN(n5832) );
  OR2_X1 U7438 ( .A1(n5753), .A2(n6798), .ZN(n5831) );
  OR2_X1 U7439 ( .A1(n8518), .A2(n10286), .ZN(n8238) );
  NAND2_X1 U7440 ( .A1(n8518), .A2(n10286), .ZN(n8227) );
  NAND2_X1 U7441 ( .A1(n8238), .A2(n8227), .ZN(n8157) );
  INV_X1 U7442 ( .A(n10286), .ZN(n5834) );
  NAND2_X1 U7443 ( .A1(n8518), .A2(n5834), .ZN(n5835) );
  NAND2_X1 U7444 ( .A1(n5744), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5842) );
  INV_X1 U7445 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6592) );
  OR2_X1 U7446 ( .A1(n5745), .A2(n6592), .ZN(n5841) );
  OR2_X1 U7447 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  AND2_X1 U7448 ( .A1(n5856), .A2(n5838), .ZN(n7425) );
  OR2_X1 U7449 ( .A1(n5746), .A2(n7425), .ZN(n5840) );
  INV_X1 U7450 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7426) );
  OR2_X1 U7451 ( .A1(n5914), .A2(n7426), .ZN(n5839) );
  NAND2_X1 U7452 ( .A1(n6810), .A2(n8142), .ZN(n5849) );
  NOR2_X1 U7453 ( .A1(n5843), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5865) );
  OR2_X1 U7454 ( .A1(n5865), .A2(n7988), .ZN(n5846) );
  INV_X1 U7455 ( .A(n5846), .ZN(n5844) );
  NAND2_X1 U7456 ( .A1(n5844), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5847) );
  INV_X1 U7457 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7458 ( .A1(n5846), .A2(n5845), .ZN(n5852) );
  AND2_X1 U7459 ( .A1(n5847), .A2(n5852), .ZN(n6593) );
  AOI22_X1 U7460 ( .A1(n5962), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5961), .B2(
        n6593), .ZN(n5848) );
  NAND2_X1 U7461 ( .A1(n7451), .A2(n10291), .ZN(n5850) );
  INV_X1 U7462 ( .A(n7451), .ZN(n8517) );
  INV_X1 U7463 ( .A(n10291), .ZN(n7428) );
  NAND2_X1 U7464 ( .A1(n8517), .A2(n7428), .ZN(n5851) );
  NAND2_X1 U7465 ( .A1(n5852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5853) );
  XNOR2_X1 U7466 ( .A(n5853), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U7467 ( .A1(n5962), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5961), .B2(
        n10135), .ZN(n5854) );
  INV_X1 U7468 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7469 ( .A1(n5745), .A2(n5855), .ZN(n5861) );
  NAND2_X1 U7470 ( .A1(n5856), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5857) );
  AND2_X1 U7471 ( .A1(n5875), .A2(n5857), .ZN(n7715) );
  OR2_X1 U7472 ( .A1(n5746), .A2(n7715), .ZN(n5860) );
  INV_X1 U7473 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7452) );
  OR2_X1 U7474 ( .A1(n5914), .A2(n7452), .ZN(n5859) );
  NAND2_X1 U7475 ( .A1(n5744), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5858) );
  NAND4_X1 U7476 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n8516)
         );
  AND2_X1 U7477 ( .A1(n7714), .A2(n8516), .ZN(n5863) );
  OAI21_X1 U7478 ( .B1(n7449), .B2(n5863), .A(n5862), .ZN(n7471) );
  NAND2_X1 U7479 ( .A1(n6866), .A2(n8142), .ZN(n5872) );
  NOR2_X1 U7480 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5864) );
  AND2_X1 U7481 ( .A1(n5865), .A2(n5864), .ZN(n5869) );
  NOR2_X1 U7482 ( .A1(n5869), .A2(n7988), .ZN(n5866) );
  MUX2_X1 U7483 ( .A(n7988), .B(n5866), .S(P2_IR_REG_11__SCAN_IN), .Z(n5867)
         );
  INV_X1 U7484 ( .A(n5867), .ZN(n5870) );
  INV_X1 U7485 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7486 ( .A1(n5869), .A2(n5868), .ZN(n5893) );
  AND2_X1 U7487 ( .A1(n5870), .A2(n5893), .ZN(n10153) );
  AOI22_X1 U7488 ( .A1(n5962), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5961), .B2(
        n10153), .ZN(n5871) );
  NAND2_X1 U7489 ( .A1(n5872), .A2(n5871), .ZN(n7476) );
  NAND2_X1 U7490 ( .A1(n5744), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5880) );
  INV_X1 U7491 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5873) );
  OR2_X1 U7492 ( .A1(n5745), .A2(n5873), .ZN(n5879) );
  INV_X1 U7493 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5874) );
  OR2_X1 U7494 ( .A1(n5914), .A2(n5874), .ZN(n5878) );
  NAND2_X1 U7495 ( .A1(n5875), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5876) );
  AND2_X1 U7496 ( .A1(n5885), .A2(n5876), .ZN(n7477) );
  OR2_X1 U7497 ( .A1(n5746), .A2(n7477), .ZN(n5877) );
  NAND2_X1 U7498 ( .A1(n7476), .A2(n7827), .ZN(n8248) );
  AND2_X2 U7499 ( .A1(n8253), .A2(n8248), .ZN(n8162) );
  INV_X1 U7500 ( .A(n7827), .ZN(n8515) );
  NAND2_X1 U7501 ( .A1(n7476), .A2(n8515), .ZN(n5881) );
  NAND2_X1 U7502 ( .A1(n6986), .A2(n8142), .ZN(n5884) );
  NAND2_X1 U7503 ( .A1(n5893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U7504 ( .A(n5882), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U7505 ( .A1(n5962), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5961), .B2(
        n10168), .ZN(n5883) );
  INV_X1 U7506 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6519) );
  OR2_X1 U7507 ( .A1(n5745), .A2(n6519), .ZN(n5890) );
  AND2_X1 U7508 ( .A1(n5885), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5886) );
  NOR2_X1 U7509 ( .A1(n5899), .A2(n5886), .ZN(n7830) );
  OR2_X1 U7510 ( .A1(n5746), .A2(n7830), .ZN(n5889) );
  INV_X1 U7511 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7737) );
  OR2_X1 U7512 ( .A1(n5914), .A2(n7737), .ZN(n5888) );
  NAND2_X1 U7513 ( .A1(n5744), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5887) );
  NAND4_X1 U7514 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n8514)
         );
  OR2_X1 U7515 ( .A1(n10313), .A2(n8514), .ZN(n5891) );
  NAND2_X1 U7516 ( .A1(n10313), .A2(n8514), .ZN(n5892) );
  NAND2_X1 U7517 ( .A1(n7049), .A2(n8142), .ZN(n5896) );
  NAND2_X1 U7518 ( .A1(n5894), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5907) );
  XNOR2_X1 U7519 ( .A(n5907), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U7520 ( .A1(n5962), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5961), .B2(
        n10185), .ZN(n5895) );
  INV_X1 U7521 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10194) );
  OR2_X1 U7522 ( .A1(n5745), .A2(n10194), .ZN(n5904) );
  INV_X1 U7523 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5897) );
  OR2_X1 U7524 ( .A1(n5914), .A2(n5897), .ZN(n5903) );
  OR2_X1 U7525 ( .A1(n5899), .A2(n5898), .ZN(n5900) );
  AND2_X1 U7526 ( .A1(n5900), .A2(n5911), .ZN(n7816) );
  OR2_X1 U7527 ( .A1(n5746), .A2(n7816), .ZN(n5902) );
  NAND2_X1 U7528 ( .A1(n5744), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5901) );
  NAND4_X1 U7529 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n8513)
         );
  NAND2_X1 U7530 ( .A1(n7807), .A2(n7805), .ZN(n5905) );
  NAND2_X1 U7531 ( .A1(n7815), .A2(n8513), .ZN(n7804) );
  NAND2_X1 U7532 ( .A1(n5905), .A2(n7804), .ZN(n7882) );
  NAND2_X1 U7533 ( .A1(n7111), .A2(n8142), .ZN(n5910) );
  INV_X1 U7534 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7535 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U7536 ( .A1(n5908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7537 ( .A(n5922), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U7538 ( .A1(n5962), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5961), .B2(
        n10202), .ZN(n5909) );
  INV_X1 U7539 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9853) );
  OR2_X1 U7540 ( .A1(n5745), .A2(n9853), .ZN(n5918) );
  NAND2_X1 U7541 ( .A1(n5911), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5912) );
  AND2_X1 U7542 ( .A1(n5927), .A2(n5912), .ZN(n7891) );
  OR2_X1 U7543 ( .A1(n5746), .A2(n7891), .ZN(n5917) );
  INV_X1 U7544 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7545 ( .A1(n5914), .A2(n5913), .ZN(n5916) );
  NAND2_X1 U7546 ( .A1(n5744), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5915) );
  NAND4_X1 U7547 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n8512)
         );
  NAND2_X1 U7548 ( .A1(n7882), .A2(n5919), .ZN(n5921) );
  NAND2_X1 U7549 ( .A1(n7890), .A2(n8512), .ZN(n5920) );
  NAND2_X1 U7550 ( .A1(n5921), .A2(n5920), .ZN(n7951) );
  NAND2_X1 U7551 ( .A1(n5922), .A2(n5675), .ZN(n5923) );
  NAND2_X1 U7552 ( .A1(n5923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  XNOR2_X1 U7553 ( .A(n5924), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8555) );
  AOI22_X1 U7554 ( .A1(n5962), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5961), .B2(
        n8555), .ZN(n5925) );
  INV_X1 U7555 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9899) );
  OR2_X1 U7556 ( .A1(n5745), .A2(n9899), .ZN(n5933) );
  AND2_X1 U7557 ( .A1(n5927), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5928) );
  NOR2_X1 U7558 ( .A1(n5929), .A2(n5928), .ZN(n7959) );
  OR2_X1 U7559 ( .A1(n5746), .A2(n7959), .ZN(n5932) );
  INV_X1 U7560 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9868) );
  OR2_X1 U7561 ( .A1(n5914), .A2(n9868), .ZN(n5931) );
  NAND2_X1 U7562 ( .A1(n5744), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5930) );
  NAND4_X1 U7563 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n8511)
         );
  AND2_X1 U7564 ( .A1(n7961), .A2(n8511), .ZN(n7947) );
  NAND2_X1 U7565 ( .A1(n8048), .A2(n8720), .ZN(n8274) );
  NAND2_X1 U7566 ( .A1(n7153), .A2(n8142), .ZN(n5936) );
  NAND2_X1 U7567 ( .A1(n5941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7568 ( .A(n5934), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U7569 ( .A1(n5962), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5961), .B2(
        n10218), .ZN(n5935) );
  NAND2_X1 U7570 ( .A1(n5744), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5940) );
  INV_X1 U7571 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10231) );
  OR2_X1 U7572 ( .A1(n5745), .A2(n10231), .ZN(n5939) );
  INV_X1 U7573 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10226) );
  OR2_X1 U7574 ( .A1(n5914), .A2(n10226), .ZN(n5938) );
  XNOR2_X1 U7575 ( .A(n5949), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8025) );
  OR2_X1 U7576 ( .A1(n5746), .A2(n8025), .ZN(n5937) );
  NAND2_X1 U7577 ( .A1(n8829), .A2(n8708), .ZN(n8286) );
  NAND2_X1 U7578 ( .A1(n7116), .A2(n8142), .ZN(n5948) );
  INV_X1 U7579 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5942) );
  INV_X1 U7580 ( .A(n6058), .ZN(n5943) );
  NAND2_X1 U7581 ( .A1(n5943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7582 ( .A1(n5945), .A2(n5944), .ZN(n5958) );
  OR2_X1 U7583 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  AND2_X1 U7584 ( .A1(n5958), .A2(n5946), .ZN(n8595) );
  AOI22_X1 U7585 ( .A1(n5962), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5961), .B2(
        n8595), .ZN(n5947) );
  INV_X1 U7586 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9761) );
  OR2_X1 U7587 ( .A1(n6022), .A2(n9761), .ZN(n5955) );
  INV_X1 U7588 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U7589 ( .A1(n5949), .A2(n10240), .ZN(n5950) );
  NAND2_X1 U7590 ( .A1(n5950), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5951) );
  AND2_X1 U7591 ( .A1(n5951), .A2(n5965), .ZN(n8712) );
  OR2_X1 U7592 ( .A1(n5746), .A2(n8712), .ZN(n5954) );
  NAND2_X1 U7593 ( .A1(n6051), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7594 ( .A1(n6174), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5952) );
  NAND4_X1 U7595 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n8725)
         );
  NOR2_X1 U7596 ( .A1(n8764), .A2(n8725), .ZN(n5957) );
  INV_X1 U7597 ( .A(n8764), .ZN(n5956) );
  NAND2_X1 U7598 ( .A1(n7183), .A2(n8142), .ZN(n5964) );
  NAND2_X1 U7599 ( .A1(n5958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5960) );
  INV_X1 U7600 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5959) );
  INV_X1 U7601 ( .A(n8360), .ZN(n6610) );
  AOI22_X1 U7602 ( .A1(n5962), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6610), .B2(
        n5961), .ZN(n5963) );
  NAND2_X1 U7603 ( .A1(n5744), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5970) );
  INV_X1 U7604 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8761) );
  OR2_X1 U7605 ( .A1(n5745), .A2(n8761), .ZN(n5969) );
  INV_X1 U7606 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8699) );
  OR2_X1 U7607 ( .A1(n5914), .A2(n8699), .ZN(n5968) );
  NAND2_X1 U7608 ( .A1(n5965), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5966) );
  AND2_X1 U7609 ( .A1(n5973), .A2(n5966), .ZN(n8698) );
  OR2_X1 U7610 ( .A1(n5746), .A2(n8698), .ZN(n5967) );
  NAND2_X1 U7611 ( .A1(n8760), .A2(n8709), .ZN(n8304) );
  INV_X1 U7612 ( .A(n8709), .ZN(n8681) );
  NAND2_X1 U7613 ( .A1(n7227), .A2(n8142), .ZN(n5972) );
  OR2_X1 U7614 ( .A1(n5753), .A2(n7228), .ZN(n5971) );
  NAND2_X1 U7615 ( .A1(n5744), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7616 ( .A1(n6051), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5977) );
  AND2_X1 U7617 ( .A1(n5973), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5974) );
  OR2_X1 U7618 ( .A1(n5974), .A2(n5982), .ZN(n8686) );
  NAND2_X1 U7619 ( .A1(n5824), .A2(n8686), .ZN(n5976) );
  NAND2_X1 U7620 ( .A1(n6174), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5975) );
  NAND4_X1 U7621 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n8672)
         );
  NAND2_X1 U7622 ( .A1(n8108), .A2(n8672), .ZN(n8187) );
  NAND2_X1 U7623 ( .A1(n8680), .A2(n8679), .ZN(n8666) );
  NAND2_X1 U7624 ( .A1(n8108), .A2(n8697), .ZN(n8667) );
  NAND2_X1 U7625 ( .A1(n7275), .A2(n8142), .ZN(n5980) );
  OR2_X1 U7626 ( .A1(n5753), .A2(n7300), .ZN(n5979) );
  OR2_X1 U7627 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  NAND2_X1 U7628 ( .A1(n5992), .A2(n5983), .ZN(n8675) );
  NAND2_X1 U7629 ( .A1(n5824), .A2(n8675), .ZN(n5987) );
  INV_X1 U7630 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8808) );
  OR2_X1 U7631 ( .A1(n6022), .A2(n8808), .ZN(n5986) );
  INV_X1 U7632 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8753) );
  OR2_X1 U7633 ( .A1(n5745), .A2(n8753), .ZN(n5985) );
  INV_X1 U7634 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8674) );
  OR2_X1 U7635 ( .A1(n5914), .A2(n8674), .ZN(n5984) );
  NAND2_X1 U7636 ( .A1(n8809), .A2(n8111), .ZN(n8306) );
  AOI21_X1 U7637 ( .B1(n8666), .B2(n8667), .A(n8668), .ZN(n8652) );
  NOR2_X1 U7638 ( .A1(n8809), .A2(n8682), .ZN(n8654) );
  NAND2_X1 U7639 ( .A1(n7347), .A2(n8142), .ZN(n5989) );
  OR2_X1 U7640 ( .A1(n5753), .A2(n7348), .ZN(n5988) );
  NAND2_X1 U7641 ( .A1(n5744), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7642 ( .A1(n6051), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5990) );
  AND2_X1 U7643 ( .A1(n5991), .A2(n5990), .ZN(n5997) );
  NAND2_X1 U7644 ( .A1(n5992), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7645 ( .A1(n5994), .A2(n5993), .ZN(n8660) );
  NAND2_X1 U7646 ( .A1(n8660), .A2(n5824), .ZN(n5996) );
  NAND2_X1 U7647 ( .A1(n6174), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7648 ( .A1(n8803), .A2(n8642), .ZN(n8302) );
  NAND2_X1 U7649 ( .A1(n8309), .A2(n8302), .ZN(n8653) );
  OAI21_X1 U7650 ( .B1(n8652), .B2(n8654), .A(n8653), .ZN(n8656) );
  NAND2_X1 U7651 ( .A1(n8656), .A2(n5998), .ZN(n8640) );
  OAI21_X1 U7652 ( .B1(n8797), .B2(n8627), .A(n8640), .ZN(n5999) );
  NAND2_X1 U7653 ( .A1(n7468), .A2(n8142), .ZN(n6001) );
  OR2_X1 U7654 ( .A1(n5753), .A2(n8416), .ZN(n6000) );
  INV_X1 U7655 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6006) );
  AND2_X1 U7656 ( .A1(n6002), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6003) );
  NOR2_X2 U7657 ( .A1(n6002), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6011) );
  OR2_X1 U7658 ( .A1(n6003), .A2(n6011), .ZN(n8630) );
  NAND2_X1 U7659 ( .A1(n8630), .A2(n5824), .ZN(n6005) );
  AOI22_X1 U7660 ( .A1(n5744), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n6051), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n6004) );
  OAI211_X1 U7661 ( .C1(n5914), .C2(n6006), .A(n6005), .B(n6004), .ZN(n8508)
         );
  NOR2_X1 U7662 ( .A1(n8469), .A2(n8508), .ZN(n6007) );
  NAND2_X1 U7663 ( .A1(n7515), .A2(n8142), .ZN(n6009) );
  OR2_X1 U7664 ( .A1(n5753), .A2(n9822), .ZN(n6008) );
  INV_X1 U7665 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6010) );
  NOR2_X1 U7666 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  INV_X1 U7667 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7668 ( .A1(n6051), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7669 ( .A1(n5744), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6013) );
  OAI211_X1 U7670 ( .C1(n5914), .C2(n6015), .A(n6014), .B(n6013), .ZN(n6016)
         );
  NAND2_X1 U7671 ( .A1(n8461), .A2(n8628), .ZN(n8321) );
  NAND2_X1 U7672 ( .A1(n7723), .A2(n8142), .ZN(n6019) );
  OR2_X1 U7673 ( .A1(n5753), .A2(n6017), .ZN(n6018) );
  INV_X1 U7674 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8494) );
  NOR2_X1 U7675 ( .A1(n6020), .A2(n8494), .ZN(n6021) );
  NAND2_X1 U7676 ( .A1(n8614), .A2(n5824), .ZN(n6027) );
  INV_X1 U7677 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U7678 ( .A1(n6051), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6024) );
  INV_X1 U7679 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9772) );
  OR2_X1 U7680 ( .A1(n6022), .A2(n9772), .ZN(n6023) );
  OAI211_X1 U7681 ( .C1(n8613), .C2(n5914), .A(n6024), .B(n6023), .ZN(n6025)
         );
  INV_X1 U7682 ( .A(n6025), .ZN(n6026) );
  NAND2_X1 U7683 ( .A1(n6027), .A2(n6026), .ZN(n8507) );
  AND2_X1 U7684 ( .A1(n8786), .A2(n8507), .ZN(n6040) );
  NAND2_X1 U7685 ( .A1(n7727), .A2(n8142), .ZN(n6030) );
  OR2_X1 U7686 ( .A1(n5753), .A2(n6028), .ZN(n6029) );
  INV_X1 U7687 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7688 ( .A1(n6032), .A2(n6031), .ZN(n6049) );
  OR2_X1 U7689 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  NAND2_X1 U7690 ( .A1(n6049), .A2(n6033), .ZN(n8426) );
  NAND2_X1 U7691 ( .A1(n8426), .A2(n5824), .ZN(n6038) );
  NAND2_X1 U7692 ( .A1(n6051), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7693 ( .A1(n5744), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6034) );
  OAI211_X1 U7694 ( .C1(n5914), .C2(n6459), .A(n6035), .B(n6034), .ZN(n6036)
         );
  INV_X1 U7695 ( .A(n6036), .ZN(n6037) );
  NAND2_X1 U7696 ( .A1(n6038), .A2(n6037), .ZN(n8607) );
  AND2_X1 U7697 ( .A1(n8122), .A2(n8607), .ZN(n6045) );
  OR2_X1 U7698 ( .A1(n8122), .A2(n8607), .ZN(n6043) );
  INV_X1 U7699 ( .A(n8461), .ZN(n8619) );
  NAND2_X1 U7700 ( .A1(n8619), .A2(n8628), .ZN(n8603) );
  OR2_X1 U7701 ( .A1(n6040), .A2(n8603), .ZN(n6042) );
  INV_X1 U7702 ( .A(n8786), .ZN(n8504) );
  NAND2_X1 U7703 ( .A1(n8504), .A2(n8459), .ZN(n6041) );
  AND2_X1 U7704 ( .A1(n6043), .A2(n6433), .ZN(n6044) );
  NAND2_X1 U7705 ( .A1(n7741), .A2(n8142), .ZN(n6048) );
  OR2_X1 U7706 ( .A1(n5753), .A2(n6046), .ZN(n6047) );
  NAND2_X1 U7707 ( .A1(n6049), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7708 ( .A1(n8097), .A2(n6050), .ZN(n8126) );
  NAND2_X1 U7709 ( .A1(n8126), .A2(n5824), .ZN(n6056) );
  NAND2_X1 U7710 ( .A1(n6051), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7711 ( .A1(n5744), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6052) );
  OAI211_X1 U7712 ( .C1(n6118), .C2(n5914), .A(n6053), .B(n6052), .ZN(n6054)
         );
  INV_X1 U7713 ( .A(n6054), .ZN(n6055) );
  NOR2_X1 U7714 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6057) );
  INV_X1 U7715 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7716 ( .A1(n6062), .A2(n6059), .ZN(n6065) );
  OR2_X1 U7717 ( .A1(n6065), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7718 ( .A1(n6098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6060) );
  XNOR2_X1 U7719 ( .A(n6060), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U7720 ( .A1(n8364), .A2(n6610), .ZN(n6154) );
  INV_X1 U7721 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7722 ( .A1(n6063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6064) );
  MUX2_X1 U7723 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6064), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6066) );
  NAND2_X1 U7724 ( .A1(n6066), .A2(n6065), .ZN(n8359) );
  NAND2_X1 U7725 ( .A1(n8184), .A2(n6678), .ZN(n6067) );
  NAND2_X1 U7726 ( .A1(n6154), .A2(n6067), .ZN(n8684) );
  INV_X1 U7727 ( .A(n8097), .ZN(n6068) );
  NAND2_X1 U7728 ( .A1(n6068), .A2(n5824), .ZN(n7212) );
  INV_X1 U7729 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U7730 ( .A1(n5744), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6070) );
  INV_X1 U7731 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9644) );
  OR2_X1 U7732 ( .A1(n5745), .A2(n9644), .ZN(n6069) );
  OAI211_X1 U7733 ( .C1(n9837), .C2(n5914), .A(n6070), .B(n6069), .ZN(n6071)
         );
  INV_X1 U7734 ( .A(n6071), .ZN(n6072) );
  INV_X1 U7735 ( .A(n6167), .ZN(n8506) );
  INV_X1 U7736 ( .A(n6073), .ZN(n6530) );
  NAND2_X1 U7737 ( .A1(n6530), .A2(n6531), .ZN(n6075) );
  NAND2_X1 U7738 ( .A1(n6497), .A2(n6075), .ZN(n6748) );
  NAND2_X1 U7740 ( .A1(n6748), .A2(n8354), .ZN(n8710) );
  NAND2_X1 U7741 ( .A1(n8506), .A2(n10247), .ZN(n6078) );
  INV_X1 U7742 ( .A(n6748), .ZN(n6076) );
  NAND2_X1 U7743 ( .A1(n6088), .A2(n6081), .ZN(n6085) );
  OAI21_X1 U7744 ( .B1(n6088), .B2(n7988), .A(P2_IR_REG_24__SCAN_IN), .ZN(
        n6083) );
  NAND2_X1 U7745 ( .A1(n6085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7746 ( .A(n6086), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6095) );
  INV_X1 U7747 ( .A(n6095), .ZN(n7518) );
  INV_X1 U7748 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6789) );
  INV_X1 U7749 ( .A(n6097), .ZN(n6091) );
  INV_X1 U7750 ( .A(n6786), .ZN(n6092) );
  AND2_X1 U7751 ( .A1(n8364), .A2(n8360), .ZN(n6135) );
  NAND2_X1 U7752 ( .A1(n6135), .A2(n6678), .ZN(n6093) );
  INV_X1 U7753 ( .A(n6090), .ZN(n6094) );
  AND2_X1 U7754 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7755 ( .A1(n6097), .A2(n6096), .ZN(n6731) );
  AND2_X1 U7756 ( .A1(n6731), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7757 ( .B1(n6098), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6100) );
  INV_X1 U7758 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7759 ( .A(n6100), .B(n6099), .ZN(n6787) );
  NAND2_X1 U7760 ( .A1(n8359), .A2(n8360), .ZN(n6682) );
  NAND2_X1 U7761 ( .A1(n8354), .A2(n6682), .ZN(n6732) );
  NOR2_X1 U7762 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .ZN(
        n9648) );
  NOR4_X1 U7763 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6104) );
  NOR4_X1 U7764 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6103) );
  NOR4_X1 U7765 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6102) );
  NAND4_X1 U7766 ( .A1(n9648), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n6111)
         );
  NOR4_X1 U7767 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6108) );
  NOR4_X1 U7768 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6107) );
  NOR4_X1 U7769 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6106) );
  NOR4_X1 U7770 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6105) );
  NAND4_X1 U7771 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n6110)
         );
  OAI21_X1 U7772 ( .B1(n6111), .B2(n6110), .A(n6109), .ZN(n6733) );
  AND3_X1 U7773 ( .A1(n6785), .A2(n6732), .A3(n6733), .ZN(n6115) );
  INV_X1 U7774 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7775 ( .A1(n6109), .A2(n6112), .ZN(n6114) );
  NAND2_X1 U7776 ( .A1(n6091), .A2(n7518), .ZN(n6113) );
  AND2_X1 U7777 ( .A1(n6114), .A2(n6113), .ZN(n6774) );
  NAND2_X1 U7778 ( .A1(n6677), .A2(n6774), .ZN(n6735) );
  AND2_X1 U7779 ( .A1(n6115), .A2(n6735), .ZN(n6454) );
  INV_X1 U7780 ( .A(n6774), .ZN(n6449) );
  NAND2_X1 U7781 ( .A1(n6448), .A2(n6449), .ZN(n6116) );
  OAI211_X1 U7782 ( .C1(n6677), .C2(n6448), .A(n6454), .B(n6116), .ZN(n6140)
         );
  INV_X1 U7783 ( .A(n8364), .ZN(n7349) );
  AND2_X1 U7784 ( .A1(n8359), .A2(n6610), .ZN(n6160) );
  NAND2_X1 U7785 ( .A1(n10314), .A2(n6160), .ZN(n6446) );
  INV_X1 U7786 ( .A(n6446), .ZN(n6117) );
  NAND2_X1 U7787 ( .A1(n6117), .A2(n6785), .ZN(n8711) );
  INV_X1 U7789 ( .A(n6943), .ZN(n6119) );
  NAND2_X1 U7790 ( .A1(n6119), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U7791 ( .A1(n6944), .A2(n8197), .ZN(n10243) );
  INV_X1 U7792 ( .A(n6120), .ZN(n8148) );
  NAND2_X1 U7793 ( .A1(n10243), .A2(n8148), .ZN(n10242) );
  INV_X1 U7794 ( .A(n10265), .ZN(n6121) );
  NAND2_X1 U7795 ( .A1(n10246), .A2(n6121), .ZN(n8217) );
  NAND2_X1 U7796 ( .A1(n6123), .A2(n6122), .ZN(n8210) );
  NAND2_X1 U7797 ( .A1(n7199), .A2(n7157), .ZN(n8213) );
  NAND2_X1 U7798 ( .A1(n7160), .A2(n7030), .ZN(n7103) );
  AND2_X1 U7799 ( .A1(n8213), .A2(n7103), .ZN(n8218) );
  NAND2_X1 U7800 ( .A1(n7009), .A2(n8218), .ZN(n6124) );
  NAND2_X1 U7801 ( .A1(n8521), .A2(n10277), .ZN(n8221) );
  NAND2_X1 U7802 ( .A1(n6707), .A2(n7123), .ZN(n8223) );
  NAND2_X1 U7803 ( .A1(n8520), .A2(n10281), .ZN(n8225) );
  NAND2_X1 U7804 ( .A1(n8223), .A2(n8225), .ZN(n7119) );
  INV_X1 U7805 ( .A(n8230), .ZN(n8159) );
  INV_X1 U7806 ( .A(n7308), .ZN(n8239) );
  NAND2_X1 U7807 ( .A1(n8519), .A2(n8239), .ZN(n7317) );
  AND2_X1 U7808 ( .A1(n8227), .A2(n7317), .ZN(n8233) );
  NAND2_X1 U7809 ( .A1(n7219), .A2(n8233), .ZN(n6125) );
  NAND2_X1 U7810 ( .A1(n6125), .A2(n8238), .ZN(n7418) );
  NAND2_X1 U7811 ( .A1(n7451), .A2(n7428), .ZN(n8242) );
  NAND2_X1 U7812 ( .A1(n8517), .A2(n10291), .ZN(n8236) );
  NAND2_X1 U7813 ( .A1(n8242), .A2(n8236), .ZN(n7421) );
  INV_X1 U7814 ( .A(n8516), .ZN(n7770) );
  NAND2_X1 U7815 ( .A1(n7714), .A2(n7770), .ZN(n8243) );
  AND2_X1 U7816 ( .A1(n8248), .A2(n8243), .ZN(n8255) );
  XNOR2_X1 U7817 ( .A(n10313), .B(n8514), .ZN(n8250) );
  NAND2_X1 U7818 ( .A1(n6126), .A2(n8250), .ZN(n7733) );
  INV_X1 U7819 ( .A(n8514), .ZN(n8252) );
  OR2_X1 U7820 ( .A1(n10313), .A2(n8252), .ZN(n6127) );
  INV_X1 U7821 ( .A(n8513), .ZN(n7736) );
  NAND2_X1 U7822 ( .A1(n7815), .A2(n7736), .ZN(n8262) );
  NAND2_X1 U7823 ( .A1(n7806), .A2(n8262), .ZN(n6128) );
  OR2_X1 U7824 ( .A1(n7815), .A2(n7736), .ZN(n8261) );
  NAND2_X1 U7825 ( .A1(n6128), .A2(n8261), .ZN(n7881) );
  INV_X1 U7826 ( .A(n8512), .ZN(n7834) );
  NAND2_X1 U7827 ( .A1(n7890), .A2(n7834), .ZN(n8269) );
  OR2_X1 U7828 ( .A1(n7890), .A2(n7834), .ZN(n8266) );
  INV_X1 U7829 ( .A(n8511), .ZN(n7965) );
  NAND2_X1 U7830 ( .A1(n7961), .A2(n7965), .ZN(n8270) );
  AND2_X1 U7831 ( .A1(n8274), .A2(n8270), .ZN(n8279) );
  NAND2_X1 U7832 ( .A1(n8031), .A2(n8279), .ZN(n6129) );
  NAND2_X1 U7833 ( .A1(n8764), .A2(n8696), .ZN(n8283) );
  NAND2_X1 U7834 ( .A1(n8703), .A2(n8276), .ZN(n8690) );
  INV_X1 U7835 ( .A(n8693), .ZN(n8689) );
  NAND2_X1 U7836 ( .A1(n8690), .A2(n8689), .ZN(n8692) );
  AND2_X1 U7837 ( .A1(n8306), .A2(n8663), .ZN(n8188) );
  NAND2_X1 U7838 ( .A1(n6130), .A2(n8300), .ZN(n8650) );
  NAND2_X1 U7839 ( .A1(n8650), .A2(n8302), .ZN(n6131) );
  NAND2_X1 U7840 ( .A1(n8469), .A2(n8643), .ZN(n8316) );
  NAND2_X1 U7841 ( .A1(n8647), .A2(n8627), .ZN(n8633) );
  INV_X1 U7842 ( .A(n8312), .ZN(n6132) );
  OR2_X1 U7843 ( .A1(n8469), .A2(n8643), .ZN(n8311) );
  OAI21_X2 U7844 ( .B1(n8602), .B2(n8147), .A(n8324), .ZN(n6440) );
  NAND2_X1 U7845 ( .A1(n8122), .A2(n8497), .ZN(n8331) );
  NAND2_X1 U7846 ( .A1(n6440), .A2(n8331), .ZN(n6134) );
  NAND2_X1 U7847 ( .A1(n6134), .A2(n8330), .ZN(n6170) );
  OR2_X1 U7848 ( .A1(n8349), .A2(n6682), .ZN(n6746) );
  INV_X1 U7849 ( .A(n6135), .ZN(n6136) );
  NAND2_X1 U7850 ( .A1(n6136), .A2(n6682), .ZN(n6137) );
  NAND3_X1 U7851 ( .A1(n6746), .A2(n10303), .A3(n6137), .ZN(n10244) );
  NAND2_X1 U7852 ( .A1(n6160), .A2(n8184), .ZN(n10255) );
  NAND2_X1 U7853 ( .A1(n10244), .A2(n10255), .ZN(n6138) );
  NAND2_X1 U7854 ( .A1(n8714), .A2(n6138), .ZN(n8731) );
  INV_X1 U7855 ( .A(n6160), .ZN(n6139) );
  NAND2_X1 U7856 ( .A1(n10314), .A2(n6139), .ZN(n10254) );
  OR2_X1 U7857 ( .A1(n6140), .A2(n10254), .ZN(n8601) );
  INV_X1 U7858 ( .A(n8711), .ZN(n10257) );
  AOI22_X1 U7859 ( .A1(n8781), .A2(n8728), .B1(n10257), .B2(n8126), .ZN(n6141)
         );
  INV_X1 U7860 ( .A(n6142), .ZN(n6143) );
  INV_X1 U7861 ( .A(n6432), .ZN(n6146) );
  INV_X1 U7862 ( .A(n8318), .ZN(n6145) );
  INV_X1 U7863 ( .A(n8684), .ZN(n10252) );
  INV_X1 U7864 ( .A(n10248), .ZN(n8719) );
  OAI22_X1 U7865 ( .A1(n8459), .A2(n8710), .B1(n8719), .B2(n8643), .ZN(n6149)
         );
  INV_X1 U7866 ( .A(n6149), .ZN(n6150) );
  INV_X1 U7867 ( .A(n6677), .ZN(n6152) );
  AND3_X1 U7868 ( .A1(n6152), .A2(n6449), .A3(n6733), .ZN(n6741) );
  AND2_X1 U7869 ( .A1(n6741), .A2(n6785), .ZN(n6750) );
  NAND2_X1 U7870 ( .A1(n8196), .A2(n6678), .ZN(n6153) );
  OR2_X1 U7871 ( .A1(n6154), .A2(n6153), .ZN(n6739) );
  NAND3_X1 U7872 ( .A1(n8349), .A2(n10303), .A3(n6739), .ZN(n6720) );
  NAND2_X1 U7873 ( .A1(n6720), .A2(n10254), .ZN(n6734) );
  NAND2_X1 U7874 ( .A1(n6750), .A2(n6734), .ZN(n6157) );
  INV_X1 U7875 ( .A(n6746), .ZN(n6890) );
  INV_X1 U7876 ( .A(n6739), .ZN(n6719) );
  NAND2_X1 U7877 ( .A1(n6785), .A2(n6733), .ZN(n6155) );
  NOR2_X1 U7878 ( .A1(n6735), .A2(n6155), .ZN(n6729) );
  OAI21_X1 U7879 ( .B1(n6890), .B2(n6719), .A(n6729), .ZN(n6156) );
  INV_X2 U7880 ( .A(n10317), .ZN(n10315) );
  MUX2_X1 U7881 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8621), .S(n10315), .Z(n6158) );
  INV_X1 U7882 ( .A(n6158), .ZN(n6163) );
  XNOR2_X1 U7883 ( .A(n6159), .B(n8318), .ZN(n8624) );
  NAND2_X1 U7884 ( .A1(n7349), .A2(n6160), .ZN(n10292) );
  NAND2_X1 U7885 ( .A1(n10244), .A2(n10292), .ZN(n10306) );
  INV_X1 U7886 ( .A(n10306), .ZN(n10309) );
  OR2_X1 U7887 ( .A1(n10317), .A2(n10303), .ZN(n8796) );
  OAI22_X1 U7888 ( .A1(n8624), .A2(n8832), .B1(n8619), .B2(n8796), .ZN(n6161)
         );
  INV_X1 U7889 ( .A(n6161), .ZN(n6162) );
  NAND2_X1 U7890 ( .A1(n6163), .A2(n6162), .ZN(P2_U3452) );
  NOR2_X1 U7891 ( .A1(n8340), .A2(n8337), .ZN(n6164) );
  OAI22_X1 U7892 ( .A1(n6165), .A2(n6164), .B1(n4603), .B2(n8781), .ZN(n6168)
         );
  INV_X1 U7893 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7926) );
  OR2_X1 U7894 ( .A1(n5753), .A2(n7926), .ZN(n6166) );
  NAND2_X1 U7895 ( .A1(n8099), .A2(n6167), .ZN(n8181) );
  XNOR2_X1 U7896 ( .A(n6168), .B(n8335), .ZN(n6182) );
  NAND2_X1 U7897 ( .A1(n8781), .A2(n8337), .ZN(n6169) );
  NAND2_X1 U7898 ( .A1(n6170), .A2(n6169), .ZN(n6172) );
  NAND2_X1 U7899 ( .A1(n6172), .A2(n6171), .ZN(n8178) );
  XOR2_X1 U7900 ( .A(n8178), .B(n8173), .Z(n6173) );
  INV_X1 U7901 ( .A(n6173), .ZN(n6183) );
  INV_X1 U7902 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U7903 ( .A1(n5744), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7904 ( .A1(n6174), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6175) );
  OAI211_X1 U7905 ( .C1(n5745), .C2(n9735), .A(n6176), .B(n6175), .ZN(n6177)
         );
  INV_X1 U7906 ( .A(n6177), .ZN(n6178) );
  NAND2_X1 U7907 ( .A1(n7212), .A2(n6178), .ZN(n8505) );
  AND2_X1 U7908 ( .A1(n6497), .A2(P2_B_REG_SCAN_IN), .ZN(n6179) );
  NOR2_X1 U7909 ( .A1(n8710), .A2(n6179), .ZN(n8000) );
  AOI22_X1 U7910 ( .A1(n8505), .A2(n8000), .B1(n4603), .B2(n10248), .ZN(n6180)
         );
  OAI21_X1 U7911 ( .B1(n6183), .B2(n10244), .A(n6180), .ZN(n6181) );
  INV_X1 U7912 ( .A(n10292), .ZN(n6184) );
  INV_X1 U7913 ( .A(n8099), .ZN(n6674) );
  NOR2_X1 U7914 ( .A1(n6674), .A2(n8796), .ZN(n6186) );
  NAND2_X1 U7915 ( .A1(n6188), .A2(n6187), .ZN(P2_U3456) );
  NAND2_X1 U7916 ( .A1(n6792), .A2(n6189), .ZN(n6253) );
  INV_X4 U7917 ( .A(n6253), .ZN(n6397) );
  AOI22_X1 U7918 ( .A1(n7577), .A2(n6397), .B1(n6392), .B2(n9202), .ZN(n6248)
         );
  AND2_X1 U7919 ( .A1(n6792), .A2(n6192), .ZN(n6193) );
  NAND2_X2 U7920 ( .A1(n6191), .A2(n6193), .ZN(n6196) );
  NAND2_X1 U7921 ( .A1(n7577), .A2(n6387), .ZN(n6195) );
  NAND2_X1 U7922 ( .A1(n9202), .A2(n6397), .ZN(n6194) );
  NAND2_X1 U7923 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  XNOR2_X1 U7924 ( .A(n6197), .B(n6196), .ZN(n6247) );
  AND2_X1 U7925 ( .A1(n6199), .A2(n6397), .ZN(n6198) );
  AOI21_X1 U7926 ( .B1(n9207), .B2(n6392), .A(n6198), .ZN(n6225) );
  NAND2_X1 U7927 ( .A1(n6387), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7928 ( .A1(n9207), .A2(n6397), .ZN(n6200) );
  NAND2_X1 U7929 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  XNOR2_X1 U7930 ( .A(n6202), .B(n6388), .ZN(n6224) );
  AND2_X1 U7931 ( .A1(n7682), .A2(n6397), .ZN(n6203) );
  AOI21_X1 U7932 ( .B1(n9208), .B2(n6392), .A(n6203), .ZN(n6222) );
  AOI22_X1 U7933 ( .A1(n9208), .A2(n6397), .B1(n7682), .B2(n6214), .ZN(n6204)
         );
  XNOR2_X1 U7934 ( .A(n6204), .B(n6388), .ZN(n6223) );
  XOR2_X1 U7935 ( .A(n6222), .B(n6223), .Z(n7043) );
  INV_X1 U7936 ( .A(n6792), .ZN(n6205) );
  AOI222_X1 U7937 ( .A1(n8073), .A2(n6392), .B1(n7511), .B2(n6397), .C1(n6205), 
        .C2(P1_IR_REG_0__SCAN_IN), .ZN(n6898) );
  AOI21_X1 U7938 ( .B1(n6205), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6206), .ZN(
        n6897) );
  OAI21_X1 U7939 ( .B1(n6898), .B2(n6897), .A(n6207), .ZN(n7131) );
  NAND2_X1 U7940 ( .A1(n9211), .A2(n6397), .ZN(n6208) );
  OAI21_X1 U7941 ( .B1(n6213), .B2(n5123), .A(n6208), .ZN(n6209) );
  XNOR2_X1 U7942 ( .A(n6209), .B(n6395), .ZN(n6212) );
  AND2_X1 U7943 ( .A1(n7133), .A2(n6397), .ZN(n6210) );
  AOI21_X1 U7944 ( .B1(n9211), .B2(n6392), .A(n6210), .ZN(n6211) );
  NOR2_X1 U7945 ( .A1(n6212), .A2(n6211), .ZN(n7129) );
  NOR2_X1 U7946 ( .A1(n7131), .A2(n7129), .ZN(n7127) );
  AND2_X1 U7947 ( .A1(n6212), .A2(n6211), .ZN(n7128) );
  NOR2_X1 U7948 ( .A1(n7127), .A2(n7128), .ZN(n7145) );
  AOI22_X1 U7949 ( .A1(n9209), .A2(n6392), .B1(n6397), .B2(n7645), .ZN(n6218)
         );
  INV_X1 U7950 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7951 ( .A1(n9209), .A2(n6397), .ZN(n6215) );
  NAND2_X1 U7952 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  INV_X1 U7953 ( .A(n6218), .ZN(n6219) );
  XNOR2_X1 U7954 ( .A(n6224), .B(n6225), .ZN(n7061) );
  AOI22_X1 U7955 ( .A1(n9206), .A2(n6397), .B1(n7664), .B2(n6387), .ZN(n6226)
         );
  XOR2_X1 U7956 ( .A(n6196), .B(n6226), .Z(n6227) );
  AOI22_X1 U7957 ( .A1(n9206), .A2(n6392), .B1(n6397), .B2(n7664), .ZN(n7260)
         );
  NAND2_X1 U7958 ( .A1(n9205), .A2(n6397), .ZN(n6229) );
  NAND2_X1 U7959 ( .A1(n6387), .A2(n7436), .ZN(n6228) );
  NAND2_X1 U7960 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  XNOR2_X1 U7961 ( .A(n6230), .B(n6395), .ZN(n6233) );
  AND2_X1 U7962 ( .A1(n7436), .A2(n6397), .ZN(n6231) );
  AOI21_X1 U7963 ( .B1(n9205), .B2(n6392), .A(n6231), .ZN(n6232) );
  NOR2_X1 U7964 ( .A1(n6233), .A2(n6232), .ZN(n7291) );
  NAND2_X1 U7965 ( .A1(n6233), .A2(n6232), .ZN(n7289) );
  NAND2_X1 U7966 ( .A1(n9204), .A2(n6397), .ZN(n6235) );
  NAND2_X1 U7967 ( .A1(n7639), .A2(n6387), .ZN(n6234) );
  NAND2_X1 U7968 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  XNOR2_X1 U7969 ( .A(n6236), .B(n6395), .ZN(n6237) );
  AOI22_X1 U7970 ( .A1(n9204), .A2(n6392), .B1(n7639), .B2(n6397), .ZN(n6238)
         );
  AND2_X1 U7971 ( .A1(n6237), .A2(n6238), .ZN(n7380) );
  INV_X1 U7972 ( .A(n6237), .ZN(n6240) );
  INV_X1 U7973 ( .A(n6238), .ZN(n6239) );
  NAND2_X1 U7974 ( .A1(n6240), .A2(n6239), .ZN(n7379) );
  OAI21_X2 U7975 ( .B1(n7383), .B2(n7380), .A(n7379), .ZN(n7399) );
  NAND2_X1 U7976 ( .A1(n7585), .A2(n6387), .ZN(n6242) );
  NAND2_X1 U7977 ( .A1(n9203), .A2(n6397), .ZN(n6241) );
  NAND2_X1 U7978 ( .A1(n6242), .A2(n6241), .ZN(n6243) );
  XNOR2_X1 U7979 ( .A(n6243), .B(n6388), .ZN(n6244) );
  AOI22_X1 U7980 ( .A1(n7585), .A2(n6397), .B1(n6392), .B2(n9203), .ZN(n6245)
         );
  XNOR2_X1 U7981 ( .A(n6244), .B(n6245), .ZN(n7398) );
  NAND2_X1 U7982 ( .A1(n7399), .A2(n7398), .ZN(n7397) );
  INV_X1 U7983 ( .A(n6244), .ZN(n6246) );
  NAND2_X1 U7984 ( .A1(n7397), .A2(n4907), .ZN(n7483) );
  XNOR2_X1 U7985 ( .A(n6247), .B(n6248), .ZN(n7482) );
  NAND2_X1 U7986 ( .A1(n10008), .A2(n6387), .ZN(n6250) );
  NAND2_X1 U7987 ( .A1(n9200), .A2(n6397), .ZN(n6249) );
  NAND2_X1 U7988 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  XNOR2_X1 U7989 ( .A(n6251), .B(n6196), .ZN(n7848) );
  OAI22_X1 U7990 ( .A1(n10079), .A2(n6253), .B1(n8965), .B2(n6252), .ZN(n7847)
         );
  NAND2_X1 U7991 ( .A1(n7848), .A2(n7847), .ZN(n7846) );
  INV_X1 U7992 ( .A(n7846), .ZN(n6260) );
  NAND2_X1 U7993 ( .A1(n7759), .A2(n6387), .ZN(n6255) );
  NAND2_X1 U7994 ( .A1(n9201), .A2(n6397), .ZN(n6254) );
  NAND2_X1 U7995 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  XNOR2_X1 U7996 ( .A(n6256), .B(n6395), .ZN(n7850) );
  NAND2_X1 U7997 ( .A1(n7759), .A2(n6397), .ZN(n6258) );
  NAND2_X1 U7998 ( .A1(n9201), .A2(n6392), .ZN(n6257) );
  INV_X1 U7999 ( .A(n7847), .ZN(n6262) );
  AOI21_X1 U8000 ( .B1(n7850), .B2(n7752), .A(n6262), .ZN(n6261) );
  NAND3_X1 U8001 ( .A1(n6262), .A2(n7752), .A3(n7850), .ZN(n6263) );
  NAND2_X1 U8002 ( .A1(n5606), .A2(n6387), .ZN(n6267) );
  NAND2_X1 U8003 ( .A1(n9984), .A2(n6397), .ZN(n6266) );
  NAND2_X1 U8004 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  XNOR2_X1 U8005 ( .A(n6268), .B(n6196), .ZN(n6272) );
  NAND2_X1 U8006 ( .A1(n5606), .A2(n6397), .ZN(n6270) );
  NAND2_X1 U8007 ( .A1(n9984), .A2(n6392), .ZN(n6269) );
  NAND2_X1 U8008 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  AOI21_X1 U8009 ( .B1(n6272), .B2(n6271), .A(n6273), .ZN(n7779) );
  INV_X1 U8010 ( .A(n6273), .ZN(n6274) );
  NAND2_X1 U8011 ( .A1(n7777), .A2(n6274), .ZN(n7858) );
  NAND2_X1 U8012 ( .A1(n9969), .A2(n6387), .ZN(n6276) );
  NAND2_X1 U8013 ( .A1(n9199), .A2(n6397), .ZN(n6275) );
  NAND2_X1 U8014 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  XNOR2_X1 U8015 ( .A(n6277), .B(n6196), .ZN(n6280) );
  AOI22_X1 U8016 ( .A1(n9969), .A2(n6397), .B1(n6392), .B2(n9199), .ZN(n6278)
         );
  XNOR2_X1 U8017 ( .A(n6280), .B(n6278), .ZN(n7859) );
  INV_X1 U8018 ( .A(n6278), .ZN(n6279) );
  NAND2_X1 U8019 ( .A1(n7857), .A2(n6281), .ZN(n6286) );
  INV_X1 U8020 ( .A(n6286), .ZN(n6284) );
  AOI22_X1 U8021 ( .A1(n7794), .A2(n6387), .B1(n6397), .B2(n9983), .ZN(n6282)
         );
  XNOR2_X1 U8022 ( .A(n6282), .B(n6196), .ZN(n6285) );
  INV_X1 U8023 ( .A(n6285), .ZN(n6283) );
  NAND2_X1 U8024 ( .A1(n6284), .A2(n6283), .ZN(n6287) );
  NAND2_X1 U8025 ( .A1(n6286), .A2(n6285), .ZN(n6288) );
  AOI22_X1 U8026 ( .A1(n7794), .A2(n6397), .B1(n6392), .B2(n9983), .ZN(n8053)
         );
  NAND2_X1 U8027 ( .A1(n8052), .A2(n6288), .ZN(n6292) );
  AOI22_X1 U8028 ( .A1(n9623), .A2(n6387), .B1(n6397), .B2(n9198), .ZN(n6289)
         );
  XNOR2_X1 U8029 ( .A(n6289), .B(n6196), .ZN(n6291) );
  INV_X1 U8030 ( .A(n6291), .ZN(n6290) );
  AOI22_X1 U8031 ( .A1(n9623), .A2(n6397), .B1(n6392), .B2(n9198), .ZN(n8916)
         );
  NAND2_X1 U8032 ( .A1(n8915), .A2(n6293), .ZN(n8858) );
  NAND2_X1 U8033 ( .A1(n7908), .A2(n6387), .ZN(n6295) );
  NAND2_X1 U8034 ( .A1(n9197), .A2(n6397), .ZN(n6294) );
  NAND2_X1 U8035 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  XNOR2_X1 U8036 ( .A(n6296), .B(n6196), .ZN(n6297) );
  AOI22_X1 U8037 ( .A1(n7908), .A2(n6397), .B1(n6392), .B2(n9197), .ZN(n6298)
         );
  XNOR2_X1 U8038 ( .A(n6297), .B(n6298), .ZN(n8860) );
  NAND2_X1 U8039 ( .A1(n8858), .A2(n8860), .ZN(n8859) );
  INV_X1 U8040 ( .A(n6297), .ZN(n6299) );
  NAND2_X1 U8041 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  NAND2_X1 U8042 ( .A1(n8859), .A2(n6300), .ZN(n8869) );
  NAND2_X1 U8043 ( .A1(n9619), .A2(n6214), .ZN(n6302) );
  NAND2_X1 U8044 ( .A1(n9196), .A2(n6397), .ZN(n6301) );
  NAND2_X1 U8045 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  XNOR2_X1 U8046 ( .A(n6303), .B(n6388), .ZN(n6306) );
  NAND2_X1 U8047 ( .A1(n9619), .A2(n6397), .ZN(n6305) );
  NAND2_X1 U8048 ( .A1(n9196), .A2(n6392), .ZN(n6304) );
  NAND2_X1 U8049 ( .A1(n6305), .A2(n6304), .ZN(n6307) );
  NAND2_X1 U8050 ( .A1(n6306), .A2(n6307), .ZN(n8871) );
  NAND2_X1 U8051 ( .A1(n8869), .A2(n8871), .ZN(n6310) );
  INV_X1 U8052 ( .A(n6306), .ZN(n6309) );
  INV_X1 U8053 ( .A(n6307), .ZN(n6308) );
  NAND2_X1 U8054 ( .A1(n6309), .A2(n6308), .ZN(n8870) );
  NAND2_X1 U8055 ( .A1(n8910), .A2(n6387), .ZN(n6312) );
  NAND2_X1 U8056 ( .A1(n9195), .A2(n6397), .ZN(n6311) );
  NAND2_X1 U8057 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  XNOR2_X1 U8058 ( .A(n6313), .B(n6196), .ZN(n8901) );
  NAND2_X1 U8059 ( .A1(n8910), .A2(n6397), .ZN(n6315) );
  NAND2_X1 U8060 ( .A1(n9195), .A2(n6392), .ZN(n6314) );
  NAND2_X1 U8061 ( .A1(n6315), .A2(n6314), .ZN(n8900) );
  NOR2_X1 U8062 ( .A1(n8901), .A2(n8900), .ZN(n6318) );
  INV_X1 U8063 ( .A(n8901), .ZN(n6317) );
  INV_X1 U8064 ( .A(n8900), .ZN(n6316) );
  NAND2_X1 U8065 ( .A1(n9608), .A2(n6387), .ZN(n6320) );
  NAND2_X1 U8066 ( .A1(n9523), .A2(n6397), .ZN(n6319) );
  NAND2_X1 U8067 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  XNOR2_X1 U8068 ( .A(n6321), .B(n6395), .ZN(n6324) );
  AND2_X1 U8069 ( .A1(n9523), .A2(n6392), .ZN(n6322) );
  AOI21_X1 U8070 ( .B1(n9608), .B2(n6397), .A(n6322), .ZN(n6323) );
  NOR2_X1 U8071 ( .A1(n6324), .A2(n6323), .ZN(n8838) );
  NAND2_X1 U8072 ( .A1(n6324), .A2(n6323), .ZN(n8836) );
  NAND2_X1 U8073 ( .A1(n8835), .A2(n8836), .ZN(n8848) );
  NAND2_X1 U8074 ( .A1(n9530), .A2(n6214), .ZN(n6326) );
  NAND2_X1 U8075 ( .A1(n9511), .A2(n6397), .ZN(n6325) );
  NAND2_X1 U8076 ( .A1(n6326), .A2(n6325), .ZN(n6327) );
  XNOR2_X1 U8077 ( .A(n6327), .B(n6388), .ZN(n6337) );
  AOI22_X1 U8078 ( .A1(n9530), .A2(n6397), .B1(n6392), .B2(n9511), .ZN(n6338)
         );
  XNOR2_X1 U8079 ( .A(n6337), .B(n6338), .ZN(n8882) );
  NAND2_X1 U8080 ( .A1(n9597), .A2(n6214), .ZN(n6329) );
  NAND2_X1 U8081 ( .A1(n9524), .A2(n6397), .ZN(n6328) );
  NAND2_X1 U8082 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  XNOR2_X1 U8083 ( .A(n6330), .B(n6388), .ZN(n6333) );
  INV_X1 U8084 ( .A(n6333), .ZN(n6331) );
  AOI22_X1 U8085 ( .A1(n9597), .A2(n6397), .B1(n6392), .B2(n9524), .ZN(n6332)
         );
  NAND2_X1 U8086 ( .A1(n6331), .A2(n6332), .ZN(n6340) );
  INV_X1 U8087 ( .A(n6340), .ZN(n6334) );
  XNOR2_X1 U8088 ( .A(n6333), .B(n6332), .ZN(n8851) );
  NAND2_X1 U8089 ( .A1(n8848), .A2(n6335), .ZN(n6344) );
  INV_X1 U8090 ( .A(n6336), .ZN(n6342) );
  INV_X1 U8091 ( .A(n6337), .ZN(n6339) );
  NAND2_X1 U8092 ( .A1(n6339), .A2(n6338), .ZN(n8849) );
  AND2_X1 U8093 ( .A1(n8849), .A2(n6340), .ZN(n6341) );
  NAND2_X1 U8094 ( .A1(n9588), .A2(n6214), .ZN(n6346) );
  NAND2_X1 U8095 ( .A1(n9489), .A2(n6397), .ZN(n6345) );
  NAND2_X1 U8096 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  XNOR2_X1 U8097 ( .A(n6347), .B(n6395), .ZN(n8374) );
  AOI22_X1 U8098 ( .A1(n9588), .A2(n6397), .B1(n6392), .B2(n9489), .ZN(n8373)
         );
  NAND2_X1 U8099 ( .A1(n9494), .A2(n6387), .ZN(n6349) );
  NAND2_X1 U8100 ( .A1(n9512), .A2(n6397), .ZN(n6348) );
  NAND2_X1 U8101 ( .A1(n6349), .A2(n6348), .ZN(n6350) );
  NAND2_X1 U8102 ( .A1(n9494), .A2(n6397), .ZN(n6352) );
  NAND2_X1 U8103 ( .A1(n9512), .A2(n6392), .ZN(n6351) );
  NAND2_X1 U8104 ( .A1(n6352), .A2(n6351), .ZN(n8368) );
  NAND2_X1 U8105 ( .A1(n8370), .A2(n8368), .ZN(n6353) );
  INV_X1 U8106 ( .A(n8373), .ZN(n6356) );
  OAI21_X1 U8107 ( .B1(n8370), .B2(n8368), .A(n6356), .ZN(n6358) );
  NOR3_X1 U8108 ( .A1(n6356), .A2(n8370), .A3(n8368), .ZN(n6357) );
  AOI21_X1 U8109 ( .B1(n8374), .B2(n6358), .A(n6357), .ZN(n6465) );
  AND2_X1 U8110 ( .A1(n8403), .A2(n6392), .ZN(n6359) );
  AOI21_X1 U8111 ( .B1(n9430), .B2(n6397), .A(n6359), .ZN(n6384) );
  NAND2_X1 U8112 ( .A1(n9430), .A2(n6214), .ZN(n6361) );
  NAND2_X1 U8113 ( .A1(n8403), .A2(n6397), .ZN(n6360) );
  NAND2_X1 U8114 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  XNOR2_X1 U8115 ( .A(n6362), .B(n6388), .ZN(n6386) );
  XOR2_X1 U8116 ( .A(n6384), .B(n6386), .Z(n6470) );
  INV_X1 U8117 ( .A(n6470), .ZN(n6377) );
  NAND2_X1 U8118 ( .A1(n9575), .A2(n6214), .ZN(n6364) );
  NAND2_X1 U8119 ( .A1(n9458), .A2(n6397), .ZN(n6363) );
  NAND2_X1 U8120 ( .A1(n6364), .A2(n6363), .ZN(n6365) );
  XNOR2_X1 U8121 ( .A(n6365), .B(n6196), .ZN(n6368) );
  INV_X1 U8122 ( .A(n6368), .ZN(n6366) );
  AOI22_X1 U8123 ( .A1(n9575), .A2(n6397), .B1(n6392), .B2(n9458), .ZN(n6367)
         );
  NAND2_X1 U8124 ( .A1(n6366), .A2(n6367), .ZN(n6374) );
  INV_X1 U8125 ( .A(n6374), .ZN(n6369) );
  XNOR2_X1 U8126 ( .A(n6368), .B(n6367), .ZN(n8134) );
  INV_X1 U8127 ( .A(n6382), .ZN(n6376) );
  NAND2_X1 U8128 ( .A1(n9464), .A2(n6387), .ZN(n6371) );
  NAND2_X1 U8129 ( .A1(n9194), .A2(n6397), .ZN(n6370) );
  NAND2_X1 U8130 ( .A1(n6371), .A2(n6370), .ZN(n6372) );
  XNOR2_X1 U8131 ( .A(n6372), .B(n6196), .ZN(n6381) );
  INV_X1 U8132 ( .A(n6381), .ZN(n6373) );
  AOI22_X1 U8133 ( .A1(n9464), .A2(n6397), .B1(n6392), .B2(n9194), .ZN(n6380)
         );
  NAND2_X1 U8134 ( .A1(n6373), .A2(n6380), .ZN(n8132) );
  AND2_X1 U8135 ( .A1(n8132), .A2(n6374), .ZN(n6375) );
  AND2_X1 U8136 ( .A1(n6465), .A2(n6379), .ZN(n6378) );
  INV_X1 U8137 ( .A(n6379), .ZN(n6383) );
  XNOR2_X1 U8138 ( .A(n6381), .B(n6380), .ZN(n8382) );
  INV_X1 U8139 ( .A(n6384), .ZN(n6385) );
  NAND2_X1 U8140 ( .A1(n6386), .A2(n6385), .ZN(n6481) );
  AOI22_X1 U8141 ( .A1(n9564), .A2(n6387), .B1(n6397), .B2(n9427), .ZN(n6389)
         );
  XNOR2_X1 U8142 ( .A(n6389), .B(n6388), .ZN(n6405) );
  AOI22_X1 U8143 ( .A1(n9564), .A2(n6397), .B1(n6392), .B2(n9427), .ZN(n6404)
         );
  XNOR2_X1 U8144 ( .A(n6405), .B(n6404), .ZN(n6485) );
  INV_X1 U8145 ( .A(n6485), .ZN(n6390) );
  AND2_X1 U8146 ( .A1(n6481), .A2(n6390), .ZN(n6391) );
  NAND2_X1 U8147 ( .A1(n9026), .A2(n6397), .ZN(n6394) );
  NAND2_X1 U8148 ( .A1(n9193), .A2(n6392), .ZN(n6393) );
  NAND2_X1 U8149 ( .A1(n6394), .A2(n6393), .ZN(n6396) );
  XNOR2_X1 U8150 ( .A(n6396), .B(n6395), .ZN(n6399) );
  AOI22_X1 U8151 ( .A1(n9026), .A2(n6214), .B1(n6397), .B2(n9193), .ZN(n6398)
         );
  XNOR2_X1 U8152 ( .A(n6399), .B(n6398), .ZN(n6425) );
  INV_X1 U8153 ( .A(n6425), .ZN(n6403) );
  NOR2_X1 U8154 ( .A1(n6401), .A2(n6400), .ZN(n6631) );
  NOR2_X1 U8155 ( .A1(n6632), .A2(n6631), .ZN(n6402) );
  AND2_X1 U8156 ( .A1(n6402), .A2(n9941), .ZN(n6413) );
  INV_X1 U8157 ( .A(n9940), .ZN(n7037) );
  NAND2_X1 U8158 ( .A1(n6190), .A2(n6939), .ZN(n10095) );
  AND2_X1 U8159 ( .A1(n10095), .A2(n9115), .ZN(n6414) );
  NAND2_X1 U8160 ( .A1(n6403), .A2(n8917), .ZN(n6430) );
  NAND2_X1 U8161 ( .A1(n6405), .A2(n6404), .ZN(n6424) );
  NOR2_X1 U8162 ( .A1(n9940), .A2(n9988), .ZN(n6407) );
  NAND2_X1 U8163 ( .A1(n6413), .A2(n6407), .ZN(n6408) );
  NAND2_X1 U8164 ( .A1(n6408), .A2(n9994), .ZN(n8909) );
  NAND2_X1 U8165 ( .A1(n9192), .A2(n9982), .ZN(n6410) );
  NAND2_X1 U8166 ( .A1(n9427), .A2(n9985), .ZN(n6409) );
  AND2_X1 U8167 ( .A1(n6410), .A2(n6409), .ZN(n6625) );
  NOR2_X1 U8168 ( .A1(n9940), .A2(n6190), .ZN(n6411) );
  NAND2_X1 U8169 ( .A1(n6413), .A2(n6411), .ZN(n8862) );
  INV_X1 U8170 ( .A(n6412), .ZN(n9411) );
  INV_X1 U8171 ( .A(n6413), .ZN(n6420) );
  INV_X1 U8172 ( .A(n6414), .ZN(n6417) );
  OR2_X1 U8173 ( .A1(n6415), .A2(P1_U3086), .ZN(n7204) );
  NAND3_X1 U8174 ( .A1(n6417), .A2(n6416), .A3(n7204), .ZN(n6419) );
  AOI21_X1 U8175 ( .B1(n6420), .B2(n6419), .A(n6418), .ZN(n7038) );
  INV_X1 U8176 ( .A(n7395), .ZN(n6421) );
  NAND3_X1 U8177 ( .A1(n7038), .A2(n6421), .A3(n6792), .ZN(n6422) );
  AOI22_X1 U8178 ( .A1(n9411), .A2(n8924), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6423) );
  OAI21_X1 U8179 ( .B1(n6625), .B2(n8862), .A(n6423), .ZN(n6427) );
  INV_X1 U8180 ( .A(n8917), .ZN(n8912) );
  NOR3_X1 U8181 ( .A1(n6425), .A2(n8912), .A3(n6424), .ZN(n6426) );
  AOI211_X1 U8182 ( .C1(n9026), .C2(n8909), .A(n6427), .B(n6426), .ZN(n6428)
         );
  OAI211_X1 U8183 ( .C1(n6488), .C2(n6430), .A(n6429), .B(n6428), .ZN(P1_U3220) );
  OR2_X1 U8184 ( .A1(n6432), .A2(n6431), .ZN(n6434) );
  NAND2_X1 U8185 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  XNOR2_X1 U8186 ( .A(n6435), .B(n8327), .ZN(n6439) );
  XNOR2_X1 U8187 ( .A(n6440), .B(n8327), .ZN(n6616) );
  INV_X1 U8188 ( .A(n8122), .ZN(n8432) );
  OAI22_X1 U8189 ( .A1(n6616), .A2(n8832), .B1(n8432), .B2(n8796), .ZN(n6441)
         );
  INV_X1 U8190 ( .A(n6441), .ZN(n6443) );
  NAND2_X1 U8191 ( .A1(n10317), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8192 ( .A1(n6446), .A2(n6677), .ZN(n6447) );
  NAND2_X1 U8193 ( .A1(n6448), .A2(n6447), .ZN(n6452) );
  INV_X1 U8194 ( .A(n6448), .ZN(n6450) );
  NAND2_X1 U8195 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  AND2_X1 U8196 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  AND2_X2 U8197 ( .A1(n6454), .A2(n6453), .ZN(n10333) );
  MUX2_X1 U8198 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8621), .S(n10333), .Z(n6455) );
  INV_X1 U8199 ( .A(n6455), .ZN(n6458) );
  NAND2_X1 U8200 ( .A1(n10333), .A2(n10306), .ZN(n8770) );
  NAND2_X1 U8201 ( .A1(n10333), .A2(n10314), .ZN(n8747) );
  OAI22_X1 U8202 ( .A1(n8624), .A2(n8770), .B1(n8619), .B2(n8747), .ZN(n6456)
         );
  INV_X1 U8203 ( .A(n6456), .ZN(n6457) );
  NAND2_X1 U8204 ( .A1(n6458), .A2(n6457), .ZN(P2_U3484) );
  NAND2_X1 U8205 ( .A1(n6613), .A2(n8714), .ZN(n6464) );
  AOI22_X1 U8206 ( .A1(n8122), .A2(n8728), .B1(n10257), .B2(n8426), .ZN(n6460)
         );
  NAND2_X1 U8207 ( .A1(n6464), .A2(n6463), .ZN(P2_U3206) );
  NAND2_X1 U8208 ( .A1(n8383), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U8209 ( .A1(n6469), .A2(n6468), .ZN(n6471) );
  NAND2_X1 U8210 ( .A1(n6473), .A2(n6472), .ZN(n6480) );
  INV_X1 U8211 ( .A(n9430), .ZN(n9638) );
  INV_X1 U8212 ( .A(n9982), .ZN(n9551) );
  OR2_X1 U8213 ( .A1(n8862), .A2(n9551), .ZN(n8843) );
  INV_X1 U8214 ( .A(n8843), .ZN(n8919) );
  INV_X1 U8215 ( .A(n9431), .ZN(n6475) );
  INV_X1 U8216 ( .A(n8924), .ZN(n8907) );
  INV_X1 U8217 ( .A(n9985), .ZN(n9549) );
  OR2_X1 U8218 ( .A1(n8862), .A2(n9549), .ZN(n8921) );
  INV_X1 U8219 ( .A(n8921), .ZN(n8903) );
  AOI22_X1 U8220 ( .A1(n9458), .A2(n8903), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n6474) );
  OAI21_X1 U8221 ( .B1(n6475), .B2(n8907), .A(n6474), .ZN(n6476) );
  AOI21_X1 U8222 ( .B1(n8919), .B2(n9427), .A(n6476), .ZN(n6477) );
  OAI21_X1 U8223 ( .B1(n9638), .B2(n8928), .A(n6477), .ZN(n6478) );
  NAND2_X1 U8224 ( .A1(n6480), .A2(n6479), .ZN(P1_U3240) );
  AND2_X1 U8225 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  NAND2_X1 U8226 ( .A1(n6484), .A2(n6483), .ZN(n6486) );
  NAND2_X1 U8227 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  NAND2_X1 U8228 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  NAND2_X1 U8229 ( .A1(n6489), .A2(n8917), .ZN(n6495) );
  AOI22_X1 U8230 ( .A1(n8403), .A2(n8903), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6490) );
  OAI21_X1 U8231 ( .B1(n8395), .B2(n8907), .A(n6490), .ZN(n6491) );
  AOI21_X1 U8232 ( .B1(n8919), .B2(n9193), .A(n6491), .ZN(n6492) );
  INV_X1 U8233 ( .A(n6493), .ZN(n6494) );
  NAND2_X1 U8234 ( .A1(n6495), .A2(n6494), .ZN(P1_U3214) );
  NOR2_X1 U8235 ( .A1(n6731), .A2(P2_U3151), .ZN(n6496) );
  AND2_X1 U8236 ( .A1(n6496), .A2(n6787), .ZN(P2_U3893) );
  INV_X1 U8237 ( .A(n6731), .ZN(n6560) );
  OAI21_X1 U8238 ( .B1(n8354), .B2(n6560), .A(n6787), .ZN(n6558) );
  NAND2_X1 U8239 ( .A1(n6558), .A2(n6497), .ZN(n6498) );
  NAND2_X1 U8240 ( .A1(n6498), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8241 ( .A(n10202), .ZN(n7115) );
  INV_X1 U8242 ( .A(n10168), .ZN(n7007) );
  INV_X1 U8243 ( .A(n10135), .ZN(n6833) );
  OAI21_X1 U8244 ( .B1(n6760), .B2(n6500), .A(n6499), .ZN(n8533) );
  AND2_X1 U8245 ( .A1(n4645), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U8246 ( .A1(n5725), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6502) );
  OAI21_X1 U8247 ( .B1(n6830), .B2(n6501), .A(n6502), .ZN(n6816) );
  NAND2_X1 U8248 ( .A1(n8533), .A2(n8532), .ZN(n8531) );
  NAND2_X1 U8249 ( .A1(n6760), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8250 ( .A1(n8531), .A2(n6503), .ZN(n6504) );
  NAND2_X1 U8251 ( .A1(n6504), .A2(n6762), .ZN(n6879) );
  OAI21_X1 U8252 ( .B1(n6504), .B2(n6762), .A(n6879), .ZN(n10116) );
  INV_X1 U8253 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U8254 ( .A1(n6878), .A2(n6879), .ZN(n6505) );
  INV_X1 U8255 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10321) );
  MUX2_X1 U8256 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10321), .S(n6889), .Z(n6881)
         );
  NAND2_X1 U8257 ( .A1(n6505), .A2(n6881), .ZN(n6877) );
  NAND2_X1 U8258 ( .A1(n6889), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8259 ( .A1(n6877), .A2(n6506), .ZN(n6507) );
  INV_X1 U8260 ( .A(n6770), .ZN(n6997) );
  XNOR2_X1 U8261 ( .A(n6507), .B(n6997), .ZN(n6996) );
  NAND2_X1 U8262 ( .A1(n6996), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8263 ( .A1(n6507), .A2(n6770), .ZN(n6508) );
  INV_X1 U8264 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10325) );
  MUX2_X1 U8265 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10325), .S(n7081), .Z(n7075)
         );
  INV_X1 U8266 ( .A(n7283), .ZN(n6511) );
  AOI21_X1 U8267 ( .B1(n6512), .B2(n6511), .A(n6513), .ZN(n7279) );
  NAND2_X1 U8268 ( .A1(n7279), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7338) );
  INV_X1 U8269 ( .A(n6513), .ZN(n7336) );
  XNOR2_X1 U8270 ( .A(n6800), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7337) );
  XNOR2_X1 U8271 ( .A(n6514), .B(n4853), .ZN(n7411) );
  INV_X1 U8272 ( .A(n6514), .ZN(n6515) );
  NAND2_X1 U8273 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6833), .ZN(n6516) );
  OAI21_X1 U8274 ( .B1(n6833), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6516), .ZN(
        n10146) );
  NOR2_X1 U8275 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  NOR2_X1 U8276 ( .A1(n10153), .A2(n6517), .ZN(n6518) );
  MUX2_X1 U8277 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6519), .S(n10168), .Z(
        n10179) );
  AOI21_X1 U8278 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7007), .A(n10178), .ZN(
        n6520) );
  XNOR2_X1 U8279 ( .A(n10185), .B(n6520), .ZN(n10195) );
  XNOR2_X1 U8280 ( .A(n10202), .B(n9853), .ZN(n10212) );
  XNOR2_X1 U8281 ( .A(n8555), .B(n6521), .ZN(n8551) );
  NOR2_X1 U8282 ( .A1(n8555), .A2(n6521), .ZN(n6522) );
  NAND2_X1 U8283 ( .A1(n7102), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6523) );
  OAI21_X1 U8284 ( .B1(n7102), .B2(P2_REG1_REG_16__SCAN_IN), .A(n6523), .ZN(
        n8562) );
  INV_X1 U8285 ( .A(n6525), .ZN(n6524) );
  NOR2_X1 U8286 ( .A1(n10218), .A2(n6524), .ZN(n6526) );
  INV_X1 U8287 ( .A(n10218), .ZN(n7192) );
  INV_X1 U8288 ( .A(n8595), .ZN(n8585) );
  NAND2_X1 U8289 ( .A1(n8585), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6527) );
  OAI21_X1 U8290 ( .B1(n8585), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6527), .ZN(
        n8579) );
  INV_X1 U8291 ( .A(n6527), .ZN(n6528) );
  XNOR2_X1 U8292 ( .A(n8360), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6563) );
  XNOR2_X1 U8293 ( .A(n6529), .B(n6563), .ZN(n6532) );
  INV_X1 U8294 ( .A(n6530), .ZN(n8362) );
  NOR2_X1 U8295 ( .A1(n8362), .A2(P2_U3151), .ZN(n7742) );
  AND2_X1 U8296 ( .A1(n6558), .A2(n7742), .ZN(n6557) );
  INV_X2 U8297 ( .A(n6531), .ZN(n8361) );
  AND2_X1 U8298 ( .A1(n6557), .A2(n8361), .ZN(n10117) );
  NAND2_X1 U8299 ( .A1(n6532), .A2(n10117), .ZN(n6612) );
  NAND2_X1 U8300 ( .A1(n10202), .A2(n5913), .ZN(n10201) );
  INV_X1 U8301 ( .A(n10185), .ZN(n7052) );
  AOI22_X1 U8302 ( .A1(n10168), .A2(n7737), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n7007), .ZN(n10171) );
  INV_X1 U8303 ( .A(n10153), .ZN(n6868) );
  INV_X1 U8304 ( .A(n7081), .ZN(n6588) );
  INV_X1 U8305 ( .A(n6760), .ZN(n8539) );
  INV_X1 U8306 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U8307 ( .A1(n5725), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8308 ( .A1(n6830), .A2(n6537), .ZN(n6536) );
  NAND2_X1 U8309 ( .A1(n4645), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6534) );
  OR2_X1 U8310 ( .A1(n6534), .A2(n5725), .ZN(n6535) );
  NAND2_X1 U8311 ( .A1(n6536), .A2(n6535), .ZN(n6820) );
  NAND2_X1 U8312 ( .A1(n6820), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8313 ( .A1(n6538), .A2(n6537), .ZN(n8528) );
  NAND2_X1 U8314 ( .A1(n8529), .A2(n8528), .ZN(n8527) );
  OAI21_X1 U8315 ( .B1(n8539), .B2(n10259), .A(n8527), .ZN(n6539) );
  INV_X1 U8316 ( .A(n6762), .ZN(n10131) );
  XNOR2_X1 U8317 ( .A(n6539), .B(n10131), .ZN(n10115) );
  AOI22_X1 U8318 ( .A1(n10115), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n6762), .B2(
        n6539), .ZN(n6875) );
  MUX2_X1 U8319 ( .A(n7014), .B(P2_REG2_REG_4__SCAN_IN), .S(n6889), .Z(n6876)
         );
  OAI22_X1 U8320 ( .A1(n6997), .A2(n6540), .B1(n6992), .B2(n7107), .ZN(n7072)
         );
  MUX2_X1 U8321 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6541), .S(n7081), .Z(n7073)
         );
  INV_X1 U8322 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6542) );
  MUX2_X1 U8323 ( .A(n6542), .B(P2_REG2_REG_8__SCAN_IN), .S(n6800), .Z(n7329)
         );
  AOI22_X1 U8324 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6833), .B1(n10135), .B2(
        n7452), .ZN(n10140) );
  NAND2_X1 U8325 ( .A1(n6868), .A2(n6545), .ZN(n6546) );
  XNOR2_X1 U8326 ( .A(n6545), .B(n10153), .ZN(n10155) );
  NAND2_X1 U8327 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n10155), .ZN(n10154) );
  NAND2_X1 U8328 ( .A1(n6546), .A2(n10154), .ZN(n10170) );
  NAND2_X1 U8329 ( .A1(n10171), .A2(n10170), .ZN(n10169) );
  NAND2_X1 U8330 ( .A1(n7052), .A2(n6547), .ZN(n6548) );
  NOR2_X1 U8331 ( .A1(n8555), .A2(n6549), .ZN(n6550) );
  XNOR2_X1 U8332 ( .A(n8555), .B(n6549), .ZN(n8546) );
  NOR2_X1 U8333 ( .A1(n9868), .A2(n8546), .ZN(n8545) );
  NAND2_X1 U8334 ( .A1(n7102), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6551) );
  OAI21_X1 U8335 ( .B1(n7102), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6551), .ZN(
        n8569) );
  NOR2_X1 U8336 ( .A1(n10218), .A2(n6552), .ZN(n6553) );
  NOR2_X1 U8337 ( .A1(n10226), .A2(n10225), .ZN(n10224) );
  NAND2_X1 U8338 ( .A1(n8585), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6554) );
  OAI21_X1 U8339 ( .B1(n8585), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6554), .ZN(
        n8591) );
  INV_X1 U8340 ( .A(n6554), .ZN(n6555) );
  NOR2_X1 U8341 ( .A1(n8590), .A2(n6555), .ZN(n6556) );
  MUX2_X1 U8342 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8699), .S(n8360), .Z(n6565)
         );
  INV_X1 U8343 ( .A(n6557), .ZN(n6801) );
  OR2_X1 U8344 ( .A1(n6801), .A2(n8361), .ZN(n10227) );
  NOR2_X1 U8345 ( .A1(n8361), .A2(P2_U3151), .ZN(n7728) );
  AND2_X1 U8346 ( .A1(n6558), .A2(n7728), .ZN(n6559) );
  MUX2_X1 U8347 ( .A(P2_U3893), .B(n6559), .S(n8362), .Z(n10219) );
  AND2_X1 U8348 ( .A1(n6787), .A2(n6560), .ZN(n6561) );
  OR2_X1 U8349 ( .A1(P2_U3150), .A2(n6561), .ZN(n10134) );
  NAND2_X1 U8350 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n6562) );
  OAI21_X1 U8351 ( .B1(n10134), .B2(n4581), .A(n6562), .ZN(n6609) );
  INV_X1 U8352 ( .A(n6563), .ZN(n6564) );
  MUX2_X1 U8353 ( .A(n6565), .B(n6564), .S(n8361), .Z(n6607) );
  MUX2_X1 U8354 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8361), .Z(n6603) );
  XNOR2_X1 U8355 ( .A(n6603), .B(n10218), .ZN(n10223) );
  MUX2_X1 U8356 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8361), .Z(n6566) );
  OR2_X1 U8357 ( .A1(n6566), .A2(n7102), .ZN(n6602) );
  XNOR2_X1 U8358 ( .A(n6566), .B(n8566), .ZN(n8565) );
  MUX2_X1 U8359 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8361), .Z(n6568) );
  INV_X1 U8360 ( .A(n6568), .ZN(n6567) );
  NAND2_X1 U8361 ( .A1(n8555), .A2(n6567), .ZN(n6601) );
  XNOR2_X1 U8362 ( .A(n6568), .B(n8555), .ZN(n8549) );
  MUX2_X1 U8363 ( .A(n5913), .B(n9853), .S(n8361), .Z(n6569) );
  NAND2_X1 U8364 ( .A1(n10202), .A2(n6569), .ZN(n6600) );
  XNOR2_X1 U8365 ( .A(n6569), .B(n7115), .ZN(n10207) );
  MUX2_X1 U8366 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8361), .Z(n6570) );
  OR2_X1 U8367 ( .A1(n6570), .A2(n7052), .ZN(n6599) );
  XNOR2_X1 U8368 ( .A(n6570), .B(n10185), .ZN(n10190) );
  MUX2_X1 U8369 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8361), .Z(n6571) );
  OR2_X1 U8370 ( .A1(n6571), .A2(n7007), .ZN(n6598) );
  XNOR2_X1 U8371 ( .A(n6571), .B(n10168), .ZN(n10174) );
  MUX2_X1 U8372 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8361), .Z(n6572) );
  OR2_X1 U8373 ( .A1(n6572), .A2(n6868), .ZN(n6597) );
  XNOR2_X1 U8374 ( .A(n6572), .B(n10153), .ZN(n10158) );
  MUX2_X1 U8375 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8361), .Z(n6573) );
  OR2_X1 U8376 ( .A1(n6573), .A2(n6833), .ZN(n6596) );
  XNOR2_X1 U8377 ( .A(n6573), .B(n10135), .ZN(n10137) );
  MUX2_X1 U8378 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8361), .Z(n6586) );
  INV_X1 U8379 ( .A(n6586), .ZN(n6587) );
  MUX2_X1 U8380 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8361), .Z(n6584) );
  INV_X1 U8381 ( .A(n6584), .ZN(n6585) );
  INV_X1 U8382 ( .A(n6889), .ZN(n6583) );
  MUX2_X1 U8383 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8361), .Z(n6581) );
  INV_X1 U8384 ( .A(n6581), .ZN(n6582) );
  MUX2_X1 U8385 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8361), .Z(n6579) );
  INV_X1 U8386 ( .A(n6579), .ZN(n6580) );
  MUX2_X1 U8387 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8361), .Z(n6577) );
  INV_X1 U8388 ( .A(n6577), .ZN(n6578) );
  INV_X1 U8389 ( .A(n6830), .ZN(n6576) );
  MUX2_X1 U8390 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8361), .Z(n6574) );
  INV_X1 U8391 ( .A(n6574), .ZN(n6575) );
  XOR2_X1 U8392 ( .A(n6830), .B(n6574), .Z(n6827) );
  NAND2_X1 U8393 ( .A1(n6827), .A2(n6826), .ZN(n6825) );
  OAI21_X1 U8394 ( .B1(n6576), .B2(n6575), .A(n6825), .ZN(n8526) );
  XOR2_X1 U8395 ( .A(n6760), .B(n6577), .Z(n8525) );
  NAND2_X1 U8396 ( .A1(n8526), .A2(n8525), .ZN(n8524) );
  OAI21_X1 U8397 ( .B1(n8539), .B2(n6578), .A(n8524), .ZN(n10125) );
  XNOR2_X1 U8398 ( .A(n6579), .B(n6762), .ZN(n10126) );
  NOR2_X1 U8399 ( .A1(n10125), .A2(n10126), .ZN(n10124) );
  AOI21_X1 U8400 ( .B1(n10131), .B2(n6580), .A(n10124), .ZN(n6873) );
  XOR2_X1 U8401 ( .A(n6889), .B(n6581), .Z(n6872) );
  NAND2_X1 U8402 ( .A1(n6873), .A2(n6872), .ZN(n6871) );
  OAI21_X1 U8403 ( .B1(n6583), .B2(n6582), .A(n6871), .ZN(n6995) );
  XOR2_X1 U8404 ( .A(n6770), .B(n6584), .Z(n6994) );
  NAND2_X1 U8405 ( .A1(n6995), .A2(n6994), .ZN(n6993) );
  XNOR2_X1 U8406 ( .A(n6586), .B(n7081), .ZN(n7070) );
  MUX2_X1 U8407 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8361), .Z(n6589) );
  XNOR2_X1 U8408 ( .A(n6589), .B(n7283), .ZN(n7277) );
  MUX2_X1 U8409 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8361), .Z(n6590) );
  XOR2_X1 U8410 ( .A(n6800), .B(n6590), .Z(n7330) );
  INV_X1 U8411 ( .A(n6800), .ZN(n7343) );
  INV_X1 U8412 ( .A(n6590), .ZN(n6591) );
  AOI22_X1 U8413 ( .A1(n7331), .A2(n7330), .B1(n7343), .B2(n6591), .ZN(n7406)
         );
  MUX2_X1 U8414 ( .A(n7426), .B(n6592), .S(n8361), .Z(n6594) );
  XNOR2_X1 U8415 ( .A(n6594), .B(n6593), .ZN(n7407) );
  INV_X1 U8416 ( .A(n6594), .ZN(n6595) );
  OAI22_X1 U8417 ( .A1(n7406), .A2(n7407), .B1(n6595), .B2(n4853), .ZN(n10138)
         );
  NAND2_X1 U8418 ( .A1(n10137), .A2(n10138), .ZN(n10136) );
  NAND2_X1 U8419 ( .A1(n6596), .A2(n10136), .ZN(n10157) );
  NAND2_X1 U8420 ( .A1(n10158), .A2(n10157), .ZN(n10156) );
  NAND2_X1 U8421 ( .A1(n6597), .A2(n10156), .ZN(n10173) );
  NAND2_X1 U8422 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U8423 ( .A1(n6598), .A2(n10172), .ZN(n10189) );
  NAND2_X1 U8424 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  NAND2_X1 U8425 ( .A1(n6599), .A2(n10188), .ZN(n10206) );
  NAND2_X1 U8426 ( .A1(n10207), .A2(n10206), .ZN(n10205) );
  NAND2_X1 U8427 ( .A1(n6600), .A2(n10205), .ZN(n8548) );
  NAND2_X1 U8428 ( .A1(n8549), .A2(n8548), .ZN(n8547) );
  NAND2_X1 U8429 ( .A1(n6601), .A2(n8547), .ZN(n8564) );
  NAND2_X1 U8430 ( .A1(n8565), .A2(n8564), .ZN(n8563) );
  INV_X1 U8431 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8713) );
  INV_X1 U8432 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8765) );
  MUX2_X1 U8433 ( .A(n8713), .B(n8765), .S(n8361), .Z(n6604) );
  NAND2_X1 U8434 ( .A1(n6605), .A2(n6604), .ZN(n8581) );
  AOI21_X1 U8435 ( .B1(n8585), .B2(n8581), .A(n8580), .ZN(n6606) );
  XOR2_X1 U8436 ( .A(n6607), .B(n6606), .Z(n6608) );
  NAND2_X1 U8437 ( .A1(P2_U3893), .A2(n8362), .ZN(n10127) );
  NAND2_X1 U8438 ( .A1(n6612), .A2(n6611), .ZN(P2_U3201) );
  NAND2_X1 U8439 ( .A1(n6613), .A2(n10333), .ZN(n6615) );
  NAND2_X1 U8440 ( .A1(n6615), .A2(n6614), .ZN(n6618) );
  OAI22_X1 U8441 ( .A1(n6616), .A2(n8770), .B1(n8432), .B2(n8747), .ZN(n6617)
         );
  OR2_X1 U8442 ( .A1(n6618), .A2(n6617), .ZN(P2_U3486) );
  INV_X1 U8443 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6637) );
  INV_X1 U8444 ( .A(n10084), .ZN(n6621) );
  INV_X1 U8445 ( .A(n6622), .ZN(n9072) );
  XNOR2_X1 U8446 ( .A(n6623), .B(n9072), .ZN(n6624) );
  NAND2_X1 U8447 ( .A1(n6624), .A2(n9980), .ZN(n6626) );
  AOI21_X1 U8448 ( .B1(n8392), .B2(n9026), .A(n9968), .ZN(n6628) );
  NAND2_X1 U8449 ( .A1(n10084), .A2(n9132), .ZN(n6635) );
  NOR2_X1 U8450 ( .A1(n6631), .A2(n9940), .ZN(n6633) );
  NAND4_X1 U8451 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6639)
         );
  INV_X1 U8452 ( .A(n9941), .ZN(n6636) );
  INV_X2 U8453 ( .A(n10110), .ZN(n10113) );
  MUX2_X1 U8454 ( .A(n6637), .B(n6640), .S(n10113), .Z(n6638) );
  INV_X1 U8455 ( .A(n9026), .ZN(n9414) );
  INV_X1 U8456 ( .A(n10095), .ZN(n9624) );
  NAND2_X1 U8457 ( .A1(n10113), .A2(n9624), .ZN(n9616) );
  NAND2_X1 U8458 ( .A1(n6638), .A2(n4914), .ZN(P1_U3550) );
  INV_X1 U8459 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6641) );
  INV_X2 U8460 ( .A(n10099), .ZN(n10101) );
  MUX2_X1 U8461 ( .A(n6641), .B(n6640), .S(n10101), .Z(n6642) );
  NAND2_X1 U8462 ( .A1(n10101), .A2(n9624), .ZN(n9936) );
  NAND2_X1 U8463 ( .A1(n6642), .A2(n4906), .ZN(P1_U3518) );
  INV_X1 U8464 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6665) );
  INV_X1 U8465 ( .A(n6643), .ZN(n6644) );
  MUX2_X1 U8466 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6763), .Z(n6652) );
  XNOR2_X1 U8467 ( .A(n6652), .B(SI_30_), .ZN(n6653) );
  NAND2_X1 U8468 ( .A1(n8091), .A2(n6648), .ZN(n6651) );
  INV_X1 U8469 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8093) );
  OR2_X1 U8470 ( .A1(n6649), .A2(n8093), .ZN(n6650) );
  NAND2_X1 U8471 ( .A1(n9401), .A2(n9632), .ZN(n9402) );
  INV_X1 U8472 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6655) );
  INV_X1 U8473 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8144) );
  MUX2_X1 U8474 ( .A(n6655), .B(n8144), .S(n6763), .Z(n6656) );
  XNOR2_X1 U8475 ( .A(n6656), .B(SI_31_), .ZN(n6657) );
  NAND2_X1 U8476 ( .A1(n5174), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6663) );
  INV_X1 U8477 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8411) );
  OR2_X1 U8478 ( .A1(n5125), .A2(n8411), .ZN(n6662) );
  OR2_X1 U8479 ( .A1(n5340), .A2(n6665), .ZN(n6661) );
  AND3_X1 U8480 ( .A1(n6663), .A2(n6662), .A3(n6661), .ZN(n9035) );
  NOR2_X1 U8481 ( .A1(n9035), .A2(n6664), .ZN(n9555) );
  NOR2_X1 U8482 ( .A1(n8410), .A2(n9555), .ZN(n6668) );
  MUX2_X1 U8483 ( .A(n6665), .B(n6668), .S(n10101), .Z(n6667) );
  NAND2_X1 U8484 ( .A1(n6667), .A2(n6666), .ZN(P1_U3521) );
  INV_X1 U8485 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6669) );
  MUX2_X1 U8486 ( .A(n6669), .B(n6668), .S(n10113), .Z(n6671) );
  NAND2_X1 U8487 ( .A1(n6671), .A2(n6670), .ZN(P1_U3553) );
  INV_X1 U8488 ( .A(n10333), .ZN(n6673) );
  NAND2_X1 U8489 ( .A1(n6673), .A2(n9644), .ZN(n6672) );
  NAND2_X1 U8490 ( .A1(n6675), .A2(n4915), .ZN(P2_U3488) );
  OR2_X1 U8491 ( .A1(n6792), .A2(P1_U3086), .ZN(n6676) );
  OR2_X2 U8492 ( .A1(n6676), .A2(n7395), .ZN(n9210) );
  INV_X1 U8493 ( .A(n9210), .ZN(P1_U3973) );
  NAND2_X1 U8494 ( .A1(n6677), .A2(n8196), .ZN(n6679) );
  NAND2_X1 U8495 ( .A1(n6679), .A2(n6678), .ZN(n6681) );
  NAND2_X1 U8496 ( .A1(n6681), .A2(n6680), .ZN(n6683) );
  XNOR2_X1 U8497 ( .A(n10291), .B(n6685), .ZN(n7687) );
  XNOR2_X1 U8498 ( .A(n7687), .B(n8517), .ZN(n6728) );
  INV_X1 U8499 ( .A(n6688), .ZN(n6686) );
  NAND2_X1 U8500 ( .A1(n6686), .A2(n6982), .ZN(n6691) );
  NAND2_X1 U8501 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  INV_X1 U8502 ( .A(n6979), .ZN(n6864) );
  NAND2_X1 U8503 ( .A1(n7690), .A2(n6864), .ZN(n6690) );
  NAND2_X1 U8504 ( .A1(n6690), .A2(n8195), .ZN(n6916) );
  NAND2_X1 U8505 ( .A1(n6915), .A2(n6691), .ZN(n6923) );
  XNOR2_X1 U8506 ( .A(n5757), .B(n6685), .ZN(n6692) );
  XNOR2_X1 U8507 ( .A(n6692), .B(n6949), .ZN(n6924) );
  NAND2_X1 U8508 ( .A1(n6923), .A2(n6924), .ZN(n6922) );
  INV_X1 U8509 ( .A(n6692), .ZN(n6693) );
  NAND2_X1 U8510 ( .A1(n6693), .A2(n6949), .ZN(n6694) );
  NAND2_X1 U8511 ( .A1(n6922), .A2(n6694), .ZN(n6931) );
  INV_X1 U8512 ( .A(n6931), .ZN(n6697) );
  XNOR2_X1 U8513 ( .A(n6695), .B(n6698), .ZN(n6930) );
  NAND2_X1 U8514 ( .A1(n6697), .A2(n6696), .ZN(n6932) );
  INV_X1 U8515 ( .A(n6698), .ZN(n6699) );
  NAND2_X1 U8516 ( .A1(n6699), .A2(n10246), .ZN(n6700) );
  XNOR2_X1 U8517 ( .A(n7030), .B(n6685), .ZN(n6701) );
  NAND2_X1 U8518 ( .A1(n6701), .A2(n7160), .ZN(n7162) );
  INV_X1 U8519 ( .A(n6701), .ZN(n6702) );
  NAND2_X1 U8520 ( .A1(n8522), .A2(n6702), .ZN(n6703) );
  AND2_X1 U8521 ( .A1(n7162), .A2(n6703), .ZN(n7026) );
  XNOR2_X1 U8522 ( .A(n6685), .B(n10277), .ZN(n6704) );
  XNOR2_X1 U8523 ( .A(n6704), .B(n7199), .ZN(n7161) );
  INV_X1 U8524 ( .A(n6704), .ZN(n6705) );
  NAND2_X1 U8525 ( .A1(n6705), .A2(n7199), .ZN(n6706) );
  NAND2_X1 U8526 ( .A1(n7165), .A2(n6706), .ZN(n7194) );
  XNOR2_X1 U8527 ( .A(n6685), .B(n7123), .ZN(n6712) );
  XNOR2_X1 U8528 ( .A(n6707), .B(n6712), .ZN(n7193) );
  INV_X1 U8529 ( .A(n7193), .ZN(n6708) );
  INV_X1 U8530 ( .A(n8519), .ZN(n7374) );
  XNOR2_X1 U8531 ( .A(n6685), .B(n7308), .ZN(n6709) );
  NAND2_X1 U8532 ( .A1(n7374), .A2(n6709), .ZN(n7366) );
  INV_X1 U8533 ( .A(n6709), .ZN(n6710) );
  NAND2_X1 U8534 ( .A1(n6710), .A2(n8519), .ZN(n6711) );
  AND2_X1 U8535 ( .A1(n7366), .A2(n6711), .ZN(n7305) );
  INV_X1 U8536 ( .A(n6712), .ZN(n6713) );
  NAND2_X1 U8537 ( .A1(n6713), .A2(n8520), .ZN(n7302) );
  AND2_X1 U8538 ( .A1(n7305), .A2(n7302), .ZN(n6714) );
  XNOR2_X1 U8539 ( .A(n10286), .B(n6685), .ZN(n6716) );
  INV_X1 U8540 ( .A(n8518), .ZN(n6753) );
  XNOR2_X1 U8541 ( .A(n6716), .B(n6753), .ZN(n7367) );
  NAND2_X1 U8542 ( .A1(n6715), .A2(n7367), .ZN(n7369) );
  INV_X1 U8543 ( .A(n6716), .ZN(n6717) );
  NAND2_X1 U8544 ( .A1(n6717), .A2(n6753), .ZN(n6718) );
  NAND2_X1 U8545 ( .A1(n7369), .A2(n6718), .ZN(n6727) );
  NAND2_X1 U8546 ( .A1(n6750), .A2(n6719), .ZN(n6723) );
  INV_X1 U8547 ( .A(n6720), .ZN(n6721) );
  NAND2_X1 U8548 ( .A1(n6729), .A2(n6721), .ZN(n6722) );
  INV_X1 U8549 ( .A(n6727), .ZN(n6725) );
  INV_X1 U8550 ( .A(n6728), .ZN(n6724) );
  NAND2_X1 U8551 ( .A1(n6725), .A2(n6724), .ZN(n7689) );
  INV_X1 U8552 ( .A(n7689), .ZN(n6726) );
  AOI211_X1 U8553 ( .C1(n6728), .C2(n6727), .A(n8488), .B(n6726), .ZN(n6757)
         );
  NAND2_X1 U8554 ( .A1(n6729), .A2(n10314), .ZN(n6730) );
  NAND2_X1 U8555 ( .A1(n6730), .A2(n8711), .ZN(n8486) );
  INV_X1 U8556 ( .A(n8486), .ZN(n8503) );
  NOR2_X1 U8557 ( .A1(n8503), .A2(n10291), .ZN(n6756) );
  AND2_X1 U8558 ( .A1(n6732), .A2(n6731), .ZN(n6738) );
  INV_X1 U8559 ( .A(n6733), .ZN(n6736) );
  OAI21_X1 U8560 ( .B1(n6736), .B2(n6735), .A(n6734), .ZN(n6737) );
  OAI211_X1 U8561 ( .C1(n6741), .C2(n6739), .A(n6738), .B(n6737), .ZN(n6740)
         );
  NAND2_X1 U8562 ( .A1(n6740), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8563 ( .A1(n6890), .A2(n6785), .ZN(n8363) );
  OR2_X1 U8564 ( .A1(n6787), .A2(P2_U3151), .ZN(n8367) );
  OAI21_X1 U8565 ( .B1(n6741), .B2(n8363), .A(n8367), .ZN(n6742) );
  INV_X1 U8566 ( .A(n6742), .ZN(n6743) );
  NAND2_X1 U8567 ( .A1(n6744), .A2(n6743), .ZN(n8500) );
  INV_X1 U8568 ( .A(n7425), .ZN(n6745) );
  AND2_X1 U8569 ( .A1(n8500), .A2(n6745), .ZN(n6755) );
  NOR2_X1 U8570 ( .A1(n6748), .A2(n6746), .ZN(n6747) );
  NAND2_X1 U8571 ( .A1(n6750), .A2(n6747), .ZN(n8495) );
  AND2_X1 U8572 ( .A1(n6748), .A2(n6890), .ZN(n6749) );
  NAND2_X1 U8573 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7410) );
  INV_X1 U8574 ( .A(n7410), .ZN(n6751) );
  AOI21_X1 U8575 ( .B1(n8474), .B2(n8516), .A(n6751), .ZN(n6752) );
  OAI21_X1 U8576 ( .B1(n6753), .B2(n8495), .A(n6752), .ZN(n6754) );
  OR4_X1 U8577 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(P2_U3171)
         );
  AND2_X1 U8578 ( .A1(n6763), .A2(P2_U3151), .ZN(n7390) );
  INV_X2 U8579 ( .A(n7390), .ZN(n8418) );
  NOR2_X1 U8580 ( .A1(n6763), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7991) );
  INV_X2 U8581 ( .A(n7991), .ZN(n8415) );
  OAI222_X1 U8582 ( .A1(n6830), .A2(P2_U3151), .B1(n8418), .B2(n6764), .C1(
        n6758), .C2(n8415), .ZN(P2_U3294) );
  OAI222_X1 U8583 ( .A1(n6760), .A2(P2_U3151), .B1(n8418), .B2(n6771), .C1(
        n6759), .C2(n8415), .ZN(P2_U3293) );
  OAI222_X1 U8584 ( .A1(n6762), .A2(P2_U3151), .B1(n8418), .B2(n6765), .C1(
        n6761), .C2(n8415), .ZN(P2_U3292) );
  NAND2_X1 U8585 ( .A1(n6763), .A2(P1_U3086), .ZN(n8422) );
  AND2_X1 U8586 ( .A1(n4401), .A2(P1_U3086), .ZN(n7393) );
  INV_X2 U8587 ( .A(n7393), .ZN(n8420) );
  OAI222_X1 U8588 ( .A1(n8422), .A2(n4929), .B1(n8420), .B2(n6764), .C1(
        P1_U3086), .C2(n9219), .ZN(P1_U3354) );
  OAI222_X1 U8589 ( .A1(n8422), .A2(n6766), .B1(n8420), .B2(n6765), .C1(
        P1_U3086), .C2(n9227), .ZN(P1_U3352) );
  OAI222_X1 U8590 ( .A1(n8422), .A2(n6767), .B1(n8420), .B2(n6769), .C1(
        P1_U3086), .C2(n6914), .ZN(P1_U3351) );
  OAI222_X1 U8591 ( .A1(n6889), .A2(P2_U3151), .B1(n8418), .B2(n6769), .C1(
        n6768), .C2(n8415), .ZN(P2_U3291) );
  OAI222_X1 U8592 ( .A1(n6770), .A2(P2_U3151), .B1(n8418), .B2(n6772), .C1(
        n9803), .C2(n8415), .ZN(P2_U3290) );
  CLKBUF_X1 U8593 ( .A(n8422), .Z(n7801) );
  OAI222_X1 U8594 ( .A1(n7801), .A2(n9797), .B1(n8420), .B2(n6771), .C1(
        P1_U3086), .C2(n9955), .ZN(P1_U3353) );
  OAI222_X1 U8595 ( .A1(n7801), .A2(n6773), .B1(n8420), .B2(n6772), .C1(
        P1_U3086), .C2(n6958), .ZN(P1_U3350) );
  NAND2_X1 U8596 ( .A1(n6785), .A2(n6774), .ZN(n6775) );
  OAI21_X1 U8597 ( .B1(n6785), .B2(n6112), .A(n6775), .ZN(P2_U3377) );
  OAI222_X1 U8598 ( .A1(n7081), .A2(P2_U3151), .B1(n8418), .B2(n6777), .C1(
        n6776), .C2(n8415), .ZN(P2_U3289) );
  OAI222_X1 U8599 ( .A1(n7801), .A2(n6778), .B1(n8420), .B2(n6777), .C1(
        P1_U3086), .C2(n9240), .ZN(P1_U3349) );
  INV_X1 U8600 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U8601 ( .A1(n6919), .A2(P2_U3893), .ZN(n6779) );
  OAI21_X1 U8602 ( .B1(P2_U3893), .B2(n6780), .A(n6779), .ZN(P2_U3491) );
  OAI222_X1 U8603 ( .A1(n7283), .A2(P2_U3151), .B1(n8418), .B2(n6782), .C1(
        n6781), .C2(n8415), .ZN(P2_U3288) );
  INV_X1 U8604 ( .A(n6966), .ZN(n9254) );
  OAI222_X1 U8605 ( .A1(n8422), .A2(n6783), .B1(n8420), .B2(n6782), .C1(
        P1_U3086), .C2(n9254), .ZN(P1_U3348) );
  INV_X1 U8606 ( .A(n6109), .ZN(n6784) );
  NAND2_X1 U8607 ( .A1(n6785), .A2(n6784), .ZN(n6790) );
  AND2_X1 U8608 ( .A1(n6790), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8609 ( .A1(n6790), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8610 ( .A1(n6790), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8611 ( .A1(n6790), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8612 ( .A1(n6790), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8613 ( .A1(n6790), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8614 ( .A1(n6790), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8615 ( .A1(n6790), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8616 ( .A1(n6790), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8617 ( .A1(n6790), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8618 ( .A1(n6790), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8619 ( .A1(n6790), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8620 ( .A1(n6790), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8621 ( .A1(n6790), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8622 ( .A1(n6790), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8623 ( .A1(n6790), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8624 ( .A1(n6790), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8625 ( .A1(n6790), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8626 ( .A1(n6790), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8627 ( .A1(n6790), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8628 ( .A1(n6790), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  NOR2_X1 U8629 ( .A1(n6786), .A2(P2_U3151), .ZN(n6788) );
  AOI22_X1 U8630 ( .A1(n6790), .A2(n6789), .B1(n6788), .B2(n6787), .ZN(
        P2_U3376) );
  INV_X1 U8631 ( .A(n6790), .ZN(n6791) );
  INV_X1 U8632 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9786) );
  NOR2_X1 U8633 ( .A1(n6791), .A2(n9786), .ZN(P2_U3255) );
  INV_X1 U8634 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9721) );
  NOR2_X1 U8635 ( .A1(n6791), .A2(n9721), .ZN(P2_U3251) );
  INV_X1 U8636 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9706) );
  NOR2_X1 U8637 ( .A1(n6791), .A2(n9706), .ZN(P2_U3246) );
  INV_X1 U8638 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U8639 ( .A1(n6791), .A2(n9823), .ZN(P2_U3244) );
  INV_X1 U8640 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9850) );
  NOR2_X1 U8641 ( .A1(n6791), .A2(n9850), .ZN(P2_U3242) );
  INV_X1 U8642 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9696) );
  NOR2_X1 U8643 ( .A1(n6791), .A2(n9696), .ZN(P2_U3240) );
  INV_X1 U8644 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9886) );
  NOR2_X1 U8645 ( .A1(n6791), .A2(n9886), .ZN(P2_U3234) );
  INV_X1 U8646 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9846) );
  NOR2_X1 U8647 ( .A1(n6791), .A2(n9846), .ZN(P2_U3237) );
  INV_X1 U8648 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U8649 ( .A1(n6791), .A2(n9851), .ZN(P2_U3239) );
  OR2_X1 U8650 ( .A1(n7395), .A2(n6792), .ZN(n6793) );
  AND2_X1 U8651 ( .A1(n6793), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6835) );
  OR2_X1 U8652 ( .A1(n7395), .A2(n9115), .ZN(n6795) );
  NAND2_X1 U8653 ( .A1(n6795), .A2(n6794), .ZN(n6834) );
  NAND2_X1 U8654 ( .A1(n6835), .A2(n6834), .ZN(n9337) );
  INV_X1 U8655 ( .A(n9337), .ZN(n9950) );
  NOR2_X1 U8656 ( .A1(n9950), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8657 ( .A(n6796), .ZN(n6799) );
  INV_X1 U8658 ( .A(n6968), .ZN(n9267) );
  OAI222_X1 U8659 ( .A1(n7801), .A2(n6797), .B1(n8420), .B2(n6799), .C1(
        P1_U3086), .C2(n9267), .ZN(P1_U3347) );
  OAI222_X1 U8660 ( .A1(n6800), .A2(P2_U3151), .B1(n8418), .B2(n6799), .C1(
        n6798), .C2(n8415), .ZN(P2_U3287) );
  INV_X1 U8661 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U8662 ( .A1(n6801), .A2(n10127), .ZN(n6803) );
  AOI22_X1 U8663 ( .A1(n6803), .A2(n6802), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6805) );
  OAI211_X1 U8664 ( .C1(n10134), .C2(n6806), .A(n6805), .B(n6804), .ZN(
        P2_U3182) );
  NAND2_X1 U8665 ( .A1(n8073), .A2(P1_U3973), .ZN(n6807) );
  OAI21_X1 U8666 ( .B1(P1_U3973), .B2(n5738), .A(n6807), .ZN(P1_U3554) );
  INV_X1 U8667 ( .A(n9035), .ZN(n9108) );
  NAND2_X1 U8668 ( .A1(n9108), .A2(P1_U3973), .ZN(n6808) );
  OAI21_X1 U8669 ( .B1(P1_U3973), .B2(n8144), .A(n6808), .ZN(P1_U3585) );
  INV_X1 U8670 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9820) );
  INV_X1 U8671 ( .A(n9075), .ZN(n9074) );
  NAND2_X1 U8672 ( .A1(n9074), .A2(P1_U3973), .ZN(n6809) );
  OAI21_X1 U8673 ( .B1(n9820), .B2(P1_U3973), .A(n6809), .ZN(P1_U3584) );
  INV_X1 U8674 ( .A(n6810), .ZN(n6812) );
  OAI222_X1 U8675 ( .A1(n8415), .A2(n6811), .B1(n8418), .B2(n6812), .C1(n4853), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8676 ( .A(n7089), .ZN(n6973) );
  OAI222_X1 U8677 ( .A1(n7801), .A2(n6813), .B1(n8420), .B2(n6812), .C1(
        P1_U3086), .C2(n6973), .ZN(P1_U3346) );
  INV_X1 U8678 ( .A(n6814), .ZN(n6832) );
  INV_X1 U8679 ( .A(n7351), .ZN(n7355) );
  OAI222_X1 U8680 ( .A1(n8420), .A2(n6832), .B1(n7355), .B2(P1_U3086), .C1(
        n6815), .C2(n8422), .ZN(P1_U3345) );
  INV_X1 U8681 ( .A(n10219), .ZN(n8583) );
  NAND2_X1 U8682 ( .A1(n6816), .A2(n5729), .ZN(n6817) );
  NAND2_X1 U8683 ( .A1(n6818), .A2(n6817), .ZN(n6824) );
  XNOR2_X1 U8684 ( .A(n6820), .B(n6819), .ZN(n6821) );
  OAI22_X1 U8685 ( .A1(n10227), .A2(n6821), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7139), .ZN(n6823) );
  INV_X1 U8686 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10336) );
  NOR2_X1 U8687 ( .A1(n10134), .A2(n10336), .ZN(n6822) );
  AOI211_X1 U8688 ( .C1(n10117), .C2(n6824), .A(n6823), .B(n6822), .ZN(n6829)
         );
  INV_X1 U8689 ( .A(n10127), .ZN(n10237) );
  OAI211_X1 U8690 ( .C1(n6827), .C2(n6826), .A(n6825), .B(n10237), .ZN(n6828)
         );
  OAI211_X1 U8691 ( .C1(n8583), .C2(n6830), .A(n6829), .B(n6828), .ZN(P2_U3183) );
  OAI222_X1 U8692 ( .A1(P2_U3151), .A2(n6833), .B1(n8418), .B2(n6832), .C1(
        n6831), .C2(n8415), .ZN(P2_U3285) );
  INV_X1 U8693 ( .A(n6834), .ZN(n6836) );
  NAND2_X1 U8694 ( .A1(n6836), .A2(n6835), .ZN(n9948) );
  OR2_X1 U8695 ( .A1(n9948), .A2(n6899), .ZN(n9956) );
  INV_X1 U8696 ( .A(n6914), .ZN(n6842) );
  INV_X1 U8697 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6837) );
  MUX2_X1 U8698 ( .A(n6837), .B(P1_REG2_REG_4__SCAN_IN), .S(n6914), .Z(n6838)
         );
  INV_X1 U8699 ( .A(n6838), .ZN(n6908) );
  INV_X1 U8700 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6839) );
  MUX2_X1 U8701 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6839), .S(n6848), .Z(n9954)
         );
  INV_X1 U8702 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9700) );
  MUX2_X1 U8703 ( .A(n9700), .B(P1_REG2_REG_1__SCAN_IN), .S(n9219), .Z(n9217)
         );
  AND2_X1 U8704 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9216) );
  NAND2_X1 U8705 ( .A1(n9217), .A2(n9216), .ZN(n9215) );
  INV_X1 U8706 ( .A(n9219), .ZN(n9214) );
  NAND2_X1 U8707 ( .A1(n9214), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8708 ( .A1(n9215), .A2(n6840), .ZN(n9953) );
  NAND2_X1 U8709 ( .A1(n6847), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6841) );
  OAI21_X1 U8710 ( .B1(n6847), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6841), .ZN(
        n9231) );
  NOR2_X1 U8711 ( .A1(n9232), .A2(n9231), .ZN(n9230) );
  AOI21_X1 U8712 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6847), .A(n9230), .ZN(
        n6909) );
  NOR2_X1 U8713 ( .A1(n6908), .A2(n6909), .ZN(n6907) );
  INV_X1 U8714 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U8715 ( .A1(n6963), .A2(n6843), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n6958), .ZN(n6844) );
  OR2_X1 U8716 ( .A1(n5554), .A2(n5558), .ZN(n9189) );
  OR2_X1 U8717 ( .A1(n9948), .A2(n9189), .ZN(n9958) );
  AOI211_X1 U8718 ( .C1(n6845), .C2(n6844), .A(n6962), .B(n9958), .ZN(n6859)
         );
  NOR2_X2 U8719 ( .A1(n9948), .A2(n6846), .ZN(n9961) );
  INV_X1 U8720 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7255) );
  MUX2_X1 U8721 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7255), .S(n6914), .Z(n6904)
         );
  INV_X1 U8722 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10103) );
  MUX2_X1 U8723 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10103), .S(n6847), .Z(n9235)
         );
  INV_X1 U8724 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7180) );
  MUX2_X1 U8725 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7180), .S(n6848), .Z(n9962)
         );
  INV_X1 U8726 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9220) );
  MUX2_X1 U8727 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9220), .S(n9219), .Z(n6849)
         );
  INV_X1 U8728 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9945) );
  OR3_X1 U8729 ( .A1(n6849), .A2(n9945), .A3(n9218), .ZN(n9221) );
  OAI21_X1 U8730 ( .B1(n9219), .B2(n9220), .A(n9221), .ZN(n9963) );
  NAND2_X1 U8731 ( .A1(n9962), .A2(n9963), .ZN(n9960) );
  OAI21_X1 U8732 ( .B1(n7180), .B2(n9955), .A(n9960), .ZN(n9236) );
  NAND2_X1 U8733 ( .A1(n9235), .A2(n9236), .ZN(n9234) );
  OAI21_X1 U8734 ( .B1(n10103), .B2(n9227), .A(n9234), .ZN(n6850) );
  INV_X1 U8735 ( .A(n6850), .ZN(n6905) );
  NOR2_X1 U8736 ( .A1(n6904), .A2(n6905), .ZN(n6903) );
  NOR2_X1 U8737 ( .A1(n6914), .A2(n7255), .ZN(n6853) );
  INV_X1 U8738 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6851) );
  MUX2_X1 U8739 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6851), .S(n6963), .Z(n6852)
         );
  OAI21_X1 U8740 ( .B1(n6903), .B2(n6853), .A(n6852), .ZN(n6957) );
  INV_X1 U8741 ( .A(n6903), .ZN(n6856) );
  INV_X1 U8742 ( .A(n6853), .ZN(n6855) );
  MUX2_X1 U8743 ( .A(n6851), .B(P1_REG1_REG_5__SCAN_IN), .S(n6963), .Z(n6854)
         );
  NAND3_X1 U8744 ( .A1(n6856), .A2(n6855), .A3(n6854), .ZN(n6857) );
  AND3_X1 U8745 ( .A1(n9961), .A2(n6957), .A3(n6857), .ZN(n6858) );
  NOR2_X1 U8746 ( .A1(n6859), .A2(n6858), .ZN(n6862) );
  NOR2_X1 U8747 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9739), .ZN(n6860) );
  AOI21_X1 U8748 ( .B1(n9950), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6860), .ZN(
        n6861) );
  OAI211_X1 U8749 ( .C1(n6958), .C2(n9956), .A(n6862), .B(n6861), .ZN(P1_U3248) );
  NAND2_X1 U8750 ( .A1(n6919), .A2(n6864), .ZN(n8193) );
  AND2_X1 U8751 ( .A1(n8195), .A2(n8193), .ZN(n8149) );
  INV_X1 U8752 ( .A(n8149), .ZN(n6984) );
  OAI21_X1 U8753 ( .B1(n8684), .B2(n10306), .A(n6984), .ZN(n6863) );
  NAND2_X1 U8754 ( .A1(n6687), .A2(n10247), .ZN(n6891) );
  OAI211_X1 U8755 ( .C1(n10303), .C2(n6864), .A(n6863), .B(n6891), .ZN(n6952)
         );
  NAND2_X1 U8756 ( .A1(n6952), .A2(n10333), .ZN(n6865) );
  OAI21_X1 U8757 ( .B1(n10333), .B2(n5736), .A(n6865), .ZN(P2_U3459) );
  INV_X1 U8758 ( .A(n6866), .ZN(n6869) );
  OAI222_X1 U8759 ( .A1(n6868), .A2(P2_U3151), .B1(n8418), .B2(n6869), .C1(
        n6867), .C2(n8415), .ZN(P2_U3284) );
  INV_X1 U8760 ( .A(n7357), .ZN(n9281) );
  OAI222_X1 U8761 ( .A1(n8422), .A2(n6870), .B1(n8420), .B2(n6869), .C1(
        P1_U3086), .C2(n9281), .ZN(P1_U3344) );
  OAI211_X1 U8762 ( .C1(n6873), .C2(n6872), .A(n6871), .B(n10237), .ZN(n6888)
         );
  INV_X1 U8763 ( .A(n10134), .ZN(n10220) );
  AOI21_X1 U8764 ( .B1(n6876), .B2(n6875), .A(n6874), .ZN(n6885) );
  INV_X1 U8765 ( .A(n6877), .ZN(n6883) );
  INV_X1 U8766 ( .A(n6878), .ZN(n10119) );
  INV_X1 U8767 ( .A(n6879), .ZN(n6880) );
  NOR3_X1 U8768 ( .A1(n10119), .A2(n6881), .A3(n6880), .ZN(n6882) );
  OAI21_X1 U8769 ( .B1(n6883), .B2(n6882), .A(n10117), .ZN(n6884) );
  NAND2_X1 U8770 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7028) );
  OAI211_X1 U8771 ( .C1(n6885), .C2(n10227), .A(n6884), .B(n7028), .ZN(n6886)
         );
  AOI21_X1 U8772 ( .B1(n10220), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6886), .ZN(
        n6887) );
  OAI211_X1 U8773 ( .C1(n8583), .C2(n6889), .A(n6888), .B(n6887), .ZN(P2_U3186) );
  NOR3_X1 U8774 ( .A1(n8149), .A2(n6890), .A3(n10314), .ZN(n6893) );
  INV_X1 U8775 ( .A(n6891), .ZN(n6892) );
  OAI21_X1 U8776 ( .B1(n6893), .B2(n6892), .A(n8714), .ZN(n6895) );
  AOI22_X1 U8777 ( .A1(n8728), .A2(n6979), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10257), .ZN(n6894) );
  OAI211_X1 U8778 ( .C1(n8714), .C2(n6896), .A(n6895), .B(n6894), .ZN(P2_U3233) );
  XNOR2_X1 U8779 ( .A(n6898), .B(n6897), .ZN(n7041) );
  NAND3_X1 U8780 ( .A1(n7041), .A2(n6899), .A3(n5558), .ZN(n6902) );
  OAI21_X1 U8781 ( .B1(n5558), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6899), .ZN(
        n9944) );
  INV_X1 U8782 ( .A(n9189), .ZN(n6900) );
  AOI22_X1 U8783 ( .A1(n9218), .A2(n9944), .B1(n6900), .B2(n9216), .ZN(n6901)
         );
  NAND3_X1 U8784 ( .A1(n6902), .A2(P1_U3973), .A3(n6901), .ZN(n9965) );
  INV_X1 U8785 ( .A(n9961), .ZN(n9348) );
  AOI211_X1 U8786 ( .C1(n6905), .C2(n6904), .A(n6903), .B(n9348), .ZN(n6912)
         );
  AND2_X1 U8787 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7065) );
  INV_X1 U8788 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6906) );
  NOR2_X1 U8789 ( .A1(n9337), .A2(n6906), .ZN(n6911) );
  AOI211_X1 U8790 ( .C1(n6909), .C2(n6908), .A(n6907), .B(n9958), .ZN(n6910)
         );
  NOR4_X1 U8791 ( .A1(n6912), .A2(n7065), .A3(n6911), .A4(n6910), .ZN(n6913)
         );
  OAI211_X1 U8792 ( .C1(n9956), .C2(n6914), .A(n9965), .B(n6913), .ZN(P1_U3247) );
  INV_X1 U8793 ( .A(n8500), .ZN(n8444) );
  NAND2_X1 U8794 ( .A1(n8444), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6978) );
  INV_X1 U8795 ( .A(n6978), .ZN(n6929) );
  INV_X1 U8796 ( .A(n8488), .ZN(n8492) );
  NAND2_X1 U8797 ( .A1(n6917), .A2(n8492), .ZN(n6921) );
  INV_X1 U8798 ( .A(n8495), .ZN(n8482) );
  INV_X1 U8799 ( .A(n8474), .ZN(n8496) );
  OAI22_X1 U8800 ( .A1(n8496), .A2(n6949), .B1(n6684), .B2(n8503), .ZN(n6918)
         );
  AOI21_X1 U8801 ( .B1(n8482), .B2(n6919), .A(n6918), .ZN(n6920) );
  OAI211_X1 U8802 ( .C1(n6929), .C2(n7139), .A(n6921), .B(n6920), .ZN(P2_U3162) );
  OAI21_X1 U8803 ( .B1(n6924), .B2(n6923), .A(n6922), .ZN(n6925) );
  NAND2_X1 U8804 ( .A1(n6925), .A2(n8492), .ZN(n6928) );
  OAI22_X1 U8805 ( .A1(n8496), .A2(n6695), .B1(n5757), .B2(n8503), .ZN(n6926)
         );
  AOI21_X1 U8806 ( .B1(n8482), .B2(n6687), .A(n6926), .ZN(n6927) );
  OAI211_X1 U8807 ( .C1(n6929), .C2(n8537), .A(n6928), .B(n6927), .ZN(P2_U3177) );
  AOI21_X1 U8808 ( .B1(n6931), .B2(n6930), .A(n8488), .ZN(n6933) );
  NAND2_X1 U8809 ( .A1(n6933), .A2(n6932), .ZN(n6936) );
  AND2_X1 U8810 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10120) );
  OAI22_X1 U8811 ( .A1(n8496), .A2(n7160), .B1(n6949), .B2(n8495), .ZN(n6934)
         );
  AOI211_X1 U8812 ( .C1(n10265), .C2(n8486), .A(n10120), .B(n6934), .ZN(n6935)
         );
  OAI211_X1 U8813 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8444), .A(n6936), .B(
        n6935), .ZN(P2_U3158) );
  NOR2_X1 U8814 ( .A1(n7148), .A2(n9551), .ZN(n7507) );
  INV_X1 U8815 ( .A(n6937), .ZN(n8074) );
  NAND2_X1 U8816 ( .A1(n8073), .A2(n8082), .ZN(n9130) );
  AND2_X1 U8817 ( .A1(n8074), .A2(n9130), .ZN(n9050) );
  AOI21_X1 U8818 ( .B1(n9627), .B2(n10002), .A(n9050), .ZN(n6938) );
  AOI211_X1 U8819 ( .C1(n6939), .C2(n7511), .A(n7507), .B(n6938), .ZN(n6942)
         );
  NAND2_X1 U8820 ( .A1(n10110), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6940) );
  OAI21_X1 U8821 ( .B1(n6942), .B2(n10110), .A(n6940), .ZN(P1_U3522) );
  NAND2_X1 U8822 ( .A1(n10099), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6941) );
  OAI21_X1 U8823 ( .B1(n6942), .B2(n10099), .A(n6941), .ZN(P1_U3453) );
  OAI21_X1 U8824 ( .B1(n6119), .B2(n6945), .A(n6944), .ZN(n7143) );
  XNOR2_X1 U8825 ( .A(n6946), .B(n6119), .ZN(n6947) );
  OAI222_X1 U8826 ( .A1(n8710), .A2(n6949), .B1(n8719), .B2(n6948), .C1(n10252), .C2(n6947), .ZN(n7140) );
  AOI21_X1 U8827 ( .B1(n10306), .B2(n7143), .A(n7140), .ZN(n6991) );
  AOI22_X1 U8828 ( .A1(n8767), .A2(n6950), .B1(n6673), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n6951) );
  OAI21_X1 U8829 ( .B1(n6991), .B2(n6673), .A(n6951), .ZN(P2_U3460) );
  INV_X1 U8830 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8831 ( .A1(n6952), .A2(n10315), .ZN(n6953) );
  OAI21_X1 U8832 ( .B1(n6954), .B2(n10315), .A(n6953), .ZN(P2_U3390) );
  INV_X1 U8833 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U8834 ( .A1(n7089), .A2(n6955), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6973), .ZN(n6961) );
  INV_X1 U8835 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9860) );
  MUX2_X1 U8836 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9860), .S(n6968), .Z(n9275)
         );
  INV_X1 U8837 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U8838 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10105), .S(n6966), .Z(n9262)
         );
  NAND2_X1 U8839 ( .A1(n6965), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6959) );
  INV_X1 U8840 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6956) );
  MUX2_X1 U8841 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6956), .S(n6965), .Z(n9248)
         );
  OAI21_X1 U8842 ( .B1(n6851), .B2(n6958), .A(n6957), .ZN(n9249) );
  NAND2_X1 U8843 ( .A1(n9248), .A2(n9249), .ZN(n9247) );
  NAND2_X1 U8844 ( .A1(n6959), .A2(n9247), .ZN(n9263) );
  NAND2_X1 U8845 ( .A1(n9262), .A2(n9263), .ZN(n9261) );
  OAI21_X1 U8846 ( .B1(n9254), .B2(n10105), .A(n9261), .ZN(n9276) );
  NAND2_X1 U8847 ( .A1(n9275), .A2(n9276), .ZN(n9274) );
  OAI21_X1 U8848 ( .B1(n9267), .B2(n9860), .A(n9274), .ZN(n6960) );
  NOR2_X1 U8849 ( .A1(n6961), .A2(n6960), .ZN(n7091) );
  AOI21_X1 U8850 ( .B1(n6961), .B2(n6960), .A(n7091), .ZN(n6977) );
  INV_X1 U8851 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7619) );
  AOI22_X1 U8852 ( .A1(n7089), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7619), .B2(
        n6973), .ZN(n6970) );
  NAND2_X1 U8853 ( .A1(n6965), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6964) );
  OAI21_X1 U8854 ( .B1(n6965), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6964), .ZN(
        n9244) );
  INV_X1 U8855 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U8856 ( .A1(n6966), .A2(n9865), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9254), .ZN(n9258) );
  NOR2_X1 U8857 ( .A1(n9259), .A2(n9258), .ZN(n9257) );
  INV_X1 U8858 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U8859 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9267), .B1(n6968), .B2(
        n6967), .ZN(n9271) );
  OAI21_X1 U8860 ( .B1(n6970), .B2(n6969), .A(n7086), .ZN(n6971) );
  INV_X1 U8861 ( .A(n9958), .ZN(n9397) );
  NAND2_X1 U8862 ( .A1(n6971), .A2(n9397), .ZN(n6976) );
  NOR2_X1 U8863 ( .A1(n6972), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7484) );
  NOR2_X1 U8864 ( .A1(n9956), .A2(n6973), .ZN(n6974) );
  AOI211_X1 U8865 ( .C1(n9950), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7484), .B(
        n6974), .ZN(n6975) );
  OAI211_X1 U8866 ( .C1(n6977), .C2(n9348), .A(n6976), .B(n6975), .ZN(P1_U3252) );
  NAND2_X1 U8867 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n6978), .ZN(n6981) );
  NAND2_X1 U8868 ( .A1(n8486), .A2(n6979), .ZN(n6980) );
  OAI211_X1 U8869 ( .C1(n8496), .C2(n6982), .A(n6981), .B(n6980), .ZN(n6983)
         );
  AOI21_X1 U8870 ( .B1(n6984), .B2(n8492), .A(n6983), .ZN(n6985) );
  INV_X1 U8871 ( .A(n6985), .ZN(P2_U3172) );
  INV_X1 U8872 ( .A(n6986), .ZN(n7006) );
  INV_X1 U8873 ( .A(n8422), .ZN(n7996) );
  AOI22_X1 U8874 ( .A1(n7493), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7996), .ZN(n6987) );
  OAI21_X1 U8875 ( .B1(n7006), .B2(n8420), .A(n6987), .ZN(P1_U3343) );
  INV_X1 U8876 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6988) );
  OAI22_X1 U8877 ( .A1(n6684), .A2(n8796), .B1(n10315), .B2(n6988), .ZN(n6989)
         );
  INV_X1 U8878 ( .A(n6989), .ZN(n6990) );
  OAI21_X1 U8879 ( .B1(n6991), .B2(n10317), .A(n6990), .ZN(P2_U3393) );
  XNOR2_X1 U8880 ( .A(n6992), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7004) );
  OAI211_X1 U8881 ( .C1(n6995), .C2(n6994), .A(n6993), .B(n10237), .ZN(n7003)
         );
  XNOR2_X1 U8882 ( .A(n6996), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7001) );
  INV_X1 U8883 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6999) );
  NAND2_X1 U8884 ( .A1(n10219), .A2(n6997), .ZN(n6998) );
  NAND2_X1 U8885 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7158) );
  OAI211_X1 U8886 ( .C1(n6999), .C2(n10134), .A(n6998), .B(n7158), .ZN(n7000)
         );
  AOI21_X1 U8887 ( .B1(n10117), .B2(n7001), .A(n7000), .ZN(n7002) );
  OAI211_X1 U8888 ( .C1(n7004), .C2(n10227), .A(n7003), .B(n7002), .ZN(
        P2_U3187) );
  OAI222_X1 U8889 ( .A1(P2_U3151), .A2(n7007), .B1(n8418), .B2(n7006), .C1(
        n7005), .C2(n8415), .ZN(P2_U3283) );
  NOR2_X1 U8890 ( .A1(n8210), .A2(n4808), .ZN(n7011) );
  INV_X1 U8891 ( .A(n7009), .ZN(n7010) );
  AOI21_X1 U8892 ( .B1(n7011), .B2(n7008), .A(n7010), .ZN(n10272) );
  XNOR2_X1 U8893 ( .A(n7012), .B(n8210), .ZN(n7013) );
  AOI222_X1 U8894 ( .A1(n8684), .A2(n7013), .B1(n10246), .B2(n10248), .C1(
        n8521), .C2(n10247), .ZN(n10270) );
  MUX2_X1 U8895 ( .A(n7014), .B(n10270), .S(n8714), .Z(n7017) );
  INV_X1 U8896 ( .A(n7033), .ZN(n7015) );
  AOI22_X1 U8897 ( .A1(n8728), .A2(n7030), .B1(n10257), .B2(n7015), .ZN(n7016)
         );
  OAI211_X1 U8898 ( .C1(n10272), .C2(n8731), .A(n7017), .B(n7016), .ZN(
        P2_U3229) );
  OAI21_X1 U8899 ( .B1(n7018), .B2(n8150), .A(n7008), .ZN(n10266) );
  INV_X1 U8900 ( .A(n10266), .ZN(n7024) );
  INV_X1 U8901 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10114) );
  XOR2_X1 U8902 ( .A(n7019), .B(n8150), .Z(n7020) );
  AOI222_X1 U8903 ( .A1(n8684), .A2(n7020), .B1(n8522), .B2(n10247), .C1(n8523), .C2(n10248), .ZN(n10268) );
  MUX2_X1 U8904 ( .A(n10114), .B(n10268), .S(n8714), .Z(n7023) );
  INV_X1 U8905 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7021) );
  AOI22_X1 U8906 ( .A1(n8728), .A2(n10265), .B1(n10257), .B2(n7021), .ZN(n7022) );
  OAI211_X1 U8907 ( .C1(n7024), .C2(n8731), .A(n7023), .B(n7022), .ZN(P2_U3230) );
  OAI21_X1 U8908 ( .B1(n7027), .B2(n7026), .A(n7025), .ZN(n7035) );
  AOI22_X1 U8909 ( .A1(n8521), .A2(n8474), .B1(n8482), .B2(n10246), .ZN(n7032)
         );
  INV_X1 U8910 ( .A(n7028), .ZN(n7029) );
  AOI21_X1 U8911 ( .B1(n7030), .B2(n8486), .A(n7029), .ZN(n7031) );
  OAI211_X1 U8912 ( .C1(n7033), .C2(n8444), .A(n7032), .B(n7031), .ZN(n7034)
         );
  AOI21_X1 U8913 ( .B1(n7035), .B2(n8492), .A(n7034), .ZN(n7036) );
  INV_X1 U8914 ( .A(n7036), .ZN(P2_U3170) );
  NAND2_X1 U8915 ( .A1(n7038), .A2(n7037), .ZN(n7150) );
  OAI22_X1 U8916 ( .A1(n8928), .A2(n8082), .B1(n8843), .B2(n7148), .ZN(n7039)
         );
  AOI21_X1 U8917 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7150), .A(n7039), .ZN(
        n7040) );
  OAI21_X1 U8918 ( .B1(n7041), .B2(n8912), .A(n7040), .ZN(P1_U3232) );
  XOR2_X1 U8919 ( .A(n7043), .B(n7042), .Z(n7048) );
  OAI22_X1 U8920 ( .A1(n8928), .A2(n10067), .B1(n8921), .B2(n7044), .ZN(n7046)
         );
  MUX2_X1 U8921 ( .A(n8924), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n7045) );
  AOI211_X1 U8922 ( .C1(n8919), .C2(n9207), .A(n7046), .B(n7045), .ZN(n7047)
         );
  OAI21_X1 U8923 ( .B1(n7048), .B2(n8912), .A(n7047), .ZN(P1_U3218) );
  INV_X1 U8924 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9819) );
  INV_X1 U8925 ( .A(n7049), .ZN(n7051) );
  INV_X1 U8926 ( .A(n9302), .ZN(n9298) );
  OAI222_X1 U8927 ( .A1(n8422), .A2(n9819), .B1(n8420), .B2(n7051), .C1(
        P1_U3086), .C2(n9298), .ZN(P1_U3342) );
  INV_X1 U8928 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7050) );
  OAI222_X1 U8929 ( .A1(n7052), .A2(P2_U3151), .B1(n8418), .B2(n7051), .C1(
        n7050), .C2(n8415), .ZN(P2_U3282) );
  INV_X1 U8930 ( .A(n7053), .ZN(n7101) );
  AOI22_X1 U8931 ( .A1(n9350), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7996), .ZN(n7054) );
  OAI21_X1 U8932 ( .B1(n7101), .B2(n8420), .A(n7054), .ZN(P1_U3339) );
  INV_X1 U8933 ( .A(n7055), .ZN(n7058) );
  AOI22_X1 U8934 ( .A1(n8555), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n7991), .ZN(n7056) );
  OAI21_X1 U8935 ( .B1(n7058), .B2(n8418), .A(n7056), .ZN(P2_U3280) );
  AOI22_X1 U8936 ( .A1(n9328), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7996), .ZN(n7057) );
  OAI21_X1 U8937 ( .B1(n7058), .B2(n8420), .A(n7057), .ZN(P1_U3340) );
  INV_X1 U8938 ( .A(n7059), .ZN(n7608) );
  OAI211_X1 U8939 ( .C1(n7062), .C2(n7061), .A(n7060), .B(n8917), .ZN(n7067)
         );
  OAI22_X1 U8940 ( .A1(n8928), .A2(n7609), .B1(n8921), .B2(n7063), .ZN(n7064)
         );
  AOI211_X1 U8941 ( .C1(n8919), .C2(n9206), .A(n7065), .B(n7064), .ZN(n7066)
         );
  OAI211_X1 U8942 ( .C1(n8907), .C2(n7608), .A(n7067), .B(n7066), .ZN(P1_U3230) );
  AOI21_X1 U8943 ( .B1(n7070), .B2(n7069), .A(n7068), .ZN(n7085) );
  INV_X1 U8944 ( .A(n10227), .ZN(n10209) );
  OAI21_X1 U8945 ( .B1(n7073), .B2(n7072), .A(n7071), .ZN(n7083) );
  NAND2_X1 U8946 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7197) );
  INV_X1 U8947 ( .A(n7197), .ZN(n7074) );
  AOI21_X1 U8948 ( .B1(n10220), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7074), .ZN(
        n7080) );
  NOR2_X1 U8949 ( .A1(n7076), .A2(n7075), .ZN(n7077) );
  OAI21_X1 U8950 ( .B1(n7078), .B2(n7077), .A(n10117), .ZN(n7079) );
  OAI211_X1 U8951 ( .C1(n8583), .C2(n7081), .A(n7080), .B(n7079), .ZN(n7082)
         );
  AOI21_X1 U8952 ( .B1(n10209), .B2(n7083), .A(n7082), .ZN(n7084) );
  OAI21_X1 U8953 ( .B1(n7085), .B2(n10127), .A(n7084), .ZN(P2_U3188) );
  OAI21_X1 U8954 ( .B1(n7089), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7086), .ZN(
        n7088) );
  INV_X1 U8955 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7655) );
  AOI22_X1 U8956 ( .A1(n7351), .A2(n7655), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7355), .ZN(n7087) );
  NOR2_X1 U8957 ( .A1(n7087), .A2(n7088), .ZN(n7350) );
  AOI211_X1 U8958 ( .C1(n7088), .C2(n7087), .A(n7350), .B(n9958), .ZN(n7099)
         );
  NOR2_X1 U8959 ( .A1(n7089), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7090) );
  NOR2_X1 U8960 ( .A1(n7091), .A2(n7090), .ZN(n7094) );
  INV_X1 U8961 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7092) );
  MUX2_X1 U8962 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7092), .S(n7351), .Z(n7093)
         );
  NAND2_X1 U8963 ( .A1(n7093), .A2(n7094), .ZN(n7354) );
  OAI211_X1 U8964 ( .C1(n7094), .C2(n7093), .A(n9961), .B(n7354), .ZN(n7097)
         );
  NOR2_X1 U8965 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7755), .ZN(n7095) );
  AOI21_X1 U8966 ( .B1(n9950), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7095), .ZN(
        n7096) );
  OAI211_X1 U8967 ( .C1(n7355), .C2(n9956), .A(n7097), .B(n7096), .ZN(n7098)
         );
  OR2_X1 U8968 ( .A1(n7099), .A2(n7098), .ZN(P1_U3253) );
  INV_X1 U8969 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7100) );
  OAI222_X1 U8970 ( .A1(n7102), .A2(P2_U3151), .B1(n8418), .B2(n7101), .C1(
        n7100), .C2(n8415), .ZN(P2_U3279) );
  AND2_X1 U8971 ( .A1(n8213), .A2(n8221), .ZN(n8153) );
  NAND2_X1 U8972 ( .A1(n7009), .A2(n7103), .ZN(n7104) );
  XOR2_X1 U8973 ( .A(n8153), .B(n7104), .Z(n10275) );
  XNOR2_X1 U8974 ( .A(n7105), .B(n8153), .ZN(n7106) );
  AOI222_X1 U8975 ( .A1(n8684), .A2(n7106), .B1(n8520), .B2(n10247), .C1(n8522), .C2(n10248), .ZN(n10276) );
  MUX2_X1 U8976 ( .A(n7107), .B(n10276), .S(n8714), .Z(n7110) );
  INV_X1 U8977 ( .A(n7108), .ZN(n7168) );
  AOI22_X1 U8978 ( .A1(n8728), .A2(n7157), .B1(n10257), .B2(n7168), .ZN(n7109)
         );
  OAI211_X1 U8979 ( .C1(n8731), .C2(n10275), .A(n7110), .B(n7109), .ZN(
        P2_U3228) );
  INV_X1 U8980 ( .A(n7111), .ZN(n7114) );
  OAI222_X1 U8981 ( .A1(n8422), .A2(n7112), .B1(n8420), .B2(n7114), .C1(
        P1_U3086), .C2(n9316), .ZN(P1_U3341) );
  OAI222_X1 U8982 ( .A1(n7115), .A2(P2_U3151), .B1(n8418), .B2(n7114), .C1(
        n7113), .C2(n8415), .ZN(P2_U3281) );
  INV_X1 U8983 ( .A(n7116), .ZN(n7155) );
  AOI22_X1 U8984 ( .A1(n9389), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7996), .ZN(n7117) );
  OAI21_X1 U8985 ( .B1(n7155), .B2(n8420), .A(n7117), .ZN(P1_U3337) );
  INV_X1 U8986 ( .A(n7119), .ZN(n8154) );
  XNOR2_X1 U8987 ( .A(n7118), .B(n8154), .ZN(n10282) );
  XNOR2_X1 U8988 ( .A(n7120), .B(n7119), .ZN(n7121) );
  OAI222_X1 U8989 ( .A1(n8710), .A2(n7374), .B1(n8719), .B2(n7199), .C1(n7121), 
        .C2(n10252), .ZN(n10284) );
  NAND2_X1 U8990 ( .A1(n10284), .A2(n8714), .ZN(n7125) );
  OAI22_X1 U8991 ( .A1(n8714), .A2(n6541), .B1(n7196), .B2(n8711), .ZN(n7122)
         );
  AOI21_X1 U8992 ( .B1(n8728), .B2(n7123), .A(n7122), .ZN(n7124) );
  OAI211_X1 U8993 ( .C1(n10282), .C2(n8731), .A(n7125), .B(n7124), .ZN(
        P2_U3227) );
  NAND2_X1 U8994 ( .A1(n8403), .A2(P1_U3973), .ZN(n7126) );
  OAI21_X1 U8995 ( .B1(n6017), .B2(P1_U3973), .A(n7126), .ZN(P1_U3580) );
  INV_X1 U8996 ( .A(n7128), .ZN(n7132) );
  OR2_X1 U8997 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  AOI22_X1 U8998 ( .A1(n7127), .A2(n7132), .B1(n7131), .B2(n7130), .ZN(n7138)
         );
  AOI22_X1 U8999 ( .A1(n8919), .A2(n9209), .B1(n7133), .B2(n8909), .ZN(n7134)
         );
  OAI21_X1 U9000 ( .B1(n7135), .B2(n8921), .A(n7134), .ZN(n7136) );
  AOI21_X1 U9001 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7150), .A(n7136), .ZN(
        n7137) );
  OAI21_X1 U9002 ( .B1(n7138), .B2(n8912), .A(n7137), .ZN(P1_U3222) );
  INV_X1 U9003 ( .A(n8731), .ZN(n7224) );
  OAI22_X1 U9004 ( .A1(n8601), .A2(n6684), .B1(n8711), .B2(n7139), .ZN(n7142)
         );
  MUX2_X1 U9005 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7140), .S(n8714), .Z(n7141)
         );
  AOI211_X1 U9006 ( .C1(n7224), .C2(n7143), .A(n7142), .B(n7141), .ZN(n7144)
         );
  INV_X1 U9007 ( .A(n7144), .ZN(P2_U3232) );
  XOR2_X1 U9008 ( .A(n7146), .B(n7145), .Z(n7152) );
  AOI22_X1 U9009 ( .A1(n8919), .A2(n9208), .B1(n7645), .B2(n8909), .ZN(n7147)
         );
  OAI21_X1 U9010 ( .B1(n7148), .B2(n8921), .A(n7147), .ZN(n7149) );
  AOI21_X1 U9011 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7150), .A(n7149), .ZN(
        n7151) );
  OAI21_X1 U9012 ( .B1(n7152), .B2(n8912), .A(n7151), .ZN(P1_U3237) );
  INV_X1 U9013 ( .A(n7153), .ZN(n7191) );
  AOI22_X1 U9014 ( .A1(n9367), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7996), .ZN(n7154) );
  OAI21_X1 U9015 ( .B1(n7191), .B2(n8420), .A(n7154), .ZN(P1_U3338) );
  OAI222_X1 U9016 ( .A1(n8415), .A2(n7156), .B1(n8418), .B2(n7155), .C1(
        P2_U3151), .C2(n8585), .ZN(P2_U3277) );
  AOI22_X1 U9017 ( .A1(n8474), .A2(n8520), .B1(n7157), .B2(n8486), .ZN(n7159)
         );
  OAI211_X1 U9018 ( .C1(n7160), .C2(n8495), .A(n7159), .B(n7158), .ZN(n7167)
         );
  INV_X1 U9019 ( .A(n7161), .ZN(n7163) );
  NAND3_X1 U9020 ( .A1(n7025), .A2(n7163), .A3(n7162), .ZN(n7164) );
  AOI21_X1 U9021 ( .B1(n7165), .B2(n7164), .A(n8488), .ZN(n7166) );
  AOI211_X1 U9022 ( .C1(n7168), .C2(n8500), .A(n7167), .B(n7166), .ZN(n7169)
         );
  INV_X1 U9023 ( .A(n7169), .ZN(P2_U3167) );
  OR2_X1 U9024 ( .A1(n7170), .A2(n9047), .ZN(n7171) );
  NAND2_X1 U9025 ( .A1(n7172), .A2(n7171), .ZN(n7651) );
  AOI21_X1 U9026 ( .B1(n8081), .B2(n7645), .A(n9968), .ZN(n7173) );
  NAND2_X1 U9027 ( .A1(n7173), .A2(n7677), .ZN(n7647) );
  INV_X1 U9028 ( .A(n7647), .ZN(n7179) );
  XNOR2_X1 U9029 ( .A(n7174), .B(n9047), .ZN(n7178) );
  INV_X1 U9030 ( .A(n7175), .ZN(n10005) );
  NAND2_X1 U9031 ( .A1(n7651), .A2(n10005), .ZN(n7177) );
  AOI22_X1 U9032 ( .A1(n9982), .A2(n9208), .B1(n9211), .B2(n9985), .ZN(n7176)
         );
  OAI211_X1 U9033 ( .C1(n7178), .C2(n10002), .A(n7177), .B(n7176), .ZN(n7648)
         );
  AOI211_X1 U9034 ( .C1(n10084), .C2(n7651), .A(n7179), .B(n7648), .ZN(n7189)
         );
  OAI22_X1 U9035 ( .A1(n9616), .A2(n7186), .B1(n10113), .B2(n7180), .ZN(n7181)
         );
  INV_X1 U9036 ( .A(n7181), .ZN(n7182) );
  OAI21_X1 U9037 ( .B1(n7189), .B2(n10110), .A(n7182), .ZN(P1_U3524) );
  INV_X1 U9038 ( .A(n7183), .ZN(n8419) );
  OAI222_X1 U9039 ( .A1(P2_U3151), .A2(n8360), .B1(n8418), .B2(n8419), .C1(
        n7184), .C2(n8415), .ZN(P2_U3276) );
  INV_X1 U9040 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7185) );
  OAI22_X1 U9041 ( .A1(n9936), .A2(n7186), .B1(n10101), .B2(n7185), .ZN(n7187)
         );
  INV_X1 U9042 ( .A(n7187), .ZN(n7188) );
  OAI21_X1 U9043 ( .B1(n7189), .B2(n10099), .A(n7188), .ZN(P1_U3459) );
  OAI222_X1 U9044 ( .A1(n7192), .A2(P2_U3151), .B1(n8418), .B2(n7191), .C1(
        n7190), .C2(n8415), .ZN(P2_U3278) );
  AOI21_X1 U9045 ( .B1(n7194), .B2(n7193), .A(n8488), .ZN(n7195) );
  NAND2_X1 U9046 ( .A1(n7195), .A2(n7303), .ZN(n7203) );
  INV_X1 U9047 ( .A(n7196), .ZN(n7201) );
  NAND2_X1 U9048 ( .A1(n8474), .A2(n8519), .ZN(n7198) );
  OAI211_X1 U9049 ( .C1(n7199), .C2(n8495), .A(n7198), .B(n7197), .ZN(n7200)
         );
  AOI21_X1 U9050 ( .B1(n7201), .B2(n8500), .A(n7200), .ZN(n7202) );
  OAI211_X1 U9051 ( .C1(n10281), .C2(n8503), .A(n7203), .B(n7202), .ZN(
        P2_U3179) );
  NAND2_X1 U9052 ( .A1(n7227), .A2(n7393), .ZN(n7205) );
  OAI211_X1 U9053 ( .C1(n7206), .C2(n7801), .A(n7205), .B(n7204), .ZN(P1_U3335) );
  INV_X1 U9054 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U9055 ( .A1(n5744), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7208) );
  INV_X1 U9056 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9738) );
  OR2_X1 U9057 ( .A1(n5745), .A2(n9738), .ZN(n7207) );
  OAI211_X1 U9058 ( .C1(n7209), .C2(n5914), .A(n7208), .B(n7207), .ZN(n7210)
         );
  INV_X1 U9059 ( .A(n7210), .ZN(n7211) );
  AND2_X1 U9060 ( .A1(n7212), .A2(n7211), .ZN(n8186) );
  NAND2_X1 U9061 ( .A1(n8584), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7213) );
  OAI21_X1 U9062 ( .B1(n8186), .B2(n8584), .A(n7213), .ZN(P2_U3522) );
  OAI211_X1 U9063 ( .C1(n7215), .C2(n8159), .A(n7214), .B(n8684), .ZN(n7217)
         );
  AOI22_X1 U9064 ( .A1(n10248), .A2(n8520), .B1(n8518), .B2(n10247), .ZN(n7216) );
  NAND2_X1 U9065 ( .A1(n7217), .A2(n7216), .ZN(n7268) );
  INV_X1 U9066 ( .A(n7268), .ZN(n7226) );
  INV_X1 U9067 ( .A(n7219), .ZN(n7220) );
  AOI21_X1 U9068 ( .B1(n8159), .B2(n7218), .A(n7220), .ZN(n7269) );
  INV_X1 U9069 ( .A(n7221), .ZN(n7309) );
  AOI22_X1 U9070 ( .A1(n10260), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n10257), .B2(
        n7309), .ZN(n7222) );
  OAI21_X1 U9071 ( .B1(n8239), .B2(n8601), .A(n7222), .ZN(n7223) );
  AOI21_X1 U9072 ( .B1(n7269), .B2(n7224), .A(n7223), .ZN(n7225) );
  OAI21_X1 U9073 ( .B1(n10260), .B2(n7226), .A(n7225), .ZN(P2_U3226) );
  INV_X1 U9074 ( .A(n7227), .ZN(n7229) );
  OAI222_X1 U9075 ( .A1(n8359), .A2(P2_U3151), .B1(n8418), .B2(n7229), .C1(
        n7228), .C2(n8415), .ZN(P2_U3275) );
  NAND2_X1 U9076 ( .A1(n7245), .A2(n9051), .ZN(n7244) );
  NAND2_X1 U9077 ( .A1(n7244), .A2(n7230), .ZN(n7231) );
  OAI21_X1 U9078 ( .B1(n7231), .B2(n9052), .A(n7432), .ZN(n7669) );
  INV_X1 U9079 ( .A(n7669), .ZN(n7238) );
  OAI21_X1 U9080 ( .B1(n7234), .B2(n7233), .A(n7232), .ZN(n7236) );
  OAI22_X1 U9081 ( .A1(n7235), .A2(n9549), .B1(n7385), .B2(n9551), .ZN(n7262)
         );
  AOI21_X1 U9082 ( .B1(n7236), .B2(n9980), .A(n7262), .ZN(n7671) );
  INV_X1 U9083 ( .A(n7251), .ZN(n7237) );
  OAI211_X1 U9084 ( .C1(n7237), .C2(n7264), .A(n10010), .B(n7435), .ZN(n7667)
         );
  OAI211_X1 U9085 ( .C1(n9627), .C2(n7238), .A(n7671), .B(n7667), .ZN(n7242)
         );
  OAI22_X1 U9086 ( .A1(n9616), .A2(n7264), .B1(n10113), .B2(n6851), .ZN(n7239)
         );
  AOI21_X1 U9087 ( .B1(n7242), .B2(n10113), .A(n7239), .ZN(n7240) );
  INV_X1 U9088 ( .A(n7240), .ZN(P1_U3527) );
  INV_X1 U9089 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9809) );
  OAI22_X1 U9090 ( .A1(n9936), .A2(n7264), .B1(n10101), .B2(n9809), .ZN(n7241)
         );
  AOI21_X1 U9091 ( .B1(n7242), .B2(n10101), .A(n7241), .ZN(n7243) );
  INV_X1 U9092 ( .A(n7243), .ZN(P1_U3468) );
  OAI21_X1 U9093 ( .B1(n7245), .B2(n9051), .A(n7244), .ZN(n7246) );
  INV_X1 U9094 ( .A(n7246), .ZN(n7614) );
  OAI21_X1 U9095 ( .B1(n7249), .B2(n7247), .A(n7248), .ZN(n7250) );
  AOI222_X1 U9096 ( .A1(n9980), .A2(n7250), .B1(n9208), .B2(n9985), .C1(n9206), 
        .C2(n9982), .ZN(n7606) );
  OAI211_X1 U9097 ( .C1(n7678), .C2(n7609), .A(n7251), .B(n10010), .ZN(n7607)
         );
  OAI211_X1 U9098 ( .C1(n9627), .C2(n7614), .A(n7606), .B(n7607), .ZN(n7257)
         );
  INV_X1 U9099 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7252) );
  OAI22_X1 U9100 ( .A1(n9936), .A2(n7609), .B1(n10101), .B2(n7252), .ZN(n7253)
         );
  AOI21_X1 U9101 ( .B1(n7257), .B2(n10101), .A(n7253), .ZN(n7254) );
  INV_X1 U9102 ( .A(n7254), .ZN(P1_U3465) );
  OAI22_X1 U9103 ( .A1(n9616), .A2(n7609), .B1(n10113), .B2(n7255), .ZN(n7256)
         );
  AOI21_X1 U9104 ( .B1(n7257), .B2(n10113), .A(n7256), .ZN(n7258) );
  INV_X1 U9105 ( .A(n7258), .ZN(P1_U3526) );
  NAND2_X1 U9106 ( .A1(n4465), .A2(n7259), .ZN(n7261) );
  XNOR2_X1 U9107 ( .A(n7261), .B(n7260), .ZN(n7267) );
  INV_X1 U9108 ( .A(n8862), .ZN(n7294) );
  AOI22_X1 U9109 ( .A1(n7262), .A2(n7294), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n7263) );
  OAI21_X1 U9110 ( .B1(n7264), .B2(n8928), .A(n7263), .ZN(n7265) );
  AOI21_X1 U9111 ( .B1(n7663), .B2(n8924), .A(n7265), .ZN(n7266) );
  OAI21_X1 U9112 ( .B1(n7267), .B2(n8912), .A(n7266), .ZN(P1_U3227) );
  AOI21_X1 U9113 ( .B1(n7269), .B2(n10306), .A(n7268), .ZN(n7274) );
  AOI22_X1 U9114 ( .A1(n8767), .A2(n7308), .B1(n6673), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7270) );
  OAI21_X1 U9115 ( .B1(n7274), .B2(n6673), .A(n7270), .ZN(P2_U3466) );
  INV_X1 U9116 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7271) );
  OAI22_X1 U9117 ( .A1(n8239), .A2(n8796), .B1(n10315), .B2(n7271), .ZN(n7272)
         );
  INV_X1 U9118 ( .A(n7272), .ZN(n7273) );
  OAI21_X1 U9119 ( .B1(n7274), .B2(n10317), .A(n7273), .ZN(P2_U3411) );
  INV_X1 U9120 ( .A(n7275), .ZN(n7301) );
  OAI222_X1 U9121 ( .A1(n8420), .A2(n7301), .B1(P1_U3086), .B2(n9132), .C1(
        n9902), .C2(n7801), .ZN(P1_U3334) );
  XOR2_X1 U9122 ( .A(n7277), .B(n7276), .Z(n7287) );
  XNOR2_X1 U9123 ( .A(n7278), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7285) );
  OAI21_X1 U9124 ( .B1(n7279), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7338), .ZN(
        n7280) );
  NAND2_X1 U9125 ( .A1(n7280), .A2(n10117), .ZN(n7282) );
  AND2_X1 U9126 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7307) );
  AOI21_X1 U9127 ( .B1(n10220), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7307), .ZN(
        n7281) );
  OAI211_X1 U9128 ( .C1(n8583), .C2(n7283), .A(n7282), .B(n7281), .ZN(n7284)
         );
  AOI21_X1 U9129 ( .B1(n10209), .B2(n7285), .A(n7284), .ZN(n7286) );
  OAI21_X1 U9130 ( .B1(n7287), .B2(n10127), .A(n7286), .ZN(P2_U3189) );
  INV_X1 U9131 ( .A(n7289), .ZN(n7290) );
  NOR2_X1 U9132 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  XNOR2_X1 U9133 ( .A(n7288), .B(n7292), .ZN(n7299) );
  INV_X1 U9134 ( .A(n10018), .ZN(n7296) );
  OAI22_X1 U9135 ( .A1(n7293), .A2(n9549), .B1(n7589), .B2(n9551), .ZN(n7438)
         );
  AOI22_X1 U9136 ( .A1(n7438), .A2(n7294), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7295) );
  OAI21_X1 U9137 ( .B1(n7296), .B2(n8907), .A(n7295), .ZN(n7297) );
  AOI21_X1 U9138 ( .B1(n7436), .B2(n8909), .A(n7297), .ZN(n7298) );
  OAI21_X1 U9139 ( .B1(n7299), .B2(n8912), .A(n7298), .ZN(P1_U3239) );
  OAI222_X1 U9140 ( .A1(n8196), .A2(P2_U3151), .B1(n8418), .B2(n7301), .C1(
        n7300), .C2(n8415), .ZN(P2_U3274) );
  AND2_X1 U9141 ( .A1(n7303), .A2(n7302), .ZN(n7306) );
  OAI21_X1 U9142 ( .B1(n7306), .B2(n7305), .A(n7304), .ZN(n7315) );
  AOI21_X1 U9143 ( .B1(n8482), .B2(n8520), .A(n7307), .ZN(n7313) );
  NAND2_X1 U9144 ( .A1(n8486), .A2(n7308), .ZN(n7312) );
  NAND2_X1 U9145 ( .A1(n8500), .A2(n7309), .ZN(n7311) );
  NAND2_X1 U9146 ( .A1(n8474), .A2(n8518), .ZN(n7310) );
  NAND4_X1 U9147 ( .A1(n7313), .A2(n7312), .A3(n7311), .A4(n7310), .ZN(n7314)
         );
  AOI21_X1 U9148 ( .B1(n7315), .B2(n8492), .A(n7314), .ZN(n7316) );
  INV_X1 U9149 ( .A(n7316), .ZN(P2_U3153) );
  NAND2_X1 U9150 ( .A1(n7219), .A2(n7317), .ZN(n7318) );
  XNOR2_X1 U9151 ( .A(n7318), .B(n8157), .ZN(n10289) );
  INV_X1 U9152 ( .A(n10289), .ZN(n7326) );
  OAI211_X1 U9153 ( .C1(n7320), .C2(n8157), .A(n7319), .B(n8684), .ZN(n7322)
         );
  AOI22_X1 U9154 ( .A1(n8517), .A2(n10247), .B1(n10248), .B2(n8519), .ZN(n7321) );
  NAND2_X1 U9155 ( .A1(n7322), .A2(n7321), .ZN(n10287) );
  AOI22_X1 U9156 ( .A1(n10260), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10257), .B2(
        n7376), .ZN(n7323) );
  OAI21_X1 U9157 ( .B1(n10286), .B2(n8601), .A(n7323), .ZN(n7324) );
  AOI21_X1 U9158 ( .B1(n10287), .B2(n8714), .A(n7324), .ZN(n7325) );
  OAI21_X1 U9159 ( .B1(n7326), .B2(n8731), .A(n7325), .ZN(P2_U3225) );
  AOI21_X1 U9160 ( .B1(n7329), .B2(n7328), .A(n7327), .ZN(n7346) );
  XNOR2_X1 U9161 ( .A(n7331), .B(n7330), .ZN(n7332) );
  NAND2_X1 U9162 ( .A1(n7332), .A2(n10237), .ZN(n7345) );
  INV_X1 U9163 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7334) );
  NOR2_X1 U9164 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9838), .ZN(n7372) );
  INV_X1 U9165 ( .A(n7372), .ZN(n7333) );
  OAI21_X1 U9166 ( .B1(n10134), .B2(n7334), .A(n7333), .ZN(n7342) );
  INV_X1 U9167 ( .A(n7335), .ZN(n7340) );
  NAND3_X1 U9168 ( .A1(n7338), .A2(n7337), .A3(n7336), .ZN(n7339) );
  INV_X1 U9169 ( .A(n10117), .ZN(n10232) );
  AOI21_X1 U9170 ( .B1(n7340), .B2(n7339), .A(n10232), .ZN(n7341) );
  AOI211_X1 U9171 ( .C1(n10219), .C2(n7343), .A(n7342), .B(n7341), .ZN(n7344)
         );
  OAI211_X1 U9172 ( .C1(n7346), .C2(n10227), .A(n7345), .B(n7344), .ZN(
        P2_U3190) );
  INV_X1 U9173 ( .A(n7347), .ZN(n8089) );
  OAI222_X1 U9174 ( .A1(P2_U3151), .A2(n7349), .B1(n8418), .B2(n8089), .C1(
        n7348), .C2(n8415), .ZN(P2_U3273) );
  INV_X1 U9175 ( .A(n7493), .ZN(n7496) );
  XNOR2_X1 U9176 ( .A(n7496), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7491) );
  INV_X1 U9177 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7352) );
  AOI22_X1 U9178 ( .A1(n7357), .A2(n7352), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9281), .ZN(n9288) );
  XNOR2_X1 U9179 ( .A(n7491), .B(n7490), .ZN(n7363) );
  INV_X1 U9180 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7353) );
  MUX2_X1 U9181 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7353), .S(n7357), .Z(n9285)
         );
  OAI21_X1 U9182 ( .B1(n7355), .B2(n7092), .A(n7354), .ZN(n9286) );
  NAND2_X1 U9183 ( .A1(n9285), .A2(n9286), .ZN(n9284) );
  INV_X1 U9184 ( .A(n9284), .ZN(n7356) );
  AOI21_X1 U9185 ( .B1(n7357), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7356), .ZN(
        n7361) );
  OR2_X1 U9186 ( .A1(n7493), .A2(n10108), .ZN(n7359) );
  INV_X1 U9187 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U9188 ( .A1(n7493), .A2(n10108), .ZN(n7358) );
  NAND2_X1 U9189 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  NAND2_X1 U9190 ( .A1(n7361), .A2(n7360), .ZN(n7499) );
  OAI21_X1 U9191 ( .B1(n7361), .B2(n7360), .A(n7499), .ZN(n7362) );
  AOI22_X1 U9192 ( .A1(n9397), .A2(n7363), .B1(n9961), .B2(n7362), .ZN(n7365)
         );
  NOR2_X1 U9193 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5292), .ZN(n7782) );
  AOI21_X1 U9194 ( .B1(n9950), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7782), .ZN(
        n7364) );
  OAI211_X1 U9195 ( .C1(n7496), .C2(n9956), .A(n7365), .B(n7364), .ZN(P1_U3255) );
  INV_X1 U9196 ( .A(n7304), .ZN(n7368) );
  NOR3_X1 U9197 ( .A1(n7368), .A2(n4670), .A3(n7367), .ZN(n7371) );
  INV_X1 U9198 ( .A(n7369), .ZN(n7370) );
  OAI21_X1 U9199 ( .B1(n7371), .B2(n7370), .A(n8492), .ZN(n7378) );
  AOI21_X1 U9200 ( .B1(n8517), .B2(n8474), .A(n7372), .ZN(n7373) );
  OAI21_X1 U9201 ( .B1(n7374), .B2(n8495), .A(n7373), .ZN(n7375) );
  AOI21_X1 U9202 ( .B1(n7376), .B2(n8500), .A(n7375), .ZN(n7377) );
  OAI211_X1 U9203 ( .C1(n10286), .C2(n8503), .A(n7378), .B(n7377), .ZN(
        P2_U3161) );
  INV_X1 U9204 ( .A(n7379), .ZN(n7381) );
  NOR2_X1 U9205 ( .A1(n7381), .A2(n7380), .ZN(n7382) );
  XNOR2_X1 U9206 ( .A(n7383), .B(n7382), .ZN(n7384) );
  NAND2_X1 U9207 ( .A1(n7384), .A2(n8917), .ZN(n7389) );
  NOR2_X1 U9208 ( .A1(n8921), .A2(n7385), .ZN(n7387) );
  OAI22_X1 U9209 ( .A1(n8843), .A2(n7572), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9253), .ZN(n7386) );
  AOI211_X1 U9210 ( .C1(n8924), .C2(n7638), .A(n7387), .B(n7386), .ZN(n7388)
         );
  OAI211_X1 U9211 ( .C1(n10073), .C2(n8928), .A(n7389), .B(n7388), .ZN(
        P1_U3213) );
  NAND2_X1 U9212 ( .A1(n7394), .A2(n7390), .ZN(n7391) );
  OAI211_X1 U9213 ( .C1(n7392), .C2(n8415), .A(n7391), .B(n8367), .ZN(P2_U3272) );
  NAND2_X1 U9214 ( .A1(n7394), .A2(n7393), .ZN(n7396) );
  NAND2_X1 U9215 ( .A1(n7395), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9191) );
  OAI211_X1 U9216 ( .C1(n9710), .C2(n8422), .A(n7396), .B(n9191), .ZN(P1_U3332) );
  OAI211_X1 U9217 ( .C1(n7399), .C2(n7398), .A(n7397), .B(n8917), .ZN(n7405)
         );
  NAND2_X1 U9218 ( .A1(n8924), .A2(n7598), .ZN(n7402) );
  OAI22_X1 U9219 ( .A1(n8843), .A2(n7590), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5207), .ZN(n7400) );
  INV_X1 U9220 ( .A(n7400), .ZN(n7401) );
  OAI211_X1 U9221 ( .C1(n7589), .C2(n8921), .A(n7402), .B(n7401), .ZN(n7403)
         );
  AOI21_X1 U9222 ( .B1(n7585), .B2(n8909), .A(n7403), .ZN(n7404) );
  NAND2_X1 U9223 ( .A1(n7405), .A2(n7404), .ZN(P1_U3221) );
  XOR2_X1 U9224 ( .A(n7407), .B(n7406), .Z(n7417) );
  XNOR2_X1 U9225 ( .A(n7408), .B(n7426), .ZN(n7415) );
  NAND2_X1 U9226 ( .A1(n10220), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7409) );
  OAI211_X1 U9227 ( .C1(n8583), .C2(n4853), .A(n7410), .B(n7409), .ZN(n7414)
         );
  XNOR2_X1 U9228 ( .A(n7411), .B(n6592), .ZN(n7412) );
  NOR2_X1 U9229 ( .A1(n7412), .A2(n10232), .ZN(n7413) );
  AOI211_X1 U9230 ( .C1(n10209), .C2(n7415), .A(n7414), .B(n7413), .ZN(n7416)
         );
  OAI21_X1 U9231 ( .B1(n7417), .B2(n10127), .A(n7416), .ZN(P2_U3191) );
  XNOR2_X1 U9232 ( .A(n7418), .B(n7421), .ZN(n10293) );
  INV_X1 U9233 ( .A(n10255), .ZN(n7419) );
  NAND2_X1 U9234 ( .A1(n8714), .A2(n7419), .ZN(n8100) );
  INV_X1 U9235 ( .A(n7421), .ZN(n8155) );
  XNOR2_X1 U9236 ( .A(n7420), .B(n8155), .ZN(n7422) );
  NAND2_X1 U9237 ( .A1(n7422), .A2(n8684), .ZN(n7424) );
  AOI22_X1 U9238 ( .A1(n10248), .A2(n8518), .B1(n8516), .B2(n10247), .ZN(n7423) );
  OAI211_X1 U9239 ( .C1(n10293), .C2(n10244), .A(n7424), .B(n7423), .ZN(n10295) );
  NAND2_X1 U9240 ( .A1(n10295), .A2(n8714), .ZN(n7430) );
  OAI22_X1 U9241 ( .A1(n8714), .A2(n7426), .B1(n7425), .B2(n8711), .ZN(n7427)
         );
  AOI21_X1 U9242 ( .B1(n8728), .B2(n7428), .A(n7427), .ZN(n7429) );
  OAI211_X1 U9243 ( .C1(n10293), .C2(n8100), .A(n7430), .B(n7429), .ZN(
        P2_U3224) );
  NAND2_X1 U9244 ( .A1(n7432), .A2(n7431), .ZN(n7434) );
  NAND2_X1 U9245 ( .A1(n7434), .A2(n7437), .ZN(n7433) );
  OAI21_X1 U9246 ( .B1(n7434), .B2(n7437), .A(n7433), .ZN(n10026) );
  AOI211_X1 U9247 ( .C1(n7436), .C2(n7435), .A(n9968), .B(n7637), .ZN(n10016)
         );
  XOR2_X1 U9248 ( .A(n7437), .B(n7566), .Z(n7439) );
  AOI21_X1 U9249 ( .B1(n7439), .B2(n9980), .A(n7438), .ZN(n10028) );
  INV_X1 U9250 ( .A(n10028), .ZN(n7440) );
  AOI211_X1 U9251 ( .C1(n6629), .C2(n10026), .A(n10016), .B(n7440), .ZN(n7446)
         );
  OAI22_X1 U9252 ( .A1(n9616), .A2(n10023), .B1(n10113), .B2(n6956), .ZN(n7441) );
  INV_X1 U9253 ( .A(n7441), .ZN(n7442) );
  OAI21_X1 U9254 ( .B1(n7446), .B2(n10110), .A(n7442), .ZN(P1_U3528) );
  INV_X1 U9255 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7443) );
  OAI22_X1 U9256 ( .A1(n9936), .A2(n10023), .B1(n10101), .B2(n7443), .ZN(n7444) );
  INV_X1 U9257 ( .A(n7444), .ZN(n7445) );
  OAI21_X1 U9258 ( .B1(n7446), .B2(n10099), .A(n7445), .ZN(P1_U3471) );
  INV_X1 U9259 ( .A(n8243), .ZN(n7447) );
  OR2_X1 U9260 ( .A1(n8235), .A2(n7447), .ZN(n8158) );
  XOR2_X1 U9261 ( .A(n7448), .B(n8158), .Z(n10298) );
  XNOR2_X1 U9262 ( .A(n7449), .B(n8158), .ZN(n7450) );
  OAI222_X1 U9263 ( .A1(n8710), .A2(n7827), .B1(n8719), .B2(n7451), .C1(n7450), 
        .C2(n10252), .ZN(n10300) );
  NAND2_X1 U9264 ( .A1(n10300), .A2(n8714), .ZN(n7455) );
  OAI22_X1 U9265 ( .A1(n8714), .A2(n7452), .B1(n7715), .B2(n8711), .ZN(n7453)
         );
  AOI21_X1 U9266 ( .B1(n8728), .B2(n7714), .A(n7453), .ZN(n7454) );
  OAI211_X1 U9267 ( .C1(n10298), .C2(n8731), .A(n7455), .B(n7454), .ZN(
        P2_U3223) );
  NAND2_X1 U9268 ( .A1(n7457), .A2(n7456), .ZN(n9997) );
  OAI21_X1 U9269 ( .B1(n7457), .B2(n7456), .A(n9997), .ZN(n7653) );
  AOI211_X1 U9270 ( .C1(n7759), .C2(n4566), .A(n9968), .B(n4420), .ZN(n7658)
         );
  OAI21_X1 U9271 ( .B1(n9054), .B2(n7459), .A(n7458), .ZN(n7460) );
  NAND2_X1 U9272 ( .A1(n7460), .A2(n9980), .ZN(n7463) );
  NAND2_X1 U9273 ( .A1(n9202), .A2(n9985), .ZN(n7462) );
  NAND2_X1 U9274 ( .A1(n9200), .A2(n9982), .ZN(n7461) );
  AND2_X1 U9275 ( .A1(n7462), .A2(n7461), .ZN(n7756) );
  NAND2_X1 U9276 ( .A1(n7463), .A2(n7756), .ZN(n7659) );
  AOI211_X1 U9277 ( .C1(n7653), .C2(n6629), .A(n7658), .B(n7659), .ZN(n7467)
         );
  INV_X1 U9278 ( .A(n9936), .ZN(n7464) );
  AOI22_X1 U9279 ( .A1(n7759), .A2(n7464), .B1(n10099), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n7465) );
  OAI21_X1 U9280 ( .B1(n7467), .B2(n10099), .A(n7465), .ZN(P1_U3483) );
  INV_X1 U9281 ( .A(n9616), .ZN(n7578) );
  AOI22_X1 U9282 ( .A1(n7759), .A2(n7578), .B1(n10110), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7466) );
  OAI21_X1 U9283 ( .B1(n7467), .B2(n10110), .A(n7466), .ZN(P1_U3532) );
  INV_X1 U9284 ( .A(n7468), .ZN(n8417) );
  OAI222_X1 U9285 ( .A1(n8420), .A2(n8417), .B1(n7470), .B2(P1_U3086), .C1(
        n7469), .C2(n7801), .ZN(P1_U3331) );
  AOI21_X1 U9286 ( .B1(n7471), .B2(n8162), .A(n10252), .ZN(n7473) );
  OAI22_X1 U9287 ( .A1(n8252), .A2(n8710), .B1(n7770), .B2(n8719), .ZN(n7472)
         );
  AOI21_X1 U9288 ( .B1(n7473), .B2(n4455), .A(n7472), .ZN(n10302) );
  NAND2_X1 U9289 ( .A1(n7474), .A2(n8243), .ZN(n7475) );
  XNOR2_X1 U9290 ( .A(n7475), .B(n8162), .ZN(n10307) );
  INV_X1 U9291 ( .A(n7476), .ZN(n10304) );
  INV_X1 U9292 ( .A(n7477), .ZN(n7772) );
  AOI22_X1 U9293 ( .A1(n10260), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10257), 
        .B2(n7772), .ZN(n7478) );
  OAI21_X1 U9294 ( .B1(n10304), .B2(n8601), .A(n7478), .ZN(n7479) );
  AOI21_X1 U9295 ( .B1(n10307), .B2(n7224), .A(n7479), .ZN(n7480) );
  OAI21_X1 U9296 ( .B1(n10302), .B2(n10260), .A(n7480), .ZN(P2_U3222) );
  OAI211_X1 U9297 ( .C1(n7483), .C2(n7482), .A(n7481), .B(n8917), .ZN(n7488)
         );
  AOI21_X1 U9298 ( .B1(n8919), .B2(n9201), .A(n7484), .ZN(n7485) );
  OAI21_X1 U9299 ( .B1(n7572), .B2(n8921), .A(n7485), .ZN(n7486) );
  AOI21_X1 U9300 ( .B1(n7617), .B2(n8924), .A(n7486), .ZN(n7487) );
  OAI211_X1 U9301 ( .C1(n4568), .C2(n8928), .A(n7488), .B(n7487), .ZN(P1_U3231) );
  INV_X1 U9302 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7489) );
  AOI22_X1 U9303 ( .A1(n9302), .A2(n7489), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9298), .ZN(n7495) );
  OAI21_X1 U9304 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7493), .A(n7492), .ZN(
        n7494) );
  AOI211_X1 U9305 ( .C1(n7495), .C2(n7494), .A(n9301), .B(n9958), .ZN(n7503)
         );
  INV_X1 U9306 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10111) );
  XNOR2_X1 U9307 ( .A(n9302), .B(n10111), .ZN(n7497) );
  NAND2_X1 U9308 ( .A1(n7496), .A2(n10108), .ZN(n7498) );
  NAND3_X1 U9309 ( .A1(n7499), .A2(n7497), .A3(n7498), .ZN(n9297) );
  INV_X1 U9310 ( .A(n9297), .ZN(n7501) );
  AOI21_X1 U9311 ( .B1(n7499), .B2(n7498), .A(n7497), .ZN(n7500) );
  NOR3_X1 U9312 ( .A1(n9348), .A2(n7501), .A3(n7500), .ZN(n7502) );
  NOR2_X1 U9313 ( .A1(n7503), .A2(n7502), .ZN(n7506) );
  NAND2_X1 U9314 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7861) );
  INV_X1 U9315 ( .A(n7861), .ZN(n7504) );
  AOI21_X1 U9316 ( .B1(n9950), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7504), .ZN(
        n7505) );
  OAI211_X1 U9317 ( .C1(n9298), .C2(n9956), .A(n7506), .B(n7505), .ZN(P1_U3256) );
  AOI21_X1 U9318 ( .B1(n10017), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7507), .ZN(
        n7508) );
  OAI21_X1 U9319 ( .B1(n9050), .B2(n7509), .A(n7508), .ZN(n7510) );
  NAND2_X1 U9320 ( .A1(n7510), .A2(n9989), .ZN(n7514) );
  INV_X1 U9321 ( .A(n10022), .ZN(n10007) );
  OAI21_X1 U9322 ( .B1(n7512), .B2(n10007), .A(n7511), .ZN(n7513) );
  OAI211_X1 U9323 ( .C1(n5124), .C2(n9989), .A(n7514), .B(n7513), .ZN(P1_U3293) );
  INV_X1 U9324 ( .A(n7515), .ZN(n7517) );
  OAI222_X1 U9325 ( .A1(n8420), .A2(n7517), .B1(n7516), .B2(P1_U3086), .C1(
        n9794), .C2(n8422), .ZN(P1_U3330) );
  OAI222_X1 U9326 ( .A1(n7518), .A2(P2_U3151), .B1(n8418), .B2(n7517), .C1(
        n9822), .C2(n8415), .ZN(P2_U3270) );
  NOR2_X1 U9327 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7555) );
  NOR2_X1 U9328 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n7553) );
  INV_X1 U9329 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7550) );
  INV_X1 U9330 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8553) );
  NOR2_X1 U9331 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7548) );
  NOR2_X1 U9332 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7546) );
  NOR2_X1 U9333 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7544) );
  NOR2_X1 U9334 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7542) );
  NOR2_X1 U9335 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7540) );
  NOR2_X1 U9336 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n7537) );
  NOR2_X1 U9337 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7534) );
  NOR2_X1 U9338 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7532) );
  NOR2_X1 U9339 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7530) );
  NOR2_X1 U9340 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7528) );
  NOR2_X1 U9341 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7526) );
  NAND2_X1 U9342 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7524) );
  INV_X1 U9343 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10133) );
  INV_X1 U9344 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9732) );
  AOI22_X1 U9345 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n10133), .B2(n9732), .ZN(n10370) );
  NAND2_X1 U9346 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7522) );
  AOI21_X1 U9347 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10334) );
  INV_X1 U9348 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U9349 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7519) );
  NOR2_X1 U9350 ( .A1(n9212), .A2(n7519), .ZN(n10335) );
  NOR2_X1 U9351 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10335), .ZN(n7520) );
  NOR2_X1 U9352 ( .A1(n10334), .A2(n7520), .ZN(n10368) );
  INV_X1 U9353 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8540) );
  INV_X1 U9354 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9867) );
  AOI22_X1 U9355 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n8540), .B2(n9867), .ZN(n10367) );
  NAND2_X1 U9356 ( .A1(n10368), .A2(n10367), .ZN(n7521) );
  NAND2_X1 U9357 ( .A1(n7522), .A2(n7521), .ZN(n10369) );
  NAND2_X1 U9358 ( .A1(n10370), .A2(n10369), .ZN(n7523) );
  NAND2_X1 U9359 ( .A1(n7524), .A2(n7523), .ZN(n10372) );
  XNOR2_X1 U9360 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10371) );
  NOR2_X1 U9361 ( .A1(n10372), .A2(n10371), .ZN(n7525) );
  NOR2_X1 U9362 ( .A1(n7526), .A2(n7525), .ZN(n10360) );
  XNOR2_X1 U9363 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10359) );
  NOR2_X1 U9364 ( .A1(n10360), .A2(n10359), .ZN(n7527) );
  NOR2_X1 U9365 ( .A1(n7528), .A2(n7527), .ZN(n10358) );
  XNOR2_X1 U9366 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10357) );
  NOR2_X1 U9367 ( .A1(n10358), .A2(n10357), .ZN(n7529) );
  NOR2_X1 U9368 ( .A1(n7530), .A2(n7529), .ZN(n10364) );
  XNOR2_X1 U9369 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10363) );
  NOR2_X1 U9370 ( .A1(n10364), .A2(n10363), .ZN(n7531) );
  NOR2_X1 U9371 ( .A1(n7532), .A2(n7531), .ZN(n10366) );
  XNOR2_X1 U9372 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10365) );
  NOR2_X1 U9373 ( .A1(n10366), .A2(n10365), .ZN(n7533) );
  NOR2_X1 U9374 ( .A1(n7534), .A2(n7533), .ZN(n10362) );
  INV_X1 U9375 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7535) );
  INV_X1 U9376 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U9377 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7535), .B1(
        P2_ADDR_REG_9__SCAN_IN), .B2(n9888), .ZN(n10361) );
  NOR2_X1 U9378 ( .A1(n10362), .A2(n10361), .ZN(n7536) );
  NOR2_X1 U9379 ( .A1(n7537), .A2(n7536), .ZN(n10356) );
  INV_X1 U9380 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7538) );
  INV_X1 U9381 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9653) );
  AOI22_X1 U9382 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n7538), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(n9653), .ZN(n10355) );
  NOR2_X1 U9383 ( .A1(n10356), .A2(n10355), .ZN(n7539) );
  NOR2_X1 U9384 ( .A1(n7540), .A2(n7539), .ZN(n10354) );
  XNOR2_X1 U9385 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10353) );
  NOR2_X1 U9386 ( .A1(n10354), .A2(n10353), .ZN(n7541) );
  NOR2_X1 U9387 ( .A1(n7542), .A2(n7541), .ZN(n10352) );
  XNOR2_X1 U9388 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10351) );
  NOR2_X1 U9389 ( .A1(n10352), .A2(n10351), .ZN(n7543) );
  NOR2_X1 U9390 ( .A1(n7544), .A2(n7543), .ZN(n10350) );
  XNOR2_X1 U9391 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10349) );
  NOR2_X1 U9392 ( .A1(n10350), .A2(n10349), .ZN(n7545) );
  NOR2_X1 U9393 ( .A1(n7546), .A2(n7545), .ZN(n10348) );
  XNOR2_X1 U9394 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10347) );
  NOR2_X1 U9395 ( .A1(n10348), .A2(n10347), .ZN(n7547) );
  NOR2_X1 U9396 ( .A1(n7548), .A2(n7547), .ZN(n10346) );
  AOI22_X1 U9397 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n8553), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(n7550), .ZN(n10345) );
  NOR2_X1 U9398 ( .A1(n10346), .A2(n10345), .ZN(n7549) );
  AOI21_X1 U9399 ( .B1(n7550), .B2(n8553), .A(n7549), .ZN(n10344) );
  INV_X1 U9400 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7551) );
  INV_X1 U9401 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9758) );
  AOI22_X1 U9402 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n7551), .B1(
        P2_ADDR_REG_16__SCAN_IN), .B2(n9758), .ZN(n10343) );
  NOR2_X1 U9403 ( .A1(n10344), .A2(n10343), .ZN(n7552) );
  NOR2_X1 U9404 ( .A1(n7553), .A2(n7552), .ZN(n10342) );
  XNOR2_X1 U9405 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10341) );
  NOR2_X1 U9406 ( .A1(n10342), .A2(n10341), .ZN(n7554) );
  NOR2_X1 U9407 ( .A1(n7555), .A2(n7554), .ZN(n7556) );
  NOR2_X1 U9408 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7556), .ZN(n10339) );
  AND2_X1 U9409 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7556), .ZN(n10338) );
  NOR2_X1 U9410 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10338), .ZN(n7557) );
  NOR2_X1 U9411 ( .A1(n10339), .A2(n7557), .ZN(n7559) );
  XNOR2_X1 U9412 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7558) );
  XNOR2_X1 U9413 ( .A(n7559), .B(n7558), .ZN(ADD_1068_U4) );
  OAI21_X1 U9414 ( .B1(n7561), .B2(n7570), .A(n7560), .ZN(n7615) );
  INV_X1 U9415 ( .A(n7562), .ZN(n7584) );
  OAI211_X1 U9416 ( .C1(n7584), .C2(n4568), .A(n10010), .B(n4566), .ZN(n7563)
         );
  OAI21_X1 U9417 ( .B1(n7564), .B2(n9551), .A(n7563), .ZN(n7622) );
  OAI21_X1 U9418 ( .B1(n7566), .B2(n7565), .A(n8947), .ZN(n7627) );
  NOR2_X1 U9419 ( .A1(n7627), .A2(n7628), .ZN(n7626) );
  INV_X1 U9420 ( .A(n7567), .ZN(n8943) );
  NOR3_X1 U9421 ( .A1(n7626), .A2(n8943), .A3(n7587), .ZN(n7569) );
  INV_X1 U9422 ( .A(n8951), .ZN(n7568) );
  NOR2_X1 U9423 ( .A1(n7569), .A2(n7568), .ZN(n7571) );
  XNOR2_X1 U9424 ( .A(n7571), .B(n7570), .ZN(n7573) );
  OAI22_X1 U9425 ( .A1(n7573), .A2(n10002), .B1(n7572), .B2(n9549), .ZN(n7616)
         );
  AOI211_X1 U9426 ( .C1(n6629), .C2(n7615), .A(n7622), .B(n7616), .ZN(n7580)
         );
  INV_X1 U9427 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7574) );
  OAI22_X1 U9428 ( .A1(n4568), .A2(n9936), .B1(n10101), .B2(n7574), .ZN(n7575)
         );
  INV_X1 U9429 ( .A(n7575), .ZN(n7576) );
  OAI21_X1 U9430 ( .B1(n7580), .B2(n10099), .A(n7576), .ZN(P1_U3480) );
  AOI22_X1 U9431 ( .A1(n7578), .A2(n7577), .B1(n10110), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7579) );
  OAI21_X1 U9432 ( .B1(n7580), .B2(n10110), .A(n7579), .ZN(P1_U3531) );
  OAI21_X1 U9433 ( .B1(n7582), .B2(n7587), .A(n7581), .ZN(n7596) );
  INV_X1 U9434 ( .A(n7583), .ZN(n7636) );
  AOI211_X1 U9435 ( .C1(n7585), .C2(n7636), .A(n9968), .B(n7584), .ZN(n7602)
         );
  NOR2_X1 U9436 ( .A1(n7626), .A2(n8943), .ZN(n7586) );
  XOR2_X1 U9437 ( .A(n7587), .B(n7586), .Z(n7588) );
  OAI222_X1 U9438 ( .A1(n9551), .A2(n7590), .B1(n9549), .B2(n7589), .C1(n7588), 
        .C2(n10002), .ZN(n7597) );
  AOI211_X1 U9439 ( .C1(n6629), .C2(n7596), .A(n7602), .B(n7597), .ZN(n7595)
         );
  OAI22_X1 U9440 ( .A1(n9616), .A2(n7600), .B1(n10113), .B2(n9860), .ZN(n7591)
         );
  INV_X1 U9441 ( .A(n7591), .ZN(n7592) );
  OAI21_X1 U9442 ( .B1(n7595), .B2(n10110), .A(n7592), .ZN(P1_U3530) );
  INV_X1 U9443 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9804) );
  OAI22_X1 U9444 ( .A1(n9936), .A2(n7600), .B1(n10101), .B2(n9804), .ZN(n7593)
         );
  INV_X1 U9445 ( .A(n7593), .ZN(n7594) );
  OAI21_X1 U9446 ( .B1(n7595), .B2(n10099), .A(n7594), .ZN(P1_U3477) );
  INV_X1 U9447 ( .A(n7596), .ZN(n7605) );
  NAND2_X1 U9448 ( .A1(n7597), .A2(n9989), .ZN(n7604) );
  AOI22_X1 U9449 ( .A1(n10019), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7598), .B2(
        n10017), .ZN(n7599) );
  OAI21_X1 U9450 ( .B1(n10022), .B2(n7600), .A(n7599), .ZN(n7601) );
  AOI21_X1 U9451 ( .B1(n7602), .B2(n10015), .A(n7601), .ZN(n7603) );
  OAI211_X1 U9452 ( .C1(n7605), .C2(n9554), .A(n7604), .B(n7603), .ZN(P1_U3285) );
  MUX2_X1 U9453 ( .A(n6837), .B(n7606), .S(n9989), .Z(n7613) );
  INV_X1 U9454 ( .A(n7607), .ZN(n7611) );
  OAI22_X1 U9455 ( .A1(n10022), .A2(n7609), .B1(n7608), .B2(n9994), .ZN(n7610)
         );
  AOI21_X1 U9456 ( .B1(n7611), .B2(n10015), .A(n7610), .ZN(n7612) );
  OAI211_X1 U9457 ( .C1(n7614), .C2(n9554), .A(n7613), .B(n7612), .ZN(P1_U3289) );
  INV_X1 U9458 ( .A(n7615), .ZN(n7625) );
  NAND2_X1 U9459 ( .A1(n7616), .A2(n9989), .ZN(n7624) );
  NOR2_X1 U9460 ( .A1(n4568), .A2(n10022), .ZN(n7621) );
  INV_X1 U9461 ( .A(n7617), .ZN(n7618) );
  OAI22_X1 U9462 ( .A1(n9989), .A2(n7619), .B1(n7618), .B2(n9994), .ZN(n7620)
         );
  AOI211_X1 U9463 ( .C1(n7622), .C2(n10015), .A(n7621), .B(n7620), .ZN(n7623)
         );
  OAI211_X1 U9464 ( .C1(n7625), .C2(n9554), .A(n7624), .B(n7623), .ZN(P1_U3284) );
  AOI21_X1 U9465 ( .B1(n7628), .B2(n7627), .A(n7626), .ZN(n7634) );
  AOI22_X1 U9466 ( .A1(n9985), .A2(n9205), .B1(n9203), .B2(n9982), .ZN(n7633)
         );
  OR2_X1 U9467 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  NAND2_X1 U9468 ( .A1(n7631), .A2(n7630), .ZN(n10076) );
  NAND2_X1 U9469 ( .A1(n10076), .A2(n10005), .ZN(n7632) );
  OAI211_X1 U9470 ( .C1(n7634), .C2(n10002), .A(n7633), .B(n7632), .ZN(n10074)
         );
  INV_X1 U9471 ( .A(n10074), .ZN(n7644) );
  OR2_X1 U9472 ( .A1(n5604), .A2(n7635), .ZN(n7799) );
  INV_X1 U9473 ( .A(n7799), .ZN(n10012) );
  OAI211_X1 U9474 ( .C1(n10073), .C2(n7637), .A(n7636), .B(n10010), .ZN(n10072) );
  AOI22_X1 U9475 ( .A1(n10019), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7638), .B2(
        n10017), .ZN(n7641) );
  NAND2_X1 U9476 ( .A1(n10007), .A2(n7639), .ZN(n7640) );
  OAI211_X1 U9477 ( .C1(n10072), .C2(n9467), .A(n7641), .B(n7640), .ZN(n7642)
         );
  AOI21_X1 U9478 ( .B1(n10076), .B2(n10012), .A(n7642), .ZN(n7643) );
  OAI21_X1 U9479 ( .B1(n7644), .B2(n5604), .A(n7643), .ZN(P1_U3286) );
  AOI22_X1 U9480 ( .A1(n10007), .A2(n7645), .B1(n10017), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7646) );
  OAI21_X1 U9481 ( .B1(n9467), .B2(n7647), .A(n7646), .ZN(n7650) );
  MUX2_X1 U9482 ( .A(n7648), .B(P1_REG2_REG_2__SCAN_IN), .S(n5604), .Z(n7649)
         );
  AOI211_X1 U9483 ( .C1(n10012), .C2(n7651), .A(n7650), .B(n7649), .ZN(n7652)
         );
  INV_X1 U9484 ( .A(n7652), .ZN(P1_U3291) );
  INV_X1 U9485 ( .A(n7653), .ZN(n7662) );
  NOR2_X1 U9486 ( .A1(n5658), .A2(n10022), .ZN(n7657) );
  INV_X1 U9487 ( .A(n7758), .ZN(n7654) );
  OAI22_X1 U9488 ( .A1(n9989), .A2(n7655), .B1(n7654), .B2(n9994), .ZN(n7656)
         );
  AOI211_X1 U9489 ( .C1(n7658), .C2(n10015), .A(n7657), .B(n7656), .ZN(n7661)
         );
  NAND2_X1 U9490 ( .A1(n7659), .A2(n9989), .ZN(n7660) );
  OAI211_X1 U9491 ( .C1(n7662), .C2(n9554), .A(n7661), .B(n7660), .ZN(P1_U3283) );
  INV_X1 U9492 ( .A(n9554), .ZN(n10025) );
  AOI22_X1 U9493 ( .A1(n5604), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7663), .B2(
        n10017), .ZN(n7666) );
  NAND2_X1 U9494 ( .A1(n10007), .A2(n7664), .ZN(n7665) );
  OAI211_X1 U9495 ( .C1(n7667), .C2(n9467), .A(n7666), .B(n7665), .ZN(n7668)
         );
  AOI21_X1 U9496 ( .B1(n7669), .B2(n10025), .A(n7668), .ZN(n7670) );
  OAI21_X1 U9497 ( .B1(n7671), .B2(n5604), .A(n7670), .ZN(P1_U3288) );
  OAI21_X1 U9498 ( .B1(n9049), .B2(n7673), .A(n7672), .ZN(n7674) );
  AOI222_X1 U9499 ( .A1(n9980), .A2(n7674), .B1(n9209), .B2(n9985), .C1(n9207), 
        .C2(n9982), .ZN(n10068) );
  OAI21_X1 U9500 ( .B1(n7676), .B2(n8936), .A(n7675), .ZN(n10071) );
  INV_X1 U9501 ( .A(n7677), .ZN(n7680) );
  INV_X1 U9502 ( .A(n7678), .ZN(n7679) );
  OAI211_X1 U9503 ( .C1(n10067), .C2(n7680), .A(n7679), .B(n10010), .ZN(n10066) );
  AOI22_X1 U9504 ( .A1(n10019), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10017), .B2(
        n7681), .ZN(n7684) );
  NAND2_X1 U9505 ( .A1(n10007), .A2(n7682), .ZN(n7683) );
  OAI211_X1 U9506 ( .C1(n10066), .C2(n9467), .A(n7684), .B(n7683), .ZN(n7685)
         );
  AOI21_X1 U9507 ( .B1(n10071), .B2(n10025), .A(n7685), .ZN(n7686) );
  OAI21_X1 U9508 ( .B1(n10068), .B2(n5604), .A(n7686), .ZN(P1_U3290) );
  NAND2_X1 U9509 ( .A1(n7687), .A2(n8517), .ZN(n7688) );
  XNOR2_X1 U9510 ( .A(n8162), .B(n7690), .ZN(n7824) );
  XNOR2_X1 U9511 ( .A(n4403), .B(n6685), .ZN(n7712) );
  OR2_X1 U9512 ( .A1(n7824), .A2(n4904), .ZN(n7698) );
  NOR3_X1 U9513 ( .A1(n4403), .A2(n7690), .A3(n8516), .ZN(n7692) );
  INV_X1 U9514 ( .A(n8162), .ZN(n7691) );
  AOI211_X1 U9515 ( .C1(n7827), .C2(n7690), .A(n7692), .B(n7691), .ZN(n7695)
         );
  NOR3_X1 U9516 ( .A1(n7714), .A2(n8516), .A3(n6685), .ZN(n7693) );
  AOI211_X1 U9517 ( .C1(n7827), .C2(n6685), .A(n7693), .B(n8162), .ZN(n7694)
         );
  XNOR2_X1 U9518 ( .A(n10313), .B(n6685), .ZN(n7699) );
  XNOR2_X1 U9519 ( .A(n7699), .B(n8514), .ZN(n7826) );
  OAI21_X1 U9520 ( .B1(n7695), .B2(n7694), .A(n7826), .ZN(n7696) );
  INV_X1 U9521 ( .A(n7696), .ZN(n7697) );
  OAI21_X1 U9522 ( .B1(n7763), .B2(n7698), .A(n7697), .ZN(n7701) );
  OR2_X1 U9523 ( .A1(n7699), .A2(n8252), .ZN(n7700) );
  NAND2_X1 U9524 ( .A1(n7701), .A2(n7700), .ZN(n7746) );
  XNOR2_X1 U9525 ( .A(n7815), .B(n6685), .ZN(n7702) );
  NOR2_X1 U9526 ( .A1(n7702), .A2(n7736), .ZN(n7744) );
  NAND2_X1 U9527 ( .A1(n7702), .A2(n7736), .ZN(n7745) );
  INV_X1 U9528 ( .A(n7745), .ZN(n7703) );
  NOR2_X1 U9529 ( .A1(n7744), .A2(n7703), .ZN(n7704) );
  XNOR2_X1 U9530 ( .A(n7746), .B(n7704), .ZN(n7710) );
  NAND2_X1 U9531 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10198) );
  INV_X1 U9532 ( .A(n10198), .ZN(n7706) );
  NOR2_X1 U9533 ( .A1(n8252), .A2(n8495), .ZN(n7705) );
  AOI211_X1 U9534 ( .C1(n8474), .C2(n8512), .A(n7706), .B(n7705), .ZN(n7707)
         );
  OAI21_X1 U9535 ( .B1(n7816), .B2(n8444), .A(n7707), .ZN(n7708) );
  AOI21_X1 U9536 ( .B1(n7815), .B2(n8486), .A(n7708), .ZN(n7709) );
  OAI21_X1 U9537 ( .B1(n7710), .B2(n8488), .A(n7709), .ZN(P2_U3174) );
  XNOR2_X1 U9538 ( .A(n7763), .B(n8516), .ZN(n7711) );
  NOR2_X1 U9539 ( .A1(n7711), .A2(n7712), .ZN(n7765) );
  AOI21_X1 U9540 ( .B1(n7712), .B2(n7711), .A(n7765), .ZN(n7722) );
  INV_X1 U9541 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7713) );
  NOR2_X1 U9542 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7713), .ZN(n10144) );
  AOI21_X1 U9543 ( .B1(n8515), .B2(n8474), .A(n10144), .ZN(n7720) );
  NAND2_X1 U9544 ( .A1(n7714), .A2(n8486), .ZN(n7719) );
  INV_X1 U9545 ( .A(n7715), .ZN(n7716) );
  NAND2_X1 U9546 ( .A1(n8500), .A2(n7716), .ZN(n7718) );
  NAND2_X1 U9547 ( .A1(n8517), .A2(n8482), .ZN(n7717) );
  AND4_X1 U9548 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n7721)
         );
  OAI21_X1 U9549 ( .B1(n7722), .B2(n8488), .A(n7721), .ZN(P2_U3157) );
  INV_X1 U9550 ( .A(n7723), .ZN(n7725) );
  OAI222_X1 U9551 ( .A1(P2_U3151), .A2(n6091), .B1(n8418), .B2(n7725), .C1(
        n8415), .C2(n6017), .ZN(P2_U3269) );
  OAI222_X1 U9552 ( .A1(n8422), .A2(n7726), .B1(n8420), .B2(n7725), .C1(
        P1_U3086), .C2(n7724), .ZN(P1_U3329) );
  INV_X1 U9553 ( .A(n7727), .ZN(n7776) );
  AOI21_X1 U9554 ( .B1(n7991), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7728), .ZN(
        n7729) );
  OAI21_X1 U9555 ( .B1(n7776), .B2(n8418), .A(n7729), .ZN(P2_U3268) );
  INV_X1 U9556 ( .A(n8250), .ZN(n7730) );
  NAND3_X1 U9557 ( .A1(n7731), .A2(n7730), .A3(n8253), .ZN(n7732) );
  NAND2_X1 U9558 ( .A1(n7733), .A2(n7732), .ZN(n10310) );
  XOR2_X1 U9559 ( .A(n7734), .B(n8250), .Z(n7735) );
  OAI222_X1 U9560 ( .A1(n8719), .A2(n7827), .B1(n8710), .B2(n7736), .C1(n10252), .C2(n7735), .ZN(n10311) );
  NAND2_X1 U9561 ( .A1(n10311), .A2(n8714), .ZN(n7740) );
  OAI22_X1 U9562 ( .A1(n8714), .A2(n7737), .B1(n7830), .B2(n8711), .ZN(n7738)
         );
  AOI21_X1 U9563 ( .B1(n10313), .B2(n8728), .A(n7738), .ZN(n7739) );
  OAI211_X1 U9564 ( .C1(n8731), .C2(n10310), .A(n7740), .B(n7739), .ZN(
        P2_U3221) );
  INV_X1 U9565 ( .A(n7741), .ZN(n7803) );
  AOI21_X1 U9566 ( .B1(n7991), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7742), .ZN(
        n7743) );
  OAI21_X1 U9567 ( .B1(n7803), .B2(n8418), .A(n7743), .ZN(P2_U3267) );
  XNOR2_X1 U9568 ( .A(n7890), .B(n6685), .ZN(n7835) );
  XNOR2_X1 U9569 ( .A(n7835), .B(n8512), .ZN(n7837) );
  XOR2_X1 U9570 ( .A(n7837), .B(n7838), .Z(n7751) );
  INV_X1 U9571 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9893) );
  OAI22_X1 U9572 ( .A1(n8496), .A2(n7965), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9893), .ZN(n7747) );
  AOI21_X1 U9573 ( .B1(n8482), .B2(n8513), .A(n7747), .ZN(n7748) );
  OAI21_X1 U9574 ( .B1(n7891), .B2(n8444), .A(n7748), .ZN(n7749) );
  AOI21_X1 U9575 ( .B1(n7890), .B2(n8486), .A(n7749), .ZN(n7750) );
  OAI21_X1 U9576 ( .B1(n7751), .B2(n8488), .A(n7750), .ZN(P2_U3155) );
  INV_X1 U9577 ( .A(n7752), .ZN(n7754) );
  XNOR2_X1 U9578 ( .A(n4453), .B(n7850), .ZN(n7753) );
  NOR2_X1 U9579 ( .A1(n7753), .A2(n7754), .ZN(n7849) );
  AOI21_X1 U9580 ( .B1(n7754), .B2(n7753), .A(n7849), .ZN(n7762) );
  OAI22_X1 U9581 ( .A1(n7756), .A2(n8862), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7755), .ZN(n7757) );
  AOI21_X1 U9582 ( .B1(n7758), .B2(n8924), .A(n7757), .ZN(n7761) );
  NAND2_X1 U9583 ( .A1(n7759), .A2(n8909), .ZN(n7760) );
  OAI211_X1 U9584 ( .C1(n7762), .C2(n8912), .A(n7761), .B(n7760), .ZN(P1_U3217) );
  NOR2_X1 U9585 ( .A1(n7763), .A2(n8516), .ZN(n7764) );
  NOR3_X1 U9586 ( .A1(n7765), .A2(n7764), .A3(n7824), .ZN(n7823) );
  INV_X1 U9587 ( .A(n7823), .ZN(n7767) );
  OAI21_X1 U9588 ( .B1(n7765), .B2(n7764), .A(n7824), .ZN(n7766) );
  NAND3_X1 U9589 ( .A1(n7767), .A2(n8492), .A3(n7766), .ZN(n7774) );
  NAND2_X1 U9590 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10165) );
  INV_X1 U9591 ( .A(n10165), .ZN(n7768) );
  AOI21_X1 U9592 ( .B1(n8474), .B2(n8514), .A(n7768), .ZN(n7769) );
  OAI21_X1 U9593 ( .B1(n7770), .B2(n8495), .A(n7769), .ZN(n7771) );
  AOI21_X1 U9594 ( .B1(n7772), .B2(n8500), .A(n7771), .ZN(n7773) );
  OAI211_X1 U9595 ( .C1(n10304), .C2(n8503), .A(n7774), .B(n7773), .ZN(
        P2_U3176) );
  OAI222_X1 U9596 ( .A1(n8420), .A2(n7776), .B1(P1_U3086), .B2(n5558), .C1(
        n7775), .C2(n7801), .ZN(P1_U3328) );
  OAI21_X1 U9597 ( .B1(n7779), .B2(n7778), .A(n7777), .ZN(n7780) );
  NAND2_X1 U9598 ( .A1(n7780), .A2(n8917), .ZN(n7784) );
  AOI22_X1 U9599 ( .A1(n9982), .A2(n9199), .B1(n9200), .B2(n9985), .ZN(n7873)
         );
  NOR2_X1 U9600 ( .A1(n7873), .A2(n8862), .ZN(n7781) );
  AOI211_X1 U9601 ( .C1(n8924), .C2(n7875), .A(n7782), .B(n7781), .ZN(n7783)
         );
  OAI211_X1 U9602 ( .C1(n10087), .C2(n8928), .A(n7784), .B(n7783), .ZN(
        P1_U3224) );
  NAND2_X1 U9603 ( .A1(n7786), .A2(n7785), .ZN(n7787) );
  XOR2_X1 U9604 ( .A(n9060), .B(n7787), .Z(n7916) );
  INV_X1 U9605 ( .A(n7916), .ZN(n7800) );
  INV_X1 U9606 ( .A(n7788), .ZN(n7789) );
  AOI21_X1 U9607 ( .B1(n9060), .B2(n7790), .A(n7789), .ZN(n7793) );
  NAND2_X1 U9608 ( .A1(n7916), .A2(n10005), .ZN(n7792) );
  AOI22_X1 U9609 ( .A1(n9985), .A2(n9199), .B1(n9198), .B2(n9982), .ZN(n7791)
         );
  OAI211_X1 U9610 ( .C1(n10002), .C2(n7793), .A(n7792), .B(n7791), .ZN(n7914)
         );
  NAND2_X1 U9611 ( .A1(n7914), .A2(n9989), .ZN(n7798) );
  AOI211_X1 U9612 ( .C1(n7794), .C2(n9971), .A(n9968), .B(n7936), .ZN(n7915)
         );
  INV_X1 U9613 ( .A(n7794), .ZN(n8061) );
  AOI22_X1 U9614 ( .A1(n10019), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8058), .B2(
        n10017), .ZN(n7795) );
  OAI21_X1 U9615 ( .B1(n8061), .B2(n10022), .A(n7795), .ZN(n7796) );
  AOI21_X1 U9616 ( .B1(n7915), .B2(n10015), .A(n7796), .ZN(n7797) );
  OAI211_X1 U9617 ( .C1(n7800), .C2(n7799), .A(n7798), .B(n7797), .ZN(P1_U3279) );
  OAI222_X1 U9618 ( .A1(n8420), .A2(n7803), .B1(P1_U3086), .B2(n5554), .C1(
        n7802), .C2(n7801), .ZN(P1_U3327) );
  NAND2_X1 U9619 ( .A1(n7805), .A2(n7804), .ZN(n8259) );
  XNOR2_X1 U9620 ( .A(n7806), .B(n8259), .ZN(n7822) );
  XNOR2_X1 U9621 ( .A(n7807), .B(n8259), .ZN(n7808) );
  AOI222_X1 U9622 ( .A1(n8684), .A2(n7808), .B1(n8512), .B2(n10247), .C1(n8514), .C2(n10248), .ZN(n7814) );
  MUX2_X1 U9623 ( .A(n10194), .B(n7814), .S(n10333), .Z(n7810) );
  NAND2_X1 U9624 ( .A1(n7815), .A2(n8767), .ZN(n7809) );
  OAI211_X1 U9625 ( .C1(n8770), .C2(n7822), .A(n7810), .B(n7809), .ZN(P2_U3472) );
  INV_X1 U9626 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7811) );
  MUX2_X1 U9627 ( .A(n7811), .B(n7814), .S(n10315), .Z(n7813) );
  INV_X1 U9628 ( .A(n8796), .ZN(n8828) );
  NAND2_X1 U9629 ( .A1(n7815), .A2(n8828), .ZN(n7812) );
  OAI211_X1 U9630 ( .C1(n7822), .C2(n8832), .A(n7813), .B(n7812), .ZN(P2_U3429) );
  INV_X1 U9631 ( .A(n7814), .ZN(n7819) );
  INV_X1 U9632 ( .A(n7815), .ZN(n7817) );
  OAI22_X1 U9633 ( .A1(n7817), .A2(n10254), .B1(n7816), .B2(n8711), .ZN(n7818)
         );
  OAI21_X1 U9634 ( .B1(n7819), .B2(n7818), .A(n8714), .ZN(n7821) );
  NAND2_X1 U9635 ( .A1(n10260), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7820) );
  OAI211_X1 U9636 ( .C1(n7822), .C2(n8731), .A(n7821), .B(n7820), .ZN(P2_U3220) );
  AOI21_X1 U9637 ( .B1(n8515), .B2(n7824), .A(n7823), .ZN(n7825) );
  XOR2_X1 U9638 ( .A(n7826), .B(n7825), .Z(n7833) );
  INV_X1 U9639 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9736) );
  NOR2_X1 U9640 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9736), .ZN(n10177) );
  NOR2_X1 U9641 ( .A1(n7827), .A2(n8495), .ZN(n7828) );
  AOI211_X1 U9642 ( .C1(n8474), .C2(n8513), .A(n10177), .B(n7828), .ZN(n7829)
         );
  OAI21_X1 U9643 ( .B1(n7830), .B2(n8444), .A(n7829), .ZN(n7831) );
  AOI21_X1 U9644 ( .B1(n10313), .B2(n8486), .A(n7831), .ZN(n7832) );
  OAI21_X1 U9645 ( .B1(n7833), .B2(n8488), .A(n7832), .ZN(P2_U3164) );
  INV_X1 U9646 ( .A(n7961), .ZN(n7845) );
  AND2_X1 U9647 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  AOI21_X1 U9648 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7840) );
  XNOR2_X1 U9649 ( .A(n7961), .B(n6685), .ZN(n7966) );
  XNOR2_X1 U9650 ( .A(n7966), .B(n8511), .ZN(n7839) );
  OAI211_X1 U9651 ( .C1(n7840), .C2(n7839), .A(n7968), .B(n8492), .ZN(n7844)
         );
  NAND2_X1 U9652 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8552) );
  OAI21_X1 U9653 ( .B1(n8496), .B2(n8720), .A(n8552), .ZN(n7842) );
  NOR2_X1 U9654 ( .A1(n8444), .A2(n7959), .ZN(n7841) );
  AOI211_X1 U9655 ( .C1(n8482), .C2(n8512), .A(n7842), .B(n7841), .ZN(n7843)
         );
  OAI211_X1 U9656 ( .C1(n7845), .C2(n8503), .A(n7844), .B(n7843), .ZN(P2_U3181) );
  OAI21_X1 U9657 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n7852) );
  AOI21_X1 U9658 ( .B1(n7850), .B2(n4453), .A(n7849), .ZN(n7851) );
  XOR2_X1 U9659 ( .A(n7852), .B(n7851), .Z(n7856) );
  AOI22_X1 U9660 ( .A1(n9985), .A2(n9201), .B1(n9984), .B2(n9982), .ZN(n10001)
         );
  OAI22_X1 U9661 ( .A1(n10001), .A2(n8862), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9280), .ZN(n7854) );
  NOR2_X1 U9662 ( .A1(n10079), .A2(n8928), .ZN(n7853) );
  AOI211_X1 U9663 ( .C1(n8924), .C2(n10006), .A(n7854), .B(n7853), .ZN(n7855)
         );
  OAI21_X1 U9664 ( .B1(n7856), .B2(n8912), .A(n7855), .ZN(P1_U3236) );
  INV_X1 U9665 ( .A(n9969), .ZN(n10096) );
  OAI21_X1 U9666 ( .B1(n7859), .B2(n7858), .A(n7857), .ZN(n7860) );
  NAND2_X1 U9667 ( .A1(n7860), .A2(n8917), .ZN(n7866) );
  NAND2_X1 U9668 ( .A1(n8903), .A2(n9984), .ZN(n7862) );
  OAI211_X1 U9669 ( .C1(n8922), .C2(n8843), .A(n7862), .B(n7861), .ZN(n7863)
         );
  AOI21_X1 U9670 ( .B1(n7864), .B2(n8924), .A(n7863), .ZN(n7865) );
  OAI211_X1 U9671 ( .C1(n10096), .C2(n8928), .A(n7866), .B(n7865), .ZN(
        P1_U3234) );
  OAI222_X1 U9672 ( .A1(n8420), .A2(n7927), .B1(n7868), .B2(P1_U3086), .C1(
        n7867), .C2(n8422), .ZN(P1_U3326) );
  AND2_X1 U9673 ( .A1(n4462), .A2(n7870), .ZN(n7871) );
  XNOR2_X1 U9674 ( .A(n7871), .B(n9059), .ZN(n10090) );
  INV_X1 U9675 ( .A(n10090), .ZN(n7880) );
  XNOR2_X1 U9676 ( .A(n7872), .B(n9059), .ZN(n7874) );
  OAI21_X1 U9677 ( .B1(n7874), .B2(n10002), .A(n7873), .ZN(n10089) );
  OAI211_X1 U9678 ( .C1(n10009), .C2(n10087), .A(n9970), .B(n10010), .ZN(
        n10086) );
  AOI22_X1 U9679 ( .A1(n10019), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7875), .B2(
        n10017), .ZN(n7877) );
  NAND2_X1 U9680 ( .A1(n5606), .A2(n10007), .ZN(n7876) );
  OAI211_X1 U9681 ( .C1(n10086), .C2(n9467), .A(n7877), .B(n7876), .ZN(n7878)
         );
  AOI21_X1 U9682 ( .B1(n10089), .B2(n9989), .A(n7878), .ZN(n7879) );
  OAI21_X1 U9683 ( .B1(n7880), .B2(n9554), .A(n7879), .ZN(P1_U3281) );
  NAND2_X1 U9684 ( .A1(n8266), .A2(n8269), .ZN(n8164) );
  XNOR2_X1 U9685 ( .A(n7881), .B(n8264), .ZN(n7897) );
  XNOR2_X1 U9686 ( .A(n7882), .B(n8264), .ZN(n7883) );
  AOI222_X1 U9687 ( .A1(n8684), .A2(n7883), .B1(n8511), .B2(n10247), .C1(n8513), .C2(n10248), .ZN(n7889) );
  MUX2_X1 U9688 ( .A(n9853), .B(n7889), .S(n10333), .Z(n7885) );
  NAND2_X1 U9689 ( .A1(n7890), .A2(n8767), .ZN(n7884) );
  OAI211_X1 U9690 ( .C1(n7897), .C2(n8770), .A(n7885), .B(n7884), .ZN(P2_U3473) );
  INV_X1 U9691 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7886) );
  MUX2_X1 U9692 ( .A(n7886), .B(n7889), .S(n10315), .Z(n7888) );
  NAND2_X1 U9693 ( .A1(n7890), .A2(n8828), .ZN(n7887) );
  OAI211_X1 U9694 ( .C1(n7897), .C2(n8832), .A(n7888), .B(n7887), .ZN(P2_U3432) );
  INV_X1 U9695 ( .A(n7889), .ZN(n7894) );
  INV_X1 U9696 ( .A(n7890), .ZN(n7892) );
  OAI22_X1 U9697 ( .A1(n7892), .A2(n10254), .B1(n7891), .B2(n8711), .ZN(n7893)
         );
  OAI21_X1 U9698 ( .B1(n7894), .B2(n7893), .A(n8714), .ZN(n7896) );
  NAND2_X1 U9699 ( .A1(n10260), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7895) );
  OAI211_X1 U9700 ( .C1(n7897), .C2(n8731), .A(n7896), .B(n7895), .ZN(P2_U3219) );
  INV_X1 U9701 ( .A(n7898), .ZN(n7899) );
  AOI21_X1 U9702 ( .B1(n9063), .B2(n7900), .A(n7899), .ZN(n7922) );
  INV_X1 U9703 ( .A(n7922), .ZN(n7913) );
  NAND2_X1 U9704 ( .A1(n7901), .A2(n9980), .ZN(n7905) );
  AOI21_X1 U9705 ( .B1(n7940), .B2(n8977), .A(n9063), .ZN(n7904) );
  NAND2_X1 U9706 ( .A1(n9198), .A2(n9985), .ZN(n7903) );
  NAND2_X1 U9707 ( .A1(n9196), .A2(n9982), .ZN(n7902) );
  AND2_X1 U9708 ( .A1(n7903), .A2(n7902), .ZN(n8863) );
  OAI21_X1 U9709 ( .B1(n7905), .B2(n7904), .A(n8863), .ZN(n7920) );
  INV_X1 U9710 ( .A(n7937), .ZN(n7907) );
  INV_X1 U9711 ( .A(n7983), .ZN(n7906) );
  AOI211_X1 U9712 ( .C1(n7908), .C2(n7907), .A(n9968), .B(n7906), .ZN(n7921)
         );
  NAND2_X1 U9713 ( .A1(n7921), .A2(n10015), .ZN(n7910) );
  AOI22_X1 U9714 ( .A1(n10019), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8865), .B2(
        n10017), .ZN(n7909) );
  OAI211_X1 U9715 ( .C1(n8868), .C2(n10022), .A(n7910), .B(n7909), .ZN(n7911)
         );
  AOI21_X1 U9716 ( .B1(n7920), .B2(n9989), .A(n7911), .ZN(n7912) );
  OAI21_X1 U9717 ( .B1(n7913), .B2(n9554), .A(n7912), .ZN(P1_U3277) );
  INV_X1 U9718 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9312) );
  AOI211_X1 U9719 ( .C1(n7916), .C2(n10084), .A(n7915), .B(n7914), .ZN(n7918)
         );
  MUX2_X1 U9720 ( .A(n9312), .B(n7918), .S(n10113), .Z(n7917) );
  OAI21_X1 U9721 ( .B1(n8061), .B2(n9616), .A(n7917), .ZN(P1_U3536) );
  INV_X1 U9722 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9730) );
  MUX2_X1 U9723 ( .A(n9730), .B(n7918), .S(n10101), .Z(n7919) );
  OAI21_X1 U9724 ( .B1(n8061), .B2(n9936), .A(n7919), .ZN(P1_U3495) );
  INV_X1 U9725 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9748) );
  AOI211_X1 U9726 ( .C1(n7922), .C2(n6629), .A(n7921), .B(n7920), .ZN(n7924)
         );
  MUX2_X1 U9727 ( .A(n9748), .B(n7924), .S(n10113), .Z(n7923) );
  OAI21_X1 U9728 ( .B1(n8868), .B2(n9616), .A(n7923), .ZN(P1_U3538) );
  MUX2_X1 U9729 ( .A(n9762), .B(n7924), .S(n10101), .Z(n7925) );
  OAI21_X1 U9730 ( .B1(n8868), .B2(n9936), .A(n7925), .ZN(P1_U3501) );
  OAI222_X1 U9731 ( .A1(P2_U3151), .A2(n5698), .B1(n8418), .B2(n7927), .C1(
        n7926), .C2(n8415), .ZN(P2_U3266) );
  INV_X1 U9732 ( .A(n7928), .ZN(n7932) );
  OR2_X1 U9733 ( .A1(n7929), .A2(n7932), .ZN(n7930) );
  OR2_X1 U9734 ( .A1(n9974), .A2(n7930), .ZN(n7934) );
  OR2_X1 U9735 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U9736 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  XOR2_X1 U9737 ( .A(n9062), .B(n7935), .Z(n9628) );
  INV_X1 U9738 ( .A(n7936), .ZN(n7938) );
  AOI211_X1 U9739 ( .C1(n9623), .C2(n7938), .A(n9968), .B(n7937), .ZN(n9622)
         );
  AOI22_X1 U9740 ( .A1(n10019), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8925), .B2(
        n10017), .ZN(n7939) );
  OAI21_X1 U9741 ( .B1(n8929), .B2(n10022), .A(n7939), .ZN(n7944) );
  OAI21_X1 U9742 ( .B1(n9062), .B2(n7941), .A(n7940), .ZN(n7942) );
  AOI222_X1 U9743 ( .A1(n9980), .A2(n7942), .B1(n9983), .B2(n9985), .C1(n9197), 
        .C2(n9982), .ZN(n9626) );
  NOR2_X1 U9744 ( .A1(n9626), .A2(n10019), .ZN(n7943) );
  AOI211_X1 U9745 ( .C1(n9622), .C2(n10015), .A(n7944), .B(n7943), .ZN(n7945)
         );
  OAI21_X1 U9746 ( .B1(n9554), .B2(n9628), .A(n7945), .ZN(P1_U3278) );
  INV_X1 U9747 ( .A(n7947), .ZN(n7949) );
  AND2_X1 U9748 ( .A1(n7949), .A2(n7948), .ZN(n8165) );
  INV_X1 U9749 ( .A(n8165), .ZN(n7950) );
  XNOR2_X1 U9750 ( .A(n7946), .B(n7950), .ZN(n7964) );
  INV_X1 U9751 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7953) );
  XOR2_X1 U9752 ( .A(n7951), .B(n8165), .Z(n7952) );
  AOI222_X1 U9753 ( .A1(n8684), .A2(n7952), .B1(n8510), .B2(n10247), .C1(n8512), .C2(n10248), .ZN(n7958) );
  MUX2_X1 U9754 ( .A(n7953), .B(n7958), .S(n10315), .Z(n7955) );
  NAND2_X1 U9755 ( .A1(n7961), .A2(n8828), .ZN(n7954) );
  OAI211_X1 U9756 ( .C1(n7964), .C2(n8832), .A(n7955), .B(n7954), .ZN(P2_U3435) );
  MUX2_X1 U9757 ( .A(n9899), .B(n7958), .S(n10333), .Z(n7957) );
  NAND2_X1 U9758 ( .A1(n7961), .A2(n8767), .ZN(n7956) );
  OAI211_X1 U9759 ( .C1(n8770), .C2(n7964), .A(n7957), .B(n7956), .ZN(P2_U3474) );
  OAI21_X1 U9760 ( .B1(n7959), .B2(n8711), .A(n7958), .ZN(n7960) );
  NAND2_X1 U9761 ( .A1(n7960), .A2(n8714), .ZN(n7963) );
  AOI22_X1 U9762 ( .A1(n7961), .A2(n8728), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n10260), .ZN(n7962) );
  OAI211_X1 U9763 ( .C1(n7964), .C2(n8731), .A(n7963), .B(n7962), .ZN(P2_U3218) );
  XNOR2_X1 U9764 ( .A(n8048), .B(n6685), .ZN(n8018) );
  XNOR2_X1 U9765 ( .A(n8018), .B(n8720), .ZN(n7970) );
  OR2_X1 U9766 ( .A1(n7966), .A2(n7965), .ZN(n7967) );
  AOI21_X1 U9767 ( .B1(n7970), .B2(n7969), .A(n8022), .ZN(n7976) );
  NAND2_X1 U9768 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8567) );
  OAI21_X1 U9769 ( .B1(n8496), .B2(n8708), .A(n8567), .ZN(n7971) );
  AOI21_X1 U9770 ( .B1(n8482), .B2(n8511), .A(n7971), .ZN(n7972) );
  OAI21_X1 U9771 ( .B1(n7973), .B2(n8444), .A(n7972), .ZN(n7974) );
  AOI21_X1 U9772 ( .B1(n8048), .B2(n8486), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9773 ( .B1(n7976), .B2(n8488), .A(n7975), .ZN(P2_U3166) );
  XNOR2_X1 U9774 ( .A(n7977), .B(n9065), .ZN(n9621) );
  INV_X1 U9775 ( .A(n7978), .ZN(n7979) );
  AOI21_X1 U9776 ( .B1(n9065), .B2(n7980), .A(n7979), .ZN(n7981) );
  OAI222_X1 U9777 ( .A1(n9549), .A2(n8877), .B1(n9551), .B2(n9548), .C1(n10002), .C2(n7981), .ZN(n9617) );
  INV_X1 U9778 ( .A(n8006), .ZN(n7982) );
  AOI211_X1 U9779 ( .C1(n9619), .C2(n7983), .A(n9968), .B(n7982), .ZN(n9618)
         );
  NAND2_X1 U9780 ( .A1(n9618), .A2(n10015), .ZN(n7985) );
  AOI22_X1 U9781 ( .A1(n10019), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8874), .B2(
        n10017), .ZN(n7984) );
  OAI211_X1 U9782 ( .C1(n4570), .C2(n10022), .A(n7985), .B(n7984), .ZN(n7986)
         );
  AOI21_X1 U9783 ( .B1(n9617), .B2(n9989), .A(n7986), .ZN(n7987) );
  OAI21_X1 U9784 ( .B1(n9554), .B2(n9621), .A(n7987), .ZN(P1_U3276) );
  INV_X1 U9785 ( .A(n8143), .ZN(n7998) );
  NOR4_X1 U9786 ( .A1(n7989), .A2(n7988), .A3(P2_U3151), .A4(
        P2_IR_REG_30__SCAN_IN), .ZN(n7990) );
  AOI21_X1 U9787 ( .B1(n7991), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n7990), .ZN(
        n7992) );
  OAI21_X1 U9788 ( .B1(n7998), .B2(n8418), .A(n7992), .ZN(P2_U3264) );
  NOR4_X1 U9789 ( .A1(n7994), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n7993), .ZN(n7995) );
  AOI21_X1 U9790 ( .B1(n7996), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n7995), .ZN(
        n7997) );
  OAI21_X1 U9791 ( .B1(n7998), .B2(n8420), .A(n7997), .ZN(P1_U3324) );
  NOR2_X1 U9792 ( .A1(n5753), .A2(n9820), .ZN(n7999) );
  INV_X1 U9793 ( .A(n8000), .ZN(n8001) );
  OR2_X1 U9794 ( .A1(n8186), .A2(n8001), .ZN(n8771) );
  NOR2_X1 U9795 ( .A1(n8771), .A2(n6673), .ZN(n8732) );
  AOI21_X1 U9796 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n6673), .A(n8732), .ZN(
        n8002) );
  OAI21_X1 U9797 ( .B1(n8180), .B2(n8747), .A(n8002), .ZN(P2_U3489) );
  OAI22_X1 U9798 ( .A1(n10260), .A2(n8771), .B1(n8097), .B2(n8711), .ZN(n8599)
         );
  AOI21_X1 U9799 ( .B1(n10260), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8599), .ZN(
        n8003) );
  OAI21_X1 U9800 ( .B1(n8180), .B2(n8601), .A(n8003), .ZN(P2_U3203) );
  OAI21_X1 U9801 ( .B1(n8005), .B2(n9066), .A(n8004), .ZN(n9613) );
  INV_X1 U9802 ( .A(n9613), .ZN(n8017) );
  AOI211_X1 U9803 ( .C1(n8910), .C2(n8006), .A(n9968), .B(n9538), .ZN(n9612)
         );
  NOR2_X1 U9804 ( .A1(n4569), .A2(n10022), .ZN(n8008) );
  INV_X1 U9805 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9377) );
  OAI22_X1 U9806 ( .A1(n9989), .A2(n9377), .B1(n8906), .B2(n9994), .ZN(n8007)
         );
  AOI211_X1 U9807 ( .C1(n9612), .C2(n10015), .A(n8008), .B(n8007), .ZN(n8016)
         );
  OAI21_X1 U9808 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8012) );
  NAND2_X1 U9809 ( .A1(n8012), .A2(n9980), .ZN(n8014) );
  AOI22_X1 U9810 ( .A1(n9523), .A2(n9982), .B1(n9985), .B2(n9196), .ZN(n8013)
         );
  NAND2_X1 U9811 ( .A1(n8014), .A2(n8013), .ZN(n9611) );
  NAND2_X1 U9812 ( .A1(n9611), .A2(n9989), .ZN(n8015) );
  OAI211_X1 U9813 ( .C1(n8017), .C2(n9554), .A(n8016), .B(n8015), .ZN(P1_U3275) );
  INV_X1 U9814 ( .A(n8829), .ZN(n8030) );
  INV_X1 U9815 ( .A(n8018), .ZN(n8019) );
  NOR2_X1 U9816 ( .A1(n8019), .A2(n8510), .ZN(n8021) );
  XNOR2_X1 U9817 ( .A(n8829), .B(n6685), .ZN(n8062) );
  XNOR2_X1 U9818 ( .A(n8062), .B(n8509), .ZN(n8020) );
  INV_X1 U9819 ( .A(n8064), .ZN(n8024) );
  NOR3_X1 U9820 ( .A1(n8022), .A2(n8021), .A3(n8020), .ZN(n8023) );
  OAI21_X1 U9821 ( .B1(n8024), .B2(n8023), .A(n8492), .ZN(n8029) );
  INV_X1 U9822 ( .A(n8025), .ZN(n8727) );
  AOI22_X1 U9823 ( .A1(n8474), .A2(n8725), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8026) );
  OAI21_X1 U9824 ( .B1(n8720), .B2(n8495), .A(n8026), .ZN(n8027) );
  AOI21_X1 U9825 ( .B1(n8727), .B2(n8500), .A(n8027), .ZN(n8028) );
  OAI211_X1 U9826 ( .C1(n8030), .C2(n8503), .A(n8029), .B(n8028), .ZN(P2_U3168) );
  NAND2_X1 U9827 ( .A1(n8031), .A2(n8270), .ZN(n8032) );
  INV_X1 U9828 ( .A(n8033), .ZN(n8166) );
  XNOR2_X1 U9829 ( .A(n8032), .B(n8166), .ZN(n8051) );
  NAND2_X1 U9830 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  NAND2_X1 U9831 ( .A1(n8035), .A2(n8684), .ZN(n8036) );
  OR2_X1 U9832 ( .A1(n8037), .A2(n8036), .ZN(n8039) );
  AOI22_X1 U9833 ( .A1(n8509), .A2(n10247), .B1(n10248), .B2(n8511), .ZN(n8038) );
  MUX2_X1 U9834 ( .A(n8047), .B(n8040), .S(n10317), .Z(n8042) );
  NAND2_X1 U9835 ( .A1(n8048), .A2(n8828), .ZN(n8041) );
  OAI211_X1 U9836 ( .C1(n8051), .C2(n8832), .A(n8042), .B(n8041), .ZN(P2_U3438) );
  INV_X1 U9837 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8043) );
  MUX2_X1 U9838 ( .A(n8047), .B(n8043), .S(n10260), .Z(n8046) );
  AOI22_X1 U9839 ( .A1(n8048), .A2(n8728), .B1(n10257), .B2(n8044), .ZN(n8045)
         );
  OAI211_X1 U9840 ( .C1(n8051), .C2(n8731), .A(n8046), .B(n8045), .ZN(P2_U3217) );
  MUX2_X1 U9841 ( .A(n9771), .B(n8047), .S(n10333), .Z(n8050) );
  NAND2_X1 U9842 ( .A1(n8048), .A2(n8767), .ZN(n8049) );
  OAI211_X1 U9843 ( .C1(n8770), .C2(n8051), .A(n8050), .B(n8049), .ZN(P2_U3475) );
  NAND2_X1 U9844 ( .A1(n8054), .A2(n8917), .ZN(n8060) );
  AND2_X1 U9845 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9295) );
  AOI21_X1 U9846 ( .B1(n8919), .B2(n9198), .A(n9295), .ZN(n8055) );
  OAI21_X1 U9847 ( .B1(n8056), .B2(n8921), .A(n8055), .ZN(n8057) );
  AOI21_X1 U9848 ( .B1(n8058), .B2(n8924), .A(n8057), .ZN(n8059) );
  OAI211_X1 U9849 ( .C1(n8061), .C2(n8928), .A(n8060), .B(n8059), .ZN(P1_U3215) );
  NAND2_X1 U9850 ( .A1(n8062), .A2(n8708), .ZN(n8063) );
  XNOR2_X1 U9851 ( .A(n8764), .B(n6685), .ZN(n8103) );
  XNOR2_X1 U9852 ( .A(n8103), .B(n8725), .ZN(n8104) );
  XOR2_X1 U9853 ( .A(n8105), .B(n8104), .Z(n8069) );
  NAND2_X1 U9854 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8587) );
  OAI21_X1 U9855 ( .B1(n8496), .B2(n8709), .A(n8587), .ZN(n8065) );
  AOI21_X1 U9856 ( .B1(n8482), .B2(n8509), .A(n8065), .ZN(n8066) );
  OAI21_X1 U9857 ( .B1(n8712), .B2(n8444), .A(n8066), .ZN(n8067) );
  AOI21_X1 U9858 ( .B1(n8764), .B2(n8486), .A(n8067), .ZN(n8068) );
  OAI21_X1 U9859 ( .B1(n8069), .B2(n8488), .A(n8068), .ZN(P2_U3178) );
  OR2_X1 U9860 ( .A1(n5607), .A2(n8070), .ZN(n8072) );
  NAND2_X1 U9861 ( .A1(n8072), .A2(n8071), .ZN(n10065) );
  NAND2_X1 U9862 ( .A1(n10065), .A2(n10005), .ZN(n8080) );
  AOI22_X1 U9863 ( .A1(n8073), .A2(n9985), .B1(n9982), .B2(n9209), .ZN(n8079)
         );
  NAND2_X1 U9864 ( .A1(n8074), .A2(n5607), .ZN(n8076) );
  NAND2_X1 U9865 ( .A1(n8076), .A2(n8075), .ZN(n8077) );
  NAND2_X1 U9866 ( .A1(n8077), .A2(n9980), .ZN(n8078) );
  NAND3_X1 U9867 ( .A1(n8080), .A2(n8079), .A3(n8078), .ZN(n10063) );
  MUX2_X1 U9868 ( .A(n10063), .B(P1_REG2_REG_1__SCAN_IN), .S(n5604), .Z(n8087)
         );
  OAI211_X1 U9869 ( .C1(n10062), .C2(n8082), .A(n10010), .B(n8081), .ZN(n10061) );
  NAND2_X1 U9870 ( .A1(n10065), .A2(n10012), .ZN(n8085) );
  INV_X1 U9871 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9890) );
  OAI22_X1 U9872 ( .A1(n10022), .A2(n10062), .B1(n9890), .B2(n9994), .ZN(n8083) );
  INV_X1 U9873 ( .A(n8083), .ZN(n8084) );
  OAI211_X1 U9874 ( .C1(n9467), .C2(n10061), .A(n8085), .B(n8084), .ZN(n8086)
         );
  OR2_X1 U9875 ( .A1(n8087), .A2(n8086), .ZN(P1_U3292) );
  OAI222_X1 U9876 ( .A1(n8422), .A2(n8090), .B1(n8420), .B2(n8089), .C1(n8088), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U9877 ( .A(n8091), .ZN(n8095) );
  OAI222_X1 U9878 ( .A1(n8422), .A2(n8093), .B1(n8420), .B2(n8095), .C1(
        P1_U3086), .C2(n8092), .ZN(P1_U3325) );
  OAI222_X1 U9879 ( .A1(n8094), .A2(P2_U3151), .B1(n8418), .B2(n8095), .C1(
        n8415), .C2(n9820), .ZN(P2_U3265) );
  OAI22_X1 U9880 ( .A1(n8097), .A2(n8711), .B1(n9837), .B2(n8714), .ZN(n8098)
         );
  AOI21_X1 U9881 ( .B1(n8099), .B2(n8728), .A(n8098), .ZN(n8102) );
  OR2_X1 U9882 ( .A1(n6183), .A2(n8100), .ZN(n8101) );
  OAI211_X1 U9883 ( .C1(n8096), .C2(n10260), .A(n8102), .B(n8101), .ZN(
        P2_U3204) );
  AOI22_X2 U9884 ( .A1(n8105), .A2(n8104), .B1(n8696), .B2(n8103), .ZN(n8441)
         );
  XNOR2_X1 U9885 ( .A(n8760), .B(n6685), .ZN(n8106) );
  XNOR2_X1 U9886 ( .A(n8106), .B(n8709), .ZN(n8440) );
  INV_X1 U9887 ( .A(n8106), .ZN(n8107) );
  XNOR2_X1 U9888 ( .A(n8108), .B(n6685), .ZN(n8109) );
  XNOR2_X1 U9889 ( .A(n8109), .B(n8697), .ZN(n8473) );
  INV_X1 U9890 ( .A(n8109), .ZN(n8110) );
  XNOR2_X1 U9891 ( .A(n8809), .B(n6685), .ZN(n8112) );
  XNOR2_X1 U9892 ( .A(n8112), .B(n8111), .ZN(n8449) );
  INV_X1 U9893 ( .A(n8112), .ZN(n8113) );
  XNOR2_X1 U9894 ( .A(n8803), .B(n6685), .ZN(n8114) );
  XNOR2_X1 U9895 ( .A(n8114), .B(n8671), .ZN(n8481) );
  XNOR2_X1 U9896 ( .A(n8797), .B(n6685), .ZN(n8115) );
  OAI21_X2 U9897 ( .B1(n8433), .B2(n8657), .A(n4920), .ZN(n8464) );
  XNOR2_X1 U9898 ( .A(n8469), .B(n6685), .ZN(n8117) );
  XNOR2_X1 U9899 ( .A(n8117), .B(n8508), .ZN(n8465) );
  AOI21_X2 U9900 ( .B1(n8464), .B2(n8465), .A(n8118), .ZN(n8455) );
  XNOR2_X1 U9901 ( .A(n8461), .B(n6685), .ZN(n8119) );
  XNOR2_X1 U9902 ( .A(n8119), .B(n8628), .ZN(n8456) );
  INV_X1 U9903 ( .A(n8119), .ZN(n8120) );
  INV_X1 U9904 ( .A(n8628), .ZN(n8608) );
  OAI22_X2 U9905 ( .A1(n8455), .A2(n8456), .B1(n8120), .B2(n8608), .ZN(n8490)
         );
  XNOR2_X1 U9906 ( .A(n8786), .B(n6685), .ZN(n8121) );
  XNOR2_X1 U9907 ( .A(n8121), .B(n8507), .ZN(n8491) );
  XNOR2_X1 U9908 ( .A(n8122), .B(n6685), .ZN(n8123) );
  NOR2_X1 U9909 ( .A1(n8123), .A2(n8497), .ZN(n8124) );
  AOI21_X1 U9910 ( .B1(n8497), .B2(n8123), .A(n8124), .ZN(n8424) );
  XNOR2_X1 U9911 ( .A(n8171), .B(n6685), .ZN(n8125) );
  AOI22_X1 U9912 ( .A1(n8506), .A2(n8474), .B1(n8126), .B2(n8500), .ZN(n8128)
         );
  NAND2_X1 U9913 ( .A1(P2_U3151), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8127) );
  OAI211_X1 U9914 ( .C1(n8497), .C2(n8495), .A(n8128), .B(n8127), .ZN(n8129)
         );
  AOI21_X1 U9915 ( .B1(n8781), .B2(n8486), .A(n8129), .ZN(n8130) );
  OAI21_X1 U9916 ( .B1(n8131), .B2(n8488), .A(n8130), .ZN(P2_U3160) );
  NAND2_X1 U9917 ( .A1(n8383), .A2(n8382), .ZN(n8133) );
  NAND2_X1 U9918 ( .A1(n8133), .A2(n8132), .ZN(n8136) );
  INV_X1 U9919 ( .A(n8134), .ZN(n8135) );
  XNOR2_X1 U9920 ( .A(n8136), .B(n8135), .ZN(n8141) );
  OAI22_X1 U9921 ( .A1(n9442), .A2(n8921), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9904), .ZN(n8137) );
  AOI21_X1 U9922 ( .B1(n8919), .B2(n8403), .A(n8137), .ZN(n8138) );
  OAI21_X1 U9923 ( .B1(n9445), .B2(n8907), .A(n8138), .ZN(n8139) );
  AOI21_X1 U9924 ( .B1(n9575), .B2(n8909), .A(n8139), .ZN(n8140) );
  OAI21_X1 U9925 ( .B1(n8141), .B2(n8912), .A(n8140), .ZN(P1_U3225) );
  NAND2_X1 U9926 ( .A1(n8143), .A2(n8142), .ZN(n8146) );
  OR2_X1 U9927 ( .A1(n5753), .A2(n8144), .ZN(n8145) );
  OR2_X1 U9928 ( .A1(n8598), .A2(n8186), .ZN(n8179) );
  INV_X1 U9929 ( .A(n8179), .ZN(n8355) );
  INV_X1 U9930 ( .A(n8147), .ZN(n8325) );
  NAND2_X1 U9931 ( .A1(n8311), .A2(n8316), .ZN(n8636) );
  AND2_X1 U9932 ( .A1(n8632), .A2(n8633), .ZN(n8639) );
  INV_X1 U9933 ( .A(n8653), .ZN(n8651) );
  NAND3_X1 U9934 ( .A1(n8148), .A2(n8149), .A3(n8210), .ZN(n8152) );
  NAND2_X1 U9935 ( .A1(n6119), .A2(n8150), .ZN(n8151) );
  NOR2_X1 U9936 ( .A1(n8152), .A2(n8151), .ZN(n8156) );
  NAND4_X1 U9937 ( .A1(n8156), .A2(n8155), .A3(n8154), .A4(n8153), .ZN(n8160)
         );
  NOR4_X1 U9938 ( .A1(n8160), .A2(n8159), .A3(n8158), .A4(n8157), .ZN(n8161)
         );
  NAND4_X1 U9939 ( .A1(n8259), .A2(n8162), .A3(n8161), .A4(n8250), .ZN(n8163)
         );
  NOR4_X1 U9940 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n8167)
         );
  NAND4_X1 U9941 ( .A1(n8722), .A2(n8167), .A3(n8276), .A4(n8283), .ZN(n8168)
         );
  NOR3_X1 U9942 ( .A1(n8679), .A2(n8693), .A3(n8168), .ZN(n8169) );
  NAND4_X1 U9943 ( .A1(n8639), .A2(n8651), .A3(n8668), .A4(n8169), .ZN(n8170)
         );
  NOR4_X1 U9944 ( .A1(n8605), .A2(n6145), .A3(n8636), .A4(n8170), .ZN(n8172)
         );
  NAND4_X1 U9945 ( .A1(n8173), .A2(n8327), .A3(n8172), .A4(n8171), .ZN(n8176)
         );
  INV_X1 U9946 ( .A(n8180), .ZN(n8774) );
  INV_X1 U9947 ( .A(n8505), .ZN(n8174) );
  NAND2_X1 U9948 ( .A1(n8774), .A2(n8174), .ZN(n8351) );
  INV_X1 U9949 ( .A(n8351), .ZN(n8175) );
  NOR4_X1 U9950 ( .A1(n8355), .A2(n8176), .A3(n8353), .A4(n8175), .ZN(n8185)
         );
  INV_X1 U9951 ( .A(n8342), .ZN(n8177) );
  OAI21_X1 U9952 ( .B1(n8180), .B2(n8598), .A(n8179), .ZN(n8182) );
  NAND2_X1 U9953 ( .A1(n8351), .A2(n8181), .ZN(n8338) );
  NOR2_X1 U9954 ( .A1(n8182), .A2(n8338), .ZN(n8183) );
  NAND2_X1 U9955 ( .A1(n8598), .A2(n8186), .ZN(n8347) );
  NAND2_X1 U9956 ( .A1(n8300), .A2(n8187), .ZN(n8190) );
  INV_X1 U9957 ( .A(n8188), .ZN(n8189) );
  MUX2_X1 U9958 ( .A(n8190), .B(n8189), .S(n8349), .Z(n8308) );
  NAND2_X1 U9959 ( .A1(n8198), .A2(n8193), .ZN(n8192) );
  INV_X1 U9960 ( .A(n8197), .ZN(n8191) );
  MUX2_X1 U9961 ( .A(n8192), .B(n8191), .S(n8349), .Z(n8201) );
  NAND2_X1 U9962 ( .A1(n8193), .A2(n8349), .ZN(n8194) );
  AOI21_X1 U9963 ( .B1(n8196), .B2(n8195), .A(n8194), .ZN(n8200) );
  MUX2_X1 U9964 ( .A(n8198), .B(n8197), .S(n8354), .Z(n8199) );
  OAI211_X1 U9965 ( .C1(n8201), .C2(n8200), .A(n8148), .B(n8199), .ZN(n8209)
         );
  NAND2_X1 U9966 ( .A1(n8203), .A2(n8202), .ZN(n8206) );
  NAND2_X1 U9967 ( .A1(n8217), .A2(n8204), .ZN(n8205) );
  MUX2_X1 U9968 ( .A(n8206), .B(n8205), .S(n8354), .Z(n8207) );
  INV_X1 U9969 ( .A(n8207), .ZN(n8208) );
  NAND2_X1 U9970 ( .A1(n8209), .A2(n8208), .ZN(n8211) );
  NAND2_X1 U9971 ( .A1(n8211), .A2(n8210), .ZN(n8220) );
  NAND2_X1 U9972 ( .A1(n8522), .A2(n10271), .ZN(n8212) );
  OAI211_X1 U9973 ( .C1(n8220), .C2(n4808), .A(n8212), .B(n8221), .ZN(n8214)
         );
  NAND3_X1 U9974 ( .A1(n8214), .A2(n8223), .A3(n8213), .ZN(n8215) );
  NAND2_X1 U9975 ( .A1(n8215), .A2(n8225), .ZN(n8216) );
  NAND3_X1 U9976 ( .A1(n8242), .A2(n8349), .A3(n8238), .ZN(n8229) );
  NAND2_X1 U9977 ( .A1(n8216), .A2(n8229), .ZN(n8232) );
  INV_X1 U9978 ( .A(n8217), .ZN(n8219) );
  OAI21_X1 U9979 ( .B1(n8220), .B2(n8219), .A(n8218), .ZN(n8222) );
  NAND2_X1 U9980 ( .A1(n8222), .A2(n8221), .ZN(n8224) );
  NAND2_X1 U9981 ( .A1(n8224), .A2(n8223), .ZN(n8226) );
  NAND3_X1 U9982 ( .A1(n8226), .A2(n8349), .A3(n8225), .ZN(n8231) );
  NAND3_X1 U9983 ( .A1(n8236), .A2(n8227), .A3(n8354), .ZN(n8228) );
  NAND2_X1 U9984 ( .A1(n8229), .A2(n8228), .ZN(n8241) );
  NAND4_X1 U9985 ( .A1(n8232), .A2(n8231), .A3(n8241), .A4(n8230), .ZN(n8246)
         );
  INV_X1 U9986 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U9987 ( .A1(n8241), .A2(n8234), .ZN(n8237) );
  INV_X1 U9988 ( .A(n8235), .ZN(n8247) );
  OAI21_X1 U9989 ( .B1(n8239), .B2(n8519), .A(n8238), .ZN(n8240) );
  NAND2_X1 U9990 ( .A1(n8241), .A2(n8240), .ZN(n8244) );
  NAND3_X1 U9991 ( .A1(n8244), .A2(n8243), .A3(n8242), .ZN(n8245) );
  NAND3_X1 U9992 ( .A1(n8256), .A2(n8247), .A3(n8253), .ZN(n8249) );
  NAND3_X1 U9993 ( .A1(n8249), .A2(n8354), .A3(n8248), .ZN(n8251) );
  NAND3_X1 U9994 ( .A1(n10313), .A2(n8354), .A3(n8252), .ZN(n8258) );
  NAND2_X1 U9995 ( .A1(n8253), .A2(n8349), .ZN(n8254) );
  AOI21_X1 U9996 ( .B1(n8256), .B2(n8255), .A(n8254), .ZN(n8257) );
  NAND2_X1 U9997 ( .A1(n8514), .A2(n8349), .ZN(n8260) );
  OAI21_X1 U9998 ( .B1(n10313), .B2(n8260), .A(n8259), .ZN(n8265) );
  MUX2_X1 U9999 ( .A(n8262), .B(n8261), .S(n8354), .Z(n8263) );
  INV_X1 U10000 ( .A(n8266), .ZN(n8267) );
  NOR2_X1 U10001 ( .A1(n8272), .A2(n8267), .ZN(n8268) );
  INV_X1 U10002 ( .A(n8272), .ZN(n8273) );
  NAND2_X1 U10003 ( .A1(n8280), .A2(n4926), .ZN(n8275) );
  NAND2_X1 U10004 ( .A1(n8275), .A2(n8274), .ZN(n8278) );
  AND2_X1 U10005 ( .A1(n8722), .A2(n8354), .ZN(n8277) );
  NAND4_X1 U10006 ( .A1(n8278), .A2(n8277), .A3(n8292), .A4(n8276), .ZN(n8296)
         );
  NAND2_X1 U10007 ( .A1(n8280), .A2(n8279), .ZN(n8282) );
  NAND2_X1 U10008 ( .A1(n8282), .A2(n8281), .ZN(n8284) );
  NAND4_X1 U10009 ( .A1(n8284), .A2(n8349), .A3(n8286), .A4(n8283), .ZN(n8295)
         );
  NOR2_X1 U10010 ( .A1(n8286), .A2(n8725), .ZN(n8285) );
  OR3_X1 U10011 ( .A1(n8285), .A2(n8764), .A3(n8349), .ZN(n8291) );
  OAI211_X1 U10012 ( .C1(n8287), .C2(n8696), .A(n8764), .B(n8349), .ZN(n8290)
         );
  NAND3_X1 U10013 ( .A1(n8286), .A2(n8354), .A3(n8725), .ZN(n8289) );
  NAND3_X1 U10014 ( .A1(n8287), .A2(n8696), .A3(n8349), .ZN(n8288) );
  NAND4_X1 U10015 ( .A1(n8291), .A2(n8290), .A3(n8289), .A4(n8288), .ZN(n8293)
         );
  INV_X1 U10016 ( .A(n8292), .ZN(n8298) );
  NAND3_X1 U10017 ( .A1(n8296), .A2(n8295), .A3(n8294), .ZN(n8297) );
  NOR2_X1 U10018 ( .A1(n8679), .A2(n8298), .ZN(n8299) );
  AND2_X1 U10019 ( .A1(n8305), .A2(n8299), .ZN(n8301) );
  OAI211_X1 U10020 ( .C1(n8308), .C2(n8301), .A(n8651), .B(n8300), .ZN(n8303)
         );
  OAI211_X1 U10021 ( .C1(n8308), .C2(n8307), .A(n8651), .B(n8306), .ZN(n8310)
         );
  AND2_X1 U10022 ( .A1(n8311), .A2(n8632), .ZN(n8313) );
  MUX2_X1 U10023 ( .A(n8313), .B(n8312), .S(n8354), .Z(n8314) );
  MUX2_X1 U10024 ( .A(n8316), .B(n8315), .S(n8354), .Z(n8317) );
  NAND2_X1 U10025 ( .A1(n8319), .A2(n8318), .ZN(n8323) );
  MUX2_X1 U10026 ( .A(n8321), .B(n8320), .S(n8354), .Z(n8322) );
  AOI21_X1 U10027 ( .B1(n8323), .B2(n8322), .A(n8605), .ZN(n8329) );
  MUX2_X1 U10028 ( .A(n8325), .B(n8324), .S(n8354), .Z(n8326) );
  NAND2_X1 U10029 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  NOR2_X1 U10030 ( .A1(n8329), .A2(n8328), .ZN(n8334) );
  MUX2_X1 U10031 ( .A(n8331), .B(n8330), .S(n8349), .Z(n8332) );
  INV_X1 U10032 ( .A(n8332), .ZN(n8333) );
  MUX2_X1 U10033 ( .A(n8337), .B(n8340), .S(n8349), .Z(n8343) );
  OR2_X1 U10034 ( .A1(n8335), .A2(n8343), .ZN(n8336) );
  INV_X1 U10035 ( .A(n8338), .ZN(n8339) );
  INV_X1 U10036 ( .A(n8353), .ZN(n8341) );
  NOR2_X1 U10037 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  INV_X1 U10038 ( .A(n8347), .ZN(n8348) );
  AOI21_X1 U10039 ( .B1(n8350), .B2(n8349), .A(n8348), .ZN(n8357) );
  INV_X1 U10040 ( .A(n8350), .ZN(n8352) );
  OAI211_X1 U10041 ( .C1(n8354), .C2(n8353), .A(n8352), .B(n8351), .ZN(n8356)
         );
  AOI21_X1 U10042 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8358) );
  NOR3_X1 U10043 ( .A1(n8363), .A2(n6531), .A3(n8362), .ZN(n8366) );
  OAI21_X1 U10044 ( .B1(n8367), .B2(n8364), .A(P2_B_REG_SCAN_IN), .ZN(n8365)
         );
  INV_X1 U10045 ( .A(n8368), .ZN(n8892) );
  INV_X1 U10046 ( .A(n8370), .ZN(n8371) );
  NAND2_X1 U10047 ( .A1(n8890), .A2(n8372), .ZN(n8376) );
  XNOR2_X1 U10048 ( .A(n8374), .B(n8373), .ZN(n8375) );
  XNOR2_X1 U10049 ( .A(n8376), .B(n8375), .ZN(n8381) );
  AOI22_X1 U10050 ( .A1(n9194), .A2(n9982), .B1(n9985), .B2(n9512), .ZN(n9475)
         );
  INV_X1 U10051 ( .A(n8377), .ZN(n9478) );
  AOI22_X1 U10052 ( .A1(n9478), .A2(n8924), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8378) );
  OAI21_X1 U10053 ( .B1(n9475), .B2(n8862), .A(n8378), .ZN(n8379) );
  AOI21_X1 U10054 ( .B1(n9588), .B2(n8909), .A(n8379), .ZN(n8380) );
  OAI21_X1 U10055 ( .B1(n8381), .B2(n8912), .A(n8380), .ZN(P1_U3216) );
  XOR2_X1 U10056 ( .A(n8383), .B(n8382), .Z(n8389) );
  OAI22_X1 U10057 ( .A1(n8384), .A2(n8921), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9862), .ZN(n8385) );
  AOI21_X1 U10058 ( .B1(n8919), .B2(n9458), .A(n8385), .ZN(n8386) );
  OAI21_X1 U10059 ( .B1(n9462), .B2(n8907), .A(n8386), .ZN(n8387) );
  AOI21_X1 U10060 ( .B1(n9464), .B2(n8909), .A(n8387), .ZN(n8388) );
  OAI21_X1 U10061 ( .B1(n8389), .B2(n8912), .A(n8388), .ZN(P1_U3229) );
  XOR2_X1 U10062 ( .A(n9070), .B(n8390), .Z(n9567) );
  INV_X1 U10063 ( .A(n8391), .ZN(n8394) );
  INV_X1 U10064 ( .A(n8392), .ZN(n8393) );
  AOI211_X1 U10065 ( .C1(n9564), .C2(n8394), .A(n9968), .B(n8393), .ZN(n9563)
         );
  INV_X1 U10066 ( .A(n8395), .ZN(n8396) );
  AOI22_X1 U10067 ( .A1(n8396), .A2(n10017), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10019), .ZN(n8397) );
  OAI21_X1 U10068 ( .B1(n9025), .B2(n10022), .A(n8397), .ZN(n8408) );
  NAND2_X1 U10069 ( .A1(n9425), .A2(n9094), .ZN(n8401) );
  NAND2_X1 U10070 ( .A1(n8401), .A2(n9070), .ZN(n8400) );
  OAI21_X1 U10071 ( .B1(n9070), .B2(n8401), .A(n8400), .ZN(n8402) );
  NAND2_X1 U10072 ( .A1(n8402), .A2(n9980), .ZN(n8406) );
  NOR2_X1 U10073 ( .A1(n9566), .A2(n10019), .ZN(n8407) );
  AOI211_X1 U10074 ( .C1(n9563), .C2(n10015), .A(n8408), .B(n8407), .ZN(n8409)
         );
  OAI21_X1 U10075 ( .B1(n9567), .B2(n9554), .A(n8409), .ZN(P1_U3266) );
  INV_X1 U10076 ( .A(n8410), .ZN(n8414) );
  NAND2_X1 U10077 ( .A1(n9989), .A2(n9555), .ZN(n9406) );
  OAI21_X1 U10078 ( .B1(n9989), .B2(n8411), .A(n9406), .ZN(n8412) );
  AOI21_X1 U10079 ( .B1(n8931), .B2(n10007), .A(n8412), .ZN(n8413) );
  OAI21_X1 U10080 ( .B1(n8414), .B2(n9467), .A(n8413), .ZN(P1_U3263) );
  OAI222_X1 U10081 ( .A1(n6090), .A2(P2_U3151), .B1(n8418), .B2(n8417), .C1(
        n8416), .C2(n8415), .ZN(P2_U3271) );
  OAI222_X1 U10082 ( .A1(n8422), .A2(n8421), .B1(n8420), .B2(n8419), .C1(
        P1_U3086), .C2(n5654), .ZN(P1_U3336) );
  OAI211_X1 U10083 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n8492), .ZN(n8431)
         );
  NAND2_X1 U10084 ( .A1(P2_U3151), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10085 ( .A1(n8426), .A2(n8500), .ZN(n8427) );
  OAI211_X1 U10086 ( .C1(n8459), .C2(n8495), .A(n8428), .B(n8427), .ZN(n8429)
         );
  AOI21_X1 U10087 ( .B1(n4603), .B2(n8474), .A(n8429), .ZN(n8430) );
  OAI211_X1 U10088 ( .C1(n8432), .C2(n8503), .A(n8431), .B(n8430), .ZN(
        P2_U3154) );
  XNOR2_X1 U10089 ( .A(n8433), .B(n8657), .ZN(n8434) );
  NAND2_X1 U10090 ( .A1(n8434), .A2(n8492), .ZN(n8439) );
  INV_X1 U10091 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8435) );
  OAI22_X1 U10092 ( .A1(n8642), .A2(n8495), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8435), .ZN(n8437) );
  NOR2_X1 U10093 ( .A1(n8643), .A2(n8496), .ZN(n8436) );
  AOI211_X1 U10094 ( .C1(n8646), .C2(n8500), .A(n8437), .B(n8436), .ZN(n8438)
         );
  OAI211_X1 U10095 ( .C1(n8797), .C2(n8503), .A(n8439), .B(n8438), .ZN(
        P2_U3156) );
  XOR2_X1 U10096 ( .A(n8441), .B(n8440), .Z(n8447) );
  AOI22_X1 U10097 ( .A1(n8474), .A2(n8672), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8443) );
  NAND2_X1 U10098 ( .A1(n8482), .A2(n8725), .ZN(n8442) );
  OAI211_X1 U10099 ( .C1(n8444), .C2(n8698), .A(n8443), .B(n8442), .ZN(n8445)
         );
  AOI21_X1 U10100 ( .B1(n8760), .B2(n8486), .A(n8445), .ZN(n8446) );
  OAI21_X1 U10101 ( .B1(n8447), .B2(n8488), .A(n8446), .ZN(P2_U3159) );
  XOR2_X1 U10102 ( .A(n8449), .B(n8448), .Z(n8454) );
  AOI22_X1 U10103 ( .A1(n8671), .A2(n8474), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8451) );
  NAND2_X1 U10104 ( .A1(n8500), .A2(n8675), .ZN(n8450) );
  OAI211_X1 U10105 ( .C1(n8697), .C2(n8495), .A(n8451), .B(n8450), .ZN(n8452)
         );
  AOI21_X1 U10106 ( .B1(n8809), .B2(n8486), .A(n8452), .ZN(n8453) );
  OAI21_X1 U10107 ( .B1(n8454), .B2(n8488), .A(n8453), .ZN(P2_U3163) );
  XOR2_X1 U10108 ( .A(n8456), .B(n8455), .Z(n8463) );
  AOI22_X1 U10109 ( .A1(n8508), .A2(n8482), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8458) );
  NAND2_X1 U10110 ( .A1(n8617), .A2(n8500), .ZN(n8457) );
  OAI211_X1 U10111 ( .C1(n8459), .C2(n8496), .A(n8458), .B(n8457), .ZN(n8460)
         );
  AOI21_X1 U10112 ( .B1(n8461), .B2(n8486), .A(n8460), .ZN(n8462) );
  OAI21_X1 U10113 ( .B1(n8463), .B2(n8488), .A(n8462), .ZN(P2_U3165) );
  XOR2_X1 U10114 ( .A(n8465), .B(n8464), .Z(n8471) );
  AOI22_X1 U10115 ( .A1(n8608), .A2(n8474), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8467) );
  NAND2_X1 U10116 ( .A1(n8630), .A2(n8500), .ZN(n8466) );
  OAI211_X1 U10117 ( .C1(n8627), .C2(n8495), .A(n8467), .B(n8466), .ZN(n8468)
         );
  AOI21_X1 U10118 ( .B1(n8469), .B2(n8486), .A(n8468), .ZN(n8470) );
  OAI21_X1 U10119 ( .B1(n8471), .B2(n8488), .A(n8470), .ZN(P2_U3169) );
  XOR2_X1 U10120 ( .A(n8473), .B(n8472), .Z(n8479) );
  AOI22_X1 U10121 ( .A1(n8682), .A2(n8474), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8476) );
  NAND2_X1 U10122 ( .A1(n8500), .A2(n8686), .ZN(n8475) );
  OAI211_X1 U10123 ( .C1(n8709), .C2(n8495), .A(n8476), .B(n8475), .ZN(n8477)
         );
  AOI21_X1 U10124 ( .B1(n8815), .B2(n8486), .A(n8477), .ZN(n8478) );
  OAI21_X1 U10125 ( .B1(n8479), .B2(n8488), .A(n8478), .ZN(P2_U3173) );
  XOR2_X1 U10126 ( .A(n8481), .B(n8480), .Z(n8489) );
  AOI22_X1 U10127 ( .A1(n8682), .A2(n8482), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8484) );
  NAND2_X1 U10128 ( .A1(n8500), .A2(n8660), .ZN(n8483) );
  OAI211_X1 U10129 ( .C1(n8627), .C2(n8496), .A(n8484), .B(n8483), .ZN(n8485)
         );
  AOI21_X1 U10130 ( .B1(n8803), .B2(n8486), .A(n8485), .ZN(n8487) );
  OAI21_X1 U10131 ( .B1(n8489), .B2(n8488), .A(n8487), .ZN(P2_U3175) );
  XNOR2_X1 U10132 ( .A(n8490), .B(n8491), .ZN(n8493) );
  NAND2_X1 U10133 ( .A1(n8493), .A2(n8492), .ZN(n8502) );
  OAI22_X1 U10134 ( .A1(n8628), .A2(n8495), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8494), .ZN(n8499) );
  NOR2_X1 U10135 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  AOI211_X1 U10136 ( .C1(n8614), .C2(n8500), .A(n8499), .B(n8498), .ZN(n8501)
         );
  OAI211_X1 U10137 ( .C1(n8504), .C2(n8503), .A(n8502), .B(n8501), .ZN(
        P2_U3180) );
  MUX2_X1 U10138 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8505), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8506), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10140 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n4603), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10141 ( .A(n8607), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8584), .Z(
        P2_U3518) );
  MUX2_X1 U10142 ( .A(n8507), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8584), .Z(
        P2_U3517) );
  MUX2_X1 U10143 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8608), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10144 ( .A(n8508), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8584), .Z(
        P2_U3515) );
  MUX2_X1 U10145 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8657), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8671), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8682), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10148 ( .A(n8672), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8584), .Z(
        P2_U3511) );
  MUX2_X1 U10149 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8681), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10150 ( .A(n8725), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8584), .Z(
        P2_U3509) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8509), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10152 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8510), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10153 ( .A(n8511), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8584), .Z(
        P2_U3506) );
  MUX2_X1 U10154 ( .A(n8512), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8584), .Z(
        P2_U3505) );
  MUX2_X1 U10155 ( .A(n8513), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8584), .Z(
        P2_U3504) );
  MUX2_X1 U10156 ( .A(n8514), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8584), .Z(
        P2_U3503) );
  MUX2_X1 U10157 ( .A(n8515), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8584), .Z(
        P2_U3502) );
  MUX2_X1 U10158 ( .A(n8516), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8584), .Z(
        P2_U3501) );
  MUX2_X1 U10159 ( .A(n8517), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8584), .Z(
        P2_U3500) );
  MUX2_X1 U10160 ( .A(n8518), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8584), .Z(
        P2_U3499) );
  MUX2_X1 U10161 ( .A(n8519), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8584), .Z(
        P2_U3498) );
  MUX2_X1 U10162 ( .A(n8520), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8584), .Z(
        P2_U3497) );
  MUX2_X1 U10163 ( .A(n8521), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8584), .Z(
        P2_U3496) );
  MUX2_X1 U10164 ( .A(n8522), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8584), .Z(
        P2_U3495) );
  MUX2_X1 U10165 ( .A(n10246), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8584), .Z(
        P2_U3494) );
  MUX2_X1 U10166 ( .A(n8523), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8584), .Z(
        P2_U3493) );
  MUX2_X1 U10167 ( .A(n6687), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8584), .Z(
        P2_U3492) );
  OAI211_X1 U10168 ( .C1(n8526), .C2(n8525), .A(n8524), .B(n10237), .ZN(n8544)
         );
  OAI21_X1 U10169 ( .B1(n8529), .B2(n8528), .A(n8527), .ZN(n8530) );
  NAND2_X1 U10170 ( .A1(n10209), .A2(n8530), .ZN(n8536) );
  OAI21_X1 U10171 ( .B1(n8533), .B2(n8532), .A(n8531), .ZN(n8534) );
  NAND2_X1 U10172 ( .A1(n10117), .A2(n8534), .ZN(n8535) );
  OAI211_X1 U10173 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8537), .A(n8536), .B(
        n8535), .ZN(n8538) );
  INV_X1 U10174 ( .A(n8538), .ZN(n8543) );
  NAND2_X1 U10175 ( .A1(n10219), .A2(n8539), .ZN(n8542) );
  OR2_X1 U10176 ( .A1(n10134), .A2(n8540), .ZN(n8541) );
  NAND4_X1 U10177 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(
        P2_U3184) );
  AOI21_X1 U10178 ( .B1(n9868), .B2(n8546), .A(n8545), .ZN(n8561) );
  OAI21_X1 U10179 ( .B1(n8549), .B2(n8548), .A(n8547), .ZN(n8559) );
  AOI21_X1 U10180 ( .B1(n8551), .B2(n9899), .A(n8550), .ZN(n8557) );
  OAI21_X1 U10181 ( .B1(n10134), .B2(n8553), .A(n8552), .ZN(n8554) );
  AOI21_X1 U10182 ( .B1(n8555), .B2(n10219), .A(n8554), .ZN(n8556) );
  OAI21_X1 U10183 ( .B1(n8557), .B2(n10232), .A(n8556), .ZN(n8558) );
  AOI21_X1 U10184 ( .B1(n10237), .B2(n8559), .A(n8558), .ZN(n8560) );
  OAI21_X1 U10185 ( .B1(n8561), .B2(n10227), .A(n8560), .ZN(P2_U3197) );
  AOI21_X1 U10186 ( .B1(n4450), .B2(n8562), .A(n4414), .ZN(n8577) );
  OAI21_X1 U10187 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8575) );
  NAND2_X1 U10188 ( .A1(n10219), .A2(n8566), .ZN(n8568) );
  OAI211_X1 U10189 ( .C1(n10134), .C2(n7551), .A(n8568), .B(n8567), .ZN(n8574)
         );
  NAND2_X1 U10190 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  AOI21_X1 U10191 ( .B1(n8572), .B2(n8571), .A(n10227), .ZN(n8573) );
  AOI211_X1 U10192 ( .C1(n10237), .C2(n8575), .A(n8574), .B(n8573), .ZN(n8576)
         );
  OAI21_X1 U10193 ( .B1(n8577), .B2(n10232), .A(n8576), .ZN(P2_U3198) );
  AOI21_X1 U10194 ( .B1(n4430), .B2(n8579), .A(n8578), .ZN(n8597) );
  INV_X1 U10195 ( .A(n8580), .ZN(n8582) );
  NAND2_X1 U10196 ( .A1(n8582), .A2(n8581), .ZN(n8586) );
  OAI21_X1 U10197 ( .B1(n8586), .B2(n8584), .A(n8583), .ZN(n8594) );
  INV_X1 U10198 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8589) );
  NAND3_X1 U10199 ( .A1(n8586), .A2(n10237), .A3(n8585), .ZN(n8588) );
  OAI211_X1 U10200 ( .C1(n10134), .C2(n8589), .A(n8588), .B(n8587), .ZN(n8593)
         );
  OAI21_X1 U10201 ( .B1(n8597), .B2(n10232), .A(n8596), .ZN(P2_U3200) );
  AOI21_X1 U10202 ( .B1(n10260), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8599), .ZN(
        n8600) );
  OAI21_X1 U10203 ( .B1(n8773), .B2(n8601), .A(n8600), .ZN(P2_U3202) );
  XNOR2_X1 U10204 ( .A(n8602), .B(n8605), .ZN(n8789) );
  NAND2_X1 U10205 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  XNOR2_X1 U10206 ( .A(n8606), .B(n8605), .ZN(n8612) );
  NAND2_X1 U10207 ( .A1(n8607), .A2(n10247), .ZN(n8610) );
  AOI21_X1 U10208 ( .B1(n8612), .B2(n8684), .A(n8611), .ZN(n8785) );
  MUX2_X1 U10209 ( .A(n8613), .B(n8785), .S(n8714), .Z(n8616) );
  AOI22_X1 U10210 ( .A1(n8786), .A2(n8728), .B1(n10257), .B2(n8614), .ZN(n8615) );
  OAI211_X1 U10211 ( .C1(n8789), .C2(n8731), .A(n8616), .B(n8615), .ZN(
        P2_U3207) );
  INV_X1 U10212 ( .A(n8617), .ZN(n8618) );
  OAI22_X1 U10213 ( .A1(n8619), .A2(n10254), .B1(n8618), .B2(n8711), .ZN(n8620) );
  OAI21_X1 U10214 ( .B1(n8621), .B2(n8620), .A(n8714), .ZN(n8623) );
  NAND2_X1 U10215 ( .A1(n10260), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8622) );
  OAI211_X1 U10216 ( .C1(n8624), .C2(n8731), .A(n8623), .B(n8622), .ZN(
        P2_U3208) );
  NOR2_X1 U10217 ( .A1(n8791), .A2(n10254), .ZN(n8629) );
  XOR2_X1 U10218 ( .A(n8636), .B(n8625), .Z(n8626) );
  OAI222_X1 U10219 ( .A1(n8710), .A2(n8628), .B1(n8719), .B2(n8627), .C1(
        n10252), .C2(n8626), .ZN(n8790) );
  AOI211_X1 U10220 ( .C1(n10257), .C2(n8630), .A(n8629), .B(n8790), .ZN(n8638)
         );
  INV_X1 U10221 ( .A(n8632), .ZN(n8634) );
  OAI21_X1 U10222 ( .B1(n8631), .B2(n8634), .A(n8633), .ZN(n8635) );
  XOR2_X1 U10223 ( .A(n8636), .B(n8635), .Z(n8744) );
  AOI22_X1 U10224 ( .A1(n8744), .A2(n7224), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10260), .ZN(n8637) );
  OAI21_X1 U10225 ( .B1(n8638), .B2(n10260), .A(n8637), .ZN(P2_U3209) );
  XNOR2_X1 U10226 ( .A(n8631), .B(n8639), .ZN(n8798) );
  INV_X1 U10227 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8645) );
  XNOR2_X1 U10228 ( .A(n8640), .B(n8639), .ZN(n8641) );
  OAI222_X1 U10229 ( .A1(n8710), .A2(n8643), .B1(n8719), .B2(n8642), .C1(
        n10252), .C2(n8641), .ZN(n8795) );
  INV_X1 U10230 ( .A(n8795), .ZN(n8644) );
  MUX2_X1 U10231 ( .A(n8645), .B(n8644), .S(n8714), .Z(n8649) );
  AOI22_X1 U10232 ( .A1(n8647), .A2(n8728), .B1(n10257), .B2(n8646), .ZN(n8648) );
  OAI211_X1 U10233 ( .C1(n8798), .C2(n8731), .A(n8649), .B(n8648), .ZN(
        P2_U3210) );
  XNOR2_X1 U10234 ( .A(n8650), .B(n8651), .ZN(n8806) );
  INV_X1 U10235 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8659) );
  OR3_X1 U10236 ( .A1(n8652), .A2(n8654), .A3(n8653), .ZN(n8655) );
  NAND2_X1 U10237 ( .A1(n8656), .A2(n8655), .ZN(n8658) );
  AOI222_X1 U10238 ( .A1(n8684), .A2(n8658), .B1(n8657), .B2(n10247), .C1(
        n8682), .C2(n10248), .ZN(n8801) );
  MUX2_X1 U10239 ( .A(n8659), .B(n8801), .S(n8714), .Z(n8662) );
  AOI22_X1 U10240 ( .A1(n8803), .A2(n8728), .B1(n10257), .B2(n8660), .ZN(n8661) );
  OAI211_X1 U10241 ( .C1(n8806), .C2(n8731), .A(n8662), .B(n8661), .ZN(
        P2_U3211) );
  NAND2_X1 U10242 ( .A1(n8664), .A2(n8663), .ZN(n8665) );
  XOR2_X1 U10243 ( .A(n8668), .B(n8665), .Z(n8812) );
  INV_X1 U10244 ( .A(n8652), .ZN(n8670) );
  NAND3_X1 U10245 ( .A1(n8666), .A2(n8668), .A3(n8667), .ZN(n8669) );
  NAND2_X1 U10246 ( .A1(n8670), .A2(n8669), .ZN(n8673) );
  AOI222_X1 U10247 ( .A1(n8684), .A2(n8673), .B1(n8672), .B2(n10248), .C1(
        n8671), .C2(n10247), .ZN(n8807) );
  MUX2_X1 U10248 ( .A(n8674), .B(n8807), .S(n8714), .Z(n8677) );
  AOI22_X1 U10249 ( .A1(n8809), .A2(n8728), .B1(n10257), .B2(n8675), .ZN(n8676) );
  OAI211_X1 U10250 ( .C1(n8812), .C2(n8731), .A(n8677), .B(n8676), .ZN(
        P2_U3212) );
  XOR2_X1 U10251 ( .A(n8678), .B(n8679), .Z(n8818) );
  INV_X1 U10252 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8685) );
  OAI21_X1 U10253 ( .B1(n8680), .B2(n8679), .A(n8666), .ZN(n8683) );
  AOI222_X1 U10254 ( .A1(n8684), .A2(n8683), .B1(n8682), .B2(n10247), .C1(
        n8681), .C2(n10248), .ZN(n8813) );
  MUX2_X1 U10255 ( .A(n8685), .B(n8813), .S(n8714), .Z(n8688) );
  AOI22_X1 U10256 ( .A1(n8815), .A2(n8728), .B1(n10257), .B2(n8686), .ZN(n8687) );
  OAI211_X1 U10257 ( .C1(n8818), .C2(n8731), .A(n8688), .B(n8687), .ZN(
        P2_U3213) );
  OR2_X1 U10258 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  NAND2_X1 U10259 ( .A1(n8692), .A2(n8691), .ZN(n8822) );
  XNOR2_X1 U10260 ( .A(n8694), .B(n8693), .ZN(n8695) );
  OAI222_X1 U10261 ( .A1(n8710), .A2(n8697), .B1(n8719), .B2(n8696), .C1(n8695), .C2(n10252), .ZN(n8759) );
  NAND2_X1 U10262 ( .A1(n8759), .A2(n8714), .ZN(n8702) );
  OAI22_X1 U10263 ( .A1(n8714), .A2(n8699), .B1(n8698), .B2(n8711), .ZN(n8700)
         );
  AOI21_X1 U10264 ( .B1(n8760), .B2(n8728), .A(n8700), .ZN(n8701) );
  OAI211_X1 U10265 ( .C1(n8822), .C2(n8731), .A(n8702), .B(n8701), .ZN(
        P2_U3214) );
  OAI21_X1 U10266 ( .B1(n8704), .B2(n8705), .A(n8703), .ZN(n8825) );
  XNOR2_X1 U10267 ( .A(n8706), .B(n8705), .ZN(n8707) );
  OAI222_X1 U10268 ( .A1(n8710), .A2(n8709), .B1(n8719), .B2(n8708), .C1(n8707), .C2(n10252), .ZN(n8763) );
  NAND2_X1 U10269 ( .A1(n8763), .A2(n8714), .ZN(n8717) );
  OAI22_X1 U10270 ( .A1(n8714), .A2(n8713), .B1(n8712), .B2(n8711), .ZN(n8715)
         );
  AOI21_X1 U10271 ( .B1(n8764), .B2(n8728), .A(n8715), .ZN(n8716) );
  OAI211_X1 U10272 ( .C1(n8825), .C2(n8731), .A(n8717), .B(n8716), .ZN(
        P2_U3215) );
  XNOR2_X1 U10273 ( .A(n8718), .B(n8722), .ZN(n8833) );
  NOR2_X1 U10274 ( .A1(n8720), .A2(n8719), .ZN(n8724) );
  AOI211_X1 U10275 ( .C1(n8722), .C2(n8721), .A(n10252), .B(n4883), .ZN(n8723)
         );
  AOI211_X1 U10276 ( .C1(n10247), .C2(n8725), .A(n8724), .B(n8723), .ZN(n8826)
         );
  MUX2_X1 U10277 ( .A(n10226), .B(n8826), .S(n8714), .Z(n8730) );
  AOI22_X1 U10278 ( .A1(n8829), .A2(n8728), .B1(n10257), .B2(n8727), .ZN(n8729) );
  OAI211_X1 U10279 ( .C1(n8833), .C2(n8731), .A(n8730), .B(n8729), .ZN(
        P2_U3216) );
  AOI21_X1 U10280 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n6673), .A(n8732), .ZN(
        n8733) );
  OAI21_X1 U10281 ( .B1(n8773), .B2(n8747), .A(n8733), .ZN(P2_U3490) );
  INV_X1 U10282 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10283 ( .A1(n6673), .A2(n8734), .ZN(n8735) );
  NAND2_X1 U10284 ( .A1(n8781), .A2(n8767), .ZN(n8737) );
  OAI211_X1 U10285 ( .C1(n8784), .C2(n8770), .A(n8738), .B(n8737), .ZN(
        P2_U3487) );
  INV_X1 U10286 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U10287 ( .A1(n6673), .A2(n8739), .ZN(n8740) );
  NAND2_X1 U10288 ( .A1(n8786), .A2(n8767), .ZN(n8742) );
  OAI211_X1 U10289 ( .C1(n8770), .C2(n8789), .A(n8743), .B(n8742), .ZN(
        P2_U3485) );
  MUX2_X1 U10290 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8790), .S(n10333), .Z(
        n8746) );
  INV_X1 U10291 ( .A(n8744), .ZN(n8792) );
  OAI22_X1 U10292 ( .A1(n8792), .A2(n8770), .B1(n8791), .B2(n8747), .ZN(n8745)
         );
  OR2_X1 U10293 ( .A1(n8746), .A2(n8745), .ZN(P2_U3483) );
  MUX2_X1 U10294 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8795), .S(n10333), .Z(
        n8749) );
  OAI22_X1 U10295 ( .A1(n8798), .A2(n8770), .B1(n8797), .B2(n8747), .ZN(n8748)
         );
  OR2_X1 U10296 ( .A1(n8749), .A2(n8748), .ZN(P2_U3482) );
  INV_X1 U10297 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8750) );
  MUX2_X1 U10298 ( .A(n8750), .B(n8801), .S(n10333), .Z(n8752) );
  NAND2_X1 U10299 ( .A1(n8803), .A2(n8767), .ZN(n8751) );
  OAI211_X1 U10300 ( .C1(n8806), .C2(n8770), .A(n8752), .B(n8751), .ZN(
        P2_U3481) );
  MUX2_X1 U10301 ( .A(n8753), .B(n8807), .S(n10333), .Z(n8755) );
  NAND2_X1 U10302 ( .A1(n8809), .A2(n8767), .ZN(n8754) );
  OAI211_X1 U10303 ( .C1(n8770), .C2(n8812), .A(n8755), .B(n8754), .ZN(
        P2_U3480) );
  INV_X1 U10304 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8756) );
  MUX2_X1 U10305 ( .A(n8756), .B(n8813), .S(n10333), .Z(n8758) );
  NAND2_X1 U10306 ( .A1(n8815), .A2(n8767), .ZN(n8757) );
  OAI211_X1 U10307 ( .C1(n8818), .C2(n8770), .A(n8758), .B(n8757), .ZN(
        P2_U3479) );
  AOI21_X1 U10308 ( .B1(n10314), .B2(n8760), .A(n8759), .ZN(n8819) );
  MUX2_X1 U10309 ( .A(n8761), .B(n8819), .S(n10333), .Z(n8762) );
  OAI21_X1 U10310 ( .B1(n8770), .B2(n8822), .A(n8762), .ZN(P2_U3478) );
  AOI21_X1 U10311 ( .B1(n10314), .B2(n8764), .A(n8763), .ZN(n8823) );
  MUX2_X1 U10312 ( .A(n8765), .B(n8823), .S(n10333), .Z(n8766) );
  OAI21_X1 U10313 ( .B1(n8770), .B2(n8825), .A(n8766), .ZN(P2_U3477) );
  MUX2_X1 U10314 ( .A(n10231), .B(n8826), .S(n10333), .Z(n8769) );
  NAND2_X1 U10315 ( .A1(n8829), .A2(n8767), .ZN(n8768) );
  OAI211_X1 U10316 ( .C1(n8833), .C2(n8770), .A(n8769), .B(n8768), .ZN(
        P2_U3476) );
  NOR2_X1 U10317 ( .A1(n8771), .A2(n10317), .ZN(n8775) );
  AOI21_X1 U10318 ( .B1(n10317), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8775), .ZN(
        n8772) );
  OAI21_X1 U10319 ( .B1(n8773), .B2(n8796), .A(n8772), .ZN(P2_U3458) );
  INV_X1 U10320 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U10321 ( .A1(n8774), .A2(n8828), .ZN(n8777) );
  INV_X1 U10322 ( .A(n8775), .ZN(n8776) );
  OAI211_X1 U10323 ( .C1(n8778), .C2(n10315), .A(n8777), .B(n8776), .ZN(
        P2_U3457) );
  INV_X1 U10324 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U10325 ( .A1(n8781), .A2(n8828), .ZN(n8782) );
  OAI211_X1 U10326 ( .C1(n8784), .C2(n8832), .A(n8783), .B(n8782), .ZN(
        P2_U3455) );
  MUX2_X1 U10327 ( .A(n9772), .B(n8785), .S(n10315), .Z(n8788) );
  NAND2_X1 U10328 ( .A1(n8786), .A2(n8828), .ZN(n8787) );
  OAI211_X1 U10329 ( .C1(n8789), .C2(n8832), .A(n8788), .B(n8787), .ZN(
        P2_U3453) );
  MUX2_X1 U10330 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8790), .S(n10315), .Z(
        n8794) );
  OAI22_X1 U10331 ( .A1(n8792), .A2(n8832), .B1(n8791), .B2(n8796), .ZN(n8793)
         );
  OR2_X1 U10332 ( .A1(n8794), .A2(n8793), .ZN(P2_U3451) );
  MUX2_X1 U10333 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8795), .S(n10315), .Z(
        n8800) );
  OAI22_X1 U10334 ( .A1(n8798), .A2(n8832), .B1(n8797), .B2(n8796), .ZN(n8799)
         );
  OR2_X1 U10335 ( .A1(n8800), .A2(n8799), .ZN(P2_U3450) );
  INV_X1 U10336 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10337 ( .A(n8802), .B(n8801), .S(n10315), .Z(n8805) );
  NAND2_X1 U10338 ( .A1(n8803), .A2(n8828), .ZN(n8804) );
  OAI211_X1 U10339 ( .C1(n8806), .C2(n8832), .A(n8805), .B(n8804), .ZN(
        P2_U3449) );
  MUX2_X1 U10340 ( .A(n8808), .B(n8807), .S(n10315), .Z(n8811) );
  NAND2_X1 U10341 ( .A1(n8809), .A2(n8828), .ZN(n8810) );
  OAI211_X1 U10342 ( .C1(n8812), .C2(n8832), .A(n8811), .B(n8810), .ZN(
        P2_U3448) );
  INV_X1 U10343 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8814) );
  MUX2_X1 U10344 ( .A(n8814), .B(n8813), .S(n10315), .Z(n8817) );
  NAND2_X1 U10345 ( .A1(n8815), .A2(n8828), .ZN(n8816) );
  OAI211_X1 U10346 ( .C1(n8818), .C2(n8832), .A(n8817), .B(n8816), .ZN(
        P2_U3447) );
  INV_X1 U10347 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8820) );
  MUX2_X1 U10348 ( .A(n8820), .B(n8819), .S(n10315), .Z(n8821) );
  OAI21_X1 U10349 ( .B1(n8822), .B2(n8832), .A(n8821), .ZN(P2_U3446) );
  MUX2_X1 U10350 ( .A(n9761), .B(n8823), .S(n10315), .Z(n8824) );
  OAI21_X1 U10351 ( .B1(n8825), .B2(n8832), .A(n8824), .ZN(P2_U3444) );
  INV_X1 U10352 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8827) );
  MUX2_X1 U10353 ( .A(n8827), .B(n8826), .S(n10315), .Z(n8831) );
  NAND2_X1 U10354 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  OAI211_X1 U10355 ( .C1(n8833), .C2(n8832), .A(n8831), .B(n8830), .ZN(
        P2_U3441) );
  INV_X1 U10356 ( .A(n8836), .ZN(n8840) );
  OAI21_X1 U10357 ( .B1(n8838), .B2(n8840), .A(n8837), .ZN(n8839) );
  OAI21_X1 U10358 ( .B1(n8835), .B2(n8840), .A(n8839), .ZN(n8841) );
  NAND2_X1 U10359 ( .A1(n8841), .A2(n8917), .ZN(n8847) );
  OAI22_X1 U10360 ( .A1(n9550), .A2(n8843), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8842), .ZN(n8845) );
  NOR2_X1 U10361 ( .A1(n8907), .A2(n9542), .ZN(n8844) );
  AOI211_X1 U10362 ( .C1(n8903), .C2(n9195), .A(n8845), .B(n8844), .ZN(n8846)
         );
  OAI211_X1 U10363 ( .C1(n9541), .C2(n8928), .A(n8847), .B(n8846), .ZN(
        P1_U3219) );
  NAND2_X1 U10364 ( .A1(n8848), .A2(n8882), .ZN(n8881) );
  NAND2_X1 U10365 ( .A1(n8881), .A2(n8849), .ZN(n8850) );
  XOR2_X1 U10366 ( .A(n8851), .B(n8850), .Z(n8857) );
  OAI22_X1 U10367 ( .A1(n9550), .A2(n8921), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8852), .ZN(n8853) );
  AOI21_X1 U10368 ( .B1(n8919), .B2(n9512), .A(n8853), .ZN(n8854) );
  OAI21_X1 U10369 ( .B1(n9504), .B2(n8907), .A(n8854), .ZN(n8855) );
  AOI21_X1 U10370 ( .B1(n9597), .B2(n8909), .A(n8855), .ZN(n8856) );
  OAI21_X1 U10371 ( .B1(n8857), .B2(n8912), .A(n8856), .ZN(P1_U3223) );
  OAI21_X1 U10372 ( .B1(n8860), .B2(n8858), .A(n8859), .ZN(n8861) );
  NAND2_X1 U10373 ( .A1(n8861), .A2(n8917), .ZN(n8867) );
  NAND2_X1 U10374 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9336) );
  OAI21_X1 U10375 ( .B1(n8863), .B2(n8862), .A(n9336), .ZN(n8864) );
  AOI21_X1 U10376 ( .B1(n8865), .B2(n8924), .A(n8864), .ZN(n8866) );
  OAI211_X1 U10377 ( .C1(n8868), .C2(n8928), .A(n8867), .B(n8866), .ZN(
        P1_U3226) );
  NAND2_X1 U10378 ( .A1(n8871), .A2(n8870), .ZN(n8872) );
  XNOR2_X1 U10379 ( .A(n8869), .B(n8872), .ZN(n8880) );
  NOR2_X1 U10380 ( .A1(n8873), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9356) );
  AOI21_X1 U10381 ( .B1(n8919), .B2(n9195), .A(n9356), .ZN(n8876) );
  NAND2_X1 U10382 ( .A1(n8924), .A2(n8874), .ZN(n8875) );
  OAI211_X1 U10383 ( .C1(n8877), .C2(n8921), .A(n8876), .B(n8875), .ZN(n8878)
         );
  AOI21_X1 U10384 ( .B1(n9619), .B2(n8909), .A(n8878), .ZN(n8879) );
  OAI21_X1 U10385 ( .B1(n8880), .B2(n8912), .A(n8879), .ZN(P1_U3228) );
  OAI21_X1 U10386 ( .B1(n8882), .B2(n8848), .A(n8881), .ZN(n8883) );
  NAND2_X1 U10387 ( .A1(n8883), .A2(n8917), .ZN(n8889) );
  INV_X1 U10388 ( .A(n8884), .ZN(n9531) );
  AOI22_X1 U10389 ( .A1(n9524), .A2(n8919), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8885) );
  OAI21_X1 U10390 ( .B1(n8886), .B2(n8921), .A(n8885), .ZN(n8887) );
  AOI21_X1 U10391 ( .B1(n9531), .B2(n8924), .A(n8887), .ZN(n8888) );
  OAI211_X1 U10392 ( .C1(n9931), .C2(n8928), .A(n8889), .B(n8888), .ZN(
        P1_U3233) );
  OAI21_X1 U10393 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n8893) );
  NAND2_X1 U10394 ( .A1(n8893), .A2(n8917), .ZN(n8898) );
  AOI22_X1 U10395 ( .A1(n9489), .A2(n8919), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8894) );
  OAI21_X1 U10396 ( .B1(n8895), .B2(n8921), .A(n8894), .ZN(n8896) );
  AOI21_X1 U10397 ( .B1(n9495), .B2(n8924), .A(n8896), .ZN(n8897) );
  OAI211_X1 U10398 ( .C1(n4571), .C2(n8928), .A(n8898), .B(n8897), .ZN(
        P1_U3235) );
  XNOR2_X1 U10399 ( .A(n8901), .B(n8900), .ZN(n8902) );
  XNOR2_X1 U10400 ( .A(n8899), .B(n8902), .ZN(n8913) );
  AOI22_X1 U10401 ( .A1(n8903), .A2(n9196), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8905) );
  NAND2_X1 U10402 ( .A1(n8919), .A2(n9523), .ZN(n8904) );
  OAI211_X1 U10403 ( .C1(n8907), .C2(n8906), .A(n8905), .B(n8904), .ZN(n8908)
         );
  AOI21_X1 U10404 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8911) );
  OAI21_X1 U10405 ( .B1(n8913), .B2(n8912), .A(n8911), .ZN(P1_U3238) );
  OAI21_X1 U10406 ( .B1(n8914), .B2(n8916), .A(n8915), .ZN(n8918) );
  NAND2_X1 U10407 ( .A1(n8918), .A2(n8917), .ZN(n8927) );
  NOR2_X1 U10408 ( .A1(n9733), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9323) );
  AOI21_X1 U10409 ( .B1(n8919), .B2(n9197), .A(n9323), .ZN(n8920) );
  OAI21_X1 U10410 ( .B1(n8922), .B2(n8921), .A(n8920), .ZN(n8923) );
  AOI21_X1 U10411 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8926) );
  OAI211_X1 U10412 ( .C1(n8929), .C2(n8928), .A(n8927), .B(n8926), .ZN(
        P1_U3241) );
  AOI211_X1 U10413 ( .C1(n9182), .C2(n5401), .A(n5653), .B(n8930), .ZN(n9188)
         );
  INV_X1 U10414 ( .A(n9125), .ZN(n9044) );
  INV_X1 U10415 ( .A(n8932), .ZN(n8989) );
  NAND2_X1 U10416 ( .A1(n9002), .A2(n8989), .ZN(n8933) );
  NAND2_X1 U10417 ( .A1(n8933), .A2(n9003), .ZN(n9085) );
  NAND2_X1 U10418 ( .A1(n8977), .A2(n8934), .ZN(n9163) );
  INV_X1 U10419 ( .A(n8935), .ZN(n9133) );
  AOI211_X1 U10420 ( .C1(n7174), .C2(n9135), .A(n9133), .B(n8936), .ZN(n8938)
         );
  INV_X1 U10421 ( .A(n9134), .ZN(n8937) );
  INV_X1 U10422 ( .A(n8940), .ZN(n9138) );
  NOR3_X1 U10423 ( .A1(n8938), .A2(n8937), .A3(n9138), .ZN(n8942) );
  INV_X1 U10424 ( .A(n8946), .ZN(n8939) );
  MUX2_X1 U10425 ( .A(n8942), .B(n8941), .S(n9125), .Z(n8948) );
  NOR2_X1 U10426 ( .A1(n8943), .A2(n9044), .ZN(n8944) );
  NAND2_X1 U10427 ( .A1(n8946), .A2(n8945), .ZN(n9142) );
  INV_X1 U10428 ( .A(n8950), .ZN(n8953) );
  NAND2_X1 U10429 ( .A1(n8951), .A2(n8955), .ZN(n8952) );
  MUX2_X1 U10430 ( .A(n8953), .B(n8952), .S(n9125), .Z(n8954) );
  AOI21_X1 U10431 ( .B1(n8956), .B2(n8955), .A(n8954), .ZN(n8961) );
  NAND2_X1 U10432 ( .A1(n8962), .A2(n8957), .ZN(n8958) );
  MUX2_X1 U10433 ( .A(n8959), .B(n8958), .S(n9125), .Z(n8960) );
  NOR2_X1 U10434 ( .A1(n8961), .A2(n8960), .ZN(n8970) );
  INV_X1 U10435 ( .A(n8962), .ZN(n8963) );
  OAI21_X1 U10436 ( .B1(n8970), .B2(n8963), .A(n9146), .ZN(n8964) );
  NAND3_X1 U10437 ( .A1(n8964), .A2(n9151), .A3(n9153), .ZN(n8966) );
  OR2_X1 U10438 ( .A1(n10008), .A2(n8965), .ZN(n9149) );
  NAND2_X1 U10439 ( .A1(n8966), .A2(n4923), .ZN(n8967) );
  INV_X1 U10440 ( .A(n8968), .ZN(n8969) );
  OAI21_X1 U10441 ( .B1(n8970), .B2(n8969), .A(n9151), .ZN(n8971) );
  NAND3_X1 U10442 ( .A1(n8971), .A2(n9146), .A3(n9149), .ZN(n8972) );
  NAND2_X1 U10443 ( .A1(n8972), .A2(n4922), .ZN(n8973) );
  XNOR2_X1 U10444 ( .A(n9969), .B(n9199), .ZN(n9978) );
  INV_X1 U10445 ( .A(n9159), .ZN(n8974) );
  MUX2_X1 U10446 ( .A(n8975), .B(n8974), .S(n9125), .Z(n8976) );
  AOI21_X1 U10447 ( .B1(n9125), .B2(n9162), .A(n9062), .ZN(n8981) );
  INV_X1 U10448 ( .A(n9162), .ZN(n8979) );
  INV_X1 U10449 ( .A(n9160), .ZN(n8978) );
  OAI211_X1 U10450 ( .C1(n8979), .C2(n8978), .A(n9044), .B(n8977), .ZN(n8980)
         );
  OAI21_X1 U10451 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n8986) );
  NAND2_X1 U10452 ( .A1(n8987), .A2(n9165), .ZN(n8984) );
  INV_X1 U10453 ( .A(n9169), .ZN(n8983) );
  MUX2_X1 U10454 ( .A(n8984), .B(n8983), .S(n9125), .Z(n8985) );
  AOI21_X1 U10455 ( .B1(n8986), .B2(n9063), .A(n8985), .ZN(n8996) );
  NAND2_X1 U10456 ( .A1(n9170), .A2(n8987), .ZN(n9166) );
  AOI21_X1 U10457 ( .B1(n8996), .B2(n8994), .A(n9166), .ZN(n8988) );
  NOR4_X1 U10458 ( .A1(n8988), .A2(n4839), .A3(n4835), .A4(n9044), .ZN(n8993)
         );
  INV_X1 U10459 ( .A(n9002), .ZN(n8992) );
  NOR2_X1 U10460 ( .A1(n8989), .A2(n9125), .ZN(n8998) );
  OAI21_X1 U10461 ( .B1(n8989), .B2(n9608), .A(n9044), .ZN(n8990) );
  AOI22_X1 U10462 ( .A1(n8998), .A2(n9523), .B1(n8990), .B2(n9001), .ZN(n8991)
         );
  NOR3_X1 U10463 ( .A1(n8993), .A2(n8992), .A3(n8991), .ZN(n9000) );
  NAND2_X1 U10464 ( .A1(n8995), .A2(n8994), .ZN(n9172) );
  OAI211_X1 U10465 ( .C1(n8996), .C2(n9172), .A(n9044), .B(n9170), .ZN(n8997)
         );
  MUX2_X1 U10466 ( .A(n8998), .B(n8997), .S(n9171), .Z(n8999) );
  NAND2_X1 U10467 ( .A1(n9000), .A2(n8999), .ZN(n9006) );
  NAND2_X1 U10468 ( .A1(n9002), .A2(n9001), .ZN(n9096) );
  INV_X1 U10469 ( .A(n9003), .ZN(n9004) );
  NAND2_X1 U10470 ( .A1(n9452), .A2(n9007), .ZN(n9084) );
  OR2_X1 U10471 ( .A1(n9494), .A2(n9008), .ZN(n9009) );
  NAND2_X1 U10472 ( .A1(n9010), .A2(n9009), .ZN(n9080) );
  MUX2_X1 U10473 ( .A(n9084), .B(n9080), .S(n9125), .Z(n9013) );
  INV_X1 U10474 ( .A(n9454), .ZN(n9012) );
  MUX2_X1 U10475 ( .A(n9010), .B(n9452), .S(n9125), .Z(n9011) );
  MUX2_X1 U10476 ( .A(n9088), .B(n9081), .S(n9125), .Z(n9014) );
  OAI211_X1 U10477 ( .C1(n9023), .C2(n9420), .A(n9045), .B(n9094), .ZN(n9016)
         );
  INV_X1 U10478 ( .A(n9079), .ZN(n9018) );
  NOR2_X1 U10479 ( .A1(n9018), .A2(n9125), .ZN(n9019) );
  INV_X1 U10480 ( .A(n9045), .ZN(n9022) );
  INV_X1 U10481 ( .A(n9420), .ZN(n9021) );
  NOR3_X1 U10482 ( .A1(n9414), .A2(n9125), .A3(n9193), .ZN(n9032) );
  NAND2_X1 U10483 ( .A1(n9193), .A2(n9125), .ZN(n9028) );
  NAND3_X1 U10484 ( .A1(n9025), .A2(n9125), .A3(n9427), .ZN(n9027) );
  AOI21_X1 U10485 ( .B1(n9028), .B2(n9027), .A(n9026), .ZN(n9031) );
  NOR3_X1 U10486 ( .A1(n9564), .A2(n9029), .A3(n9028), .ZN(n9030) );
  NOR3_X1 U10487 ( .A1(n9032), .A2(n9031), .A3(n9030), .ZN(n9033) );
  NOR2_X1 U10488 ( .A1(n9075), .A2(n9035), .ZN(n9112) );
  NOR3_X1 U10489 ( .A1(n9182), .A2(n9112), .A3(n9405), .ZN(n9037) );
  AOI211_X1 U10490 ( .C1(n9125), .C2(n9632), .A(n9075), .B(n9036), .ZN(n9041)
         );
  OAI21_X1 U10491 ( .B1(n9044), .B2(n9110), .A(n9405), .ZN(n9040) );
  AOI211_X1 U10492 ( .C1(n9632), .C2(n9110), .A(n9112), .B(n9044), .ZN(n9038)
         );
  AOI211_X1 U10493 ( .C1(n9041), .C2(n9040), .A(n9039), .B(n9038), .ZN(n9042)
         );
  NAND2_X1 U10494 ( .A1(n9043), .A2(n9042), .ZN(n9077) );
  OAI21_X1 U10495 ( .B1(n9183), .B2(n9044), .A(n9077), .ZN(n9187) );
  OR2_X1 U10496 ( .A1(n9420), .A2(n9022), .ZN(n9437) );
  INV_X1 U10497 ( .A(n9437), .ZN(n9439) );
  INV_X1 U10498 ( .A(n9046), .ZN(n9999) );
  INV_X1 U10499 ( .A(n9147), .ZN(n9057) );
  INV_X1 U10500 ( .A(n9047), .ZN(n9048) );
  NAND4_X1 U10501 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9132), .ZN(n9053)
         );
  NOR4_X1 U10502 ( .A1(n9053), .A2(n5607), .A3(n9052), .A4(n9051), .ZN(n9055)
         );
  NAND4_X1 U10503 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9058)
         );
  NOR4_X1 U10504 ( .A1(n9060), .A2(n9999), .A3(n9059), .A4(n9058), .ZN(n9061)
         );
  NAND4_X1 U10505 ( .A1(n9063), .A2(n9062), .A3(n9061), .A4(n9978), .ZN(n9064)
         );
  NOR3_X1 U10506 ( .A1(n9066), .A2(n9065), .A3(n9064), .ZN(n9067) );
  NAND4_X1 U10507 ( .A1(n9510), .A2(n9521), .A3(n9546), .A4(n9067), .ZN(n9068)
         );
  NOR4_X1 U10508 ( .A1(n9454), .A2(n9484), .A3(n9473), .A4(n9068), .ZN(n9069)
         );
  NAND4_X1 U10509 ( .A1(n9421), .A2(n9070), .A3(n9439), .A4(n9069), .ZN(n9071)
         );
  NOR4_X1 U10510 ( .A1(n9182), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n9118)
         );
  NOR2_X1 U10511 ( .A1(n9632), .A2(n9074), .ZN(n9109) );
  NOR2_X1 U10512 ( .A1(n9405), .A2(n9075), .ZN(n9180) );
  NOR2_X1 U10513 ( .A1(n9109), .A2(n9180), .ZN(n9119) );
  NAND3_X1 U10514 ( .A1(n9118), .A2(n9119), .A3(n9183), .ZN(n9076) );
  OAI21_X1 U10515 ( .B1(n9077), .B2(n9132), .A(n9076), .ZN(n9129) );
  NAND2_X1 U10516 ( .A1(n9079), .A2(n9078), .ZN(n9099) );
  NAND3_X1 U10517 ( .A1(n9088), .A2(n9452), .A3(n9080), .ZN(n9082) );
  NAND2_X1 U10518 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  NOR2_X1 U10519 ( .A1(n9420), .A2(n9083), .ZN(n9098) );
  INV_X1 U10520 ( .A(n9084), .ZN(n9087) );
  INV_X1 U10521 ( .A(n9085), .ZN(n9086) );
  NAND3_X1 U10522 ( .A1(n9088), .A2(n9087), .A3(n9086), .ZN(n9089) );
  AOI21_X1 U10523 ( .B1(n9098), .B2(n9089), .A(n9022), .ZN(n9090) );
  OR2_X1 U10524 ( .A1(n9099), .A2(n9090), .ZN(n9093) );
  NAND3_X1 U10525 ( .A1(n9093), .A2(n9092), .A3(n9091), .ZN(n9102) );
  INV_X1 U10526 ( .A(n9094), .ZN(n9095) );
  NOR2_X1 U10527 ( .A1(n9102), .A2(n9095), .ZN(n9176) );
  INV_X1 U10528 ( .A(n9176), .ZN(n9106) );
  INV_X1 U10529 ( .A(n9096), .ZN(n9097) );
  NAND2_X1 U10530 ( .A1(n9098), .A2(n9097), .ZN(n9105) );
  INV_X1 U10531 ( .A(n9099), .ZN(n9103) );
  OAI211_X1 U10532 ( .C1(n9103), .C2(n9102), .A(n9101), .B(n9100), .ZN(n9104)
         );
  AOI21_X1 U10533 ( .B1(n9176), .B2(n9105), .A(n9104), .ZN(n9179) );
  OAI21_X1 U10534 ( .B1(n9106), .B2(n9520), .A(n9179), .ZN(n9107) );
  OAI21_X1 U10535 ( .B1(n9632), .B2(n9108), .A(n9107), .ZN(n9114) );
  INV_X1 U10536 ( .A(n9109), .ZN(n9111) );
  NAND2_X1 U10537 ( .A1(n9111), .A2(n9110), .ZN(n9177) );
  INV_X1 U10538 ( .A(n9112), .ZN(n9113) );
  OAI22_X1 U10539 ( .A1(n9114), .A2(n9177), .B1(n9405), .B2(n9113), .ZN(n9117)
         );
  INV_X1 U10540 ( .A(n9182), .ZN(n9116) );
  AOI21_X1 U10541 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9123) );
  INV_X1 U10542 ( .A(n9118), .ZN(n9121) );
  INV_X1 U10543 ( .A(n9119), .ZN(n9120) );
  NOR2_X1 U10544 ( .A1(n9121), .A2(n9120), .ZN(n9122) );
  OAI21_X1 U10545 ( .B1(n9123), .B2(n9122), .A(n9183), .ZN(n9124) );
  NAND2_X1 U10546 ( .A1(n9124), .A2(n5654), .ZN(n9127) );
  NAND2_X1 U10547 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  INV_X1 U10548 ( .A(n9130), .ZN(n9131) );
  AOI211_X1 U10549 ( .C1(n10062), .C2(n9211), .A(n9132), .B(n9131), .ZN(n9137)
         );
  OR2_X1 U10550 ( .A1(n7174), .A2(n9133), .ZN(n9136) );
  OAI211_X1 U10551 ( .C1(n9137), .C2(n9136), .A(n9135), .B(n9134), .ZN(n9140)
         );
  AOI21_X1 U10552 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9143) );
  OAI21_X1 U10553 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9144) );
  INV_X1 U10554 ( .A(n9144), .ZN(n9148) );
  OAI211_X1 U10555 ( .C1(n9148), .C2(n9147), .A(n9146), .B(n9145), .ZN(n9152)
         );
  INV_X1 U10556 ( .A(n9149), .ZN(n9150) );
  AOI21_X1 U10557 ( .B1(n9152), .B2(n9151), .A(n9150), .ZN(n9156) );
  INV_X1 U10558 ( .A(n9153), .ZN(n9155) );
  OAI21_X1 U10559 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9158) );
  NAND3_X1 U10560 ( .A1(n9158), .A2(n9976), .A3(n9157), .ZN(n9161) );
  AND3_X1 U10561 ( .A1(n9161), .A2(n9160), .A3(n9159), .ZN(n9164) );
  OAI21_X1 U10562 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9168) );
  INV_X1 U10563 ( .A(n9165), .ZN(n9167) );
  AOI211_X1 U10564 ( .C1(n9169), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9173)
         );
  OAI211_X1 U10565 ( .C1(n9173), .C2(n9172), .A(n9171), .B(n9170), .ZN(n9174)
         );
  NAND3_X1 U10566 ( .A1(n9176), .A2(n9175), .A3(n9174), .ZN(n9178) );
  AOI21_X1 U10567 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9181) );
  NOR2_X1 U10568 ( .A1(n9181), .A2(n9180), .ZN(n9184) );
  AOI21_X1 U10569 ( .B1(n9184), .B2(n9183), .A(n9182), .ZN(n9185) );
  XNOR2_X1 U10570 ( .A(n9185), .B(n5401), .ZN(n9186) );
  OAI21_X1 U10571 ( .B1(n9191), .B2(n5653), .A(P1_B_REG_SCAN_IN), .ZN(n9190)
         );
  MUX2_X1 U10572 ( .A(n9192), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9210), .Z(
        P1_U3583) );
  MUX2_X1 U10573 ( .A(n9193), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9210), .Z(
        P1_U3582) );
  MUX2_X1 U10574 ( .A(n9427), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9210), .Z(
        P1_U3581) );
  MUX2_X1 U10575 ( .A(n9458), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9210), .Z(
        P1_U3579) );
  MUX2_X1 U10576 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9194), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10577 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9489), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10578 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9512), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10579 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9524), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10580 ( .A(n9511), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9210), .Z(
        P1_U3574) );
  MUX2_X1 U10581 ( .A(n9523), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9210), .Z(
        P1_U3573) );
  MUX2_X1 U10582 ( .A(n9195), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9210), .Z(
        P1_U3572) );
  MUX2_X1 U10583 ( .A(n9196), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9210), .Z(
        P1_U3571) );
  MUX2_X1 U10584 ( .A(n9197), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9210), .Z(
        P1_U3570) );
  MUX2_X1 U10585 ( .A(n9198), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9210), .Z(
        P1_U3569) );
  MUX2_X1 U10586 ( .A(n9983), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9210), .Z(
        P1_U3568) );
  MUX2_X1 U10587 ( .A(n9199), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9210), .Z(
        P1_U3567) );
  MUX2_X1 U10588 ( .A(n9984), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9210), .Z(
        P1_U3566) );
  MUX2_X1 U10589 ( .A(n9200), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9210), .Z(
        P1_U3565) );
  MUX2_X1 U10590 ( .A(n9201), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9210), .Z(
        P1_U3564) );
  MUX2_X1 U10591 ( .A(n9202), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9210), .Z(
        P1_U3563) );
  MUX2_X1 U10592 ( .A(n9203), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9210), .Z(
        P1_U3562) );
  MUX2_X1 U10593 ( .A(n9204), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9210), .Z(
        P1_U3561) );
  MUX2_X1 U10594 ( .A(n9205), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9210), .Z(
        P1_U3560) );
  MUX2_X1 U10595 ( .A(n9206), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9210), .Z(
        P1_U3559) );
  MUX2_X1 U10596 ( .A(n9207), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9210), .Z(
        P1_U3558) );
  MUX2_X1 U10597 ( .A(n9208), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9210), .Z(
        P1_U3557) );
  MUX2_X1 U10598 ( .A(n9209), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9210), .Z(
        P1_U3556) );
  MUX2_X1 U10599 ( .A(n9211), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9210), .Z(
        P1_U3555) );
  INV_X1 U10600 ( .A(n9956), .ZN(n9355) );
  OAI22_X1 U10601 ( .A1(n9337), .A2(n9212), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9890), .ZN(n9213) );
  AOI21_X1 U10602 ( .B1(n9355), .B2(n9214), .A(n9213), .ZN(n9226) );
  OAI211_X1 U10603 ( .C1(n9217), .C2(n9216), .A(n9397), .B(n9215), .ZN(n9225)
         );
  NOR2_X1 U10604 ( .A1(n9218), .A2(n9945), .ZN(n9223) );
  MUX2_X1 U10605 ( .A(n9220), .B(P1_REG1_REG_1__SCAN_IN), .S(n9219), .Z(n9222)
         );
  OAI211_X1 U10606 ( .C1(n9223), .C2(n9222), .A(n9961), .B(n9221), .ZN(n9224)
         );
  NAND3_X1 U10607 ( .A1(n9226), .A2(n9225), .A3(n9224), .ZN(P1_U3244) );
  AND2_X1 U10608 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9229) );
  NOR2_X1 U10609 ( .A1(n9956), .A2(n9227), .ZN(n9228) );
  AOI211_X1 U10610 ( .C1(n9950), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9229), .B(
        n9228), .ZN(n9239) );
  AOI211_X1 U10611 ( .C1(n9232), .C2(n9231), .A(n9230), .B(n9958), .ZN(n9233)
         );
  INV_X1 U10612 ( .A(n9233), .ZN(n9238) );
  OAI211_X1 U10613 ( .C1(n9236), .C2(n9235), .A(n9961), .B(n9234), .ZN(n9237)
         );
  NAND3_X1 U10614 ( .A1(n9239), .A2(n9238), .A3(n9237), .ZN(P1_U3246) );
  NOR2_X1 U10615 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5235), .ZN(n9242) );
  NOR2_X1 U10616 ( .A1(n9956), .A2(n9240), .ZN(n9241) );
  AOI211_X1 U10617 ( .C1(n9950), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9242), .B(
        n9241), .ZN(n9252) );
  AOI211_X1 U10618 ( .C1(n9245), .C2(n9244), .A(n9243), .B(n9958), .ZN(n9246)
         );
  INV_X1 U10619 ( .A(n9246), .ZN(n9251) );
  OAI211_X1 U10620 ( .C1(n9249), .C2(n9248), .A(n9961), .B(n9247), .ZN(n9250)
         );
  NAND3_X1 U10621 ( .A1(n9252), .A2(n9251), .A3(n9250), .ZN(P1_U3249) );
  NOR2_X1 U10622 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9253), .ZN(n9256) );
  NOR2_X1 U10623 ( .A1(n9956), .A2(n9254), .ZN(n9255) );
  AOI211_X1 U10624 ( .C1(n9950), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n9256), .B(
        n9255), .ZN(n9266) );
  AOI211_X1 U10625 ( .C1(n9259), .C2(n9258), .A(n9257), .B(n9958), .ZN(n9260)
         );
  INV_X1 U10626 ( .A(n9260), .ZN(n9265) );
  OAI211_X1 U10627 ( .C1(n9263), .C2(n9262), .A(n9961), .B(n9261), .ZN(n9264)
         );
  NAND3_X1 U10628 ( .A1(n9266), .A2(n9265), .A3(n9264), .ZN(P1_U3250) );
  NOR2_X1 U10629 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5207), .ZN(n9269) );
  NOR2_X1 U10630 ( .A1(n9956), .A2(n9267), .ZN(n9268) );
  AOI211_X1 U10631 ( .C1(n9950), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9269), .B(
        n9268), .ZN(n9279) );
  AOI211_X1 U10632 ( .C1(n9272), .C2(n9271), .A(n9270), .B(n9958), .ZN(n9273)
         );
  INV_X1 U10633 ( .A(n9273), .ZN(n9278) );
  OAI211_X1 U10634 ( .C1(n9276), .C2(n9275), .A(n9961), .B(n9274), .ZN(n9277)
         );
  NAND3_X1 U10635 ( .A1(n9279), .A2(n9278), .A3(n9277), .ZN(P1_U3251) );
  NOR2_X1 U10636 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9280), .ZN(n9283) );
  NOR2_X1 U10637 ( .A1(n9956), .A2(n9281), .ZN(n9282) );
  AOI211_X1 U10638 ( .C1(n9950), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9283), .B(
        n9282), .ZN(n9293) );
  OAI211_X1 U10639 ( .C1(n9286), .C2(n9285), .A(n9961), .B(n9284), .ZN(n9292)
         );
  AOI211_X1 U10640 ( .C1(n9289), .C2(n9288), .A(n9287), .B(n9958), .ZN(n9290)
         );
  INV_X1 U10641 ( .A(n9290), .ZN(n9291) );
  NAND3_X1 U10642 ( .A1(n9293), .A2(n9292), .A3(n9291), .ZN(P1_U3254) );
  NOR2_X1 U10643 ( .A1(n9956), .A2(n9316), .ZN(n9294) );
  AOI211_X1 U10644 ( .C1(n9950), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9295), .B(
        n9294), .ZN(n9310) );
  NOR2_X1 U10645 ( .A1(n9316), .A2(n9312), .ZN(n9296) );
  AOI21_X1 U10646 ( .B1(n9312), .B2(n9316), .A(n9296), .ZN(n9300) );
  OAI21_X1 U10647 ( .B1(n10111), .B2(n9298), .A(n9297), .ZN(n9299) );
  NAND2_X1 U10648 ( .A1(n9300), .A2(n9299), .ZN(n9311) );
  OAI211_X1 U10649 ( .C1(n9300), .C2(n9299), .A(n9961), .B(n9311), .ZN(n9309)
         );
  NAND2_X1 U10650 ( .A1(n9304), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9303) );
  OAI21_X1 U10651 ( .B1(n9304), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9303), .ZN(
        n9305) );
  AOI211_X1 U10652 ( .C1(n9306), .C2(n9305), .A(n9313), .B(n9958), .ZN(n9307)
         );
  INV_X1 U10653 ( .A(n9307), .ZN(n9308) );
  NAND3_X1 U10654 ( .A1(n9310), .A2(n9309), .A3(n9308), .ZN(P1_U3257) );
  INV_X1 U10655 ( .A(n9328), .ZN(n9326) );
  OAI21_X1 U10656 ( .B1(n9316), .B2(n9312), .A(n9311), .ZN(n9329) );
  XNOR2_X1 U10657 ( .A(n9329), .B(n9326), .ZN(n9327) );
  XOR2_X1 U10658 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9327), .Z(n9322) );
  INV_X1 U10659 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9320) );
  INV_X1 U10660 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9315) );
  OAI21_X1 U10661 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9318) );
  AND2_X1 U10662 ( .A1(n9318), .A2(n9328), .ZN(n9340) );
  INV_X1 U10663 ( .A(n9340), .ZN(n9317) );
  OAI21_X1 U10664 ( .B1(n9328), .B2(n9318), .A(n9317), .ZN(n9319) );
  NOR2_X1 U10665 ( .A1(n9320), .A2(n9319), .ZN(n9339) );
  AOI211_X1 U10666 ( .C1(n9320), .C2(n9319), .A(n9339), .B(n9958), .ZN(n9321)
         );
  AOI21_X1 U10667 ( .B1(n9961), .B2(n9322), .A(n9321), .ZN(n9325) );
  AOI21_X1 U10668 ( .B1(n9950), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9323), .ZN(
        n9324) );
  OAI211_X1 U10669 ( .C1(n9326), .C2(n9956), .A(n9325), .B(n9324), .ZN(
        P1_U3258) );
  NAND2_X1 U10670 ( .A1(n9327), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U10671 ( .A1(n9329), .A2(n9328), .ZN(n9330) );
  NAND2_X1 U10672 ( .A1(n9331), .A2(n9330), .ZN(n9335) );
  OR2_X1 U10673 ( .A1(n9350), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U10674 ( .A1(n9350), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U10675 ( .A1(n9358), .A2(n9332), .ZN(n9334) );
  INV_X1 U10676 ( .A(n9359), .ZN(n9333) );
  AOI21_X1 U10677 ( .B1(n9335), .B2(n9334), .A(n9333), .ZN(n9347) );
  OAI21_X1 U10678 ( .B1(n9337), .B2(n9758), .A(n9336), .ZN(n9338) );
  AOI21_X1 U10679 ( .B1(n9355), .B2(n9350), .A(n9338), .ZN(n9346) );
  INV_X1 U10680 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9341) );
  OR2_X1 U10681 ( .A1(n9350), .A2(n9341), .ZN(n9343) );
  NAND2_X1 U10682 ( .A1(n9350), .A2(n9341), .ZN(n9342) );
  NAND2_X1 U10683 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  NAND2_X1 U10684 ( .A1(n9344), .A2(n4910), .ZN(n9352) );
  OAI211_X1 U10685 ( .C1(n4910), .C2(n9344), .A(n9397), .B(n9352), .ZN(n9345)
         );
  OAI211_X1 U10686 ( .C1(n9348), .C2(n9347), .A(n9346), .B(n9345), .ZN(
        P1_U3259) );
  OR2_X1 U10687 ( .A1(n9367), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U10688 ( .A1(n9367), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9349) );
  AND2_X1 U10689 ( .A1(n9375), .A2(n9349), .ZN(n9353) );
  NAND2_X1 U10690 ( .A1(n9350), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U10691 ( .A1(n9397), .A2(n9354), .ZN(n9366) );
  NAND2_X1 U10692 ( .A1(n9355), .A2(n9367), .ZN(n9365) );
  AOI21_X1 U10693 ( .B1(n9950), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9356), .ZN(
        n9364) );
  INV_X1 U10694 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9357) );
  XNOR2_X1 U10695 ( .A(n9367), .B(n9357), .ZN(n9361) );
  NAND2_X1 U10696 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  NAND2_X1 U10697 ( .A1(n9360), .A2(n9361), .ZN(n9371) );
  OAI21_X1 U10698 ( .B1(n9361), .B2(n9360), .A(n9371), .ZN(n9362) );
  NAND2_X1 U10699 ( .A1(n9961), .A2(n9362), .ZN(n9363) );
  NAND4_X1 U10700 ( .A1(n9366), .A2(n9365), .A3(n9364), .A4(n9363), .ZN(
        P1_U3260) );
  OR2_X1 U10701 ( .A1(n9367), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9368) );
  INV_X1 U10702 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9614) );
  XNOR2_X1 U10703 ( .A(n9389), .B(n9614), .ZN(n9369) );
  AOI21_X1 U10704 ( .B1(n9371), .B2(n9368), .A(n9369), .ZN(n9385) );
  AND2_X1 U10705 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U10706 ( .A1(n9371), .A2(n9370), .ZN(n9391) );
  NAND2_X1 U10707 ( .A1(n9961), .A2(n9391), .ZN(n9384) );
  AND2_X1 U10708 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9374) );
  INV_X1 U10709 ( .A(n9389), .ZN(n9372) );
  NOR2_X1 U10710 ( .A1(n9956), .A2(n9372), .ZN(n9373) );
  AOI211_X1 U10711 ( .C1(n9950), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9374), .B(
        n9373), .ZN(n9383) );
  OR2_X1 U10712 ( .A1(n9389), .A2(n9377), .ZN(n9379) );
  NAND2_X1 U10713 ( .A1(n9389), .A2(n9377), .ZN(n9378) );
  NAND2_X1 U10714 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  NAND2_X1 U10715 ( .A1(n9381), .A2(n9380), .ZN(n9387) );
  OAI211_X1 U10716 ( .C1(n9381), .C2(n9380), .A(n9397), .B(n9387), .ZN(n9382)
         );
  OAI211_X1 U10717 ( .C1(n9385), .C2(n9384), .A(n9383), .B(n9382), .ZN(
        P1_U3261) );
  NAND2_X1 U10718 ( .A1(n9389), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U10719 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  XNOR2_X1 U10720 ( .A(n9388), .B(n9879), .ZN(n9396) );
  NAND2_X1 U10721 ( .A1(n9389), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U10722 ( .A1(n9391), .A2(n9390), .ZN(n9393) );
  INV_X1 U10723 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9392) );
  XNOR2_X1 U10724 ( .A(n9393), .B(n9392), .ZN(n9398) );
  INV_X1 U10725 ( .A(n9398), .ZN(n9394) );
  NAND2_X1 U10726 ( .A1(n9961), .A2(n9394), .ZN(n9395) );
  NAND2_X1 U10727 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9400) );
  NAND2_X1 U10728 ( .A1(n9950), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9399) );
  INV_X1 U10729 ( .A(n9401), .ZN(n9404) );
  INV_X1 U10730 ( .A(n9402), .ZN(n9403) );
  NAND2_X1 U10731 ( .A1(n5604), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9407) );
  OAI211_X1 U10732 ( .C1(n9632), .C2(n10022), .A(n9407), .B(n9406), .ZN(n9408)
         );
  AOI21_X1 U10733 ( .B1(n9556), .B2(n10015), .A(n9408), .ZN(n9409) );
  INV_X1 U10734 ( .A(n9409), .ZN(P1_U3264) );
  NAND2_X1 U10735 ( .A1(n9410), .A2(n10015), .ZN(n9413) );
  AOI22_X1 U10736 ( .A1(n9411), .A2(n10017), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10019), .ZN(n9412) );
  OAI211_X1 U10737 ( .C1(n9414), .C2(n10022), .A(n9413), .B(n9412), .ZN(n9415)
         );
  AOI21_X1 U10738 ( .B1(n9416), .B2(n9989), .A(n9415), .ZN(n9417) );
  OAI21_X1 U10739 ( .B1(n9418), .B2(n9554), .A(n9417), .ZN(P1_U3265) );
  XOR2_X1 U10740 ( .A(n9421), .B(n9419), .Z(n9570) );
  INV_X1 U10741 ( .A(n9570), .ZN(n9436) );
  OR2_X1 U10742 ( .A1(n9440), .A2(n9420), .ZN(n9423) );
  NOR2_X1 U10743 ( .A1(n9421), .A2(n9022), .ZN(n9422) );
  NAND2_X1 U10744 ( .A1(n9423), .A2(n9422), .ZN(n9424) );
  NAND2_X1 U10745 ( .A1(n9425), .A2(n9424), .ZN(n9426) );
  NAND2_X1 U10746 ( .A1(n9426), .A2(n9980), .ZN(n9429) );
  AOI22_X1 U10747 ( .A1(n9427), .A2(n9982), .B1(n9985), .B2(n9458), .ZN(n9428)
         );
  NAND2_X1 U10748 ( .A1(n9429), .A2(n9428), .ZN(n9568) );
  AOI211_X1 U10749 ( .C1(n9430), .C2(n9444), .A(n9968), .B(n8391), .ZN(n9569)
         );
  NAND2_X1 U10750 ( .A1(n9569), .A2(n10015), .ZN(n9433) );
  AOI22_X1 U10751 ( .A1(n9431), .A2(n10017), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10019), .ZN(n9432) );
  OAI211_X1 U10752 ( .C1(n9638), .C2(n10022), .A(n9433), .B(n9432), .ZN(n9434)
         );
  AOI21_X1 U10753 ( .B1(n9568), .B2(n9989), .A(n9434), .ZN(n9435) );
  OAI21_X1 U10754 ( .B1(n9436), .B2(n9554), .A(n9435), .ZN(P1_U3267) );
  XNOR2_X1 U10755 ( .A(n9438), .B(n9437), .ZN(n9577) );
  XNOR2_X1 U10756 ( .A(n9440), .B(n9439), .ZN(n9441) );
  OAI222_X1 U10757 ( .A1(n9551), .A2(n9443), .B1(n9549), .B2(n9442), .C1(
        n10002), .C2(n9441), .ZN(n9573) );
  AOI211_X1 U10758 ( .C1(n9575), .C2(n9461), .A(n9968), .B(n5659), .ZN(n9574)
         );
  NAND2_X1 U10759 ( .A1(n9574), .A2(n10015), .ZN(n9448) );
  INV_X1 U10760 ( .A(n9445), .ZN(n9446) );
  AOI22_X1 U10761 ( .A1(n9446), .A2(n10017), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10019), .ZN(n9447) );
  OAI211_X1 U10762 ( .C1(n4792), .C2(n10022), .A(n9448), .B(n9447), .ZN(n9449)
         );
  AOI21_X1 U10763 ( .B1(n9573), .B2(n9989), .A(n9449), .ZN(n9450) );
  OAI21_X1 U10764 ( .B1(n9577), .B2(n9554), .A(n9450), .ZN(P1_U3268) );
  XNOR2_X1 U10765 ( .A(n9451), .B(n9454), .ZN(n9583) );
  INV_X1 U10766 ( .A(n9583), .ZN(n9470) );
  NAND2_X1 U10767 ( .A1(n9453), .A2(n9452), .ZN(n9455) );
  NAND2_X1 U10768 ( .A1(n9455), .A2(n9454), .ZN(n9457) );
  NAND3_X1 U10769 ( .A1(n9457), .A2(n9980), .A3(n9456), .ZN(n9460) );
  AOI22_X1 U10770 ( .A1(n9458), .A2(n9982), .B1(n9985), .B2(n9489), .ZN(n9459)
         );
  NAND2_X1 U10771 ( .A1(n9460), .A2(n9459), .ZN(n9581) );
  OAI211_X1 U10772 ( .C1(n9579), .C2(n9477), .A(n10010), .B(n9461), .ZN(n9578)
         );
  INV_X1 U10773 ( .A(n9462), .ZN(n9463) );
  AOI22_X1 U10774 ( .A1(n9463), .A2(n10017), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10019), .ZN(n9466) );
  NAND2_X1 U10775 ( .A1(n9464), .A2(n10007), .ZN(n9465) );
  OAI211_X1 U10776 ( .C1(n9578), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9468)
         );
  AOI21_X1 U10777 ( .B1(n9581), .B2(n9989), .A(n9468), .ZN(n9469) );
  OAI21_X1 U10778 ( .B1(n9470), .B2(n9554), .A(n9469), .ZN(P1_U3269) );
  XNOR2_X1 U10779 ( .A(n9472), .B(n9471), .ZN(n9590) );
  XNOR2_X1 U10780 ( .A(n9474), .B(n9473), .ZN(n9476) );
  OAI21_X1 U10781 ( .B1(n9476), .B2(n10002), .A(n9475), .ZN(n9586) );
  INV_X1 U10782 ( .A(n9588), .ZN(n9481) );
  AOI211_X1 U10783 ( .C1(n9588), .C2(n9492), .A(n9968), .B(n9477), .ZN(n9587)
         );
  NAND2_X1 U10784 ( .A1(n9587), .A2(n10015), .ZN(n9480) );
  AOI22_X1 U10785 ( .A1(n9478), .A2(n10017), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10019), .ZN(n9479) );
  OAI211_X1 U10786 ( .C1(n9481), .C2(n10022), .A(n9480), .B(n9479), .ZN(n9482)
         );
  AOI21_X1 U10787 ( .B1(n9586), .B2(n9989), .A(n9482), .ZN(n9483) );
  OAI21_X1 U10788 ( .B1(n9590), .B2(n9554), .A(n9483), .ZN(P1_U3270) );
  XNOR2_X1 U10789 ( .A(n9485), .B(n9484), .ZN(n9593) );
  INV_X1 U10790 ( .A(n9593), .ZN(n9500) );
  OAI21_X1 U10791 ( .B1(n9487), .B2(n4750), .A(n9486), .ZN(n9488) );
  NAND2_X1 U10792 ( .A1(n9488), .A2(n9980), .ZN(n9491) );
  AOI22_X1 U10793 ( .A1(n9489), .A2(n9982), .B1(n9985), .B2(n9524), .ZN(n9490)
         );
  NAND2_X1 U10794 ( .A1(n9491), .A2(n9490), .ZN(n9591) );
  INV_X1 U10795 ( .A(n9492), .ZN(n9493) );
  AOI211_X1 U10796 ( .C1(n9494), .C2(n9502), .A(n9968), .B(n9493), .ZN(n9592)
         );
  NAND2_X1 U10797 ( .A1(n9592), .A2(n10015), .ZN(n9497) );
  AOI22_X1 U10798 ( .A1(n9495), .A2(n10017), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10019), .ZN(n9496) );
  OAI211_X1 U10799 ( .C1(n4571), .C2(n10022), .A(n9497), .B(n9496), .ZN(n9498)
         );
  AOI21_X1 U10800 ( .B1(n9591), .B2(n9989), .A(n9498), .ZN(n9499) );
  OAI21_X1 U10801 ( .B1(n9500), .B2(n9554), .A(n9499), .ZN(P1_U3271) );
  XNOR2_X1 U10802 ( .A(n9501), .B(n9510), .ZN(n9600) );
  INV_X1 U10803 ( .A(n9502), .ZN(n9503) );
  AOI211_X1 U10804 ( .C1(n9597), .C2(n9527), .A(n9968), .B(n9503), .ZN(n9596)
         );
  INV_X1 U10805 ( .A(n9597), .ZN(n9507) );
  INV_X1 U10806 ( .A(n9504), .ZN(n9505) );
  AOI22_X1 U10807 ( .A1(n9505), .A2(n10017), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10019), .ZN(n9506) );
  OAI21_X1 U10808 ( .B1(n9507), .B2(n10022), .A(n9506), .ZN(n9515) );
  OAI21_X1 U10809 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9513) );
  AOI222_X1 U10810 ( .A1(n9980), .A2(n9513), .B1(n9512), .B2(n9982), .C1(n9511), .C2(n9985), .ZN(n9599) );
  NOR2_X1 U10811 ( .A1(n9599), .A2(n10019), .ZN(n9514) );
  AOI211_X1 U10812 ( .C1(n9596), .C2(n10015), .A(n9515), .B(n9514), .ZN(n9516)
         );
  OAI21_X1 U10813 ( .B1(n9600), .B2(n9554), .A(n9516), .ZN(P1_U3272) );
  XNOR2_X1 U10814 ( .A(n9518), .B(n9517), .ZN(n9603) );
  INV_X1 U10815 ( .A(n9603), .ZN(n9536) );
  OAI21_X1 U10816 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9522) );
  NAND2_X1 U10817 ( .A1(n9522), .A2(n9980), .ZN(n9526) );
  AOI22_X1 U10818 ( .A1(n9524), .A2(n9982), .B1(n9985), .B2(n9523), .ZN(n9525)
         );
  NAND2_X1 U10819 ( .A1(n9526), .A2(n9525), .ZN(n9601) );
  INV_X1 U10820 ( .A(n9539), .ZN(n9529) );
  INV_X1 U10821 ( .A(n9527), .ZN(n9528) );
  AOI211_X1 U10822 ( .C1(n9530), .C2(n9529), .A(n9968), .B(n9528), .ZN(n9602)
         );
  NAND2_X1 U10823 ( .A1(n9602), .A2(n10015), .ZN(n9533) );
  AOI22_X1 U10824 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n10019), .B1(n9531), 
        .B2(n10017), .ZN(n9532) );
  OAI211_X1 U10825 ( .C1(n9931), .C2(n10022), .A(n9533), .B(n9532), .ZN(n9534)
         );
  AOI21_X1 U10826 ( .B1(n9601), .B2(n9989), .A(n9534), .ZN(n9535) );
  OAI21_X1 U10827 ( .B1(n9536), .B2(n9554), .A(n9535), .ZN(P1_U3273) );
  XNOR2_X1 U10828 ( .A(n9537), .B(n9546), .ZN(n9610) );
  INV_X1 U10829 ( .A(n9538), .ZN(n9540) );
  AOI211_X1 U10830 ( .C1(n9608), .C2(n9540), .A(n9968), .B(n9539), .ZN(n9607)
         );
  NOR2_X1 U10831 ( .A1(n9541), .A2(n10022), .ZN(n9544) );
  OAI22_X1 U10832 ( .A1(n9989), .A2(n9879), .B1(n9542), .B2(n9994), .ZN(n9543)
         );
  AOI211_X1 U10833 ( .C1(n9607), .C2(n10015), .A(n9544), .B(n9543), .ZN(n9553)
         );
  XOR2_X1 U10834 ( .A(n9546), .B(n9545), .Z(n9547) );
  OAI222_X1 U10835 ( .A1(n9551), .A2(n9550), .B1(n9549), .B2(n9548), .C1(n9547), .C2(n10002), .ZN(n9606) );
  NAND2_X1 U10836 ( .A1(n9606), .A2(n9989), .ZN(n9552) );
  OAI211_X1 U10837 ( .C1(n9610), .C2(n9554), .A(n9553), .B(n9552), .ZN(
        P1_U3274) );
  INV_X1 U10838 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9718) );
  NOR2_X1 U10839 ( .A1(n9556), .A2(n9555), .ZN(n9629) );
  MUX2_X1 U10840 ( .A(n9718), .B(n9629), .S(n10113), .Z(n9557) );
  OAI21_X1 U10841 ( .B1(n9632), .B2(n9616), .A(n9557), .ZN(P1_U3552) );
  MUX2_X1 U10842 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9633), .S(n10113), .Z(
        P1_U3551) );
  AOI21_X1 U10843 ( .B1(n9624), .B2(n9564), .A(n9563), .ZN(n9565) );
  OAI211_X1 U10844 ( .C1(n9567), .C2(n9627), .A(n9566), .B(n9565), .ZN(n9634)
         );
  MUX2_X1 U10845 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9634), .S(n10113), .Z(
        P1_U3549) );
  INV_X1 U10846 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9571) );
  MUX2_X1 U10847 ( .A(n9571), .B(n9635), .S(n10113), .Z(n9572) );
  OAI21_X1 U10848 ( .B1(n9638), .B2(n9616), .A(n9572), .ZN(P1_U3548) );
  AOI211_X1 U10849 ( .C1(n9624), .C2(n9575), .A(n9574), .B(n9573), .ZN(n9576)
         );
  OAI21_X1 U10850 ( .B1(n9627), .B2(n9577), .A(n9576), .ZN(n9639) );
  MUX2_X1 U10851 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9639), .S(n10113), .Z(
        P1_U3547) );
  INV_X1 U10852 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9584) );
  OAI21_X1 U10853 ( .B1(n9579), .B2(n10095), .A(n9578), .ZN(n9580) );
  OR2_X1 U10854 ( .A1(n9581), .A2(n9580), .ZN(n9582) );
  AOI21_X1 U10855 ( .B1(n9583), .B2(n6629), .A(n9582), .ZN(n9640) );
  MUX2_X1 U10856 ( .A(n9584), .B(n9640), .S(n10113), .Z(n9585) );
  INV_X1 U10857 ( .A(n9585), .ZN(P1_U3546) );
  AOI211_X1 U10858 ( .C1(n9624), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9589)
         );
  OAI21_X1 U10859 ( .B1(n9627), .B2(n9590), .A(n9589), .ZN(n9923) );
  MUX2_X1 U10860 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9923), .S(n10113), .Z(
        P1_U3545) );
  INV_X1 U10861 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9594) );
  AOI211_X1 U10862 ( .C1(n9593), .C2(n6629), .A(n9592), .B(n9591), .ZN(n9924)
         );
  MUX2_X1 U10863 ( .A(n9594), .B(n9924), .S(n10113), .Z(n9595) );
  OAI21_X1 U10864 ( .B1(n4571), .B2(n9616), .A(n9595), .ZN(P1_U3544) );
  AOI21_X1 U10865 ( .B1(n9624), .B2(n9597), .A(n9596), .ZN(n9598) );
  OAI211_X1 U10866 ( .C1(n9600), .C2(n9627), .A(n9599), .B(n9598), .ZN(n9927)
         );
  MUX2_X1 U10867 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9927), .S(n10113), .Z(
        P1_U3543) );
  INV_X1 U10868 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9604) );
  AOI211_X1 U10869 ( .C1(n9603), .C2(n6629), .A(n9602), .B(n9601), .ZN(n9928)
         );
  MUX2_X1 U10870 ( .A(n9604), .B(n9928), .S(n10113), .Z(n9605) );
  OAI21_X1 U10871 ( .B1(n9931), .B2(n9616), .A(n9605), .ZN(P1_U3542) );
  AOI211_X1 U10872 ( .C1(n9624), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9609)
         );
  OAI21_X1 U10873 ( .B1(n9627), .B2(n9610), .A(n9609), .ZN(n9932) );
  MUX2_X1 U10874 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9932), .S(n10113), .Z(
        P1_U3541) );
  AOI211_X1 U10875 ( .C1(n9613), .C2(n6629), .A(n9612), .B(n9611), .ZN(n9933)
         );
  MUX2_X1 U10876 ( .A(n9614), .B(n9933), .S(n10113), .Z(n9615) );
  OAI21_X1 U10877 ( .B1(n4569), .B2(n9616), .A(n9615), .ZN(P1_U3540) );
  AOI211_X1 U10878 ( .C1(n9624), .C2(n9619), .A(n9618), .B(n9617), .ZN(n9620)
         );
  OAI21_X1 U10879 ( .B1(n9627), .B2(n9621), .A(n9620), .ZN(n9937) );
  MUX2_X1 U10880 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9937), .S(n10113), .Z(
        P1_U3539) );
  AOI21_X1 U10881 ( .B1(n9624), .B2(n9623), .A(n9622), .ZN(n9625) );
  OAI211_X1 U10882 ( .C1(n9628), .C2(n9627), .A(n9626), .B(n9625), .ZN(n9938)
         );
  MUX2_X1 U10883 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9938), .S(n10113), .Z(
        P1_U3537) );
  MUX2_X1 U10884 ( .A(n9630), .B(n9629), .S(n10101), .Z(n9631) );
  OAI21_X1 U10885 ( .B1(n9632), .B2(n9936), .A(n9631), .ZN(P1_U3520) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9634), .S(n10101), .Z(
        P1_U3517) );
  INV_X1 U10887 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9636) );
  MUX2_X1 U10888 ( .A(n9636), .B(n9635), .S(n10101), .Z(n9637) );
  OAI21_X1 U10889 ( .B1(n9638), .B2(n9936), .A(n9637), .ZN(P1_U3516) );
  MUX2_X1 U10890 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9639), .S(n10101), .Z(
        P1_U3515) );
  MUX2_X1 U10891 ( .A(n9641), .B(n9640), .S(n10101), .Z(n9922) );
  NAND4_X1 U10892 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .A3(P2_ADDR_REG_1__SCAN_IN), .A4(n9888), .ZN(n9642) );
  NOR3_X1 U10893 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        n9642), .ZN(n9652) );
  NOR4_X1 U10894 ( .A1(P1_B_REG_SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), .A3(
        P1_REG3_REG_6__SCAN_IN), .A4(n10036), .ZN(n9643) );
  NAND3_X1 U10895 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9643), .A3(n10035), .ZN(
        n9650) );
  NOR4_X1 U10896 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .A3(P2_ADDR_REG_17__SCAN_IN), .A4(n9644), .ZN(n9647) );
  NOR4_X1 U10897 ( .A1(SI_19_), .A2(P2_DATAO_REG_21__SCAN_IN), .A3(n4580), 
        .A4(n9819), .ZN(n9646) );
  NOR4_X1 U10898 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(n5292), .A3(n7755), .A4(
        n9747), .ZN(n9645) );
  NAND4_X1 U10899 ( .A1(n9648), .A2(n9647), .A3(n9646), .A4(n9645), .ZN(n9649)
         );
  NOR4_X1 U10900 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(P1_U3086), .A3(n9650), 
        .A4(n9649), .ZN(n9651) );
  NAND4_X1 U10901 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(n9652), .A4(n9651), .ZN(n9664) );
  NAND4_X1 U10902 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(SI_26_), .A3(n9837), .A4(
        n5110), .ZN(n9663) );
  NAND4_X1 U10903 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_REG2_REG_21__SCAN_IN), 
        .A3(n5691), .A4(n9694), .ZN(n9662) );
  NOR4_X1 U10904 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_REG2_REG_17__SCAN_IN), 
        .A3(P1_REG2_REG_26__SCAN_IN), .A4(P2_ADDR_REG_14__SCAN_IN), .ZN(n9659)
         );
  NAND4_X1 U10905 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .A3(n9653), .A4(n9868), .ZN(n9657) );
  INV_X1 U10906 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9840) );
  NAND4_X1 U10907 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(n10325), .A3(n9840), .A4(
        n9874), .ZN(n9656) );
  NAND4_X1 U10908 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_REG2_REG_30__SCAN_IN), 
        .A3(P2_REG2_REG_0__SCAN_IN), .A4(n9735), .ZN(n9655) );
  NAND4_X1 U10909 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_REG1_REG_14__SCAN_IN), .A4(n9736), .ZN(n9654) );
  NOR4_X1 U10910 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n9658)
         );
  NAND3_X1 U10911 ( .A1(n9660), .A2(n9659), .A3(n9658), .ZN(n9661) );
  NOR4_X1 U10912 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9692)
         );
  INV_X1 U10913 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9665) );
  NAND4_X1 U10914 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(P1_REG0_REG_17__SCAN_IN), 
        .A3(n9762), .A4(n9665), .ZN(n9669) );
  NAND4_X1 U10915 ( .A1(P1_REG0_REG_22__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(P1_REG2_REG_19__SCAN_IN), .A4(P1_REG0_REG_18__SCAN_IN), .ZN(n9668)
         );
  INV_X1 U10916 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9863) );
  NAND4_X1 U10917 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_REG0_REG_0__SCAN_IN), 
        .A3(n5124), .A4(n9863), .ZN(n9667) );
  NAND4_X1 U10918 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(P1_REG1_REG_3__SCAN_IN), 
        .A3(n6851), .A4(n9809), .ZN(n9666) );
  NOR4_X1 U10919 ( .A1(n9669), .A2(n9668), .A3(n9667), .A4(n9666), .ZN(n9691)
         );
  NOR4_X1 U10920 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        n8659), .A4(n5913), .ZN(n9690) );
  NOR4_X1 U10921 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(P2_REG1_REG_31__SCAN_IN), 
        .A3(n9822), .A4(n9823), .ZN(n9670) );
  NAND3_X1 U10922 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .A3(n9670), .ZN(n9683) );
  NAND4_X1 U10923 ( .A1(n9803), .A2(n9745), .A3(P1_DATAO_REG_0__SCAN_IN), .A4(
        SI_3_), .ZN(n9672) );
  INV_X1 U10924 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9906) );
  NAND4_X1 U10925 ( .A1(n10194), .A2(n9906), .A3(P2_IR_REG_17__SCAN_IN), .A4(
        P2_IR_REG_8__SCAN_IN), .ZN(n9671) );
  NOR2_X1 U10926 ( .A1(n9672), .A2(n9671), .ZN(n9681) );
  NOR4_X1 U10927 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P1_DATAO_REG_30__SCAN_IN), 
        .A3(P1_REG1_REG_30__SCAN_IN), .A4(n9794), .ZN(n9674) );
  NOR4_X1 U10928 ( .A1(P2_D_REG_1__SCAN_IN), .A2(P1_REG2_REG_7__SCAN_IN), .A3(
        n9862), .A4(n9904), .ZN(n9673) );
  NAND2_X1 U10929 ( .A1(n9674), .A2(n9673), .ZN(n9675) );
  NOR2_X1 U10930 ( .A1(SI_23_), .A2(n9675), .ZN(n9676) );
  NAND4_X1 U10931 ( .A1(n9676), .A2(n7550), .A3(P1_REG0_REG_13__SCAN_IN), .A4(
        n10111), .ZN(n9679) );
  NAND4_X1 U10932 ( .A1(n9677), .A2(P2_DATAO_REG_2__SCAN_IN), .A3(
        P2_DATAO_REG_23__SCAN_IN), .A4(P1_DATAO_REG_6__SCAN_IN), .ZN(n9678) );
  NOR2_X1 U10933 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  NAND2_X1 U10934 ( .A1(n9681), .A2(n9680), .ZN(n9682) );
  NOR2_X1 U10935 ( .A1(n9683), .A2(n9682), .ZN(n9688) );
  NAND4_X1 U10936 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P1_REG1_REG_8__SCAN_IN), 
        .A3(P1_REG0_REG_8__SCAN_IN), .A4(n7353), .ZN(n9684) );
  NOR3_X1 U10937 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(P1_REG0_REG_14__SCAN_IN), 
        .A3(n9684), .ZN(n9687) );
  NOR4_X1 U10938 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(P2_REG2_REG_2__SCAN_IN), 
        .A3(P2_WR_REG_SCAN_IN), .A4(n9893), .ZN(n9686) );
  NOR4_X1 U10939 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_REG0_REG_26__SCAN_IN), .A4(n9771), .ZN(n9685) );
  AND4_X1 U10940 ( .A1(n9688), .A2(n9687), .A3(n9686), .A4(n9685), .ZN(n9689)
         );
  NAND4_X1 U10941 ( .A1(n9692), .A2(n9691), .A3(n9690), .A4(n9689), .ZN(n9920)
         );
  INV_X1 U10942 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U10943 ( .A1(n9694), .A2(keyinput93), .B1(n10100), .B2(keyinput54), 
        .ZN(n9693) );
  OAI221_X1 U10944 ( .B1(n9694), .B2(keyinput93), .C1(n10100), .C2(keyinput54), 
        .A(n9693), .ZN(n9704) );
  AOI22_X1 U10945 ( .A1(n4580), .A2(keyinput92), .B1(n9696), .B2(keyinput107), 
        .ZN(n9695) );
  OAI221_X1 U10946 ( .B1(n4580), .B2(keyinput92), .C1(n9696), .C2(keyinput107), 
        .A(n9695), .ZN(n9703) );
  AOI22_X1 U10947 ( .A1(n10111), .A2(keyinput70), .B1(n8659), .B2(keyinput97), 
        .ZN(n9697) );
  OAI221_X1 U10948 ( .B1(n10111), .B2(keyinput70), .C1(n8659), .C2(keyinput97), 
        .A(n9697), .ZN(n9702) );
  INV_X1 U10949 ( .A(keyinput17), .ZN(n9699) );
  AOI22_X1 U10950 ( .A1(n9700), .A2(keyinput23), .B1(P2_ADDR_REG_14__SCAN_IN), 
        .B2(n9699), .ZN(n9698) );
  OAI221_X1 U10951 ( .B1(n9700), .B2(keyinput23), .C1(n9699), .C2(
        P2_ADDR_REG_14__SCAN_IN), .A(n9698), .ZN(n9701) );
  NOR4_X1 U10952 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(n9756)
         );
  AOI22_X1 U10953 ( .A1(n9706), .A2(keyinput98), .B1(keyinput25), .B2(n8674), 
        .ZN(n9705) );
  OAI221_X1 U10954 ( .B1(n9706), .B2(keyinput98), .C1(n8674), .C2(keyinput25), 
        .A(n9705), .ZN(n9716) );
  AOI22_X1 U10955 ( .A1(n9708), .A2(keyinput127), .B1(n10035), .B2(keyinput38), 
        .ZN(n9707) );
  OAI221_X1 U10956 ( .B1(n9708), .B2(keyinput127), .C1(n10035), .C2(keyinput38), .A(n9707), .ZN(n9715) );
  AOI22_X1 U10957 ( .A1(n9710), .A2(keyinput4), .B1(keyinput74), .B2(n5576), 
        .ZN(n9709) );
  OAI221_X1 U10958 ( .B1(n9710), .B2(keyinput4), .C1(n5576), .C2(keyinput74), 
        .A(n9709), .ZN(n9714) );
  INV_X1 U10959 ( .A(P1_B_REG_SCAN_IN), .ZN(n9712) );
  AOI22_X1 U10960 ( .A1(n9712), .A2(keyinput86), .B1(n6112), .B2(keyinput83), 
        .ZN(n9711) );
  OAI221_X1 U10961 ( .B1(n9712), .B2(keyinput86), .C1(n6112), .C2(keyinput83), 
        .A(n9711), .ZN(n9713) );
  NOR4_X1 U10962 ( .A1(n9716), .A2(n9715), .A3(n9714), .A4(n9713), .ZN(n9755)
         );
  AOI22_X1 U10963 ( .A1(n9718), .A2(keyinput100), .B1(n5196), .B2(keyinput11), 
        .ZN(n9717) );
  OAI221_X1 U10964 ( .B1(n9718), .B2(keyinput100), .C1(n5196), .C2(keyinput11), 
        .A(n9717), .ZN(n9728) );
  INV_X1 U10965 ( .A(keyinput125), .ZN(n9720) );
  AOI22_X1 U10966 ( .A1(n9721), .A2(keyinput105), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n9720), .ZN(n9719) );
  OAI221_X1 U10967 ( .B1(n9721), .B2(keyinput105), .C1(n9720), .C2(
        P2_ADDR_REG_17__SCAN_IN), .A(n9719), .ZN(n9727) );
  INV_X1 U10968 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U10969 ( .A1(n5493), .A2(keyinput48), .B1(n10059), .B2(keyinput57), 
        .ZN(n9722) );
  OAI221_X1 U10970 ( .B1(n5493), .B2(keyinput48), .C1(n10059), .C2(keyinput57), 
        .A(n9722), .ZN(n9726) );
  INV_X1 U10971 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10038) );
  INV_X1 U10972 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9724) );
  AOI22_X1 U10973 ( .A1(n10038), .A2(keyinput40), .B1(n9724), .B2(keyinput28), 
        .ZN(n9723) );
  OAI221_X1 U10974 ( .B1(n10038), .B2(keyinput40), .C1(n9724), .C2(keyinput28), 
        .A(n9723), .ZN(n9725) );
  NOR4_X1 U10975 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n9754)
         );
  AOI22_X1 U10976 ( .A1(n7755), .A2(keyinput9), .B1(keyinput67), .B2(n9730), 
        .ZN(n9729) );
  OAI221_X1 U10977 ( .B1(n7755), .B2(keyinput9), .C1(n9730), .C2(keyinput67), 
        .A(n9729), .ZN(n9752) );
  AOI22_X1 U10978 ( .A1(n9733), .A2(keyinput37), .B1(keyinput10), .B2(n9732), 
        .ZN(n9731) );
  OAI221_X1 U10979 ( .B1(n9733), .B2(keyinput37), .C1(n9732), .C2(keyinput10), 
        .A(n9731), .ZN(n9742) );
  AOI22_X1 U10980 ( .A1(n9736), .A2(keyinput95), .B1(keyinput103), .B2(n9735), 
        .ZN(n9734) );
  OAI221_X1 U10981 ( .B1(n9736), .B2(keyinput95), .C1(n9735), .C2(keyinput103), 
        .A(n9734), .ZN(n9741) );
  AOI22_X1 U10982 ( .A1(n9739), .A2(keyinput68), .B1(keyinput120), .B2(n9738), 
        .ZN(n9737) );
  OAI221_X1 U10983 ( .B1(n9739), .B2(keyinput68), .C1(n9738), .C2(keyinput120), 
        .A(n9737), .ZN(n9740) );
  OR3_X1 U10984 ( .A1(n9742), .A2(n9741), .A3(n9740), .ZN(n9751) );
  AOI22_X1 U10985 ( .A1(n9745), .A2(keyinput24), .B1(keyinput43), .B2(n9744), 
        .ZN(n9743) );
  OAI221_X1 U10986 ( .B1(n9745), .B2(keyinput24), .C1(n9744), .C2(keyinput43), 
        .A(n9743), .ZN(n9750) );
  AOI22_X1 U10987 ( .A1(n9748), .A2(keyinput109), .B1(n9747), .B2(keyinput6), 
        .ZN(n9746) );
  OAI221_X1 U10988 ( .B1(n9748), .B2(keyinput109), .C1(n9747), .C2(keyinput6), 
        .A(n9746), .ZN(n9749) );
  NOR4_X1 U10989 ( .A1(n9752), .A2(n9751), .A3(n9750), .A4(n9749), .ZN(n9753)
         );
  AND4_X1 U10990 ( .A1(n9756), .A2(n9755), .A3(n9754), .A4(n9753), .ZN(n9831)
         );
  AOI22_X1 U10991 ( .A1(n5124), .A2(keyinput124), .B1(keyinput81), .B2(n9758), 
        .ZN(n9757) );
  OAI221_X1 U10992 ( .B1(n5124), .B2(keyinput124), .C1(n9758), .C2(keyinput81), 
        .A(n9757), .ZN(n9768) );
  AOI22_X1 U10993 ( .A1(n10321), .A2(keyinput62), .B1(keyinput39), .B2(n10053), 
        .ZN(n9759) );
  OAI221_X1 U10994 ( .B1(n10321), .B2(keyinput62), .C1(n10053), .C2(keyinput39), .A(n9759), .ZN(n9767) );
  AOI22_X1 U10995 ( .A1(n9762), .A2(keyinput36), .B1(n9761), .B2(keyinput110), 
        .ZN(n9760) );
  OAI221_X1 U10996 ( .B1(n9762), .B2(keyinput36), .C1(n9761), .C2(keyinput110), 
        .A(n9760), .ZN(n9766) );
  INV_X1 U10997 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U10998 ( .A1(n10050), .A2(keyinput82), .B1(keyinput29), .B2(n9764), 
        .ZN(n9763) );
  OAI221_X1 U10999 ( .B1(n10050), .B2(keyinput82), .C1(n9764), .C2(keyinput29), 
        .A(n9763), .ZN(n9765) );
  NOR4_X1 U11000 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n9830)
         );
  AOI22_X1 U11001 ( .A1(n5126), .A2(keyinput71), .B1(P1_U3086), .B2(keyinput46), .ZN(n9769) );
  OAI221_X1 U11002 ( .B1(n5126), .B2(keyinput71), .C1(P1_U3086), .C2(
        keyinput46), .A(n9769), .ZN(n9784) );
  AOI22_X1 U11003 ( .A1(n9772), .A2(keyinput90), .B1(keyinput2), .B2(n9771), 
        .ZN(n9770) );
  OAI221_X1 U11004 ( .B1(n9772), .B2(keyinput90), .C1(n9771), .C2(keyinput2), 
        .A(n9770), .ZN(n9783) );
  XNOR2_X1 U11005 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput115), .ZN(n9776)
         );
  XNOR2_X1 U11006 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput15), .ZN(n9775) );
  XNOR2_X1 U11007 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput56), .ZN(n9774) );
  XNOR2_X1 U11008 ( .A(P1_REG0_REG_22__SCAN_IN), .B(keyinput58), .ZN(n9773) );
  NAND4_X1 U11009 ( .A1(n9776), .A2(n9775), .A3(n9774), .A4(n9773), .ZN(n9782)
         );
  XNOR2_X1 U11010 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput113), .ZN(n9780) );
  XNOR2_X1 U11011 ( .A(SI_3_), .B(keyinput111), .ZN(n9779) );
  XNOR2_X1 U11012 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput126), .ZN(n9778) );
  XNOR2_X1 U11013 ( .A(P1_REG0_REG_21__SCAN_IN), .B(keyinput114), .ZN(n9777)
         );
  NAND4_X1 U11014 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n9781)
         );
  OR4_X1 U11015 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9789)
         );
  AOI22_X1 U11016 ( .A1(n7353), .A2(keyinput118), .B1(keyinput30), .B2(n10103), 
        .ZN(n9785) );
  OAI221_X1 U11017 ( .B1(n7353), .B2(keyinput118), .C1(n10103), .C2(keyinput30), .A(n9785), .ZN(n9788) );
  XNOR2_X1 U11018 ( .A(n9786), .B(keyinput33), .ZN(n9787) );
  NOR3_X1 U11019 ( .A1(n9789), .A2(n9788), .A3(n9787), .ZN(n9829) );
  XOR2_X1 U11020 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput27), .Z(n9793) );
  XOR2_X1 U11021 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput61), .Z(n9792) );
  XOR2_X1 U11022 ( .A(P1_REG1_REG_15__SCAN_IN), .B(keyinput119), .Z(n9791) );
  XOR2_X1 U11023 ( .A(P2_REG2_REG_17__SCAN_IN), .B(keyinput55), .Z(n9790) );
  NOR4_X1 U11024 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(n9817)
         );
  XNOR2_X1 U11025 ( .A(n9794), .B(keyinput32), .ZN(n9801) );
  XNOR2_X1 U11026 ( .A(n9795), .B(keyinput75), .ZN(n9800) );
  XNOR2_X1 U11027 ( .A(n9796), .B(keyinput42), .ZN(n9799) );
  XNOR2_X1 U11028 ( .A(n9797), .B(keyinput66), .ZN(n9798) );
  NOR4_X1 U11029 ( .A1(n9801), .A2(n9800), .A3(n9799), .A4(n9798), .ZN(n9816)
         );
  XOR2_X1 U11030 ( .A(P2_REG1_REG_29__SCAN_IN), .B(keyinput79), .Z(n9808) );
  XNOR2_X1 U11031 ( .A(n9802), .B(keyinput123), .ZN(n9807) );
  XNOR2_X1 U11032 ( .A(n9803), .B(keyinput44), .ZN(n9806) );
  XNOR2_X1 U11033 ( .A(keyinput51), .B(n9804), .ZN(n9805) );
  NOR4_X1 U11034 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(n9815)
         );
  XNOR2_X1 U11035 ( .A(keyinput108), .B(n5069), .ZN(n9813) );
  XNOR2_X1 U11036 ( .A(keyinput34), .B(n9677), .ZN(n9812) );
  XNOR2_X1 U11037 ( .A(keyinput89), .B(n9809), .ZN(n9811) );
  XNOR2_X1 U11038 ( .A(keyinput94), .B(n5292), .ZN(n9810) );
  NOR4_X1 U11039 ( .A1(n9813), .A2(n9812), .A3(n9811), .A4(n9810), .ZN(n9814)
         );
  NAND4_X1 U11040 ( .A1(n9817), .A2(n9816), .A3(n9815), .A4(n9814), .ZN(n9827)
         );
  AOI22_X1 U11041 ( .A1(n9820), .A2(keyinput50), .B1(n9819), .B2(keyinput7), 
        .ZN(n9818) );
  OAI221_X1 U11042 ( .B1(n9820), .B2(keyinput50), .C1(n9819), .C2(keyinput7), 
        .A(n9818), .ZN(n9826) );
  AOI22_X1 U11043 ( .A1(n9823), .A2(keyinput14), .B1(keyinput41), .B2(n9822), 
        .ZN(n9821) );
  OAI221_X1 U11044 ( .B1(n9823), .B2(keyinput14), .C1(n9822), .C2(keyinput41), 
        .A(n9821), .ZN(n9825) );
  XNOR2_X1 U11045 ( .A(n10336), .B(keyinput19), .ZN(n9824) );
  NOR4_X1 U11046 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9828)
         );
  AND4_X1 U11047 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n9918)
         );
  AOI22_X1 U11048 ( .A1(n5691), .A2(keyinput0), .B1(keyinput112), .B2(n5110), 
        .ZN(n9832) );
  OAI221_X1 U11049 ( .B1(n5691), .B2(keyinput0), .C1(n5110), .C2(keyinput112), 
        .A(n9832), .ZN(n9844) );
  AOI22_X1 U11050 ( .A1(n9835), .A2(keyinput104), .B1(n9834), .B2(keyinput102), 
        .ZN(n9833) );
  OAI221_X1 U11051 ( .B1(n9835), .B2(keyinput104), .C1(n9834), .C2(keyinput102), .A(n9833), .ZN(n9843) );
  AOI22_X1 U11052 ( .A1(n9838), .A2(keyinput20), .B1(keyinput117), .B2(n9837), 
        .ZN(n9836) );
  OAI221_X1 U11053 ( .B1(n9838), .B2(keyinput20), .C1(n9837), .C2(keyinput117), 
        .A(n9836), .ZN(n9842) );
  AOI22_X1 U11054 ( .A1(n5738), .A2(keyinput99), .B1(n9840), .B2(keyinput5), 
        .ZN(n9839) );
  OAI221_X1 U11055 ( .B1(n5738), .B2(keyinput99), .C1(n9840), .C2(keyinput5), 
        .A(n9839), .ZN(n9841) );
  NOR4_X1 U11056 ( .A1(n9844), .A2(n9843), .A3(n9842), .A4(n9841), .ZN(n9917)
         );
  AOI22_X1 U11057 ( .A1(n10036), .A2(keyinput106), .B1(n9846), .B2(keyinput12), 
        .ZN(n9845) );
  OAI221_X1 U11058 ( .B1(n10036), .B2(keyinput106), .C1(n9846), .C2(keyinput12), .A(n9845), .ZN(n9857) );
  INV_X1 U11059 ( .A(keyinput91), .ZN(n9848) );
  AOI22_X1 U11060 ( .A1(n9934), .A2(keyinput84), .B1(P2_ADDR_REG_13__SCAN_IN), 
        .B2(n9848), .ZN(n9847) );
  OAI221_X1 U11061 ( .B1(n9934), .B2(keyinput84), .C1(n9848), .C2(
        P2_ADDR_REG_13__SCAN_IN), .A(n9847), .ZN(n9856) );
  AOI22_X1 U11062 ( .A1(n9851), .A2(keyinput52), .B1(keyinput80), .B2(n9850), 
        .ZN(n9849) );
  OAI221_X1 U11063 ( .B1(n9851), .B2(keyinput52), .C1(n9850), .C2(keyinput80), 
        .A(n9849), .ZN(n9855) );
  AOI22_X1 U11064 ( .A1(n10039), .A2(keyinput53), .B1(n9853), .B2(keyinput49), 
        .ZN(n9852) );
  OAI221_X1 U11065 ( .B1(n10039), .B2(keyinput53), .C1(n9853), .C2(keyinput49), 
        .A(n9852), .ZN(n9854) );
  NOR4_X1 U11066 ( .A1(n9857), .A2(n9856), .A3(n9855), .A4(n9854), .ZN(n9916)
         );
  INV_X1 U11067 ( .A(keyinput63), .ZN(n9859) );
  AOI22_X1 U11068 ( .A1(n9860), .A2(keyinput18), .B1(P1_ADDR_REG_10__SCAN_IN), 
        .B2(n9859), .ZN(n9858) );
  OAI221_X1 U11069 ( .B1(n9860), .B2(keyinput18), .C1(n9859), .C2(
        P1_ADDR_REG_10__SCAN_IN), .A(n9858), .ZN(n9872) );
  AOI22_X1 U11070 ( .A1(n9863), .A2(keyinput16), .B1(n9862), .B2(keyinput13), 
        .ZN(n9861) );
  OAI221_X1 U11071 ( .B1(n9863), .B2(keyinput16), .C1(n9862), .C2(keyinput13), 
        .A(n9861), .ZN(n9871) );
  AOI22_X1 U11072 ( .A1(n9865), .A2(keyinput60), .B1(n10042), .B2(keyinput64), 
        .ZN(n9864) );
  OAI221_X1 U11073 ( .B1(n9865), .B2(keyinput60), .C1(n10042), .C2(keyinput64), 
        .A(n9864), .ZN(n9870) );
  AOI22_X1 U11074 ( .A1(n9868), .A2(keyinput85), .B1(keyinput116), .B2(n9867), 
        .ZN(n9866) );
  OAI221_X1 U11075 ( .B1(n9868), .B2(keyinput85), .C1(n9867), .C2(keyinput116), 
        .A(n9866), .ZN(n9869) );
  NOR4_X1 U11076 ( .A1(n9872), .A2(n9871), .A3(n9870), .A4(n9869), .ZN(n9914)
         );
  AOI22_X1 U11077 ( .A1(n10045), .A2(keyinput47), .B1(keyinput65), .B2(n9874), 
        .ZN(n9873) );
  OAI221_X1 U11078 ( .B1(n10045), .B2(keyinput47), .C1(n9874), .C2(keyinput65), 
        .A(n9873), .ZN(n9884) );
  INV_X1 U11079 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9876) );
  AOI22_X1 U11080 ( .A1(n9876), .A2(keyinput77), .B1(n10325), .B2(keyinput59), 
        .ZN(n9875) );
  OAI221_X1 U11081 ( .B1(n9876), .B2(keyinput77), .C1(n10325), .C2(keyinput59), 
        .A(n9875), .ZN(n9883) );
  AOI22_X1 U11082 ( .A1(n9879), .A2(keyinput8), .B1(n9878), .B2(keyinput96), 
        .ZN(n9877) );
  OAI221_X1 U11083 ( .B1(n9879), .B2(keyinput8), .C1(n9878), .C2(keyinput96), 
        .A(n9877), .ZN(n9882) );
  AOI22_X1 U11084 ( .A1(n6099), .A2(keyinput122), .B1(keyinput72), .B2(n8613), 
        .ZN(n9880) );
  OAI221_X1 U11085 ( .B1(n6099), .B2(keyinput122), .C1(n8613), .C2(keyinput72), 
        .A(n9880), .ZN(n9881) );
  NOR4_X1 U11086 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(n9913)
         );
  AOI22_X1 U11087 ( .A1(n5675), .A2(keyinput87), .B1(keyinput78), .B2(n9886), 
        .ZN(n9885) );
  OAI221_X1 U11088 ( .B1(n5675), .B2(keyinput87), .C1(n9886), .C2(keyinput78), 
        .A(n9885), .ZN(n9897) );
  AOI22_X1 U11089 ( .A1(n9888), .A2(keyinput88), .B1(n5913), .B2(keyinput101), 
        .ZN(n9887) );
  OAI221_X1 U11090 ( .B1(n9888), .B2(keyinput88), .C1(n5913), .C2(keyinput101), 
        .A(n9887), .ZN(n9896) );
  AOI22_X1 U11091 ( .A1(n9890), .A2(keyinput35), .B1(n5235), .B2(keyinput22), 
        .ZN(n9889) );
  OAI221_X1 U11092 ( .B1(n9890), .B2(keyinput35), .C1(n5235), .C2(keyinput22), 
        .A(n9889), .ZN(n9895) );
  INV_X1 U11093 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9892) );
  AOI22_X1 U11094 ( .A1(n9893), .A2(keyinput69), .B1(keyinput76), .B2(n9892), 
        .ZN(n9891) );
  OAI221_X1 U11095 ( .B1(n9893), .B2(keyinput69), .C1(n9892), .C2(keyinput76), 
        .A(n9891), .ZN(n9894) );
  NOR4_X1 U11096 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n9912)
         );
  AOI22_X1 U11097 ( .A1(n10259), .A2(keyinput31), .B1(keyinput121), .B2(n9899), 
        .ZN(n9898) );
  OAI221_X1 U11098 ( .B1(n10259), .B2(keyinput31), .C1(n9899), .C2(keyinput121), .A(n9898), .ZN(n9910) );
  INV_X1 U11099 ( .A(keyinput21), .ZN(n9901) );
  AOI22_X1 U11100 ( .A1(n9902), .A2(keyinput45), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n9901), .ZN(n9900) );
  OAI221_X1 U11101 ( .B1(n9902), .B2(keyinput45), .C1(n9901), .C2(
        P1_ADDR_REG_15__SCAN_IN), .A(n9900), .ZN(n9909) );
  AOI22_X1 U11102 ( .A1(n9904), .A2(keyinput1), .B1(n10194), .B2(keyinput26), 
        .ZN(n9903) );
  OAI221_X1 U11103 ( .B1(n9904), .B2(keyinput1), .C1(n10194), .C2(keyinput26), 
        .A(n9903), .ZN(n9908) );
  AOI22_X1 U11104 ( .A1(n6851), .A2(keyinput73), .B1(n9906), .B2(keyinput3), 
        .ZN(n9905) );
  OAI221_X1 U11105 ( .B1(n6851), .B2(keyinput73), .C1(n9906), .C2(keyinput3), 
        .A(n9905), .ZN(n9907) );
  NOR4_X1 U11106 ( .A1(n9910), .A2(n9909), .A3(n9908), .A4(n9907), .ZN(n9911)
         );
  AND4_X1 U11107 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(n9915)
         );
  NAND4_X1 U11108 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n9919)
         );
  XOR2_X1 U11109 ( .A(n9920), .B(n9919), .Z(n9921) );
  XNOR2_X1 U11110 ( .A(n9922), .B(n9921), .ZN(P1_U3514) );
  MUX2_X1 U11111 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9923), .S(n10101), .Z(
        P1_U3513) );
  MUX2_X1 U11112 ( .A(n9925), .B(n9924), .S(n10101), .Z(n9926) );
  OAI21_X1 U11113 ( .B1(n4571), .B2(n9936), .A(n9926), .ZN(P1_U3512) );
  MUX2_X1 U11114 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9927), .S(n10101), .Z(
        P1_U3511) );
  INV_X1 U11115 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9929) );
  MUX2_X1 U11116 ( .A(n9929), .B(n9928), .S(n10101), .Z(n9930) );
  OAI21_X1 U11117 ( .B1(n9931), .B2(n9936), .A(n9930), .ZN(P1_U3510) );
  MUX2_X1 U11118 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9932), .S(n10101), .Z(
        P1_U3509) );
  MUX2_X1 U11119 ( .A(n9934), .B(n9933), .S(n10101), .Z(n9935) );
  OAI21_X1 U11120 ( .B1(n4569), .B2(n9936), .A(n9935), .ZN(P1_U3507) );
  MUX2_X1 U11121 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9937), .S(n10101), .Z(
        P1_U3504) );
  MUX2_X1 U11122 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9938), .S(n10101), .Z(
        P1_U3498) );
  MUX2_X1 U11123 ( .A(P1_D_REG_1__SCAN_IN), .B(n9939), .S(n10060), .Z(P1_U3440) );
  MUX2_X1 U11124 ( .A(n9941), .B(P1_D_REG_0__SCAN_IN), .S(n9940), .Z(P1_U3439)
         );
  INV_X1 U11125 ( .A(n9942), .ZN(n9943) );
  MUX2_X1 U11126 ( .A(n9943), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11127 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11128 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11129 ( .B1(n5558), .B2(n9945), .A(n9944), .ZN(n9946) );
  XNOR2_X1 U11130 ( .A(n9946), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9949) );
  AOI22_X1 U11131 ( .A1(n9950), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9947) );
  OAI21_X1 U11132 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(P1_U3243) );
  AOI22_X1 U11133 ( .A1(n9950), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9967) );
  INV_X1 U11134 ( .A(n9951), .ZN(n9952) );
  OAI21_X1 U11135 ( .B1(n9954), .B2(n9953), .A(n9952), .ZN(n9957) );
  OAI22_X1 U11136 ( .A1(n9958), .A2(n9957), .B1(n9956), .B2(n9955), .ZN(n9959)
         );
  INV_X1 U11137 ( .A(n9959), .ZN(n9966) );
  OAI211_X1 U11138 ( .C1(n9963), .C2(n9962), .A(n9961), .B(n9960), .ZN(n9964)
         );
  NAND4_X1 U11139 ( .A1(n9967), .A2(n9966), .A3(n9965), .A4(n9964), .ZN(
        P1_U3245) );
  AOI21_X1 U11140 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9972) );
  NAND2_X1 U11141 ( .A1(n9972), .A2(n9971), .ZN(n10093) );
  INV_X1 U11142 ( .A(n10093), .ZN(n9973) );
  AOI22_X1 U11143 ( .A1(n9973), .A2(n10015), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n10019), .ZN(n9993) );
  XNOR2_X1 U11144 ( .A(n9974), .B(n9978), .ZN(n10092) );
  NOR2_X1 U11145 ( .A1(n10092), .A2(n9975), .ZN(n9991) );
  NAND2_X1 U11146 ( .A1(n9977), .A2(n9976), .ZN(n9979) );
  XNOR2_X1 U11147 ( .A(n9979), .B(n9978), .ZN(n9981) );
  NAND2_X1 U11148 ( .A1(n9981), .A2(n9980), .ZN(n9987) );
  AOI22_X1 U11149 ( .A1(n9985), .A2(n9984), .B1(n9983), .B2(n9982), .ZN(n9986)
         );
  AND2_X1 U11150 ( .A1(n9987), .A2(n9986), .ZN(n10094) );
  OAI21_X1 U11151 ( .B1(n10096), .B2(n9988), .A(n10094), .ZN(n9990) );
  OAI21_X1 U11152 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(n9992) );
  OAI211_X1 U11153 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(
        P1_U3280) );
  NAND2_X1 U11154 ( .A1(n9997), .A2(n9996), .ZN(n9998) );
  XNOR2_X1 U11155 ( .A(n9998), .B(n9999), .ZN(n10083) );
  XNOR2_X1 U11156 ( .A(n10000), .B(n9999), .ZN(n10003) );
  OAI21_X1 U11157 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(n10004) );
  AOI21_X1 U11158 ( .B1(n10083), .B2(n10005), .A(n10004), .ZN(n10080) );
  AOI222_X1 U11159 ( .A1(n10008), .A2(n10007), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n10019), .C1(n10006), .C2(n10017), .ZN(n10014) );
  OAI211_X1 U11160 ( .C1(n10079), .C2(n4420), .A(n4564), .B(n10010), .ZN(
        n10078) );
  INV_X1 U11161 ( .A(n10078), .ZN(n10011) );
  AOI22_X1 U11162 ( .A1(n10083), .A2(n10012), .B1(n10015), .B2(n10011), .ZN(
        n10013) );
  OAI211_X1 U11163 ( .C1(n5604), .C2(n10080), .A(n10014), .B(n10013), .ZN(
        P1_U3282) );
  NAND2_X1 U11164 ( .A1(n10016), .A2(n10015), .ZN(n10021) );
  AOI22_X1 U11165 ( .A1(n10019), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10018), 
        .B2(n10017), .ZN(n10020) );
  OAI211_X1 U11166 ( .C1(n10023), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10024) );
  AOI21_X1 U11167 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(n10027) );
  OAI21_X1 U11168 ( .B1(n5604), .B2(n10028), .A(n10027), .ZN(P1_U3287) );
  INV_X1 U11169 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U11170 ( .A1(n10060), .A2(n10029), .ZN(P1_U3294) );
  INV_X1 U11171 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U11172 ( .A1(n10060), .A2(n10030), .ZN(P1_U3295) );
  INV_X1 U11173 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U11174 ( .A1(n10060), .A2(n10031), .ZN(P1_U3296) );
  INV_X1 U11175 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U11176 ( .A1(n10044), .A2(n10032), .ZN(P1_U3297) );
  INV_X1 U11177 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10033) );
  NOR2_X1 U11178 ( .A1(n10044), .A2(n10033), .ZN(P1_U3298) );
  INV_X1 U11179 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U11180 ( .A1(n10044), .A2(n10034), .ZN(P1_U3299) );
  NOR2_X1 U11181 ( .A1(n10044), .A2(n10035), .ZN(P1_U3300) );
  NOR2_X1 U11182 ( .A1(n10044), .A2(n10036), .ZN(P1_U3301) );
  INV_X1 U11183 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U11184 ( .A1(n10044), .A2(n10037), .ZN(P1_U3302) );
  NOR2_X1 U11185 ( .A1(n10044), .A2(n10038), .ZN(P1_U3303) );
  NOR2_X1 U11186 ( .A1(n10044), .A2(n10039), .ZN(P1_U3304) );
  INV_X1 U11187 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U11188 ( .A1(n10044), .A2(n10040), .ZN(P1_U3305) );
  INV_X1 U11189 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U11190 ( .A1(n10044), .A2(n10041), .ZN(P1_U3306) );
  NOR2_X1 U11191 ( .A1(n10044), .A2(n10042), .ZN(P1_U3307) );
  INV_X1 U11192 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U11193 ( .A1(n10044), .A2(n10043), .ZN(P1_U3308) );
  NOR2_X1 U11194 ( .A1(n10060), .A2(n10045), .ZN(P1_U3309) );
  INV_X1 U11195 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U11196 ( .A1(n10060), .A2(n10046), .ZN(P1_U3310) );
  INV_X1 U11197 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U11198 ( .A1(n10060), .A2(n10047), .ZN(P1_U3311) );
  INV_X1 U11199 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U11200 ( .A1(n10060), .A2(n10048), .ZN(P1_U3312) );
  INV_X1 U11201 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U11202 ( .A1(n10060), .A2(n10049), .ZN(P1_U3313) );
  NOR2_X1 U11203 ( .A1(n10060), .A2(n10050), .ZN(P1_U3314) );
  INV_X1 U11204 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U11205 ( .A1(n10060), .A2(n10051), .ZN(P1_U3315) );
  INV_X1 U11206 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U11207 ( .A1(n10060), .A2(n10052), .ZN(P1_U3316) );
  NOR2_X1 U11208 ( .A1(n10060), .A2(n10053), .ZN(P1_U3317) );
  INV_X1 U11209 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U11210 ( .A1(n10060), .A2(n10054), .ZN(P1_U3318) );
  INV_X1 U11211 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U11212 ( .A1(n10060), .A2(n10055), .ZN(P1_U3319) );
  INV_X1 U11213 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U11214 ( .A1(n10060), .A2(n10056), .ZN(P1_U3320) );
  INV_X1 U11215 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U11216 ( .A1(n10060), .A2(n10057), .ZN(P1_U3321) );
  INV_X1 U11217 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U11218 ( .A1(n10060), .A2(n10058), .ZN(P1_U3322) );
  NOR2_X1 U11219 ( .A1(n10060), .A2(n10059), .ZN(P1_U3323) );
  OAI21_X1 U11220 ( .B1(n10062), .B2(n10095), .A(n10061), .ZN(n10064) );
  AOI211_X1 U11221 ( .C1(n10084), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10102) );
  AOI22_X1 U11222 ( .A1(n10101), .A2(n10102), .B1(n5118), .B2(n10099), .ZN(
        P1_U3456) );
  OAI21_X1 U11223 ( .B1(n10067), .B2(n10095), .A(n10066), .ZN(n10070) );
  INV_X1 U11224 ( .A(n10068), .ZN(n10069) );
  AOI211_X1 U11225 ( .C1(n6629), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        n10104) );
  AOI22_X1 U11226 ( .A1(n10101), .A2(n10104), .B1(n5151), .B2(n10099), .ZN(
        P1_U3462) );
  OAI21_X1 U11227 ( .B1(n10073), .B2(n10095), .A(n10072), .ZN(n10075) );
  AOI211_X1 U11228 ( .C1(n10084), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10106) );
  INV_X1 U11229 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U11230 ( .A1(n10101), .A2(n10106), .B1(n10077), .B2(n10099), .ZN(
        P1_U3474) );
  OAI21_X1 U11231 ( .B1(n10079), .B2(n10095), .A(n10078), .ZN(n10082) );
  INV_X1 U11232 ( .A(n10080), .ZN(n10081) );
  AOI211_X1 U11233 ( .C1(n10084), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10107) );
  INV_X1 U11234 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11235 ( .A1(n10101), .A2(n10107), .B1(n10085), .B2(n10099), .ZN(
        P1_U3486) );
  OAI21_X1 U11236 ( .B1(n10087), .B2(n10095), .A(n10086), .ZN(n10088) );
  AOI211_X1 U11237 ( .C1(n10090), .C2(n6629), .A(n10089), .B(n10088), .ZN(
        n10109) );
  INV_X1 U11238 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U11239 ( .A1(n10101), .A2(n10109), .B1(n10091), .B2(n10099), .ZN(
        P1_U3489) );
  INV_X1 U11240 ( .A(n10092), .ZN(n10098) );
  OAI211_X1 U11241 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10097) );
  AOI21_X1 U11242 ( .B1(n10098), .B2(n6629), .A(n10097), .ZN(n10112) );
  AOI22_X1 U11243 ( .A1(n10101), .A2(n10112), .B1(n10100), .B2(n10099), .ZN(
        P1_U3492) );
  AOI22_X1 U11244 ( .A1(n10113), .A2(n10102), .B1(n9220), .B2(n10110), .ZN(
        P1_U3523) );
  AOI22_X1 U11245 ( .A1(n10113), .A2(n10104), .B1(n10103), .B2(n10110), .ZN(
        P1_U3525) );
  AOI22_X1 U11246 ( .A1(n10113), .A2(n10106), .B1(n10105), .B2(n10110), .ZN(
        P1_U3529) );
  AOI22_X1 U11247 ( .A1(n10113), .A2(n10107), .B1(n7353), .B2(n10110), .ZN(
        P1_U3533) );
  AOI22_X1 U11248 ( .A1(n10113), .A2(n10109), .B1(n10108), .B2(n10110), .ZN(
        P1_U3534) );
  AOI22_X1 U11249 ( .A1(n10113), .A2(n10112), .B1(n10111), .B2(n10110), .ZN(
        P1_U3535) );
  XNOR2_X1 U11250 ( .A(n10115), .B(n10114), .ZN(n10123) );
  AND2_X1 U11251 ( .A1(n10116), .A2(n10319), .ZN(n10118) );
  OAI21_X1 U11252 ( .B1(n10119), .B2(n10118), .A(n10117), .ZN(n10122) );
  INV_X1 U11253 ( .A(n10120), .ZN(n10121) );
  OAI211_X1 U11254 ( .C1(n10123), .C2(n10227), .A(n10122), .B(n10121), .ZN(
        n10130) );
  AOI21_X1 U11255 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(n10128) );
  NOR2_X1 U11256 ( .A1(n10128), .A2(n10127), .ZN(n10129) );
  AOI211_X1 U11257 ( .C1(n10219), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10132) );
  OAI21_X1 U11258 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(P2_U3185) );
  AOI22_X1 U11259 ( .A1(n10220), .A2(P2_ADDR_REG_10__SCAN_IN), .B1(n10219), 
        .B2(n10135), .ZN(n10152) );
  OAI21_X1 U11260 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(n10143) );
  OAI21_X1 U11261 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10142) );
  AOI22_X1 U11262 ( .A1(n10143), .A2(n10237), .B1(n10209), .B2(n10142), .ZN(
        n10151) );
  INV_X1 U11263 ( .A(n10144), .ZN(n10150) );
  AOI21_X1 U11264 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(n10148) );
  OR2_X1 U11265 ( .A1(n10148), .A2(n10232), .ZN(n10149) );
  NAND4_X1 U11266 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        P2_U3192) );
  AOI22_X1 U11267 ( .A1(n10220), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10219), 
        .B2(n10153), .ZN(n10167) );
  OAI21_X1 U11268 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n10155), .A(n10154), 
        .ZN(n10160) );
  OAI21_X1 U11269 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10159) );
  AOI22_X1 U11270 ( .A1(n10160), .A2(n10209), .B1(n10237), .B2(n10159), .ZN(
        n10166) );
  AOI21_X1 U11271 ( .B1(n10162), .B2(n5873), .A(n10161), .ZN(n10163) );
  OR2_X1 U11272 ( .A1(n10232), .A2(n10163), .ZN(n10164) );
  NAND4_X1 U11273 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        P2_U3193) );
  AOI22_X1 U11274 ( .A1(n10220), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n10219), 
        .B2(n10168), .ZN(n10184) );
  OAI21_X1 U11275 ( .B1(n10171), .B2(n10170), .A(n10169), .ZN(n10176) );
  OAI21_X1 U11276 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10175) );
  AOI22_X1 U11277 ( .A1(n10176), .A2(n10209), .B1(n10237), .B2(n10175), .ZN(
        n10183) );
  INV_X1 U11278 ( .A(n10177), .ZN(n10182) );
  AOI21_X1 U11279 ( .B1(n4458), .B2(n10179), .A(n10178), .ZN(n10180) );
  OR2_X1 U11280 ( .A1(n10180), .A2(n10232), .ZN(n10181) );
  NAND4_X1 U11281 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        P2_U3194) );
  AOI22_X1 U11282 ( .A1(n10220), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(n10219), 
        .B2(n10185), .ZN(n10200) );
  OAI21_X1 U11283 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n10187), .A(n10186), 
        .ZN(n10192) );
  OAI21_X1 U11284 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(n10191) );
  AOI22_X1 U11285 ( .A1(n10192), .A2(n10209), .B1(n10237), .B2(n10191), .ZN(
        n10199) );
  AOI21_X1 U11286 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10196) );
  OR2_X1 U11287 ( .A1(n10232), .A2(n10196), .ZN(n10197) );
  NAND4_X1 U11288 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        P2_U3195) );
  AOI22_X1 U11289 ( .A1(n10220), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n10219), 
        .B2(n10202), .ZN(n10217) );
  OAI21_X1 U11290 ( .B1(n10202), .B2(n5913), .A(n10201), .ZN(n10203) );
  XOR2_X1 U11291 ( .A(n10204), .B(n10203), .Z(n10210) );
  OAI21_X1 U11292 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10208) );
  AOI22_X1 U11293 ( .A1(n10210), .A2(n10209), .B1(n10237), .B2(n10208), .ZN(
        n10216) );
  NAND2_X1 U11294 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10215)
         );
  AOI21_X1 U11295 ( .B1(n4463), .B2(n10212), .A(n10211), .ZN(n10213) );
  OR2_X1 U11296 ( .A1(n10213), .A2(n10232), .ZN(n10214) );
  NAND4_X1 U11297 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        P2_U3196) );
  AOI22_X1 U11298 ( .A1(n10220), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n10219), 
        .B2(n10218), .ZN(n10239) );
  OAI21_X1 U11299 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(n10236) );
  AOI21_X1 U11300 ( .B1(n10226), .B2(n10225), .A(n10224), .ZN(n10228) );
  NOR2_X1 U11301 ( .A1(n10228), .A2(n10227), .ZN(n10235) );
  AOI21_X1 U11302 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(n10233) );
  NOR2_X1 U11303 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  OAI211_X1 U11304 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10240), .A(n10239), .B(
        n10238), .ZN(P2_U3199) );
  XNOR2_X1 U11305 ( .A(n10241), .B(n8148), .ZN(n10251) );
  OAI21_X1 U11306 ( .B1(n10243), .B2(n8148), .A(n10242), .ZN(n10253) );
  INV_X1 U11307 ( .A(n10244), .ZN(n10245) );
  NAND2_X1 U11308 ( .A1(n10253), .A2(n10245), .ZN(n10250) );
  AOI22_X1 U11309 ( .A1(n6687), .A2(n10248), .B1(n10247), .B2(n10246), .ZN(
        n10249) );
  OAI211_X1 U11310 ( .C1(n10252), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        n10263) );
  INV_X1 U11311 ( .A(n10253), .ZN(n10261) );
  OAI22_X1 U11312 ( .A1(n10261), .A2(n10255), .B1(n5757), .B2(n10254), .ZN(
        n10256) );
  AOI211_X1 U11313 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n10257), .A(n10263), .B(
        n10256), .ZN(n10258) );
  AOI22_X1 U11314 ( .A1(n10260), .A2(n10259), .B1(n10258), .B2(n8714), .ZN(
        P2_U3231) );
  INV_X1 U11315 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10264) );
  OAI22_X1 U11316 ( .A1(n10261), .A2(n10292), .B1(n5757), .B2(n10303), .ZN(
        n10262) );
  NOR2_X1 U11317 ( .A1(n10263), .A2(n10262), .ZN(n10318) );
  AOI22_X1 U11318 ( .A1(n10317), .A2(n10264), .B1(n10318), .B2(n10315), .ZN(
        P2_U3396) );
  INV_X1 U11319 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U11320 ( .A1(n10266), .A2(n10306), .B1(n10314), .B2(n10265), .ZN(
        n10267) );
  AND2_X1 U11321 ( .A1(n10268), .A2(n10267), .ZN(n10320) );
  AOI22_X1 U11322 ( .A1(n10317), .A2(n10269), .B1(n10320), .B2(n10315), .ZN(
        P2_U3399) );
  INV_X1 U11323 ( .A(n10270), .ZN(n10274) );
  OAI22_X1 U11324 ( .A1(n10272), .A2(n10309), .B1(n10271), .B2(n10303), .ZN(
        n10273) );
  NOR2_X1 U11325 ( .A1(n10274), .A2(n10273), .ZN(n10322) );
  AOI22_X1 U11326 ( .A1(n10317), .A2(n9677), .B1(n10322), .B2(n10315), .ZN(
        P2_U3402) );
  INV_X1 U11327 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10280) );
  INV_X1 U11328 ( .A(n10275), .ZN(n10279) );
  OAI21_X1 U11329 ( .B1(n10277), .B2(n10303), .A(n10276), .ZN(n10278) );
  AOI21_X1 U11330 ( .B1(n10279), .B2(n10306), .A(n10278), .ZN(n10324) );
  AOI22_X1 U11331 ( .A1(n10317), .A2(n10280), .B1(n10324), .B2(n10315), .ZN(
        P2_U3405) );
  INV_X1 U11332 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10285) );
  OAI22_X1 U11333 ( .A1(n10282), .A2(n10309), .B1(n10281), .B2(n10303), .ZN(
        n10283) );
  NOR2_X1 U11334 ( .A1(n10284), .A2(n10283), .ZN(n10326) );
  AOI22_X1 U11335 ( .A1(n10317), .A2(n10285), .B1(n10326), .B2(n10315), .ZN(
        P2_U3408) );
  INV_X1 U11336 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10290) );
  NOR2_X1 U11337 ( .A1(n10286), .A2(n10303), .ZN(n10288) );
  AOI211_X1 U11338 ( .C1(n10306), .C2(n10289), .A(n10288), .B(n10287), .ZN(
        n10328) );
  AOI22_X1 U11339 ( .A1(n10317), .A2(n10290), .B1(n10328), .B2(n10315), .ZN(
        P2_U3414) );
  INV_X1 U11340 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10296) );
  OAI22_X1 U11341 ( .A1(n10293), .A2(n10292), .B1(n10291), .B2(n10303), .ZN(
        n10294) );
  NOR2_X1 U11342 ( .A1(n10295), .A2(n10294), .ZN(n10329) );
  AOI22_X1 U11343 ( .A1(n10317), .A2(n10296), .B1(n10329), .B2(n10315), .ZN(
        P2_U3417) );
  INV_X1 U11344 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10301) );
  OAI22_X1 U11345 ( .A1(n10298), .A2(n10309), .B1(n4403), .B2(n10303), .ZN(
        n10299) );
  NOR2_X1 U11346 ( .A1(n10300), .A2(n10299), .ZN(n10330) );
  AOI22_X1 U11347 ( .A1(n10317), .A2(n10301), .B1(n10330), .B2(n10315), .ZN(
        P2_U3420) );
  INV_X1 U11348 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10308) );
  OAI21_X1 U11349 ( .B1(n10304), .B2(n10303), .A(n10302), .ZN(n10305) );
  AOI21_X1 U11350 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(n10331) );
  AOI22_X1 U11351 ( .A1(n10317), .A2(n10308), .B1(n10331), .B2(n10315), .ZN(
        P2_U3423) );
  INV_X1 U11352 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U11353 ( .A1(n10310), .A2(n10309), .ZN(n10312) );
  AOI211_X1 U11354 ( .C1(n10314), .C2(n10313), .A(n10312), .B(n10311), .ZN(
        n10332) );
  AOI22_X1 U11355 ( .A1(n10317), .A2(n10316), .B1(n10332), .B2(n10315), .ZN(
        P2_U3426) );
  AOI22_X1 U11356 ( .A1(n10333), .A2(n10318), .B1(n6500), .B2(n6673), .ZN(
        P2_U3461) );
  AOI22_X1 U11357 ( .A1(n10333), .A2(n10320), .B1(n10319), .B2(n6673), .ZN(
        P2_U3462) );
  AOI22_X1 U11358 ( .A1(n10333), .A2(n10322), .B1(n10321), .B2(n6673), .ZN(
        P2_U3463) );
  INV_X1 U11359 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U11360 ( .A1(n10333), .A2(n10324), .B1(n10323), .B2(n6673), .ZN(
        P2_U3464) );
  AOI22_X1 U11361 ( .A1(n10333), .A2(n10326), .B1(n10325), .B2(n6673), .ZN(
        P2_U3465) );
  INV_X1 U11362 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U11363 ( .A1(n10333), .A2(n10328), .B1(n10327), .B2(n6673), .ZN(
        P2_U3467) );
  AOI22_X1 U11364 ( .A1(n10333), .A2(n10329), .B1(n6592), .B2(n6673), .ZN(
        P2_U3468) );
  AOI22_X1 U11365 ( .A1(n10333), .A2(n10330), .B1(n5855), .B2(n6673), .ZN(
        P2_U3469) );
  AOI22_X1 U11366 ( .A1(n10333), .A2(n10331), .B1(n5873), .B2(n6673), .ZN(
        P2_U3470) );
  AOI22_X1 U11367 ( .A1(n10333), .A2(n10332), .B1(n6519), .B2(n6673), .ZN(
        P2_U3471) );
  NOR2_X1 U11368 ( .A1(n10335), .A2(n10334), .ZN(n10337) );
  XNOR2_X1 U11369 ( .A(n10337), .B(n10336), .ZN(ADD_1068_U5) );
  XOR2_X1 U11370 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11371 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  XOR2_X1 U11372 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10340), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11373 ( .A(n10342), .B(n10341), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11374 ( .A(n10344), .B(n10343), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11375 ( .A(n10346), .B(n10345), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11376 ( .A(n10348), .B(n10347), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11377 ( .A(n10350), .B(n10349), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11378 ( .A(n10352), .B(n10351), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11379 ( .A(n10354), .B(n10353), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11380 ( .A(n10356), .B(n10355), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11381 ( .A(n10358), .B(n10357), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11382 ( .A(n10360), .B(n10359), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11383 ( .A(n10362), .B(n10361), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11384 ( .A(n10364), .B(n10363), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11385 ( .A(n10366), .B(n10365), .ZN(ADD_1068_U48) );
  XOR2_X1 U11386 ( .A(n10368), .B(n10367), .Z(ADD_1068_U54) );
  XOR2_X1 U11387 ( .A(n10370), .B(n10369), .Z(ADD_1068_U53) );
  XNOR2_X1 U11388 ( .A(n10372), .B(n10371), .ZN(ADD_1068_U52) );
  INV_X2 U4907 ( .A(n6395), .ZN(n6388) );
  AND2_X1 U7739 ( .A1(n8364), .A2(n8184), .ZN(n8354) );
  INV_X1 U4905 ( .A(n8354), .ZN(n8349) );
  INV_X2 U5959 ( .A(n10260), .ZN(n8714) );
endmodule

